module sparc_mul_top ( mul_exu_ack, mul_spu_ack, mul_spu_shf_ack, mul_data_out, 
        so, rclk, grst_l, arst_l, exu_mul_input_vld, exu_mul_rs1_data, 
        exu_mul_rs2_data, spu_mul_req_vld, spu_mul_acc, spu_mul_areg_shf, 
        spu_mul_areg_rst, spu_mul_op1_data, spu_mul_op2_data, 
        spu_mul_mulres_lshft, si, se );
  output [63:0] mul_data_out;
  input [63:0] exu_mul_rs1_data;
  input [63:0] exu_mul_rs2_data;
  input [63:0] spu_mul_op1_data;
  input [63:0] spu_mul_op2_data;
  input rclk, grst_l, arst_l, exu_mul_input_vld, spu_mul_req_vld, spu_mul_acc,
         spu_mul_areg_shf, spu_mul_areg_rst, spu_mul_mulres_lshft, si, se;
  output mul_exu_ack, mul_spu_ack, mul_spu_shf_ack, so;
  wire   n18338, n18339, rst_l, c0_act, byp_sel, byp_imm, acc_imm, acc_actc2,
         acc_actc3, acc_reg_enb, acc_reg_rst, acc_reg_shf, x2, rstff_n4 ,
         control_n25 , control_n24 , control_n23 , control_n22 ,
         control_n21 , control_n20 , control_n19 , control_n18 ,
         control_n17 , control_n16 , control_n15 , control_n14 ,
         control_n13 , control_n12 , control_n11 , control_n10 ,
         control_n9 , control_n8 , control_n7 , control_N11 ,
         control_N10 , control_N9 , control_N8 , control_N7 , control_N6 ,
         control_acc_actc1 , control_N5 , control_mul_ecl_ack_d ,
         control_mul_spu_ack_d , control_c3_act , control_N4 ,
         control_c2_act , control_N3 , control_N2 , control_favor_e ,
         control_acc_actc4 , control_c1_act , dpath_n1128 , dpath_n1127 ,
         dpath_n1126 , dpath_n1125 , dpath_n1124 , dpath_n1123 ,
         dpath_n1122 , dpath_n1121 , dpath_n1120 , dpath_n1119 ,
         dpath_n1118 , dpath_n1117 , dpath_n1116 , dpath_n1115 ,
         dpath_n1114 , dpath_n1113 , dpath_n1112 , dpath_n1111 ,
         dpath_n1110 , dpath_n1109 , dpath_n1108 , dpath_n1107 ,
         dpath_n1106 , dpath_n1105 , dpath_n1104 , dpath_n1103 ,
         dpath_n1102 , dpath_n1101 , dpath_n1100 , dpath_n1099 ,
         dpath_n1098 , dpath_n1097 , dpath_n1096 , dpath_n1095 ,
         dpath_n1094 , dpath_n1093 , dpath_n1092 , dpath_n1091 ,
         dpath_n1090 , dpath_n1089 , dpath_n1088 , dpath_n1087 ,
         dpath_n1086 , dpath_n1085 , dpath_n1084 , dpath_n1083 ,
         dpath_n1082 , dpath_n1081 , dpath_n1080 , dpath_n1079 ,
         dpath_n1078 , dpath_n1077 , dpath_n1076 , dpath_n1075 ,
         dpath_n1074 , dpath_n1073 , dpath_n1072 , dpath_n1071 ,
         dpath_n1070 , dpath_n1069 , dpath_n1068 , dpath_n1067 ,
         dpath_n1066 , dpath_n1065 , dpath_n1064 , dpath_n1063 ,
         dpath_n1062 , dpath_n1061 , dpath_n1060 , dpath_n1059 ,
         dpath_n1058 , dpath_n1057 , dpath_n1056 , dpath_n1055 ,
         dpath_n1054 , dpath_n1053 , dpath_n1052 , dpath_n1051 ,
         dpath_n1050 , dpath_n1049 , dpath_n1048 , dpath_n1047 ,
         dpath_n1046 , dpath_n1045 , dpath_n1044 , dpath_n1043 ,
         dpath_n1042 , dpath_n1041 , dpath_n1040 , dpath_n1039 ,
         dpath_n1038 , dpath_n1037 , dpath_n1036 , dpath_n1035 ,
         dpath_n1034 , dpath_n1033 , dpath_n1032 , dpath_n1031 ,
         dpath_n1030 , dpath_n1029 , dpath_n1028 , dpath_n1027 ,
         dpath_n1026 , dpath_n1025 , dpath_n1024 , dpath_n1023 ,
         dpath_n1022 , dpath_n1021 , dpath_n1020 , dpath_n1019 ,
         dpath_n1018 , dpath_n1017 , dpath_n1016 , dpath_n1015 ,
         dpath_n1014 , dpath_n1013 , dpath_n1012 , dpath_n1011 ,
         dpath_n1010 , dpath_n1009 , dpath_n1008 , dpath_n1007 ,
         dpath_n1006 , dpath_n1005 , dpath_n1004 , dpath_n1003 ,
         dpath_n1002 , dpath_n1001 , dpath_n1000 , dpath_n999 ,
         dpath_n998 , dpath_n997 , dpath_n996 , dpath_n995 , dpath_n994 ,
         dpath_n993 , dpath_n992 , dpath_n991 , dpath_n990 , dpath_n989 ,
         dpath_n988 , dpath_n987 , dpath_n986 , dpath_n985 , dpath_n984 ,
         dpath_n983 , dpath_n982 , dpath_n981 , dpath_n980 , dpath_n979 ,
         dpath_n978 , dpath_n977 , dpath_n976 , dpath_n975 , dpath_n974 ,
         dpath_n973 , dpath_n972 , dpath_n971 , dpath_n970 , dpath_n969 ,
         dpath_n968 , dpath_n967 , dpath_n966 , dpath_n965 , dpath_n964 ,
         dpath_n963 , dpath_n962 , dpath_n961 , dpath_n960 , dpath_n959 ,
         dpath_n958 , dpath_n957 , dpath_n956 , dpath_n955 , dpath_n954 ,
         dpath_n953 , dpath_n952 , dpath_n951 , dpath_n950 , dpath_n949 ,
         dpath_n948 , dpath_n947 , dpath_n946 , dpath_n945 , dpath_n944 ,
         dpath_n943 , dpath_n942 , dpath_n941 , dpath_n940 , dpath_n939 ,
         dpath_n938 , dpath_n937 , dpath_n936 , dpath_n935 , dpath_n934 ,
         dpath_n933 , dpath_n932 , dpath_n931 , dpath_n930 , dpath_n929 ,
         dpath_n928 , dpath_n927 , dpath_n926 , dpath_n925 , dpath_n924 ,
         dpath_n923 , dpath_n922 , dpath_n921 , dpath_n920 , dpath_n919 ,
         dpath_n918 , dpath_n917 , dpath_n916 , dpath_n915 , dpath_n914 ,
         dpath_n913 , dpath_n912 , dpath_n911 , dpath_n910 , dpath_n909 ,
         dpath_n908 , dpath_n907 , dpath_n906 , dpath_n905 , dpath_n904 ,
         dpath_n903 , dpath_n902 , dpath_n901 , dpath_n900 , dpath_n899 ,
         dpath_n898 , dpath_n897 , dpath_n896 , dpath_n895 , dpath_n894 ,
         dpath_n893 , dpath_n892 , dpath_n891 , dpath_n890 , dpath_n889 ,
         dpath_n888 , dpath_n887 , dpath_n886 , dpath_n885 , dpath_n884 ,
         dpath_n883 , dpath_n882 , dpath_n881 , dpath_n880 , dpath_n879 ,
         dpath_n878 , dpath_n877 , dpath_n876 , dpath_n875 , dpath_n874 ,
         dpath_n873 , dpath_n872 , dpath_n871 , dpath_n870 , dpath_n869 ,
         dpath_n868 , dpath_n867 , dpath_n866 , dpath_n865 , dpath_n864 ,
         dpath_n863 , dpath_n862 , dpath_n861 , dpath_n860 , dpath_n859 ,
         dpath_n858 , dpath_n857 , dpath_n856 , dpath_n855 , dpath_n854 ,
         dpath_n853 , dpath_n852 , dpath_n851 , dpath_n850 , dpath_n849 ,
         dpath_n848 , dpath_n847 , dpath_n846 , dpath_n845 , dpath_n844 ,
         dpath_n843 , dpath_n842 , dpath_n841 , dpath_n840 , dpath_n839 ,
         dpath_n838 , dpath_n837 , dpath_n836 , dpath_n835 , dpath_n834 ,
         dpath_n833 , dpath_n832 , dpath_n831 , dpath_n830 , dpath_n829 ,
         dpath_n828 , dpath_n827 , dpath_n826 , dpath_n825 , dpath_n824 ,
         dpath_n823 , dpath_n822 , dpath_n821 , dpath_n820 , dpath_n819 ,
         dpath_n818 , dpath_n817 , dpath_n816 , dpath_n815 , dpath_n814 ,
         dpath_n813 , dpath_n812 , dpath_n811 , dpath_n810 , dpath_n809 ,
         dpath_n808 , dpath_n807 , dpath_n806 , dpath_n805 , dpath_n804 ,
         dpath_n803 , dpath_n802 , dpath_n801 , dpath_n800 , dpath_n799 ,
         dpath_n798 , dpath_n797 , dpath_n796 , dpath_n795 , dpath_n794 ,
         dpath_n793 , dpath_n792 , dpath_n791 , dpath_n790 , dpath_n789 ,
         dpath_n788 , dpath_n787 , dpath_n786 , dpath_n785 , dpath_n784 ,
         dpath_n783 , dpath_n782 , dpath_n781 , dpath_n780 , dpath_n779 ,
         dpath_n778 , dpath_n777 , dpath_n776 , dpath_n775 , dpath_n774 ,
         dpath_n773 , dpath_n772 , dpath_n771 , dpath_n770 , dpath_n769 ,
         dpath_n768 , dpath_n767 , dpath_n766 , dpath_n765 , dpath_n764 ,
         dpath_n763 , dpath_n762 , dpath_n761 , dpath_n760 , dpath_n759 ,
         dpath_n758 , dpath_n757 , dpath_n756 , dpath_n755 , dpath_n754 ,
         dpath_n753 , dpath_n752 , dpath_n751 , dpath_n750 , dpath_n749 ,
         dpath_n748 , dpath_n747 , dpath_n746 , dpath_n745 , dpath_n744 ,
         dpath_n743 , dpath_n742 , dpath_n741 , dpath_n740 , dpath_n739 ,
         dpath_n738 , dpath_n737 , dpath_n736 , dpath_n735 , dpath_n734 ,
         dpath_n733 , dpath_n732 , dpath_n731 , dpath_n730 , dpath_n729 ,
         dpath_n728 , dpath_n727 , dpath_n726 , dpath_n725 , dpath_n724 ,
         dpath_n723 , dpath_n722 , dpath_n721 , dpath_n720 , dpath_n719 ,
         dpath_n718 , dpath_n717 , dpath_n716 , dpath_n715 , dpath_n714 ,
         dpath_n713 , dpath_n712 , dpath_n711 , dpath_n710 , dpath_n709 ,
         dpath_n708 , dpath_n707 , dpath_n706 , dpath_n705 , dpath_n704 ,
         dpath_n703 , dpath_n702 , dpath_n701 , dpath_n700 , dpath_n699 ,
         dpath_n698 , dpath_n697 , dpath_n696 , dpath_n695 , dpath_n694 ,
         dpath_n693 , dpath_n692 , dpath_n691 , dpath_n690 , dpath_n689 ,
         dpath_n688 , dpath_n687 , dpath_n686 , dpath_n685 , dpath_n684 ,
         dpath_n683 , dpath_n682 , dpath_n681 , dpath_n680 , dpath_n679 ,
         dpath_n678 , dpath_n677 , dpath_n676 , dpath_n675 , dpath_n674 ,
         dpath_n673 , dpath_n672 , dpath_n671 , dpath_n670 , dpath_n669 ,
         dpath_n668 , dpath_n667 , dpath_n666 , dpath_n665 , dpath_n664 ,
         dpath_n663 , dpath_n662 , dpath_n661 , dpath_n660 , dpath_n659 ,
         dpath_n658 , dpath_n657 , dpath_n656 , dpath_n655 , dpath_n654 ,
         dpath_n653 , dpath_n652 , dpath_n651 , dpath_n650 , dpath_n649 ,
         dpath_n648 , dpath_n647 , dpath_n646 , dpath_n645 , dpath_n644 ,
         dpath_n643 , dpath_n642 , dpath_n641 , dpath_n640 , dpath_n639 ,
         dpath_n638 , dpath_n637 , dpath_n636 , dpath_n635 , dpath_n634 ,
         dpath_n633 , dpath_n632 , dpath_n631 , dpath_n630 , dpath_n629 ,
         dpath_n628 , dpath_n627 , dpath_n626 , dpath_n625 , dpath_n624 ,
         dpath_n623 , dpath_n622 , dpath_n621 , dpath_n620 , dpath_n619 ,
         dpath_n618 , dpath_n617 , dpath_n616 , dpath_n615 , dpath_n614 ,
         dpath_n613 , dpath_n612 , dpath_n611 , dpath_n610 , dpath_n609 ,
         dpath_n608 , dpath_n607 , dpath_n606 , dpath_n605 , dpath_n604 ,
         dpath_n603 , dpath_n602 , dpath_n601 , dpath_n600 , dpath_n599 ,
         dpath_n598 , dpath_n597 , dpath_n596 , dpath_n595 , dpath_n594 ,
         dpath_n593 , dpath_n592 , dpath_n591 , dpath_n590 , dpath_n589 ,
         dpath_n588 , dpath_n587 , dpath_n586 , dpath_n585 , dpath_n584 ,
         dpath_n583 , dpath_n582 , dpath_n581 , dpath_n580 , dpath_n579 ,
         dpath_n578 , dpath_n577 , dpath_n576 , dpath_n575 , dpath_n574 ,
         dpath_n573 , dpath_n572 , dpath_n571 , dpath_n570 , dpath_n569 ,
         dpath_n568 , dpath_n567 , dpath_n566 , dpath_n565 , dpath_n564 ,
         dpath_n563 , dpath_n562 , dpath_n561 , dpath_n560 , dpath_n559 ,
         dpath_n558 , dpath_n557 , dpath_n556 , dpath_n555 , dpath_n554 ,
         dpath_n553 , dpath_n552 , dpath_n551 , dpath_n550 , dpath_n549 ,
         dpath_n548 , dpath_n547 , dpath_n546 , dpath_n545 , dpath_n544 ,
         dpath_n543 , dpath_n542 , dpath_n541 , dpath_n540 , dpath_n539 ,
         dpath_n538 , dpath_n537 , dpath_n536 , dpath_n535 , dpath_n534 ,
         dpath_n533 , dpath_n532 , dpath_n531 , dpath_n530 , dpath_n529 ,
         dpath_n528 , dpath_n527 , dpath_n526 , dpath_n525 , dpath_n524 ,
         dpath_n523 , dpath_n522 , dpath_n521 , dpath_n520 , dpath_n519 ,
         dpath_n518 , dpath_n517 , dpath_n516 , dpath_n515 , dpath_n514 ,
         dpath_n513 , dpath_n512 , dpath_n511 , dpath_n510 , dpath_n509 ,
         dpath_n508 , dpath_n507 , dpath_n506 , dpath_n505 , dpath_n504 ,
         dpath_n503 , dpath_n502 , dpath_n501 , dpath_n500 , dpath_n499 ,
         dpath_n498 , dpath_n497 , dpath_n496 , dpath_n495 , dpath_n494 ,
         dpath_n493 , dpath_n492 , dpath_n491 , dpath_n490 , dpath_n489 ,
         dpath_n488 , dpath_n487 , dpath_n486 , dpath_n485 , dpath_n484 ,
         dpath_n483 , dpath_n482 , dpath_n481 , dpath_n480 , dpath_n479 ,
         dpath_n478 , dpath_n477 , dpath_n476 , dpath_n475 , dpath_n474 ,
         dpath_n473 , dpath_n472 , dpath_n471 , dpath_n470 , dpath_n469 ,
         dpath_n468 , dpath_n467 , dpath_n466 , dpath_n465 , dpath_n464 ,
         dpath_n463 , dpath_n462 , dpath_n461 , dpath_n460 , dpath_n459 ,
         dpath_n458 , dpath_n457 , dpath_n456 , dpath_n455 , dpath_n454 ,
         dpath_n453 , dpath_n452 , dpath_n451 , dpath_n450 , dpath_n449 ,
         dpath_n448 , dpath_n447 , dpath_n446 , dpath_n445 , dpath_n444 ,
         dpath_n443 , dpath_n442 , dpath_n441 , dpath_n440 , dpath_n439 ,
         dpath_n438 , dpath_n437 , dpath_n436 , dpath_n435 , dpath_n434 ,
         dpath_n433 , dpath_n432 , dpath_n431 , dpath_n430 , dpath_n429 ,
         dpath_n428 , dpath_n427 , dpath_n426 , dpath_n425 , dpath_n424 ,
         dpath_n423 , dpath_n422 , dpath_n421 , dpath_n420 , dpath_n419 ,
         dpath_n418 , dpath_n417 , dpath_n416 , dpath_n415 , dpath_n414 ,
         dpath_n413 , dpath_n412 , dpath_n411 , dpath_n410 , dpath_n409 ,
         dpath_n408 , dpath_n407 , dpath_n406 , dpath_n405 , dpath_n404 ,
         dpath_n403 , dpath_n402 , dpath_n401 , dpath_n400 , dpath_n399 ,
         dpath_n398 , dpath_n397 , dpath_n396 , dpath_n395 , dpath_n394 ,
         dpath_n393 , dpath_n392 , dpath_n391 , dpath_n390 , dpath_n389 ,
         dpath_n388 , dpath_n387 , dpath_n386 , dpath_n385 , dpath_n384 ,
         dpath_n383 , dpath_n382 , dpath_n381 , dpath_n380 , dpath_n379 ,
         dpath_n378 , dpath_n377 , dpath_n376 , dpath_n375 , dpath_n374 ,
         dpath_n373 , dpath_n372 , dpath_n371 , dpath_n370 , dpath_n369 ,
         dpath_n368 , dpath_n367 , dpath_n366 , dpath_n365 , dpath_n364 ,
         dpath_n363 , dpath_n362 , dpath_n361 , dpath_n360 , dpath_n359 ,
         dpath_n358 , dpath_n357 , dpath_n356 , dpath_n355 , dpath_n354 ,
         dpath_n353 , dpath_n352 , dpath_n351 , dpath_n350 , dpath_n349 ,
         dpath_n348 , dpath_n347 , dpath_n346 , dpath_n345 , dpath_n344 ,
         dpath_n343 , dpath_n342 , dpath_n341 , dpath_n340 , dpath_n339 ,
         dpath_n338 , dpath_n337 , dpath_n336 , dpath_n335 , dpath_n334 ,
         dpath_n333 , dpath_n332 , dpath_n331 , dpath_n330 , dpath_n329 ,
         dpath_n328 , dpath_n327 , dpath_n326 , dpath_n325 , dpath_n324 ,
         dpath_n323 , dpath_n322 , dpath_n321 , dpath_n320 , dpath_n319 ,
         dpath_n318 , dpath_n317 , dpath_n316 , dpath_n315 , dpath_n314 ,
         dpath_n313 , dpath_n312 , dpath_n311 , dpath_n310 , dpath_n309 ,
         dpath_n308 , dpath_n307 , dpath_n306 , dpath_n305 , dpath_n304 ,
         dpath_n303 , dpath_n302 , dpath_n301 , dpath_n300 , dpath_n299 ,
         dpath_n298 , dpath_n297 , dpath_n296 , dpath_n295 , dpath_n294 ,
         dpath_n293 , dpath_n292 , dpath_n291 , dpath_n290 , dpath_n289 ,
         dpath_n288 , dpath_n287 , dpath_n286 , dpath_n285 , dpath_n284 ,
         dpath_n283 , dpath_n282 , dpath_n281 , dpath_n280 , dpath_n279 ,
         dpath_n278 , dpath_n277 , dpath_n276 , dpath_n275 , dpath_n274 ,
         dpath_n273 , dpath_n272 , dpath_n271 , dpath_n270 , dpath_n269 ,
         dpath_n268 , dpath_n267 , dpath_n266 , dpath_n265 , dpath_n264 ,
         dpath_n263 , dpath_n262 , dpath_n261 , dpath_n260 , dpath_n259 ,
         dpath_n258 , dpath_n257 , dpath_n256 , dpath_n255 , dpath_n254 ,
         dpath_n253 , dpath_n252 , dpath_n251 , dpath_n250 , dpath_n249 ,
         dpath_n248 , dpath_n247 , dpath_n246 , dpath_n245 , dpath_n244 ,
         dpath_n243 , dpath_n242 , dpath_n241 , dpath_n240 , dpath_n239 ,
         dpath_n238 , dpath_n237 , dpath_n236 , dpath_n235 , dpath_n234 ,
         dpath_n233 , dpath_n232 , dpath_n231 , dpath_n230 , dpath_n229 ,
         dpath_n228 , dpath_n227 , dpath_n226 , dpath_n225 , dpath_n224 ,
         dpath_n223 , dpath_n222 , dpath_n221 , dpath_n220 , dpath_n219 ,
         dpath_n218 , dpath_n217 , dpath_n216 , dpath_n215 , dpath_n214 ,
         dpath_n213 , dpath_n212 , dpath_n211 , dpath_n210 , dpath_n209 ,
         dpath_n208 , dpath_n207 , dpath_n206 , dpath_n205 , dpath_n204 ,
         dpath_n203 , dpath_n202 , dpath_n201 , dpath_n200 , dpath_n199 ,
         dpath_n198 , dpath_n197 , dpath_n196 , dpath_n195 , dpath_n194 ,
         dpath_n193 , dpath_n192 , dpath_n191 , dpath_n190 , dpath_n189 ,
         dpath_n188 , dpath_n187 , dpath_n186 , dpath_n185 , dpath_n184 ,
         dpath_n183 , dpath_n182 , dpath_n181 , dpath_n180 , dpath_n179 ,
         dpath_n178 , dpath_n177 , dpath_n176 , dpath_n175 , dpath_n174 ,
         dpath_n173 , dpath_n172 , dpath_n171 , dpath_n170 , dpath_n169 ,
         dpath_n168 , dpath_n167 , dpath_n166 , dpath_n165 , dpath_n164 ,
         dpath_n163 , dpath_n162 , dpath_n161 , dpath_n160 , dpath_n159 ,
         dpath_n158 , dpath_n157 , dpath_n156 , dpath_n155 , dpath_n154 ,
         dpath_n153 , dpath_n152 , dpath_n151 , dpath_n150 , dpath_n149 ,
         dpath_n148 , dpath_n147 , dpath_n146 , dpath_n145 , dpath_n144 ,
         dpath_n143 , dpath_n142 , dpath_n141 , dpath_n140 , dpath_n139 ,
         dpath_n138 , dpath_n137 , dpath_n136 , dpath_n135 , dpath_n134 ,
         dpath_n133 , dpath_n132 , dpath_n131 , dpath_n130 , dpath_n129 ,
         dpath_n128 , dpath_n127 , dpath_n126 , dpath_n125 , dpath_n124 ,
         dpath_n123 , dpath_n122 , dpath_n121 , dpath_n120 , dpath_n119 ,
         dpath_n118 , dpath_n117 , dpath_n116 , dpath_n115 , dpath_n114 ,
         dpath_n113 , dpath_n112 , dpath_n111 , dpath_n110 , dpath_n109 ,
         dpath_n108 , dpath_n107 , dpath_n106 , dpath_n105 , dpath_n104 ,
         dpath_n103 , dpath_n102 , dpath_n101 , dpath_n100 , dpath_n99 ,
         dpath_n98 , dpath_n97 , dpath_n96 , dpath_n95 , dpath_n94 ,
         dpath_n93 , dpath_n92 , dpath_n91 , dpath_n90 , dpath_n89 ,
         dpath_n88 , dpath_n87 , dpath_n86 , dpath_n85 , dpath_n84 ,
         dpath_n83 , dpath_n82 , dpath_n81 , dpath_n80 , dpath_n79 ,
         dpath_n78 , dpath_n77 , dpath_n76 , dpath_n75 , dpath_n74 ,
         dpath_n73 , dpath_n72 , dpath_n71 , dpath_n70 , dpath_n69 ,
         dpath_n68 , dpath_n67 , dpath_n66 , dpath_n65 , dpath_n64 ,
         dpath_n63 , dpath_n62 , dpath_n61 , dpath_n60 , dpath_n59 ,
         dpath_n58 , dpath_n57 , dpath_n56 , dpath_n55 , dpath_n54 ,
         dpath_n53 , dpath_n52 , dpath_n51 , dpath_n50 , dpath_n49 ,
         dpath_n48 , dpath_n47 , dpath_n46 , dpath_n45 , dpath_n44 ,
         dpath_n43 , dpath_n42 , dpath_n41 , dpath_n40 , dpath_n39 ,
         dpath_n38 , dpath_n37 , dpath_n36 , dpath_n35 , dpath_n34 ,
         dpath_n33 , dpath_n32 , dpath_n31 , dpath_n30 , dpath_n29 ,
         dpath_n28 , dpath_n27 , dpath_n26 , dpath_n25 , dpath_n24 ,
         dpath_n23 , dpath_n22 , dpath_n21 , dpath_n20 , dpath_n19 ,
         dpath_n18 , dpath_n17 , dpath_n16 , dpath_n15 , dpath_n14 ,
         dpath_n13 , dpath_n12 , dpath_n11 , dpath_n10 , dpath_n9 ,
         dpath_clk_enb1 , dpath_acc_reg_in[135] , dpath_acc_reg_in[134] ,
         dpath_acc_reg_in[133] , dpath_acc_reg_in[132] ,
         dpath_acc_reg_in[131] , dpath_acc_reg_in[130] ,
         dpath_acc_reg_in[129] , dpath_acc_reg_in[128] ,
         dpath_acc_reg_in[127] , dpath_acc_reg_in[126] ,
         dpath_acc_reg_in[125] , dpath_acc_reg_in[124] ,
         dpath_acc_reg_in[123] , dpath_acc_reg_in[122] ,
         dpath_acc_reg_in[121] , dpath_acc_reg_in[120] ,
         dpath_acc_reg_in[119] , dpath_acc_reg_in[118] ,
         dpath_acc_reg_in[117] , dpath_acc_reg_in[116] ,
         dpath_acc_reg_in[115] , dpath_acc_reg_in[114] ,
         dpath_acc_reg_in[113] , dpath_acc_reg_in[112] ,
         dpath_acc_reg_in[111] , dpath_acc_reg_in[110] ,
         dpath_acc_reg_in[109] , dpath_acc_reg_in[108] ,
         dpath_acc_reg_in[107] , dpath_acc_reg_in[106] ,
         dpath_acc_reg_in[105] , dpath_acc_reg_in[104] ,
         dpath_acc_reg_in[103] , dpath_acc_reg_in[102] ,
         dpath_acc_reg_in[101] , dpath_acc_reg_in[100] ,
         dpath_acc_reg_in[99] , dpath_acc_reg_in[98] ,
         dpath_acc_reg_in[97] , dpath_acc_reg_in[96] ,
         dpath_acc_reg_in[95] , dpath_acc_reg_in[94] ,
         dpath_acc_reg_in[93] , dpath_acc_reg_in[92] ,
         dpath_acc_reg_in[91] , dpath_acc_reg_in[90] ,
         dpath_acc_reg_in[89] , dpath_acc_reg_in[88] ,
         dpath_acc_reg_in[87] , dpath_acc_reg_in[86] ,
         dpath_acc_reg_in[85] , dpath_acc_reg_in[84] ,
         dpath_acc_reg_in[83] , dpath_acc_reg_in[82] ,
         dpath_acc_reg_in[81] , dpath_acc_reg_in[80] ,
         dpath_acc_reg_in[79] , dpath_acc_reg_in[78] ,
         dpath_acc_reg_in[77] , dpath_acc_reg_in[76] ,
         dpath_acc_reg_in[75] , dpath_acc_reg_in[74] ,
         dpath_acc_reg_in[73] , dpath_acc_reg_in[72] ,
         dpath_acc_reg_in[71] , dpath_acc_reg_in[70] ,
         dpath_acc_reg_in[69] , dpath_acc_reg_in[68] ,
         dpath_acc_reg_in[67] , dpath_acc_reg_in[66] ,
         dpath_acc_reg_in[65] , dpath_acc_reg_in[64] ,
         dpath_acc_reg_in[63] , dpath_acc_reg_in[62] ,
         dpath_acc_reg_in[61] , dpath_acc_reg_in[60] ,
         dpath_acc_reg_in[59] , dpath_acc_reg_in[58] ,
         dpath_acc_reg_in[57] , dpath_acc_reg_in[56] ,
         dpath_acc_reg_in[55] , dpath_acc_reg_in[54] ,
         dpath_acc_reg_in[53] , dpath_acc_reg_in[52] ,
         dpath_acc_reg_in[51] , dpath_acc_reg_in[50] ,
         dpath_acc_reg_in[49] , dpath_acc_reg_in[48] ,
         dpath_acc_reg_in[47] , dpath_acc_reg_in[46] ,
         dpath_acc_reg_in[45] , dpath_acc_reg_in[44] ,
         dpath_acc_reg_in[43] , dpath_acc_reg_in[42] ,
         dpath_acc_reg_in[41] , dpath_acc_reg_in[40] ,
         dpath_acc_reg_in[39] , dpath_acc_reg_in[38] ,
         dpath_acc_reg_in[37] , dpath_acc_reg_in[36] ,
         dpath_acc_reg_in[35] , dpath_acc_reg_in[34] ,
         dpath_acc_reg_in[33] , dpath_acc_reg_in[32] ,
         dpath_acc_reg_in[31] , dpath_acc_reg_in[30] ,
         dpath_acc_reg_in[29] , dpath_acc_reg_in[28] ,
         dpath_acc_reg_in[27] , dpath_acc_reg_in[26] ,
         dpath_acc_reg_in[25] , dpath_acc_reg_in[24] ,
         dpath_acc_reg_in[23] , dpath_acc_reg_in[22] ,
         dpath_acc_reg_in[21] , dpath_acc_reg_in[20] ,
         dpath_acc_reg_in[19] , dpath_acc_reg_in[18] ,
         dpath_acc_reg_in[17] , dpath_acc_reg_in[16] ,
         dpath_acc_reg_in[15] , dpath_acc_reg_in[14] ,
         dpath_acc_reg_in[13] , dpath_acc_reg_in[12] ,
         dpath_acc_reg_in[11] , dpath_acc_reg_in[10] , dpath_acc_reg_in[9] ,
         dpath_acc_reg_in[8] , dpath_acc_reg_in[7] , dpath_acc_reg_in[6] ,
         dpath_acc_reg_in[5] , dpath_acc_reg_in[4] , dpath_acc_reg_in[3] ,
         dpath_acc_reg_in[2] , dpath_acc_reg_in[1] , dpath_acc_reg_in[0] ,
         dpath_acc_reg_shf2 , dpath_areg[96] , dpath_areg[95] ,
         dpath_areg[94] , dpath_areg[93] , dpath_areg[92] ,
         dpath_areg[91] , dpath_areg[90] , dpath_areg[89] ,
         dpath_areg[88] , dpath_areg[87] , dpath_areg[86] ,
         dpath_areg[85] , dpath_areg[84] , dpath_areg[83] ,
         dpath_areg[82] , dpath_areg[81] , dpath_areg[80] ,
         dpath_areg[79] , dpath_areg[78] , dpath_areg[77] ,
         dpath_areg[76] , dpath_areg[75] , dpath_areg[74] ,
         dpath_areg[73] , dpath_areg[72] , dpath_areg[71] ,
         dpath_areg[70] , dpath_areg[69] , dpath_areg[68] ,
         dpath_areg[67] , dpath_areg[66] , dpath_areg[65] ,
         dpath_areg[64] , dpath_areg[63] , dpath_areg[62] ,
         dpath_areg[61] , dpath_areg[60] , dpath_areg[59] ,
         dpath_areg[58] , dpath_areg[57] , dpath_areg[56] ,
         dpath_areg[55] , dpath_areg[54] , dpath_areg[53] ,
         dpath_areg[52] , dpath_areg[51] , dpath_areg[50] ,
         dpath_areg[49] , dpath_areg[48] , dpath_areg[47] ,
         dpath_areg[46] , dpath_areg[45] , dpath_areg[44] ,
         dpath_areg[43] , dpath_areg[42] , dpath_areg[41] ,
         dpath_areg[40] , dpath_areg[39] , dpath_areg[38] ,
         dpath_areg[37] , dpath_areg[36] , dpath_areg[35] ,
         dpath_areg[34] , dpath_areg[33] , dpath_areg[32] ,
         dpath_areg[31] , dpath_areg[30] , dpath_areg[29] ,
         dpath_areg[28] , dpath_areg[27] , dpath_areg[26] ,
         dpath_areg[25] , dpath_areg[24] , dpath_areg[23] ,
         dpath_areg[22] , dpath_areg[21] , dpath_areg[20] ,
         dpath_areg[19] , dpath_areg[18] , dpath_areg[17] ,
         dpath_areg[16] , dpath_areg[15] , dpath_areg[14] ,
         dpath_areg[13] , dpath_areg[12] , dpath_areg[11] ,
         dpath_areg[10] , dpath_areg[9] , dpath_areg[8] , dpath_areg[7] ,
         dpath_areg[6] , dpath_areg[5] , dpath_areg[4] , dpath_areg[3] ,
         dpath_areg[2] , dpath_areg[1] , dpath_areg[0] , dpath_mout[0] ,
         dpath_mout[1] , dpath_mout[2] , dpath_mout[3] , dpath_mout[4] ,
         dpath_mout[5] , dpath_mout[6] , dpath_mout[7] , dpath_mout[8] ,
         dpath_mout[9] , dpath_mout[10] , dpath_mout[11] , dpath_mout[12] ,
         dpath_mout[13] , dpath_mout[14] , dpath_mout[15] ,
         dpath_mout[16] , dpath_mout[17] , dpath_mout[18] ,
         dpath_mout[19] , dpath_mout[20] , dpath_mout[21] ,
         dpath_mout[22] , dpath_mout[23] , dpath_mout[24] ,
         dpath_mout[25] , dpath_mout[26] , dpath_mout[27] ,
         dpath_mout[28] , dpath_mout[29] , dpath_mout[30] ,
         dpath_mout[31] , dpath_mout[32] , dpath_mout[33] ,
         dpath_mout[34] , dpath_mout[35] , dpath_mout[36] ,
         dpath_mout[37] , dpath_mout[38] , dpath_mout[39] ,
         dpath_mout[40] , dpath_mout[41] , dpath_mout[42] ,
         dpath_mout[43] , dpath_mout[44] , dpath_mout[45] ,
         dpath_mout[46] , dpath_mout[47] , dpath_mout[48] ,
         dpath_mout[49] , dpath_mout[50] , dpath_mout[51] ,
         dpath_mout[52] , dpath_mout[53] , dpath_mout[54] ,
         dpath_mout[55] , dpath_mout[56] , dpath_mout[57] ,
         dpath_mout[58] , dpath_mout[59] , dpath_mout[60] ,
         dpath_mout[61] , dpath_mout[62] , dpath_mout[63] ,
         dpath_mout[64] , dpath_mout[65] , dpath_mout[66] ,
         dpath_mout[67] , dpath_mout[68] , dpath_mout[69] ,
         dpath_mout[70] , dpath_mout[71] , dpath_mout[72] ,
         dpath_mout[73] , dpath_mout[74] , dpath_mout[75] ,
         dpath_mout[76] , dpath_mout[77] , dpath_mout[78] ,
         dpath_mout[79] , dpath_mout[80] , dpath_mout[81] ,
         dpath_mout[82] , dpath_mout[83] , dpath_mout[84] ,
         dpath_mout[85] , dpath_mout[86] , dpath_mout[87] ,
         dpath_mout[88] , dpath_mout[89] , dpath_mout[90] ,
         dpath_mout[91] , dpath_mout[92] , dpath_mout[93] ,
         dpath_mout[94] , dpath_mout[95] , dpath_mout[96] ,
         dpath_mout[97] , dpath_mout[98] , dpath_mout[99] ,
         dpath_mout[100] , dpath_mout[101] , dpath_mout[102] ,
         dpath_mout[103] , dpath_mout[104] , dpath_mout[105] ,
         dpath_mout[106] , dpath_mout[107] , dpath_mout[108] ,
         dpath_mout[109] , dpath_mout[110] , dpath_mout[111] ,
         dpath_mout[112] , dpath_mout[113] , dpath_mout[114] ,
         dpath_mout[115] , dpath_mout[116] , dpath_mout[117] ,
         dpath_mout[118] , dpath_mout[119] , dpath_mout[120] ,
         dpath_mout[121] , dpath_mout[122] , dpath_mout[123] ,
         dpath_mout[124] , dpath_mout[125] , dpath_mout[126] ,
         dpath_mout[127] , dpath_mout[128] , dpath_mout[129] ,
         dpath_mout[130] , dpath_mout[131] , dpath_mout[132] ,
         dpath_mout[133] , dpath_mout[134] , dpath_mout[135] ,
         dpath_acc_reg[0] , dpath_acc_reg[1] , dpath_acc_reg[2] ,
         dpath_acc_reg[3] , dpath_acc_reg[4] , dpath_acc_reg[5] ,
         dpath_acc_reg[6] , dpath_acc_reg[7] , dpath_acc_reg[8] ,
         dpath_acc_reg[9] , dpath_acc_reg[10] , dpath_acc_reg[11] ,
         dpath_acc_reg[12] , dpath_acc_reg[13] , dpath_acc_reg[14] ,
         dpath_acc_reg[15] , dpath_acc_reg[16] , dpath_acc_reg[17] ,
         dpath_acc_reg[18] , dpath_acc_reg[19] , dpath_acc_reg[20] ,
         dpath_acc_reg[21] , dpath_acc_reg[22] , dpath_acc_reg[23] ,
         dpath_acc_reg[24] , dpath_acc_reg[25] , dpath_acc_reg[26] ,
         dpath_acc_reg[27] , dpath_acc_reg[28] , dpath_acc_reg[29] ,
         dpath_acc_reg[30] , dpath_acc_reg[31] , dpath_acc_reg[32] ,
         dpath_acc_reg[33] , dpath_acc_reg[34] , dpath_acc_reg[35] ,
         dpath_acc_reg[36] , dpath_acc_reg[37] , dpath_acc_reg[38] ,
         dpath_acc_reg[39] , dpath_acc_reg[40] , dpath_acc_reg[41] ,
         dpath_acc_reg[42] , dpath_acc_reg[43] , dpath_acc_reg[44] ,
         dpath_acc_reg[45] , dpath_acc_reg[46] , dpath_acc_reg[47] ,
         dpath_acc_reg[48] , dpath_acc_reg[49] , dpath_acc_reg[50] ,
         dpath_acc_reg[51] , dpath_acc_reg[52] , dpath_acc_reg[53] ,
         dpath_acc_reg[54] , dpath_acc_reg[55] , dpath_acc_reg[56] ,
         dpath_acc_reg[57] , dpath_acc_reg[58] , dpath_acc_reg[59] ,
         dpath_acc_reg[60] , dpath_acc_reg[61] , dpath_acc_reg[62] ,
         dpath_acc_reg[63] , dpath_acc_reg[64] , dpath_acc_reg[65] ,
         dpath_acc_reg[66] , dpath_acc_reg[67] , dpath_acc_reg[68] ,
         dpath_acc_reg[69] , dpath_acc_reg[70] , dpath_acc_reg[71] ,
         dpath_acc_reg[72] , dpath_acc_reg[73] , dpath_acc_reg[74] ,
         dpath_acc_reg[75] , dpath_acc_reg[76] , dpath_acc_reg[77] ,
         dpath_acc_reg[78] , dpath_acc_reg[79] , dpath_acc_reg[80] ,
         dpath_acc_reg[81] , dpath_acc_reg[82] , dpath_acc_reg[83] ,
         dpath_acc_reg[84] , dpath_acc_reg[85] , dpath_acc_reg[86] ,
         dpath_acc_reg[87] , dpath_acc_reg[88] , dpath_acc_reg[89] ,
         dpath_acc_reg[90] , dpath_acc_reg[91] , dpath_acc_reg[92] ,
         dpath_acc_reg[93] , dpath_acc_reg[94] , dpath_acc_reg[95] ,
         dpath_acc_reg[96] , dpath_acc_reg[97] , dpath_acc_reg[98] ,
         dpath_acc_reg[99] , dpath_acc_reg[100] , dpath_acc_reg[101] ,
         dpath_acc_reg[102] , dpath_acc_reg[103] , dpath_acc_reg[104] ,
         dpath_acc_reg[105] , dpath_acc_reg[106] , dpath_acc_reg[107] ,
         dpath_acc_reg[108] , dpath_acc_reg[109] , dpath_acc_reg[110] ,
         dpath_acc_reg[111] , dpath_acc_reg[112] , dpath_acc_reg[113] ,
         dpath_acc_reg[114] , dpath_acc_reg[115] , dpath_acc_reg[116] ,
         dpath_acc_reg[117] , dpath_acc_reg[118] , dpath_acc_reg[119] ,
         dpath_acc_reg[120] , dpath_acc_reg[121] , dpath_acc_reg[122] ,
         dpath_acc_reg[123] , dpath_acc_reg[124] , dpath_acc_reg[125] ,
         dpath_acc_reg[126] , dpath_acc_reg[127] , dpath_acc_reg[128] ,
         dpath_acc_reg[129] , dpath_acc_reg[130] , dpath_acc_reg[131] ,
         dpath_acc_reg[132] , dpath_acc_reg[133] , dpath_acc_reg[134] ,
         dpath_acc_reg[135] , dpath_mul_op2_d[63] , dpath_mul_op2_d[62] ,
         dpath_mul_op2_d[61] , dpath_mul_op2_d[60] , dpath_mul_op2_d[59] ,
         dpath_mul_op2_d[58] , dpath_mul_op2_d[57] , dpath_mul_op2_d[56] ,
         dpath_mul_op2_d[55] , dpath_mul_op2_d[54] , dpath_mul_op2_d[53] ,
         dpath_mul_op2_d[52] , dpath_mul_op2_d[51] , dpath_mul_op2_d[50] ,
         dpath_mul_op2_d[49] , dpath_mul_op2_d[48] , dpath_mul_op2_d[47] ,
         dpath_mul_op2_d[46] , dpath_mul_op2_d[45] , dpath_mul_op2_d[44] ,
         dpath_mul_op2_d[43] , dpath_mul_op2_d[42] , dpath_mul_op2_d[41] ,
         dpath_mul_op2_d[40] , dpath_mul_op2_d[39] , dpath_mul_op2_d[38] ,
         dpath_mul_op2_d[37] , dpath_mul_op2_d[36] , dpath_mul_op2_d[35] ,
         dpath_mul_op2_d[34] , dpath_mul_op2_d[33] , dpath_mul_op2_d[32] ,
         dpath_mul_op2_d[30] , dpath_mul_op2_d[28] , dpath_mul_op2_d[26] ,
         dpath_mul_op2_d[24] , dpath_mul_op2_d[22] , dpath_mul_op2_d[20] ,
         dpath_mul_op2_d[18] , dpath_mul_op2_d[16] , dpath_mul_op2_d[14] ,
         dpath_mul_op2_d[12] , dpath_mul_op2_d[10] , dpath_mul_op2_d[8] ,
         dpath_mul_op2_d[6] , dpath_mul_op2_d[4] , dpath_mul_op2_d[2] ,
         dpath_mul_op2_d[0] , dpath_mulcore_add_co96 ,
         dpath_mulcore_addout[103] , dpath_mulcore_addout[102] ,
         dpath_mulcore_addout[101] , dpath_mulcore_addout[100] ,
         dpath_mulcore_addout[99] , dpath_mulcore_addout[98] ,
         dpath_mulcore_addout[97] , dpath_mulcore_addout[96] ,
         dpath_mulcore_addout[95] , dpath_mulcore_addout[94] ,
         dpath_mulcore_addout[93] , dpath_mulcore_addout[92] ,
         dpath_mulcore_addout[91] , dpath_mulcore_addout[90] ,
         dpath_mulcore_addout[89] , dpath_mulcore_addout[88] ,
         dpath_mulcore_addout[87] , dpath_mulcore_addout[86] ,
         dpath_mulcore_addout[85] , dpath_mulcore_addout[84] ,
         dpath_mulcore_addout[83] , dpath_mulcore_addout[82] ,
         dpath_mulcore_addout[81] , dpath_mulcore_addout[80] ,
         dpath_mulcore_addout[79] , dpath_mulcore_addout[78] ,
         dpath_mulcore_addout[77] , dpath_mulcore_addout[76] ,
         dpath_mulcore_addout[75] , dpath_mulcore_addout[74] ,
         dpath_mulcore_addout[73] , dpath_mulcore_addout[72] ,
         dpath_mulcore_addout[71] , dpath_mulcore_addout[70] ,
         dpath_mulcore_addout[69] , dpath_mulcore_addout[68] ,
         dpath_mulcore_addout[67] , dpath_mulcore_addout[66] ,
         dpath_mulcore_addout[65] , dpath_mulcore_addout[64] ,
         dpath_mulcore_addout[63] , dpath_mulcore_addout[62] ,
         dpath_mulcore_addout[61] , dpath_mulcore_addout[60] ,
         dpath_mulcore_addout[59] , dpath_mulcore_addout[58] ,
         dpath_mulcore_addout[57] , dpath_mulcore_addout[56] ,
         dpath_mulcore_addout[55] , dpath_mulcore_addout[54] ,
         dpath_mulcore_addout[53] , dpath_mulcore_addout[52] ,
         dpath_mulcore_addout[51] , dpath_mulcore_addout[50] ,
         dpath_mulcore_addout[49] , dpath_mulcore_addout[48] ,
         dpath_mulcore_addout[47] , dpath_mulcore_addout[46] ,
         dpath_mulcore_addout[45] , dpath_mulcore_addout[44] ,
         dpath_mulcore_addout[43] , dpath_mulcore_addout[42] ,
         dpath_mulcore_addout[41] , dpath_mulcore_addout[40] ,
         dpath_mulcore_addout[39] , dpath_mulcore_addout[38] ,
         dpath_mulcore_addout[37] , dpath_mulcore_addout[36] ,
         dpath_mulcore_addout[35] , dpath_mulcore_addout[34] ,
         dpath_mulcore_addout[33] , dpath_mulcore_addout[32] ,
         dpath_mulcore_addout[31] , dpath_mulcore_addout[30] ,
         dpath_mulcore_addout[29] , dpath_mulcore_addout[28] ,
         dpath_mulcore_addout[27] , dpath_mulcore_addout[26] ,
         dpath_mulcore_addout[25] , dpath_mulcore_addout[24] ,
         dpath_mulcore_addout[23] , dpath_mulcore_addout[22] ,
         dpath_mulcore_addout[21] , dpath_mulcore_addout[20] ,
         dpath_mulcore_addout[19] , dpath_mulcore_addout[18] ,
         dpath_mulcore_addout[17] , dpath_mulcore_addout[16] ,
         dpath_mulcore_addout[15] , dpath_mulcore_addout[14] ,
         dpath_mulcore_addout[13] , dpath_mulcore_addout[12] ,
         dpath_mulcore_addout[11] , dpath_mulcore_addout[10] ,
         dpath_mulcore_addout[9] , dpath_mulcore_addout[8] ,
         dpath_mulcore_addout[7] , dpath_mulcore_addout[6] ,
         dpath_mulcore_addout[5] , dpath_mulcore_addout[4] ,
         dpath_mulcore_addout[3] , dpath_mulcore_addout[2] ,
         dpath_mulcore_addout[1] , dpath_mulcore_addout[0] ,
         dpath_mulcore_addin_cin , dpath_mulcore_add_cin ,
         dpath_mulcore_add_co31 , dpath_mulcore_pcout_in[97] ,
         dpath_mulcore_pcout_in[96] , dpath_mulcore_pcout_in[95] ,
         dpath_mulcore_pcout_in[94] , dpath_mulcore_pcout_in[93] ,
         dpath_mulcore_pcout_in[92] , dpath_mulcore_pcout_in[91] ,
         dpath_mulcore_pcout_in[90] , dpath_mulcore_pcout_in[89] ,
         dpath_mulcore_pcout_in[88] , dpath_mulcore_pcout_in[87] ,
         dpath_mulcore_pcout_in[86] , dpath_mulcore_pcout_in[85] ,
         dpath_mulcore_pcout_in[84] , dpath_mulcore_pcout_in[83] ,
         dpath_mulcore_pcout_in[82] , dpath_mulcore_pcout_in[81] ,
         dpath_mulcore_pcout_in[80] , dpath_mulcore_pcout_in[79] ,
         dpath_mulcore_pcout_in[78] , dpath_mulcore_pcout_in[77] ,
         dpath_mulcore_pcout_in[76] , dpath_mulcore_pcout_in[75] ,
         dpath_mulcore_pcout_in[74] , dpath_mulcore_pcout_in[73] ,
         dpath_mulcore_pcout_in[72] , dpath_mulcore_pcout_in[71] ,
         dpath_mulcore_pcout_in[70] , dpath_mulcore_pcout_in[69] ,
         dpath_mulcore_pcout_in[68] , dpath_mulcore_pcout_in[67] ,
         dpath_mulcore_pcout_in[66] , dpath_mulcore_pcout_in[65] ,
         dpath_mulcore_pcout_in[64] , dpath_mulcore_pcout_in[63] ,
         dpath_mulcore_pcout_in[62] , dpath_mulcore_pcout_in[61] ,
         dpath_mulcore_pcout_in[60] , dpath_mulcore_pcout_in[59] ,
         dpath_mulcore_pcout_in[58] , dpath_mulcore_pcout_in[57] ,
         dpath_mulcore_pcout_in[56] , dpath_mulcore_pcout_in[55] ,
         dpath_mulcore_pcout_in[54] , dpath_mulcore_pcout_in[53] ,
         dpath_mulcore_pcout_in[52] , dpath_mulcore_pcout_in[51] ,
         dpath_mulcore_pcout_in[50] , dpath_mulcore_pcout_in[49] ,
         dpath_mulcore_pcout_in[48] , dpath_mulcore_pcout_in[47] ,
         dpath_mulcore_pcout_in[46] , dpath_mulcore_pcout_in[45] ,
         dpath_mulcore_pcout_in[44] , dpath_mulcore_pcout_in[43] ,
         dpath_mulcore_pcout_in[42] , dpath_mulcore_pcout_in[41] ,
         dpath_mulcore_pcout_in[40] , dpath_mulcore_pcout_in[39] ,
         dpath_mulcore_pcout_in[38] , dpath_mulcore_pcout_in[37] ,
         dpath_mulcore_pcout_in[36] , dpath_mulcore_pcout_in[35] ,
         dpath_mulcore_pcout_in[34] , dpath_mulcore_pcout_in[33] ,
         dpath_mulcore_pcout_in[32] , dpath_mulcore_pcout_in[31] ,
         dpath_mulcore_pcout_in[30] , dpath_mulcore_psum_in[98] ,
         dpath_mulcore_psum_in[97] , dpath_mulcore_psum_in[96] ,
         dpath_mulcore_psum_in[95] , dpath_mulcore_psum_in[94] ,
         dpath_mulcore_psum_in[93] , dpath_mulcore_psum_in[92] ,
         dpath_mulcore_psum_in[91] , dpath_mulcore_psum_in[90] ,
         dpath_mulcore_psum_in[89] , dpath_mulcore_psum_in[88] ,
         dpath_mulcore_psum_in[87] , dpath_mulcore_psum_in[86] ,
         dpath_mulcore_psum_in[85] , dpath_mulcore_psum_in[84] ,
         dpath_mulcore_psum_in[83] , dpath_mulcore_psum_in[82] ,
         dpath_mulcore_psum_in[81] , dpath_mulcore_psum_in[80] ,
         dpath_mulcore_psum_in[79] , dpath_mulcore_psum_in[78] ,
         dpath_mulcore_psum_in[77] , dpath_mulcore_psum_in[76] ,
         dpath_mulcore_psum_in[75] , dpath_mulcore_psum_in[74] ,
         dpath_mulcore_psum_in[73] , dpath_mulcore_psum_in[72] ,
         dpath_mulcore_psum_in[71] , dpath_mulcore_psum_in[70] ,
         dpath_mulcore_psum_in[69] , dpath_mulcore_psum_in[68] ,
         dpath_mulcore_psum_in[67] , dpath_mulcore_psum_in[66] ,
         dpath_mulcore_psum_in[65] , dpath_mulcore_psum_in[64] ,
         dpath_mulcore_psum_in[63] , dpath_mulcore_psum_in[62] ,
         dpath_mulcore_psum_in[61] , dpath_mulcore_psum_in[60] ,
         dpath_mulcore_psum_in[59] , dpath_mulcore_psum_in[58] ,
         dpath_mulcore_psum_in[57] , dpath_mulcore_psum_in[56] ,
         dpath_mulcore_psum_in[55] , dpath_mulcore_psum_in[54] ,
         dpath_mulcore_psum_in[53] , dpath_mulcore_psum_in[52] ,
         dpath_mulcore_psum_in[51] , dpath_mulcore_psum_in[50] ,
         dpath_mulcore_psum_in[49] , dpath_mulcore_psum_in[48] ,
         dpath_mulcore_psum_in[47] , dpath_mulcore_psum_in[46] ,
         dpath_mulcore_psum_in[45] , dpath_mulcore_psum_in[44] ,
         dpath_mulcore_psum_in[43] , dpath_mulcore_psum_in[42] ,
         dpath_mulcore_psum_in[41] , dpath_mulcore_psum_in[40] ,
         dpath_mulcore_psum_in[39] , dpath_mulcore_psum_in[38] ,
         dpath_mulcore_psum_in[37] , dpath_mulcore_psum_in[36] ,
         dpath_mulcore_psum_in[35] , dpath_mulcore_psum_in[34] ,
         dpath_mulcore_psum_in[33] , dpath_mulcore_psum_in[32] ,
         dpath_mulcore_psum_in[31] , dpath_mulcore_addin_sum[97] ,
         dpath_mulcore_addin_sum[96] , dpath_mulcore_addin_sum[95] ,
         dpath_mulcore_addin_sum[94] , dpath_mulcore_addin_sum[93] ,
         dpath_mulcore_addin_sum[92] , dpath_mulcore_addin_sum[91] ,
         dpath_mulcore_addin_sum[90] , dpath_mulcore_addin_sum[89] ,
         dpath_mulcore_addin_sum[88] , dpath_mulcore_addin_sum[87] ,
         dpath_mulcore_addin_sum[86] , dpath_mulcore_addin_sum[85] ,
         dpath_mulcore_addin_sum[84] , dpath_mulcore_addin_sum[83] ,
         dpath_mulcore_addin_sum[82] , dpath_mulcore_addin_sum[81] ,
         dpath_mulcore_addin_sum[80] , dpath_mulcore_addin_sum[79] ,
         dpath_mulcore_addin_sum[78] , dpath_mulcore_addin_sum[77] ,
         dpath_mulcore_addin_sum[76] , dpath_mulcore_addin_sum[75] ,
         dpath_mulcore_addin_sum[74] , dpath_mulcore_addin_sum[73] ,
         dpath_mulcore_addin_sum[72] , dpath_mulcore_addin_sum[71] ,
         dpath_mulcore_addin_sum[70] , dpath_mulcore_addin_sum[69] ,
         dpath_mulcore_addin_sum[68] , dpath_mulcore_addin_sum[67] ,
         dpath_mulcore_addin_sum[66] , dpath_mulcore_addin_sum[65] ,
         dpath_mulcore_addin_sum[64] , dpath_mulcore_addin_sum[63] ,
         dpath_mulcore_addin_sum[62] , dpath_mulcore_addin_sum[61] ,
         dpath_mulcore_addin_sum[60] , dpath_mulcore_addin_sum[59] ,
         dpath_mulcore_addin_sum[58] , dpath_mulcore_addin_sum[57] ,
         dpath_mulcore_addin_sum[56] , dpath_mulcore_addin_sum[55] ,
         dpath_mulcore_addin_sum[54] , dpath_mulcore_addin_sum[53] ,
         dpath_mulcore_addin_sum[52] , dpath_mulcore_addin_sum[51] ,
         dpath_mulcore_addin_sum[50] , dpath_mulcore_addin_sum[49] ,
         dpath_mulcore_addin_sum[48] , dpath_mulcore_addin_sum[47] ,
         dpath_mulcore_addin_sum[46] , dpath_mulcore_addin_sum[45] ,
         dpath_mulcore_addin_sum[44] , dpath_mulcore_addin_sum[43] ,
         dpath_mulcore_addin_sum[42] , dpath_mulcore_addin_sum[41] ,
         dpath_mulcore_addin_sum[40] , dpath_mulcore_addin_sum[39] ,
         dpath_mulcore_addin_sum[38] , dpath_mulcore_addin_sum[37] ,
         dpath_mulcore_addin_sum[36] , dpath_mulcore_addin_sum[35] ,
         dpath_mulcore_addin_sum[34] , dpath_mulcore_addin_sum[33] ,
         dpath_mulcore_addin_sum[32] , dpath_mulcore_addin_sum[31] ,
         dpath_mulcore_addin_sum[30] , dpath_mulcore_addin_sum[29] ,
         dpath_mulcore_addin_sum[28] , dpath_mulcore_addin_sum[27] ,
         dpath_mulcore_addin_sum[26] , dpath_mulcore_addin_sum[25] ,
         dpath_mulcore_addin_sum[24] , dpath_mulcore_addin_sum[23] ,
         dpath_mulcore_addin_sum[22] , dpath_mulcore_addin_sum[21] ,
         dpath_mulcore_addin_sum[20] , dpath_mulcore_addin_sum[19] ,
         dpath_mulcore_addin_sum[18] , dpath_mulcore_addin_sum[17] ,
         dpath_mulcore_addin_sum[16] , dpath_mulcore_addin_sum[15] ,
         dpath_mulcore_addin_sum[14] , dpath_mulcore_addin_sum[13] ,
         dpath_mulcore_addin_sum[12] , dpath_mulcore_addin_sum[11] ,
         dpath_mulcore_addin_sum[10] , dpath_mulcore_addin_sum[9] ,
         dpath_mulcore_addin_sum[8] , dpath_mulcore_addin_sum[7] ,
         dpath_mulcore_addin_sum[6] , dpath_mulcore_addin_sum[5] ,
         dpath_mulcore_addin_sum[4] , dpath_mulcore_addin_sum[3] ,
         dpath_mulcore_addin_sum[2] , dpath_mulcore_addin_sum[1] ,
         dpath_mulcore_addin_sum[0] , dpath_mulcore_ary2_sum[97] ,
         dpath_mulcore_ary2_sum[96] , dpath_mulcore_ary2_sum[95] ,
         dpath_mulcore_ary2_sum[94] , dpath_mulcore_ary2_sum[93] ,
         dpath_mulcore_ary2_sum[92] , dpath_mulcore_ary2_sum[91] ,
         dpath_mulcore_ary2_sum[90] , dpath_mulcore_ary2_sum[89] ,
         dpath_mulcore_ary2_sum[88] , dpath_mulcore_ary2_sum[87] ,
         dpath_mulcore_ary2_sum[86] , dpath_mulcore_ary2_sum[85] ,
         dpath_mulcore_ary2_sum[84] , dpath_mulcore_ary2_sum[83] ,
         dpath_mulcore_ary2_sum[82] , dpath_mulcore_ary2_sum[81] ,
         dpath_mulcore_ary2_sum[80] , dpath_mulcore_ary2_sum[79] ,
         dpath_mulcore_ary2_sum[78] , dpath_mulcore_ary2_sum[77] ,
         dpath_mulcore_ary2_sum[76] , dpath_mulcore_ary2_sum[75] ,
         dpath_mulcore_ary2_sum[74] , dpath_mulcore_ary2_sum[73] ,
         dpath_mulcore_ary2_sum[72] , dpath_mulcore_ary2_sum[71] ,
         dpath_mulcore_ary2_sum[70] , dpath_mulcore_ary2_sum[69] ,
         dpath_mulcore_ary2_sum[68] , dpath_mulcore_ary2_sum[67] ,
         dpath_mulcore_ary2_sum[66] , dpath_mulcore_ary2_sum[65] ,
         dpath_mulcore_ary2_sum[64] , dpath_mulcore_ary2_sum[63] ,
         dpath_mulcore_ary2_sum[62] , dpath_mulcore_ary2_sum[61] ,
         dpath_mulcore_ary2_sum[60] , dpath_mulcore_ary2_sum[59] ,
         dpath_mulcore_ary2_sum[58] , dpath_mulcore_ary2_sum[57] ,
         dpath_mulcore_ary2_sum[56] , dpath_mulcore_ary2_sum[55] ,
         dpath_mulcore_ary2_sum[54] , dpath_mulcore_ary2_sum[53] ,
         dpath_mulcore_ary2_sum[52] , dpath_mulcore_ary2_sum[51] ,
         dpath_mulcore_ary2_sum[50] , dpath_mulcore_ary2_sum[49] ,
         dpath_mulcore_ary2_sum[48] , dpath_mulcore_ary2_sum[47] ,
         dpath_mulcore_ary2_sum[46] , dpath_mulcore_ary2_sum[45] ,
         dpath_mulcore_ary2_sum[44] , dpath_mulcore_ary2_sum[43] ,
         dpath_mulcore_ary2_sum[42] , dpath_mulcore_ary2_sum[41] ,
         dpath_mulcore_ary2_sum[40] , dpath_mulcore_ary2_sum[39] ,
         dpath_mulcore_ary2_sum[38] , dpath_mulcore_ary2_sum[37] ,
         dpath_mulcore_ary2_sum[36] , dpath_mulcore_ary2_sum[35] ,
         dpath_mulcore_ary2_sum[34] , dpath_mulcore_ary2_sum[33] ,
         dpath_mulcore_ary2_sum[32] , dpath_mulcore_ary2_sum[31] ,
         dpath_mulcore_ary2_sum[30] , dpath_mulcore_ary2_sum[29] ,
         dpath_mulcore_ary2_sum[28] , dpath_mulcore_ary2_sum[27] ,
         dpath_mulcore_ary2_sum[26] , dpath_mulcore_ary2_sum[25] ,
         dpath_mulcore_ary2_sum[24] , dpath_mulcore_ary2_sum[23] ,
         dpath_mulcore_ary2_sum[22] , dpath_mulcore_ary2_sum[21] ,
         dpath_mulcore_ary2_sum[20] , dpath_mulcore_ary2_sum[19] ,
         dpath_mulcore_ary2_sum[18] , dpath_mulcore_ary2_sum[17] ,
         dpath_mulcore_ary2_sum[16] , dpath_mulcore_ary2_sum[15] ,
         dpath_mulcore_ary2_sum[14] , dpath_mulcore_ary2_sum[13] ,
         dpath_mulcore_ary2_sum[12] , dpath_mulcore_ary2_sum[11] ,
         dpath_mulcore_ary2_sum[10] , dpath_mulcore_ary2_sum[9] ,
         dpath_mulcore_ary2_sum[8] , dpath_mulcore_ary2_sum[7] ,
         dpath_mulcore_ary2_sum[6] , dpath_mulcore_ary2_sum[5] ,
         dpath_mulcore_ary2_sum[4] , dpath_mulcore_ary2_sum[3] ,
         dpath_mulcore_ary2_sum[2] , dpath_mulcore_ary2_sum[1] ,
         dpath_mulcore_ary2_sum[0] , dpath_mulcore_addin_cout[96] ,
         dpath_mulcore_addin_cout[95] , dpath_mulcore_addin_cout[94] ,
         dpath_mulcore_addin_cout[93] , dpath_mulcore_addin_cout[92] ,
         dpath_mulcore_addin_cout[91] , dpath_mulcore_addin_cout[90] ,
         dpath_mulcore_addin_cout[89] , dpath_mulcore_addin_cout[88] ,
         dpath_mulcore_addin_cout[87] , dpath_mulcore_addin_cout[86] ,
         dpath_mulcore_addin_cout[85] , dpath_mulcore_addin_cout[84] ,
         dpath_mulcore_addin_cout[83] , dpath_mulcore_addin_cout[82] ,
         dpath_mulcore_addin_cout[81] , dpath_mulcore_addin_cout[80] ,
         dpath_mulcore_addin_cout[79] , dpath_mulcore_addin_cout[78] ,
         dpath_mulcore_addin_cout[77] , dpath_mulcore_addin_cout[76] ,
         dpath_mulcore_addin_cout[75] , dpath_mulcore_addin_cout[74] ,
         dpath_mulcore_addin_cout[73] , dpath_mulcore_addin_cout[72] ,
         dpath_mulcore_addin_cout[71] , dpath_mulcore_addin_cout[70] ,
         dpath_mulcore_addin_cout[69] , dpath_mulcore_addin_cout[68] ,
         dpath_mulcore_addin_cout[67] , dpath_mulcore_addin_cout[66] ,
         dpath_mulcore_addin_cout[65] , dpath_mulcore_addin_cout[64] ,
         dpath_mulcore_addin_cout[63] , dpath_mulcore_addin_cout[62] ,
         dpath_mulcore_addin_cout[61] , dpath_mulcore_addin_cout[60] ,
         dpath_mulcore_addin_cout[59] , dpath_mulcore_addin_cout[58] ,
         dpath_mulcore_addin_cout[57] , dpath_mulcore_addin_cout[56] ,
         dpath_mulcore_addin_cout[55] , dpath_mulcore_addin_cout[54] ,
         dpath_mulcore_addin_cout[53] , dpath_mulcore_addin_cout[52] ,
         dpath_mulcore_addin_cout[51] , dpath_mulcore_addin_cout[50] ,
         dpath_mulcore_addin_cout[49] , dpath_mulcore_addin_cout[48] ,
         dpath_mulcore_addin_cout[47] , dpath_mulcore_addin_cout[46] ,
         dpath_mulcore_addin_cout[45] , dpath_mulcore_addin_cout[44] ,
         dpath_mulcore_addin_cout[43] , dpath_mulcore_addin_cout[42] ,
         dpath_mulcore_addin_cout[41] , dpath_mulcore_addin_cout[40] ,
         dpath_mulcore_addin_cout[39] , dpath_mulcore_addin_cout[38] ,
         dpath_mulcore_addin_cout[37] , dpath_mulcore_addin_cout[36] ,
         dpath_mulcore_addin_cout[35] , dpath_mulcore_addin_cout[34] ,
         dpath_mulcore_addin_cout[33] , dpath_mulcore_addin_cout[32] ,
         dpath_mulcore_addin_cout[31] , dpath_mulcore_addin_cout[30] ,
         dpath_mulcore_addin_cout[29] , dpath_mulcore_addin_cout[28] ,
         dpath_mulcore_addin_cout[27] , dpath_mulcore_addin_cout[26] ,
         dpath_mulcore_addin_cout[25] , dpath_mulcore_addin_cout[24] ,
         dpath_mulcore_addin_cout[23] , dpath_mulcore_addin_cout[22] ,
         dpath_mulcore_addin_cout[21] , dpath_mulcore_addin_cout[20] ,
         dpath_mulcore_addin_cout[19] , dpath_mulcore_addin_cout[18] ,
         dpath_mulcore_addin_cout[17] , dpath_mulcore_addin_cout[16] ,
         dpath_mulcore_addin_cout[15] , dpath_mulcore_addin_cout[14] ,
         dpath_mulcore_addin_cout[13] , dpath_mulcore_addin_cout[12] ,
         dpath_mulcore_addin_cout[11] , dpath_mulcore_addin_cout[10] ,
         dpath_mulcore_addin_cout[9] , dpath_mulcore_addin_cout[8] ,
         dpath_mulcore_addin_cout[7] , dpath_mulcore_addin_cout[6] ,
         dpath_mulcore_addin_cout[5] , dpath_mulcore_addin_cout[4] ,
         dpath_mulcore_addin_cout[3] , dpath_mulcore_addin_cout[2] ,
         dpath_mulcore_addin_cout[1] , dpath_mulcore_addin_cout[0] ,
         dpath_mulcore_ary2_cout[96] , dpath_mulcore_ary2_cout[95] ,
         dpath_mulcore_ary2_cout[94] , dpath_mulcore_ary2_cout[93] ,
         dpath_mulcore_ary2_cout[92] , dpath_mulcore_ary2_cout[91] ,
         dpath_mulcore_ary2_cout[90] , dpath_mulcore_ary2_cout[89] ,
         dpath_mulcore_ary2_cout[88] , dpath_mulcore_ary2_cout[87] ,
         dpath_mulcore_ary2_cout[86] , dpath_mulcore_ary2_cout[85] ,
         dpath_mulcore_ary2_cout[84] , dpath_mulcore_ary2_cout[83] ,
         dpath_mulcore_ary2_cout[82] , dpath_mulcore_ary2_cout[81] ,
         dpath_mulcore_ary2_cout[80] , dpath_mulcore_ary2_cout[79] ,
         dpath_mulcore_ary2_cout[78] , dpath_mulcore_ary2_cout[77] ,
         dpath_mulcore_ary2_cout[76] , dpath_mulcore_ary2_cout[75] ,
         dpath_mulcore_ary2_cout[74] , dpath_mulcore_ary2_cout[73] ,
         dpath_mulcore_ary2_cout[72] , dpath_mulcore_ary2_cout[71] ,
         dpath_mulcore_ary2_cout[70] , dpath_mulcore_ary2_cout[69] ,
         dpath_mulcore_ary2_cout[68] , dpath_mulcore_ary2_cout[67] ,
         dpath_mulcore_ary2_cout[66] , dpath_mulcore_ary2_cout[65] ,
         dpath_mulcore_ary2_cout[64] , dpath_mulcore_ary2_cout[63] ,
         dpath_mulcore_ary2_cout[62] , dpath_mulcore_ary2_cout[61] ,
         dpath_mulcore_ary2_cout[60] , dpath_mulcore_ary2_cout[59] ,
         dpath_mulcore_ary2_cout[58] , dpath_mulcore_ary2_cout[57] ,
         dpath_mulcore_ary2_cout[56] , dpath_mulcore_ary2_cout[55] ,
         dpath_mulcore_ary2_cout[54] , dpath_mulcore_ary2_cout[53] ,
         dpath_mulcore_ary2_cout[52] , dpath_mulcore_ary2_cout[51] ,
         dpath_mulcore_ary2_cout[50] , dpath_mulcore_ary2_cout[49] ,
         dpath_mulcore_ary2_cout[48] , dpath_mulcore_ary2_cout[47] ,
         dpath_mulcore_ary2_cout[46] , dpath_mulcore_ary2_cout[45] ,
         dpath_mulcore_ary2_cout[44] , dpath_mulcore_ary2_cout[43] ,
         dpath_mulcore_ary2_cout[42] , dpath_mulcore_ary2_cout[41] ,
         dpath_mulcore_ary2_cout[40] , dpath_mulcore_ary2_cout[39] ,
         dpath_mulcore_ary2_cout[38] , dpath_mulcore_ary2_cout[37] ,
         dpath_mulcore_ary2_cout[36] , dpath_mulcore_ary2_cout[35] ,
         dpath_mulcore_ary2_cout[34] , dpath_mulcore_ary2_cout[33] ,
         dpath_mulcore_ary2_cout[32] , dpath_mulcore_ary2_cout[31] ,
         dpath_mulcore_ary2_cout[30] , dpath_mulcore_ary2_cout[29] ,
         dpath_mulcore_ary2_cout[28] , dpath_mulcore_ary2_cout[27] ,
         dpath_mulcore_ary2_cout[26] , dpath_mulcore_ary2_cout[25] ,
         dpath_mulcore_ary2_cout[24] , dpath_mulcore_ary2_cout[23] ,
         dpath_mulcore_ary2_cout[22] , dpath_mulcore_ary2_cout[21] ,
         dpath_mulcore_ary2_cout[20] , dpath_mulcore_ary2_cout[19] ,
         dpath_mulcore_ary2_cout[18] , dpath_mulcore_ary2_cout[17] ,
         dpath_mulcore_ary2_cout[16] , dpath_mulcore_ary2_cout[15] ,
         dpath_mulcore_ary2_cout[14] , dpath_mulcore_ary2_cout[13] ,
         dpath_mulcore_ary2_cout[12] , dpath_mulcore_ary2_cout[11] ,
         dpath_mulcore_ary2_cout[10] , dpath_mulcore_ary2_cout[9] ,
         dpath_mulcore_ary2_cout[8] , dpath_mulcore_ary2_cout[7] ,
         dpath_mulcore_ary2_cout[6] , dpath_mulcore_ary2_cout[5] ,
         dpath_mulcore_ary2_cout[4] , dpath_mulcore_ary2_cout[3] ,
         dpath_mulcore_ary2_cout[2] , dpath_mulcore_ary2_cout[1] ,
         dpath_mulcore_ary2_cout[0] , dpath_mulcore_ps[98] ,
         dpath_mulcore_ps[97] , dpath_mulcore_ps[96] ,
         dpath_mulcore_ps[95] , dpath_mulcore_ps[94] ,
         dpath_mulcore_ps[93] , dpath_mulcore_ps[92] ,
         dpath_mulcore_ps[91] , dpath_mulcore_ps[90] ,
         dpath_mulcore_ps[89] , dpath_mulcore_ps[88] ,
         dpath_mulcore_ps[87] , dpath_mulcore_ps[86] ,
         dpath_mulcore_ps[85] , dpath_mulcore_ps[84] ,
         dpath_mulcore_ps[83] , dpath_mulcore_ps[82] ,
         dpath_mulcore_ps[81] , dpath_mulcore_ps[80] ,
         dpath_mulcore_ps[79] , dpath_mulcore_ps[78] ,
         dpath_mulcore_ps[77] , dpath_mulcore_ps[76] ,
         dpath_mulcore_ps[75] , dpath_mulcore_ps[74] ,
         dpath_mulcore_ps[73] , dpath_mulcore_ps[72] ,
         dpath_mulcore_ps[71] , dpath_mulcore_ps[70] ,
         dpath_mulcore_ps[69] , dpath_mulcore_ps[68] ,
         dpath_mulcore_ps[67] , dpath_mulcore_ps[66] ,
         dpath_mulcore_ps[65] , dpath_mulcore_ps[64] ,
         dpath_mulcore_ps[63] , dpath_mulcore_ps[62] ,
         dpath_mulcore_ps[61] , dpath_mulcore_ps[60] ,
         dpath_mulcore_ps[59] , dpath_mulcore_ps[58] ,
         dpath_mulcore_ps[57] , dpath_mulcore_ps[56] ,
         dpath_mulcore_ps[55] , dpath_mulcore_ps[54] ,
         dpath_mulcore_ps[53] , dpath_mulcore_ps[52] ,
         dpath_mulcore_ps[51] , dpath_mulcore_ps[50] ,
         dpath_mulcore_ps[49] , dpath_mulcore_ps[48] ,
         dpath_mulcore_ps[47] , dpath_mulcore_ps[46] ,
         dpath_mulcore_ps[45] , dpath_mulcore_ps[44] ,
         dpath_mulcore_ps[43] , dpath_mulcore_ps[42] ,
         dpath_mulcore_ps[41] , dpath_mulcore_ps[40] ,
         dpath_mulcore_ps[39] , dpath_mulcore_ps[38] ,
         dpath_mulcore_ps[37] , dpath_mulcore_ps[36] ,
         dpath_mulcore_ps[35] , dpath_mulcore_ps[34] ,
         dpath_mulcore_ps[33] , dpath_mulcore_ps[32] ,
         dpath_mulcore_ps[31] , dpath_mulcore_pc[97] ,
         dpath_mulcore_pc[96] , dpath_mulcore_pc[95] ,
         dpath_mulcore_pc[94] , dpath_mulcore_pc[93] ,
         dpath_mulcore_pc[92] , dpath_mulcore_pc[91] ,
         dpath_mulcore_pc[90] , dpath_mulcore_pc[89] ,
         dpath_mulcore_pc[88] , dpath_mulcore_pc[87] ,
         dpath_mulcore_pc[86] , dpath_mulcore_pc[85] ,
         dpath_mulcore_pc[84] , dpath_mulcore_pc[83] ,
         dpath_mulcore_pc[82] , dpath_mulcore_pc[81] ,
         dpath_mulcore_pc[80] , dpath_mulcore_pc[79] ,
         dpath_mulcore_pc[78] , dpath_mulcore_pc[77] ,
         dpath_mulcore_pc[76] , dpath_mulcore_pc[75] ,
         dpath_mulcore_pc[74] , dpath_mulcore_pc[73] ,
         dpath_mulcore_pc[72] , dpath_mulcore_pc[71] ,
         dpath_mulcore_pc[70] , dpath_mulcore_pc[69] ,
         dpath_mulcore_pc[68] , dpath_mulcore_pc[67] ,
         dpath_mulcore_pc[66] , dpath_mulcore_pc[65] ,
         dpath_mulcore_pc[64] , dpath_mulcore_pc[63] ,
         dpath_mulcore_pc[62] , dpath_mulcore_pc[61] ,
         dpath_mulcore_pc[60] , dpath_mulcore_pc[59] ,
         dpath_mulcore_pc[58] , dpath_mulcore_pc[57] ,
         dpath_mulcore_pc[56] , dpath_mulcore_pc[55] ,
         dpath_mulcore_pc[54] , dpath_mulcore_pc[53] ,
         dpath_mulcore_pc[52] , dpath_mulcore_pc[51] ,
         dpath_mulcore_pc[50] , dpath_mulcore_pc[49] ,
         dpath_mulcore_pc[48] , dpath_mulcore_pc[47] ,
         dpath_mulcore_pc[46] , dpath_mulcore_pc[45] ,
         dpath_mulcore_pc[44] , dpath_mulcore_pc[43] ,
         dpath_mulcore_pc[42] , dpath_mulcore_pc[41] ,
         dpath_mulcore_pc[40] , dpath_mulcore_pc[39] ,
         dpath_mulcore_pc[38] , dpath_mulcore_pc[37] ,
         dpath_mulcore_pc[36] , dpath_mulcore_pc[35] ,
         dpath_mulcore_pc[34] , dpath_mulcore_pc[33] ,
         dpath_mulcore_pc[32] , dpath_mulcore_pc[31] ,
         dpath_mulcore_pc[30] , dpath_mulcore_psum[0] ,
         dpath_mulcore_psum[1] , dpath_mulcore_psum[2] ,
         dpath_mulcore_psum[3] , dpath_mulcore_psum[4] ,
         dpath_mulcore_psum[5] , dpath_mulcore_psum[6] ,
         dpath_mulcore_psum[7] , dpath_mulcore_psum[8] ,
         dpath_mulcore_psum[9] , dpath_mulcore_psum[10] ,
         dpath_mulcore_psum[11] , dpath_mulcore_psum[12] ,
         dpath_mulcore_psum[13] , dpath_mulcore_psum[14] ,
         dpath_mulcore_psum[16] , dpath_mulcore_psum[17] ,
         dpath_mulcore_psum[18] , dpath_mulcore_psum[19] ,
         dpath_mulcore_psum[20] , dpath_mulcore_psum[21] ,
         dpath_mulcore_psum[22] , dpath_mulcore_psum[23] ,
         dpath_mulcore_psum[24] , dpath_mulcore_psum[25] ,
         dpath_mulcore_psum[26] , dpath_mulcore_psum[27] ,
         dpath_mulcore_psum[28] , dpath_mulcore_psum[29] ,
         dpath_mulcore_psum[30] , dpath_mulcore_psum[31] ,
         dpath_mulcore_psum[32] , dpath_mulcore_psum[33] ,
         dpath_mulcore_psum[34] , dpath_mulcore_psum[35] ,
         dpath_mulcore_psum[36] , dpath_mulcore_psum[37] ,
         dpath_mulcore_psum[38] , dpath_mulcore_psum[39] ,
         dpath_mulcore_psum[40] , dpath_mulcore_psum[41] ,
         dpath_mulcore_psum[42] , dpath_mulcore_psum[43] ,
         dpath_mulcore_psum[44] , dpath_mulcore_psum[45] ,
         dpath_mulcore_psum[46] , dpath_mulcore_psum[47] ,
         dpath_mulcore_psum[48] , dpath_mulcore_psum[49] ,
         dpath_mulcore_psum[50] , dpath_mulcore_psum[51] ,
         dpath_mulcore_psum[52] , dpath_mulcore_psum[53] ,
         dpath_mulcore_psum[54] , dpath_mulcore_psum[55] ,
         dpath_mulcore_psum[56] , dpath_mulcore_psum[57] ,
         dpath_mulcore_psum[58] , dpath_mulcore_psum[59] ,
         dpath_mulcore_psum[60] , dpath_mulcore_psum[61] ,
         dpath_mulcore_psum[62] , dpath_mulcore_psum[63] ,
         dpath_mulcore_psum[64] , dpath_mulcore_psum[65] ,
         dpath_mulcore_psum[66] , dpath_mulcore_psum[67] ,
         dpath_mulcore_psum[68] , dpath_mulcore_psum[69] ,
         dpath_mulcore_psum[70] , dpath_mulcore_psum[71] ,
         dpath_mulcore_psum[72] , dpath_mulcore_psum[73] ,
         dpath_mulcore_psum[74] , dpath_mulcore_psum[75] ,
         dpath_mulcore_psum[76] , dpath_mulcore_psum[77] ,
         dpath_mulcore_psum[78] , dpath_mulcore_psum[79] ,
         dpath_mulcore_psum[80] , dpath_mulcore_psum[81] ,
         dpath_mulcore_psum[82] , dpath_mulcore_psum[83] ,
         dpath_mulcore_psum[84] , dpath_mulcore_psum[85] ,
         dpath_mulcore_psum[86] , dpath_mulcore_psum[87] ,
         dpath_mulcore_psum[88] , dpath_mulcore_psum[89] ,
         dpath_mulcore_psum[90] , dpath_mulcore_psum[91] ,
         dpath_mulcore_psum[92] , dpath_mulcore_psum[93] ,
         dpath_mulcore_psum[94] , dpath_mulcore_psum[95] ,
         dpath_mulcore_psum[96] , dpath_mulcore_psum[97] ,
         dpath_mulcore_psum[98] , dpath_mulcore_pcout[0] ,
         dpath_mulcore_pcout[1] , dpath_mulcore_pcout[2] ,
         dpath_mulcore_pcout[3] , dpath_mulcore_pcout[4] ,
         dpath_mulcore_pcout[5] , dpath_mulcore_pcout[6] ,
         dpath_mulcore_pcout[7] , dpath_mulcore_pcout[8] ,
         dpath_mulcore_pcout[9] , dpath_mulcore_pcout[10] ,
         dpath_mulcore_pcout[11] , dpath_mulcore_pcout[12] ,
         dpath_mulcore_pcout[13] , dpath_mulcore_pcout[14] ,
         dpath_mulcore_pcout[16] , dpath_mulcore_pcout[17] ,
         dpath_mulcore_pcout[18] , dpath_mulcore_pcout[19] ,
         dpath_mulcore_pcout[20] , dpath_mulcore_pcout[21] ,
         dpath_mulcore_pcout[22] , dpath_mulcore_pcout[23] ,
         dpath_mulcore_pcout[24] , dpath_mulcore_pcout[25] ,
         dpath_mulcore_pcout[26] , dpath_mulcore_pcout[27] ,
         dpath_mulcore_pcout[28] , dpath_mulcore_pcout[29] ,
         dpath_mulcore_pcout[30] , dpath_mulcore_pcout[31] ,
         dpath_mulcore_pcout[32] , dpath_mulcore_pcout[33] ,
         dpath_mulcore_pcout[34] , dpath_mulcore_pcout[35] ,
         dpath_mulcore_pcout[36] , dpath_mulcore_pcout[37] ,
         dpath_mulcore_pcout[38] , dpath_mulcore_pcout[39] ,
         dpath_mulcore_pcout[40] , dpath_mulcore_pcout[41] ,
         dpath_mulcore_pcout[42] , dpath_mulcore_pcout[43] ,
         dpath_mulcore_pcout[44] , dpath_mulcore_pcout[45] ,
         dpath_mulcore_pcout[46] , dpath_mulcore_pcout[47] ,
         dpath_mulcore_pcout[48] , dpath_mulcore_pcout[49] ,
         dpath_mulcore_pcout[50] , dpath_mulcore_pcout[51] ,
         dpath_mulcore_pcout[52] , dpath_mulcore_pcout[53] ,
         dpath_mulcore_pcout[54] , dpath_mulcore_pcout[55] ,
         dpath_mulcore_pcout[56] , dpath_mulcore_pcout[57] ,
         dpath_mulcore_pcout[58] , dpath_mulcore_pcout[59] ,
         dpath_mulcore_pcout[60] , dpath_mulcore_pcout[61] ,
         dpath_mulcore_pcout[62] , dpath_mulcore_pcout[63] ,
         dpath_mulcore_pcout[64] , dpath_mulcore_pcout[65] ,
         dpath_mulcore_pcout[66] , dpath_mulcore_pcout[67] ,
         dpath_mulcore_pcout[68] , dpath_mulcore_pcout[69] ,
         dpath_mulcore_pcout[70] , dpath_mulcore_pcout[71] ,
         dpath_mulcore_pcout[72] , dpath_mulcore_pcout[73] ,
         dpath_mulcore_pcout[74] , dpath_mulcore_pcout[75] ,
         dpath_mulcore_pcout[76] , dpath_mulcore_pcout[77] ,
         dpath_mulcore_pcout[78] , dpath_mulcore_pcout[79] ,
         dpath_mulcore_pcout[80] , dpath_mulcore_pcout[81] ,
         dpath_mulcore_pcout[82] , dpath_mulcore_pcout[83] ,
         dpath_mulcore_pcout[84] , dpath_mulcore_pcout[85] ,
         dpath_mulcore_pcout[86] , dpath_mulcore_pcout[87] ,
         dpath_mulcore_pcout[88] , dpath_mulcore_pcout[89] ,
         dpath_mulcore_pcout[90] , dpath_mulcore_pcout[91] ,
         dpath_mulcore_pcout[92] , dpath_mulcore_pcout[93] ,
         dpath_mulcore_pcout[94] , dpath_mulcore_pcout[95] ,
         dpath_mulcore_pcout[96] , dpath_mulcore_pcout[97] ,
         dpath_mulcore_psumx2 , dpath_mulcore_pcoutx2 ,
         dpath_mulcore_a1s[81] , dpath_mulcore_a1s[80] ,
         dpath_mulcore_a1s[79] , dpath_mulcore_a1s[78] ,
         dpath_mulcore_a1s[77] , dpath_mulcore_a1s[76] ,
         dpath_mulcore_a1s[75] , dpath_mulcore_a1s[74] ,
         dpath_mulcore_a1s[73] , dpath_mulcore_a1s[72] ,
         dpath_mulcore_a1s[71] , dpath_mulcore_a1s[70] ,
         dpath_mulcore_a1s[69] , dpath_mulcore_a1s[68] ,
         dpath_mulcore_a1s[67] , dpath_mulcore_a1s[66] ,
         dpath_mulcore_a1s[65] , dpath_mulcore_a1s[64] ,
         dpath_mulcore_a1s[63] , dpath_mulcore_a1s[62] ,
         dpath_mulcore_a1s[61] , dpath_mulcore_a1s[60] ,
         dpath_mulcore_a1s[59] , dpath_mulcore_a1s[58] ,
         dpath_mulcore_a1s[57] , dpath_mulcore_a1s[56] ,
         dpath_mulcore_a1s[55] , dpath_mulcore_a1s[54] ,
         dpath_mulcore_a1s[53] , dpath_mulcore_a1s[52] ,
         dpath_mulcore_a1s[51] , dpath_mulcore_a1s[50] ,
         dpath_mulcore_a1s[49] , dpath_mulcore_a1s[48] ,
         dpath_mulcore_a1s[47] , dpath_mulcore_a1s[46] ,
         dpath_mulcore_a1s[45] , dpath_mulcore_a1s[44] ,
         dpath_mulcore_a1s[43] , dpath_mulcore_a1s[42] ,
         dpath_mulcore_a1s[41] , dpath_mulcore_a1s[40] ,
         dpath_mulcore_a1s[39] , dpath_mulcore_a1s[38] ,
         dpath_mulcore_a1s[37] , dpath_mulcore_a1s[36] ,
         dpath_mulcore_a1s[35] , dpath_mulcore_a1s[34] ,
         dpath_mulcore_a1s[33] , dpath_mulcore_a1s[32] ,
         dpath_mulcore_a1s[31] , dpath_mulcore_a1s[30] ,
         dpath_mulcore_a1s[29] , dpath_mulcore_a1s[28] ,
         dpath_mulcore_a1s[27] , dpath_mulcore_a1s[26] ,
         dpath_mulcore_a1s[25] , dpath_mulcore_a1s[24] ,
         dpath_mulcore_a1s[23] , dpath_mulcore_a1s[22] ,
         dpath_mulcore_a1s[21] , dpath_mulcore_a1s[20] ,
         dpath_mulcore_a1s[19] , dpath_mulcore_a1s[18] ,
         dpath_mulcore_a1s[17] , dpath_mulcore_a1s[16] ,
         dpath_mulcore_a1s[15] , dpath_mulcore_a1s[14] ,
         dpath_mulcore_a1s[13] , dpath_mulcore_a1s[12] ,
         dpath_mulcore_a1s[11] , dpath_mulcore_a1s[10] ,
         dpath_mulcore_a1s[9] , dpath_mulcore_a1s[8] ,
         dpath_mulcore_a1s[7] , dpath_mulcore_a1s[6] ,
         dpath_mulcore_a1s[5] , dpath_mulcore_a1s[4] ,
         dpath_mulcore_a1s[3] , dpath_mulcore_a1s[2] ,
         dpath_mulcore_a1s[1] , dpath_mulcore_a1s[0] ,
         dpath_mulcore_a1c[80] , dpath_mulcore_a1c[79] ,
         dpath_mulcore_a1c[78] , dpath_mulcore_a1c[77] ,
         dpath_mulcore_a1c[76] , dpath_mulcore_a1c[75] ,
         dpath_mulcore_a1c[74] , dpath_mulcore_a1c[73] ,
         dpath_mulcore_a1c[72] , dpath_mulcore_a1c[71] ,
         dpath_mulcore_a1c[70] , dpath_mulcore_a1c[69] ,
         dpath_mulcore_a1c[68] , dpath_mulcore_a1c[67] ,
         dpath_mulcore_a1c[66] , dpath_mulcore_a1c[65] ,
         dpath_mulcore_a1c[64] , dpath_mulcore_a1c[63] ,
         dpath_mulcore_a1c[62] , dpath_mulcore_a1c[61] ,
         dpath_mulcore_a1c[60] , dpath_mulcore_a1c[59] ,
         dpath_mulcore_a1c[58] , dpath_mulcore_a1c[57] ,
         dpath_mulcore_a1c[56] , dpath_mulcore_a1c[55] ,
         dpath_mulcore_a1c[54] , dpath_mulcore_a1c[53] ,
         dpath_mulcore_a1c[52] , dpath_mulcore_a1c[51] ,
         dpath_mulcore_a1c[50] , dpath_mulcore_a1c[49] ,
         dpath_mulcore_a1c[48] , dpath_mulcore_a1c[47] ,
         dpath_mulcore_a1c[46] , dpath_mulcore_a1c[45] ,
         dpath_mulcore_a1c[44] , dpath_mulcore_a1c[43] ,
         dpath_mulcore_a1c[42] , dpath_mulcore_a1c[41] ,
         dpath_mulcore_a1c[40] , dpath_mulcore_a1c[39] ,
         dpath_mulcore_a1c[38] , dpath_mulcore_a1c[37] ,
         dpath_mulcore_a1c[36] , dpath_mulcore_a1c[35] ,
         dpath_mulcore_a1c[34] , dpath_mulcore_a1c[33] ,
         dpath_mulcore_a1c[32] , dpath_mulcore_a1c[31] ,
         dpath_mulcore_a1c[30] , dpath_mulcore_a1c[29] ,
         dpath_mulcore_a1c[28] , dpath_mulcore_a1c[27] ,
         dpath_mulcore_a1c[26] , dpath_mulcore_a1c[25] ,
         dpath_mulcore_a1c[24] , dpath_mulcore_a1c[23] ,
         dpath_mulcore_a1c[22] , dpath_mulcore_a1c[21] ,
         dpath_mulcore_a1c[20] , dpath_mulcore_a1c[19] ,
         dpath_mulcore_a1c[18] , dpath_mulcore_a1c[17] ,
         dpath_mulcore_a1c[16] , dpath_mulcore_a1c[15] ,
         dpath_mulcore_a1c[14] , dpath_mulcore_a1c[13] ,
         dpath_mulcore_a1c[12] , dpath_mulcore_a1c[11] ,
         dpath_mulcore_a1c[10] , dpath_mulcore_a1c[9] ,
         dpath_mulcore_a1c[8] , dpath_mulcore_a1c[7] ,
         dpath_mulcore_a1c[6] , dpath_mulcore_a1c[5] ,
         dpath_mulcore_a1c[4] , dpath_mulcore_a1sum[79] ,
         dpath_mulcore_a1sum[78] , dpath_mulcore_a1sum[77] ,
         dpath_mulcore_a1sum[76] , dpath_mulcore_a1sum[75] ,
         dpath_mulcore_a1sum[74] , dpath_mulcore_a1sum[73] ,
         dpath_mulcore_a1sum[72] , dpath_mulcore_a1sum[71] ,
         dpath_mulcore_a1sum[70] , dpath_mulcore_a1sum[69] ,
         dpath_mulcore_a1sum[68] , dpath_mulcore_a1sum[67] ,
         dpath_mulcore_a1sum[66] , dpath_mulcore_a1sum[65] ,
         dpath_mulcore_a1sum[64] , dpath_mulcore_a1sum[63] ,
         dpath_mulcore_a1sum[62] , dpath_mulcore_a1sum[61] ,
         dpath_mulcore_a1sum[60] , dpath_mulcore_a1sum[59] ,
         dpath_mulcore_a1sum[58] , dpath_mulcore_a1sum[57] ,
         dpath_mulcore_a1sum[56] , dpath_mulcore_a1sum[55] ,
         dpath_mulcore_a1sum[54] , dpath_mulcore_a1sum[53] ,
         dpath_mulcore_a1sum[52] , dpath_mulcore_a1sum[51] ,
         dpath_mulcore_a1sum[50] , dpath_mulcore_a1sum[49] ,
         dpath_mulcore_a1sum[48] , dpath_mulcore_a1sum[47] ,
         dpath_mulcore_a1sum[46] , dpath_mulcore_a1sum[45] ,
         dpath_mulcore_a1sum[44] , dpath_mulcore_a1sum[43] ,
         dpath_mulcore_a1sum[42] , dpath_mulcore_a1sum[41] ,
         dpath_mulcore_a1sum[40] , dpath_mulcore_a1sum[39] ,
         dpath_mulcore_a1sum[38] , dpath_mulcore_a1sum[37] ,
         dpath_mulcore_a1sum[36] , dpath_mulcore_a1sum[35] ,
         dpath_mulcore_a1sum[34] , dpath_mulcore_a1sum[33] ,
         dpath_mulcore_a1sum[32] , dpath_mulcore_a1sum[31] ,
         dpath_mulcore_a1sum[30] , dpath_mulcore_a1sum[29] ,
         dpath_mulcore_a1sum[28] , dpath_mulcore_a1sum[27] ,
         dpath_mulcore_a1sum[26] , dpath_mulcore_a1sum[25] ,
         dpath_mulcore_a1sum[24] , dpath_mulcore_a1sum[23] ,
         dpath_mulcore_a1sum[22] , dpath_mulcore_a1sum[21] ,
         dpath_mulcore_a1sum[20] , dpath_mulcore_a1sum[19] ,
         dpath_mulcore_a1sum[18] , dpath_mulcore_a1sum[17] ,
         dpath_mulcore_a1sum[16] , dpath_mulcore_a1sum[15] ,
         dpath_mulcore_a1sum[14] , dpath_mulcore_a1sum[13] ,
         dpath_mulcore_a1sum[12] , dpath_mulcore_a1sum[10] ,
         dpath_mulcore_a1sum[9] , dpath_mulcore_a1sum[8] ,
         dpath_mulcore_a1sum[7] , dpath_mulcore_a1sum[6] ,
         dpath_mulcore_a1sum[5] , dpath_mulcore_a1sum[4] ,
         dpath_mulcore_a1sum[3] , dpath_mulcore_a1sum[2] ,
         dpath_mulcore_a1sum[1] , dpath_mulcore_a1sum[0] ,
         dpath_mulcore_a1cout[79] , dpath_mulcore_a1cout[78] ,
         dpath_mulcore_a1cout[77] , dpath_mulcore_a1cout[76] ,
         dpath_mulcore_a1cout[75] , dpath_mulcore_a1cout[74] ,
         dpath_mulcore_a1cout[73] , dpath_mulcore_a1cout[72] ,
         dpath_mulcore_a1cout[71] , dpath_mulcore_a1cout[70] ,
         dpath_mulcore_a1cout[69] , dpath_mulcore_a1cout[68] ,
         dpath_mulcore_a1cout[67] , dpath_mulcore_a1cout[66] ,
         dpath_mulcore_a1cout[65] , dpath_mulcore_a1cout[64] ,
         dpath_mulcore_a1cout[63] , dpath_mulcore_a1cout[62] ,
         dpath_mulcore_a1cout[61] , dpath_mulcore_a1cout[60] ,
         dpath_mulcore_a1cout[59] , dpath_mulcore_a1cout[58] ,
         dpath_mulcore_a1cout[57] , dpath_mulcore_a1cout[56] ,
         dpath_mulcore_a1cout[55] , dpath_mulcore_a1cout[54] ,
         dpath_mulcore_a1cout[53] , dpath_mulcore_a1cout[52] ,
         dpath_mulcore_a1cout[51] , dpath_mulcore_a1cout[50] ,
         dpath_mulcore_a1cout[49] , dpath_mulcore_a1cout[48] ,
         dpath_mulcore_a1cout[47] , dpath_mulcore_a1cout[46] ,
         dpath_mulcore_a1cout[45] , dpath_mulcore_a1cout[44] ,
         dpath_mulcore_a1cout[43] , dpath_mulcore_a1cout[42] ,
         dpath_mulcore_a1cout[41] , dpath_mulcore_a1cout[40] ,
         dpath_mulcore_a1cout[39] , dpath_mulcore_a1cout[38] ,
         dpath_mulcore_a1cout[37] , dpath_mulcore_a1cout[36] ,
         dpath_mulcore_a1cout[35] , dpath_mulcore_a1cout[34] ,
         dpath_mulcore_a1cout[33] , dpath_mulcore_a1cout[32] ,
         dpath_mulcore_a1cout[31] , dpath_mulcore_a1cout[30] ,
         dpath_mulcore_a1cout[29] , dpath_mulcore_a1cout[28] ,
         dpath_mulcore_a1cout[27] , dpath_mulcore_a1cout[26] ,
         dpath_mulcore_a1cout[25] , dpath_mulcore_a1cout[24] ,
         dpath_mulcore_a1cout[23] , dpath_mulcore_a1cout[22] ,
         dpath_mulcore_a1cout[21] , dpath_mulcore_a1cout[20] ,
         dpath_mulcore_a1cout[19] , dpath_mulcore_a1cout[18] ,
         dpath_mulcore_a1cout[17] , dpath_mulcore_a1cout[16] ,
         dpath_mulcore_a1cout[15] , dpath_mulcore_a1cout[14] ,
         dpath_mulcore_a1cout[13] , dpath_mulcore_a1cout[12] ,
         dpath_mulcore_a1cout[10] , dpath_mulcore_a1cout[9] ,
         dpath_mulcore_a1cout[8] , dpath_mulcore_a1cout[7] ,
         dpath_mulcore_a1cout[6] , dpath_mulcore_a1cout[5] ,
         dpath_mulcore_a1cout[4] , dpath_mulcore_a0s[80] ,
         dpath_mulcore_a0s[79] , dpath_mulcore_a0s[78] ,
         dpath_mulcore_a0s[77] , dpath_mulcore_a0s[76] ,
         dpath_mulcore_a0s[75] , dpath_mulcore_a0s[74] ,
         dpath_mulcore_a0s[73] , dpath_mulcore_a0s[72] ,
         dpath_mulcore_a0s[71] , dpath_mulcore_a0s[70] ,
         dpath_mulcore_a0s[69] , dpath_mulcore_a0s[68] ,
         dpath_mulcore_a0s[67] , dpath_mulcore_a0s[66] ,
         dpath_mulcore_a0s[65] , dpath_mulcore_a0s[64] ,
         dpath_mulcore_a0s[63] , dpath_mulcore_a0s[62] ,
         dpath_mulcore_a0s[61] , dpath_mulcore_a0s[60] ,
         dpath_mulcore_a0s[59] , dpath_mulcore_a0s[58] ,
         dpath_mulcore_a0s[57] , dpath_mulcore_a0s[56] ,
         dpath_mulcore_a0s[55] , dpath_mulcore_a0s[54] ,
         dpath_mulcore_a0s[53] , dpath_mulcore_a0s[52] ,
         dpath_mulcore_a0s[51] , dpath_mulcore_a0s[50] ,
         dpath_mulcore_a0s[49] , dpath_mulcore_a0s[48] ,
         dpath_mulcore_a0s[47] , dpath_mulcore_a0s[46] ,
         dpath_mulcore_a0s[45] , dpath_mulcore_a0s[44] ,
         dpath_mulcore_a0s[43] , dpath_mulcore_a0s[42] ,
         dpath_mulcore_a0s[41] , dpath_mulcore_a0s[40] ,
         dpath_mulcore_a0s[39] , dpath_mulcore_a0s[38] ,
         dpath_mulcore_a0s[37] , dpath_mulcore_a0s[36] ,
         dpath_mulcore_a0s[35] , dpath_mulcore_a0s[34] ,
         dpath_mulcore_a0s[33] , dpath_mulcore_a0s[32] ,
         dpath_mulcore_a0s[31] , dpath_mulcore_a0s[30] ,
         dpath_mulcore_a0s[29] , dpath_mulcore_a0s[28] ,
         dpath_mulcore_a0s[27] , dpath_mulcore_a0s[26] ,
         dpath_mulcore_a0s[25] , dpath_mulcore_a0s[24] ,
         dpath_mulcore_a0s[23] , dpath_mulcore_a0s[22] ,
         dpath_mulcore_a0s[21] , dpath_mulcore_a0s[20] ,
         dpath_mulcore_a0s[19] , dpath_mulcore_a0s[18] ,
         dpath_mulcore_a0s[17] , dpath_mulcore_a0s[16] ,
         dpath_mulcore_a0s[15] , dpath_mulcore_a0s[14] ,
         dpath_mulcore_a0s[13] , dpath_mulcore_a0s[12] ,
         dpath_mulcore_a0s[11] , dpath_mulcore_a0s[10] ,
         dpath_mulcore_a0s[9] , dpath_mulcore_a0s[8] ,
         dpath_mulcore_a0s[7] , dpath_mulcore_a0s[6] ,
         dpath_mulcore_a0s[5] , dpath_mulcore_a0s[4] ,
         dpath_mulcore_a0s[3] , dpath_mulcore_a0s[2] ,
         dpath_mulcore_a0s[1] , dpath_mulcore_a0s[0] ,
         dpath_mulcore_a0c[79] , dpath_mulcore_a0c[78] ,
         dpath_mulcore_a0c[77] , dpath_mulcore_a0c[76] ,
         dpath_mulcore_a0c[75] , dpath_mulcore_a0c[74] ,
         dpath_mulcore_a0c[73] , dpath_mulcore_a0c[72] ,
         dpath_mulcore_a0c[71] , dpath_mulcore_a0c[70] ,
         dpath_mulcore_a0c[69] , dpath_mulcore_a0c[68] ,
         dpath_mulcore_a0c[67] , dpath_mulcore_a0c[66] ,
         dpath_mulcore_a0c[65] , dpath_mulcore_a0c[64] ,
         dpath_mulcore_a0c[63] , dpath_mulcore_a0c[62] ,
         dpath_mulcore_a0c[61] , dpath_mulcore_a0c[60] ,
         dpath_mulcore_a0c[59] , dpath_mulcore_a0c[58] ,
         dpath_mulcore_a0c[57] , dpath_mulcore_a0c[56] ,
         dpath_mulcore_a0c[55] , dpath_mulcore_a0c[54] ,
         dpath_mulcore_a0c[53] , dpath_mulcore_a0c[52] ,
         dpath_mulcore_a0c[51] , dpath_mulcore_a0c[50] ,
         dpath_mulcore_a0c[49] , dpath_mulcore_a0c[48] ,
         dpath_mulcore_a0c[47] , dpath_mulcore_a0c[46] ,
         dpath_mulcore_a0c[45] , dpath_mulcore_a0c[44] ,
         dpath_mulcore_a0c[43] , dpath_mulcore_a0c[42] ,
         dpath_mulcore_a0c[41] , dpath_mulcore_a0c[40] ,
         dpath_mulcore_a0c[39] , dpath_mulcore_a0c[38] ,
         dpath_mulcore_a0c[37] , dpath_mulcore_a0c[36] ,
         dpath_mulcore_a0c[35] , dpath_mulcore_a0c[34] ,
         dpath_mulcore_a0c[33] , dpath_mulcore_a0c[32] ,
         dpath_mulcore_a0c[31] , dpath_mulcore_a0c[30] ,
         dpath_mulcore_a0c[29] , dpath_mulcore_a0c[28] ,
         dpath_mulcore_a0c[27] , dpath_mulcore_a0c[26] ,
         dpath_mulcore_a0c[25] , dpath_mulcore_a0c[24] ,
         dpath_mulcore_a0c[23] , dpath_mulcore_a0c[22] ,
         dpath_mulcore_a0c[21] , dpath_mulcore_a0c[20] ,
         dpath_mulcore_a0c[19] , dpath_mulcore_a0c[18] ,
         dpath_mulcore_a0c[17] , dpath_mulcore_a0c[16] ,
         dpath_mulcore_a0c[15] , dpath_mulcore_a0c[14] ,
         dpath_mulcore_a0c[13] , dpath_mulcore_a0c[12] ,
         dpath_mulcore_a0c[11] , dpath_mulcore_a0c[10] ,
         dpath_mulcore_a0c[9] , dpath_mulcore_a0c[8] ,
         dpath_mulcore_a0c[7] , dpath_mulcore_a0c[6] ,
         dpath_mulcore_a0c[5] , dpath_mulcore_a0c[4] ,
         dpath_mulcore_a0sum[79] , dpath_mulcore_a0sum[78] ,
         dpath_mulcore_a0sum[77] , dpath_mulcore_a0sum[76] ,
         dpath_mulcore_a0sum[75] , dpath_mulcore_a0sum[74] ,
         dpath_mulcore_a0sum[73] , dpath_mulcore_a0sum[72] ,
         dpath_mulcore_a0sum[71] , dpath_mulcore_a0sum[70] ,
         dpath_mulcore_a0sum[69] , dpath_mulcore_a0sum[68] ,
         dpath_mulcore_a0sum[67] , dpath_mulcore_a0sum[66] ,
         dpath_mulcore_a0sum[65] , dpath_mulcore_a0sum[64] ,
         dpath_mulcore_a0sum[63] , dpath_mulcore_a0sum[62] ,
         dpath_mulcore_a0sum[61] , dpath_mulcore_a0sum[60] ,
         dpath_mulcore_a0sum[59] , dpath_mulcore_a0sum[58] ,
         dpath_mulcore_a0sum[57] , dpath_mulcore_a0sum[56] ,
         dpath_mulcore_a0sum[55] , dpath_mulcore_a0sum[54] ,
         dpath_mulcore_a0sum[53] , dpath_mulcore_a0sum[52] ,
         dpath_mulcore_a0sum[51] , dpath_mulcore_a0sum[50] ,
         dpath_mulcore_a0sum[49] , dpath_mulcore_a0sum[48] ,
         dpath_mulcore_a0sum[47] , dpath_mulcore_a0sum[46] ,
         dpath_mulcore_a0sum[45] , dpath_mulcore_a0sum[44] ,
         dpath_mulcore_a0sum[43] , dpath_mulcore_a0sum[42] ,
         dpath_mulcore_a0sum[41] , dpath_mulcore_a0sum[40] ,
         dpath_mulcore_a0sum[39] , dpath_mulcore_a0sum[38] ,
         dpath_mulcore_a0sum[37] , dpath_mulcore_a0sum[36] ,
         dpath_mulcore_a0sum[35] , dpath_mulcore_a0sum[34] ,
         dpath_mulcore_a0sum[33] , dpath_mulcore_a0sum[32] ,
         dpath_mulcore_a0sum[31] , dpath_mulcore_a0sum[30] ,
         dpath_mulcore_a0sum[29] , dpath_mulcore_a0sum[28] ,
         dpath_mulcore_a0sum[27] , dpath_mulcore_a0sum[26] ,
         dpath_mulcore_a0sum[25] , dpath_mulcore_a0sum[24] ,
         dpath_mulcore_a0sum[23] , dpath_mulcore_a0sum[22] ,
         dpath_mulcore_a0sum[21] , dpath_mulcore_a0sum[20] ,
         dpath_mulcore_a0sum[19] , dpath_mulcore_a0sum[18] ,
         dpath_mulcore_a0sum[17] , dpath_mulcore_a0sum[16] ,
         dpath_mulcore_a0sum[15] , dpath_mulcore_a0sum[14] ,
         dpath_mulcore_a0sum[13] , dpath_mulcore_a0sum[12] ,
         dpath_mulcore_a0sum[10] , dpath_mulcore_a0sum[9] ,
         dpath_mulcore_a0sum[8] , dpath_mulcore_a0sum[7] ,
         dpath_mulcore_a0sum[6] , dpath_mulcore_a0sum[5] ,
         dpath_mulcore_a0sum[4] , dpath_mulcore_a0sum[3] ,
         dpath_mulcore_a0sum[2] , dpath_mulcore_a0sum[1] ,
         dpath_mulcore_a0sum[0] , dpath_mulcore_a0cout[79] ,
         dpath_mulcore_a0cout[78] , dpath_mulcore_a0cout[77] ,
         dpath_mulcore_a0cout[76] , dpath_mulcore_a0cout[75] ,
         dpath_mulcore_a0cout[74] , dpath_mulcore_a0cout[73] ,
         dpath_mulcore_a0cout[72] , dpath_mulcore_a0cout[71] ,
         dpath_mulcore_a0cout[70] , dpath_mulcore_a0cout[69] ,
         dpath_mulcore_a0cout[68] , dpath_mulcore_a0cout[67] ,
         dpath_mulcore_a0cout[66] , dpath_mulcore_a0cout[65] ,
         dpath_mulcore_a0cout[64] , dpath_mulcore_a0cout[63] ,
         dpath_mulcore_a0cout[62] , dpath_mulcore_a0cout[61] ,
         dpath_mulcore_a0cout[60] , dpath_mulcore_a0cout[59] ,
         dpath_mulcore_a0cout[58] , dpath_mulcore_a0cout[57] ,
         dpath_mulcore_a0cout[56] , dpath_mulcore_a0cout[55] ,
         dpath_mulcore_a0cout[54] , dpath_mulcore_a0cout[53] ,
         dpath_mulcore_a0cout[52] , dpath_mulcore_a0cout[51] ,
         dpath_mulcore_a0cout[50] , dpath_mulcore_a0cout[49] ,
         dpath_mulcore_a0cout[48] , dpath_mulcore_a0cout[47] ,
         dpath_mulcore_a0cout[46] , dpath_mulcore_a0cout[45] ,
         dpath_mulcore_a0cout[44] , dpath_mulcore_a0cout[43] ,
         dpath_mulcore_a0cout[42] , dpath_mulcore_a0cout[41] ,
         dpath_mulcore_a0cout[40] , dpath_mulcore_a0cout[39] ,
         dpath_mulcore_a0cout[38] , dpath_mulcore_a0cout[37] ,
         dpath_mulcore_a0cout[36] , dpath_mulcore_a0cout[35] ,
         dpath_mulcore_a0cout[34] , dpath_mulcore_a0cout[33] ,
         dpath_mulcore_a0cout[32] , dpath_mulcore_a0cout[31] ,
         dpath_mulcore_a0cout[30] , dpath_mulcore_a0cout[29] ,
         dpath_mulcore_a0cout[28] , dpath_mulcore_a0cout[27] ,
         dpath_mulcore_a0cout[26] , dpath_mulcore_a0cout[25] ,
         dpath_mulcore_a0cout[24] , dpath_mulcore_a0cout[23] ,
         dpath_mulcore_a0cout[22] , dpath_mulcore_a0cout[21] ,
         dpath_mulcore_a0cout[20] , dpath_mulcore_a0cout[19] ,
         dpath_mulcore_a0cout[18] , dpath_mulcore_a0cout[17] ,
         dpath_mulcore_a0cout[16] , dpath_mulcore_a0cout[15] ,
         dpath_mulcore_a0cout[14] , dpath_mulcore_a0cout[13] ,
         dpath_mulcore_a0cout[12] , dpath_mulcore_a0cout[10] ,
         dpath_mulcore_a0cout[9] , dpath_mulcore_a0cout[8] ,
         dpath_mulcore_a0cout[7] , dpath_mulcore_a0cout[6] ,
         dpath_mulcore_a0cout[5] , dpath_mulcore_a0cout[4] ,
         dpath_mulcore_b16 , dpath_mulcore_b15[2] , dpath_mulcore_b15[1] ,
         dpath_mulcore_b15[0] , dpath_mulcore_b14[2] ,
         dpath_mulcore_b14[1] , dpath_mulcore_b14[0] ,
         dpath_mulcore_b13[2] , dpath_mulcore_b13[1] ,
         dpath_mulcore_b13[0] , dpath_mulcore_b12[2] ,
         dpath_mulcore_b12[1] , dpath_mulcore_b12[0] ,
         dpath_mulcore_b11[2] , dpath_mulcore_b11[1] ,
         dpath_mulcore_b11[0] , dpath_mulcore_b10[2] ,
         dpath_mulcore_b10[1] , dpath_mulcore_b10[0] , dpath_mulcore_b9[2] ,
         dpath_mulcore_b9[1] , dpath_mulcore_b9[0] , dpath_mulcore_b8[2] ,
         dpath_mulcore_b8[1] , dpath_mulcore_b8[0] , dpath_mulcore_b7[2] ,
         dpath_mulcore_b7[1] , dpath_mulcore_b7[0] , dpath_mulcore_b6[2] ,
         dpath_mulcore_b6[1] , dpath_mulcore_b6[0] , dpath_mulcore_b5[2] ,
         dpath_mulcore_b5[1] , dpath_mulcore_b5[0] , dpath_mulcore_b4[2] ,
         dpath_mulcore_b4[1] , dpath_mulcore_b4[0] , dpath_mulcore_b3[2] ,
         dpath_mulcore_b3[1] , dpath_mulcore_b3[0] , dpath_mulcore_b2[2] ,
         dpath_mulcore_b2[1] , dpath_mulcore_b2[0] , dpath_mulcore_b1[2] ,
         dpath_mulcore_b1[1] , dpath_mulcore_b1[0] , dpath_mulcore_b0[2] ,
         dpath_mulcore_b0[1] , dpath_mulcore_b0[0] ,
         dpath_mulcore_op1_l[63] , dpath_mulcore_op1_l[62] ,
         dpath_mulcore_op1_l[61] , dpath_mulcore_op1_l[60] ,
         dpath_mulcore_op1_l[59] , dpath_mulcore_op1_l[58] ,
         dpath_mulcore_op1_l[57] , dpath_mulcore_op1_l[56] ,
         dpath_mulcore_op1_l[55] , dpath_mulcore_op1_l[54] ,
         dpath_mulcore_op1_l[53] , dpath_mulcore_op1_l[52] ,
         dpath_mulcore_op1_l[51] , dpath_mulcore_op1_l[50] ,
         dpath_mulcore_op1_l[49] , dpath_mulcore_op1_l[48] ,
         dpath_mulcore_op1_l[47] , dpath_mulcore_op1_l[46] ,
         dpath_mulcore_op1_l[45] , dpath_mulcore_op1_l[44] ,
         dpath_mulcore_op1_l[43] , dpath_mulcore_op1_l[42] ,
         dpath_mulcore_op1_l[41] , dpath_mulcore_op1_l[40] ,
         dpath_mulcore_op1_l[39] , dpath_mulcore_op1_l[38] ,
         dpath_mulcore_op1_l[37] , dpath_mulcore_op1_l[36] ,
         dpath_mulcore_op1_l[35] , dpath_mulcore_op1_l[34] ,
         dpath_mulcore_op1_l[33] , dpath_mulcore_op1_l[32] ,
         dpath_mulcore_op1_l[31] , dpath_mulcore_op1_l[30] ,
         dpath_mulcore_op1_l[29] , dpath_mulcore_op1_l[28] ,
         dpath_mulcore_op1_l[27] , dpath_mulcore_op1_l[26] ,
         dpath_mulcore_op1_l[25] , dpath_mulcore_op1_l[24] ,
         dpath_mulcore_op1_l[23] , dpath_mulcore_op1_l[22] ,
         dpath_mulcore_op1_l[21] , dpath_mulcore_op1_l[20] ,
         dpath_mulcore_op1_l[19] , dpath_mulcore_op1_l[18] ,
         dpath_mulcore_op1_l[17] , dpath_mulcore_op1_l[16] ,
         dpath_mulcore_op1_l[15] , dpath_mulcore_op1_l[14] ,
         dpath_mulcore_op1_l[13] , dpath_mulcore_op1_l[12] ,
         dpath_mulcore_op1_l[11] , dpath_mulcore_op1_l[10] ,
         dpath_mulcore_op1_l[9] , dpath_mulcore_op1_l[8] ,
         dpath_mulcore_op1_l[7] , dpath_mulcore_op1_l[6] ,
         dpath_mulcore_op1_l[5] , dpath_mulcore_op1_l[4] ,
         dpath_mulcore_op1_l[3] , dpath_mulcore_op1_l[2] ,
         dpath_mulcore_op1_l[1] , dpath_mulcore_op1_l[0] ,
         dpath_mulcore_clk_enb1 , dpath_mulcore_x2_c2c3 ,
         dpath_mulcore_x2_c3 , dpath_mulcore_x2_c2 , dpath_mulcore_x2_c1 ,
         dpath_mulcore_cyc2 , dpath_mulcore_cyc1 , dpath_mulcore_clk_enb0 ,
         dpath_mulcore_rs1_l[0] , dpath_mulcore_rs1_l[1] ,
         dpath_mulcore_rs1_l[2] , dpath_mulcore_rs1_l[3] ,
         dpath_mulcore_rs1_l[4] , dpath_mulcore_rs1_l[5] ,
         dpath_mulcore_rs1_l[6] , dpath_mulcore_rs1_l[7] ,
         dpath_mulcore_rs1_l[8] , dpath_mulcore_rs1_l[9] ,
         dpath_mulcore_rs1_l[10] , dpath_mulcore_rs1_l[11] ,
         dpath_mulcore_rs1_l[12] , dpath_mulcore_rs1_l[13] ,
         dpath_mulcore_rs1_l[14] , dpath_mulcore_rs1_l[15] ,
         dpath_mulcore_rs1_l[16] , dpath_mulcore_rs1_l[17] ,
         dpath_mulcore_rs1_l[18] , dpath_mulcore_rs1_l[19] ,
         dpath_mulcore_rs1_l[20] , dpath_mulcore_rs1_l[21] ,
         dpath_mulcore_rs1_l[22] , dpath_mulcore_rs1_l[23] ,
         dpath_mulcore_rs1_l[24] , dpath_mulcore_rs1_l[25] ,
         dpath_mulcore_rs1_l[26] , dpath_mulcore_rs1_l[27] ,
         dpath_mulcore_rs1_l[28] , dpath_mulcore_rs1_l[29] ,
         dpath_mulcore_rs1_l[30] , dpath_mulcore_rs1_l[31] ,
         dpath_mulcore_rs1_l[32] , dpath_mulcore_rs1_l[33] ,
         dpath_mulcore_rs1_l[34] , dpath_mulcore_rs1_l[35] ,
         dpath_mulcore_rs1_l[36] , dpath_mulcore_rs1_l[37] ,
         dpath_mulcore_rs1_l[38] , dpath_mulcore_rs1_l[39] ,
         dpath_mulcore_rs1_l[40] , dpath_mulcore_rs1_l[41] ,
         dpath_mulcore_rs1_l[42] , dpath_mulcore_rs1_l[43] ,
         dpath_mulcore_rs1_l[44] , dpath_mulcore_rs1_l[45] ,
         dpath_mulcore_rs1_l[46] , dpath_mulcore_rs1_l[47] ,
         dpath_mulcore_rs1_l[48] , dpath_mulcore_rs1_l[49] ,
         dpath_mulcore_rs1_l[50] , dpath_mulcore_rs1_l[51] ,
         dpath_mulcore_rs1_l[52] , dpath_mulcore_rs1_l[53] ,
         dpath_mulcore_rs1_l[54] , dpath_mulcore_rs1_l[55] ,
         dpath_mulcore_rs1_l[56] , dpath_mulcore_rs1_l[57] ,
         dpath_mulcore_rs1_l[58] , dpath_mulcore_rs1_l[59] ,
         dpath_mulcore_rs1_l[60] , dpath_mulcore_rs1_l[61] ,
         dpath_mulcore_rs1_l[62] , dpath_mulcore_rs1_l[63] ,
         dpath_dffshf_n3 , dpath_accum_n273 , dpath_accum_n271 ,
         dpath_accum_n269 , dpath_accum_n267 , dpath_accum_n265 ,
         dpath_accum_n263 , dpath_accum_n261 , dpath_accum_n259 ,
         dpath_accum_n257 , dpath_accum_n255 , dpath_accum_n253 ,
         dpath_accum_n251 , dpath_accum_n249 , dpath_accum_n247 ,
         dpath_accum_n245 , dpath_accum_n243 , dpath_accum_n241 ,
         dpath_accum_n239 , dpath_accum_n237 , dpath_accum_n235 ,
         dpath_accum_n233 , dpath_accum_n231 , dpath_accum_n229 ,
         dpath_accum_n227 , dpath_accum_n225 , dpath_accum_n223 ,
         dpath_accum_n221 , dpath_accum_n219 , dpath_accum_n217 ,
         dpath_accum_n215 , dpath_accum_n213 , dpath_accum_n211 ,
         dpath_accum_n209 , dpath_accum_n207 , dpath_accum_n205 ,
         dpath_accum_n203 , dpath_accum_n201 , dpath_accum_n199 ,
         dpath_accum_n197 , dpath_accum_n195 , dpath_accum_n193 ,
         dpath_accum_n191 , dpath_accum_n189 , dpath_accum_n187 ,
         dpath_accum_n185 , dpath_accum_n183 , dpath_accum_n181 ,
         dpath_accum_n179 , dpath_accum_n177 , dpath_accum_n175 ,
         dpath_accum_n173 , dpath_accum_n171 , dpath_accum_n169 ,
         dpath_accum_n167 , dpath_accum_n165 , dpath_accum_n163 ,
         dpath_accum_n161 , dpath_accum_n159 , dpath_accum_n157 ,
         dpath_accum_n155 , dpath_accum_n153 , dpath_accum_n151 ,
         dpath_accum_n149 , dpath_accum_n147 , dpath_accum_n145 ,
         dpath_accum_n143 , dpath_accum_n141 , dpath_accum_n139 ,
         dpath_accum_n137 , dpath_accum_n135 , dpath_accum_n133 ,
         dpath_accum_n131 , dpath_accum_n129 , dpath_accum_n127 ,
         dpath_accum_n125 , dpath_accum_n123 , dpath_accum_n121 ,
         dpath_accum_n119 , dpath_accum_n117 , dpath_accum_n115 ,
         dpath_accum_n113 , dpath_accum_n111 , dpath_accum_n109 ,
         dpath_accum_n107 , dpath_accum_n105 , dpath_accum_n103 ,
         dpath_accum_n101 , dpath_accum_n99 , dpath_accum_n97 ,
         dpath_accum_n95 , dpath_accum_n93 , dpath_accum_n91 ,
         dpath_accum_n89 , dpath_accum_n87 , dpath_accum_n85 ,
         dpath_accum_n83 , dpath_accum_n81 , dpath_accum_n79 ,
         dpath_accum_n77 , dpath_accum_n75 , dpath_accum_n73 ,
         dpath_accum_n71 , dpath_accum_n69 , dpath_accum_n67 ,
         dpath_accum_n65 , dpath_accum_n63 , dpath_accum_n61 ,
         dpath_accum_n59 , dpath_accum_n57 , dpath_accum_n55 ,
         dpath_accum_n53 , dpath_accum_n51 , dpath_accum_n49 ,
         dpath_accum_n47 , dpath_accum_n45 , dpath_accum_n43 ,
         dpath_accum_n41 , dpath_accum_n39 , dpath_accum_n37 ,
         dpath_accum_n35 , dpath_accum_n33 , dpath_accum_n31 ,
         dpath_accum_n29 , dpath_accum_n27 , dpath_accum_n25 ,
         dpath_accum_n23 , dpath_accum_n21 , dpath_accum_n19 ,
         dpath_accum_n17 , dpath_accum_n15 , dpath_accum_n13 ,
         dpath_accum_n11 , dpath_accum_n9 , dpath_accum_n7 ,
         dpath_accum_n5 , dpath_accum_n3 , dpath_accum_n2 ,
         dpath_ckbuf_1_clken , dpath_ckbuf_1_N1 , dpath_ckbuf_1_enb_l ,
         dpath_mulcore_cyc1_dff_n3 , dpath_mulcore_cyc1_dff_n2 ,
         dpath_mulcore_ffrs1_n129 , dpath_mulcore_ffrs1_n127 ,
         dpath_mulcore_ffrs1_n125 , dpath_mulcore_ffrs1_n123 ,
         dpath_mulcore_ffrs1_n121 , dpath_mulcore_ffrs1_n119 ,
         dpath_mulcore_ffrs1_n117 , dpath_mulcore_ffrs1_n115 ,
         dpath_mulcore_ffrs1_n113 , dpath_mulcore_ffrs1_n111 ,
         dpath_mulcore_ffrs1_n109 , dpath_mulcore_ffrs1_n107 ,
         dpath_mulcore_ffrs1_n105 , dpath_mulcore_ffrs1_n103 ,
         dpath_mulcore_ffrs1_n101 , dpath_mulcore_ffrs1_n99 ,
         dpath_mulcore_ffrs1_n97 , dpath_mulcore_ffrs1_n95 ,
         dpath_mulcore_ffrs1_n93 , dpath_mulcore_ffrs1_n91 ,
         dpath_mulcore_ffrs1_n89 , dpath_mulcore_ffrs1_n87 ,
         dpath_mulcore_ffrs1_n85 , dpath_mulcore_ffrs1_n83 ,
         dpath_mulcore_ffrs1_n81 , dpath_mulcore_ffrs1_n79 ,
         dpath_mulcore_ffrs1_n77 , dpath_mulcore_ffrs1_n75 ,
         dpath_mulcore_ffrs1_n73 , dpath_mulcore_ffrs1_n71 ,
         dpath_mulcore_ffrs1_n69 , dpath_mulcore_ffrs1_n67 ,
         dpath_mulcore_ffrs1_n65 , dpath_mulcore_ffrs1_n63 ,
         dpath_mulcore_ffrs1_n61 , dpath_mulcore_ffrs1_n59 ,
         dpath_mulcore_ffrs1_n57 , dpath_mulcore_ffrs1_n55 ,
         dpath_mulcore_ffrs1_n53 , dpath_mulcore_ffrs1_n51 ,
         dpath_mulcore_ffrs1_n49 , dpath_mulcore_ffrs1_n47 ,
         dpath_mulcore_ffrs1_n45 , dpath_mulcore_ffrs1_n43 ,
         dpath_mulcore_ffrs1_n41 , dpath_mulcore_ffrs1_n39 ,
         dpath_mulcore_ffrs1_n37 , dpath_mulcore_ffrs1_n35 ,
         dpath_mulcore_ffrs1_n33 , dpath_mulcore_ffrs1_n31 ,
         dpath_mulcore_ffrs1_n29 , dpath_mulcore_ffrs1_n27 ,
         dpath_mulcore_ffrs1_n25 , dpath_mulcore_ffrs1_n23 ,
         dpath_mulcore_ffrs1_n21 , dpath_mulcore_ffrs1_n19 ,
         dpath_mulcore_ffrs1_n17 , dpath_mulcore_ffrs1_n15 ,
         dpath_mulcore_ffrs1_n13 , dpath_mulcore_ffrs1_n11 ,
         dpath_mulcore_ffrs1_n9 , dpath_mulcore_ffrs1_n7 ,
         dpath_mulcore_ffrs1_n5 , dpath_mulcore_ffrs1_n3 ,
         dpath_mulcore_booth_b15_outmx[2] ,
         dpath_mulcore_booth_b15_outmx[1] ,
         dpath_mulcore_booth_b15_outmx[0] ,
         dpath_mulcore_booth_b14_outmx[2] ,
         dpath_mulcore_booth_b14_outmx[1] ,
         dpath_mulcore_booth_b14_outmx[0] ,
         dpath_mulcore_booth_b13_outmx[2] ,
         dpath_mulcore_booth_b13_outmx[1] ,
         dpath_mulcore_booth_b13_outmx[0] ,
         dpath_mulcore_booth_b12_outmx[2] ,
         dpath_mulcore_booth_b12_outmx[1] ,
         dpath_mulcore_booth_b12_outmx[0] ,
         dpath_mulcore_booth_b11_outmx[2] ,
         dpath_mulcore_booth_b11_outmx[1] ,
         dpath_mulcore_booth_b11_outmx[0] ,
         dpath_mulcore_booth_b10_outmx[2] ,
         dpath_mulcore_booth_b10_outmx[1] ,
         dpath_mulcore_booth_b10_outmx[0] , dpath_mulcore_booth_b9_outmx[2] ,
         dpath_mulcore_booth_b9_outmx[1] , dpath_mulcore_booth_b9_outmx[0] ,
         dpath_mulcore_booth_b8_outmx[2] , dpath_mulcore_booth_b8_outmx[1] ,
         dpath_mulcore_booth_b8_outmx[0] , dpath_mulcore_booth_b7_outmx[2] ,
         dpath_mulcore_booth_b7_outmx[1] , dpath_mulcore_booth_b7_outmx[0] ,
         dpath_mulcore_booth_b6_outmx[2] , dpath_mulcore_booth_b6_outmx[1] ,
         dpath_mulcore_booth_b6_outmx[0] , dpath_mulcore_booth_b5_outmx[2] ,
         dpath_mulcore_booth_b5_outmx[1] , dpath_mulcore_booth_b5_outmx[0] ,
         dpath_mulcore_booth_b4_outmx[2] , dpath_mulcore_booth_b4_outmx[1] ,
         dpath_mulcore_booth_b4_outmx[0] , dpath_mulcore_booth_b3_outmx[2] ,
         dpath_mulcore_booth_b3_outmx[1] , dpath_mulcore_booth_b3_outmx[0] ,
         dpath_mulcore_booth_b2_outmx[2] , dpath_mulcore_booth_b2_outmx[1] ,
         dpath_mulcore_booth_b2_outmx[0] , dpath_mulcore_booth_b1_outmx[2] ,
         dpath_mulcore_booth_b1_outmx[1] , dpath_mulcore_booth_b1_outmx[0] ,
         dpath_mulcore_booth_b0_outmx[2] , dpath_mulcore_booth_b0_outmx[1] ,
         dpath_mulcore_booth_b0_outmx[0] , dpath_mulcore_booth_b15_in1[2] ,
         dpath_mulcore_booth_b15_in1[1] , dpath_mulcore_booth_b15_in1[0] ,
         dpath_mulcore_booth_b14_in1[2] , dpath_mulcore_booth_b14_in1[1] ,
         dpath_mulcore_booth_b14_in1[0] , dpath_mulcore_booth_b13_in1[2] ,
         dpath_mulcore_booth_b13_in1[1] , dpath_mulcore_booth_b13_in1[0] ,
         dpath_mulcore_booth_b12_in1[2] , dpath_mulcore_booth_b12_in1[1] ,
         dpath_mulcore_booth_b12_in1[0] , dpath_mulcore_booth_b11_in1[2] ,
         dpath_mulcore_booth_b11_in1[1] , dpath_mulcore_booth_b11_in1[0] ,
         dpath_mulcore_booth_b10_in1[2] , dpath_mulcore_booth_b10_in1[1] ,
         dpath_mulcore_booth_b10_in1[0] , dpath_mulcore_booth_b9_in1[2] ,
         dpath_mulcore_booth_b9_in1[1] , dpath_mulcore_booth_b9_in1[0] ,
         dpath_mulcore_booth_b8_in1[2] , dpath_mulcore_booth_b8_in1[1] ,
         dpath_mulcore_booth_b8_in1[0] , dpath_mulcore_booth_b7_in1[2] ,
         dpath_mulcore_booth_b7_in1[1] , dpath_mulcore_booth_b7_in1[0] ,
         dpath_mulcore_booth_b6_in1[2] , dpath_mulcore_booth_b6_in1[1] ,
         dpath_mulcore_booth_b6_in1[0] , dpath_mulcore_booth_b5_in1[2] ,
         dpath_mulcore_booth_b5_in1[1] , dpath_mulcore_booth_b5_in1[0] ,
         dpath_mulcore_booth_b4_in1[2] , dpath_mulcore_booth_b4_in1[1] ,
         dpath_mulcore_booth_b4_in1[0] , dpath_mulcore_booth_b3_in1[2] ,
         dpath_mulcore_booth_b3_in1[1] , dpath_mulcore_booth_b3_in1[0] ,
         dpath_mulcore_booth_b2_in1[2] , dpath_mulcore_booth_b2_in1[1] ,
         dpath_mulcore_booth_b2_in1[0] , dpath_mulcore_booth_b1_in1[2] ,
         dpath_mulcore_booth_b1_in1[1] , dpath_mulcore_booth_b1_in1[0] ,
         dpath_mulcore_booth_b0_in1[2] , dpath_mulcore_booth_b0_in1[1] ,
         dpath_mulcore_booth_b0_in1[0] , dpath_mulcore_booth_b[31] ,
         dpath_mulcore_booth_b[32] , dpath_mulcore_booth_b[34] ,
         dpath_mulcore_booth_b[36] , dpath_mulcore_booth_b[38] ,
         dpath_mulcore_booth_b[40] , dpath_mulcore_booth_b[42] ,
         dpath_mulcore_booth_b[44] , dpath_mulcore_booth_b[46] ,
         dpath_mulcore_booth_b[48] , dpath_mulcore_booth_b[50] ,
         dpath_mulcore_booth_b[52] , dpath_mulcore_booth_b[54] ,
         dpath_mulcore_booth_b[56] , dpath_mulcore_booth_b[58] ,
         dpath_mulcore_booth_b[60] , dpath_mulcore_booth_b[62] ,
         dpath_mulcore_booth_clk_enb1 , dpath_mulcore_booth_b15_in0[2] ,
         dpath_mulcore_booth_b15_in0[1] , dpath_mulcore_booth_b15_in0[0] ,
         dpath_mulcore_booth_b14_in0[2] , dpath_mulcore_booth_b14_in0[1] ,
         dpath_mulcore_booth_b14_in0[0] , dpath_mulcore_booth_b13_in0[2] ,
         dpath_mulcore_booth_b13_in0[1] , dpath_mulcore_booth_b13_in0[0] ,
         dpath_mulcore_booth_b12_in0[2] , dpath_mulcore_booth_b12_in0[1] ,
         dpath_mulcore_booth_b12_in0[0] , dpath_mulcore_booth_b11_in0[2] ,
         dpath_mulcore_booth_b11_in0[1] , dpath_mulcore_booth_b11_in0[0] ,
         dpath_mulcore_booth_b10_in0[2] , dpath_mulcore_booth_b10_in0[1] ,
         dpath_mulcore_booth_b10_in0[0] , dpath_mulcore_booth_b9_in0[2] ,
         dpath_mulcore_booth_b9_in0[1] , dpath_mulcore_booth_b9_in0[0] ,
         dpath_mulcore_booth_b8_in0[2] , dpath_mulcore_booth_b8_in0[1] ,
         dpath_mulcore_booth_b8_in0[0] , dpath_mulcore_booth_b7_in0[2] ,
         dpath_mulcore_booth_b7_in0[1] , dpath_mulcore_booth_b7_in0[0] ,
         dpath_mulcore_booth_b6_in0[2] , dpath_mulcore_booth_b6_in0[1] ,
         dpath_mulcore_booth_b6_in0[0] , dpath_mulcore_booth_b5_in0[2] ,
         dpath_mulcore_booth_b5_in0[1] , dpath_mulcore_booth_b5_in0[0] ,
         dpath_mulcore_booth_b4_in0[2] , dpath_mulcore_booth_b4_in0[1] ,
         dpath_mulcore_booth_b4_in0[0] , dpath_mulcore_booth_b3_in0[2] ,
         dpath_mulcore_booth_b3_in0[1] , dpath_mulcore_booth_b3_in0[0] ,
         dpath_mulcore_booth_b2_in0[2] , dpath_mulcore_booth_b2_in0[1] ,
         dpath_mulcore_booth_b2_in0[0] , dpath_mulcore_booth_b1_in0[2] ,
         dpath_mulcore_booth_b1_in0[1] , dpath_mulcore_booth_b1_in0[0] ,
         dpath_mulcore_booth_b0_in0[2] , dpath_mulcore_booth_b0_in0[1] ,
         dpath_mulcore_ary1_a0_s0[67] , dpath_mulcore_ary1_a0_s0[66] ,
         dpath_mulcore_ary1_a0_s0[65] , dpath_mulcore_ary1_a0_s0[64] ,
         dpath_mulcore_ary1_a0_s0[63] , dpath_mulcore_ary1_a0_s0[62] ,
         dpath_mulcore_ary1_a0_s0[61] , dpath_mulcore_ary1_a0_s0[60] ,
         dpath_mulcore_ary1_a0_s0[59] , dpath_mulcore_ary1_a0_s0[58] ,
         dpath_mulcore_ary1_a0_s0[57] , dpath_mulcore_ary1_a0_s0[56] ,
         dpath_mulcore_ary1_a0_s0[55] , dpath_mulcore_ary1_a0_s0[54] ,
         dpath_mulcore_ary1_a0_s0[53] , dpath_mulcore_ary1_a0_s0[52] ,
         dpath_mulcore_ary1_a0_s0[51] , dpath_mulcore_ary1_a0_s0[50] ,
         dpath_mulcore_ary1_a0_s0[49] , dpath_mulcore_ary1_a0_s0[48] ,
         dpath_mulcore_ary1_a0_s0[47] , dpath_mulcore_ary1_a0_s0[46] ,
         dpath_mulcore_ary1_a0_s0[45] , dpath_mulcore_ary1_a0_s0[44] ,
         dpath_mulcore_ary1_a0_s0[43] , dpath_mulcore_ary1_a0_s0[42] ,
         dpath_mulcore_ary1_a0_s0[41] , dpath_mulcore_ary1_a0_s0[40] ,
         dpath_mulcore_ary1_a0_s0[39] , dpath_mulcore_ary1_a0_s0[38] ,
         dpath_mulcore_ary1_a0_s0[37] , dpath_mulcore_ary1_a0_s0[36] ,
         dpath_mulcore_ary1_a0_s0[35] , dpath_mulcore_ary1_a0_s0[34] ,
         dpath_mulcore_ary1_a0_s0[33] , dpath_mulcore_ary1_a0_s0[32] ,
         dpath_mulcore_ary1_a0_s0[31] , dpath_mulcore_ary1_a0_s0[30] ,
         dpath_mulcore_ary1_a0_s0[29] , dpath_mulcore_ary1_a0_s0[28] ,
         dpath_mulcore_ary1_a0_s0[27] , dpath_mulcore_ary1_a0_s0[26] ,
         dpath_mulcore_ary1_a0_s0[25] , dpath_mulcore_ary1_a0_s0[24] ,
         dpath_mulcore_ary1_a0_s0[23] , dpath_mulcore_ary1_a0_s0[22] ,
         dpath_mulcore_ary1_a0_s0[21] , dpath_mulcore_ary1_a0_s0[20] ,
         dpath_mulcore_ary1_a0_s0[19] , dpath_mulcore_ary1_a0_s0[18] ,
         dpath_mulcore_ary1_a0_s0[17] , dpath_mulcore_ary1_a0_s0[16] ,
         dpath_mulcore_ary1_a0_s0[15] , dpath_mulcore_ary1_a0_s0[14] ,
         dpath_mulcore_ary1_a0_s0[13] , dpath_mulcore_ary1_a0_s0[12] ,
         dpath_mulcore_ary1_a0_s0[11] , dpath_mulcore_ary1_a0_s0[10] ,
         dpath_mulcore_ary1_a0_s0[9] , dpath_mulcore_ary1_a0_s0[8] ,
         dpath_mulcore_ary1_a0_s0[7] , dpath_mulcore_ary1_a0_s0[6] ,
         dpath_mulcore_ary1_a0_s0[5] , dpath_mulcore_ary1_a0_s0[4] ,
         dpath_mulcore_ary1_a0_s0[3] , dpath_mulcore_ary1_a0_s0[2] ,
         dpath_mulcore_ary1_a0_c0[67] , dpath_mulcore_ary1_a0_c0[66] ,
         dpath_mulcore_ary1_a0_c0[65] , dpath_mulcore_ary1_a0_c0[64] ,
         dpath_mulcore_ary1_a0_c0[63] , dpath_mulcore_ary1_a0_c0[62] ,
         dpath_mulcore_ary1_a0_c0[61] , dpath_mulcore_ary1_a0_c0[60] ,
         dpath_mulcore_ary1_a0_c0[59] , dpath_mulcore_ary1_a0_c0[58] ,
         dpath_mulcore_ary1_a0_c0[57] , dpath_mulcore_ary1_a0_c0[56] ,
         dpath_mulcore_ary1_a0_c0[55] , dpath_mulcore_ary1_a0_c0[54] ,
         dpath_mulcore_ary1_a0_c0[53] , dpath_mulcore_ary1_a0_c0[52] ,
         dpath_mulcore_ary1_a0_c0[51] , dpath_mulcore_ary1_a0_c0[50] ,
         dpath_mulcore_ary1_a0_c0[49] , dpath_mulcore_ary1_a0_c0[48] ,
         dpath_mulcore_ary1_a0_c0[47] , dpath_mulcore_ary1_a0_c0[46] ,
         dpath_mulcore_ary1_a0_c0[45] , dpath_mulcore_ary1_a0_c0[44] ,
         dpath_mulcore_ary1_a0_c0[43] , dpath_mulcore_ary1_a0_c0[42] ,
         dpath_mulcore_ary1_a0_c0[41] , dpath_mulcore_ary1_a0_c0[40] ,
         dpath_mulcore_ary1_a0_c0[39] , dpath_mulcore_ary1_a0_c0[38] ,
         dpath_mulcore_ary1_a0_c0[37] , dpath_mulcore_ary1_a0_c0[36] ,
         dpath_mulcore_ary1_a0_c0[35] , dpath_mulcore_ary1_a0_c0[34] ,
         dpath_mulcore_ary1_a0_c0[33] , dpath_mulcore_ary1_a0_c0[32] ,
         dpath_mulcore_ary1_a0_c0[31] , dpath_mulcore_ary1_a0_c0[30] ,
         dpath_mulcore_ary1_a0_c0[29] , dpath_mulcore_ary1_a0_c0[28] ,
         dpath_mulcore_ary1_a0_c0[27] , dpath_mulcore_ary1_a0_c0[26] ,
         dpath_mulcore_ary1_a0_c0[25] , dpath_mulcore_ary1_a0_c0[24] ,
         dpath_mulcore_ary1_a0_c0[23] , dpath_mulcore_ary1_a0_c0[22] ,
         dpath_mulcore_ary1_a0_c0[21] , dpath_mulcore_ary1_a0_c0[20] ,
         dpath_mulcore_ary1_a0_c0[19] , dpath_mulcore_ary1_a0_c0[18] ,
         dpath_mulcore_ary1_a0_c0[17] , dpath_mulcore_ary1_a0_c0[16] ,
         dpath_mulcore_ary1_a0_c0[15] , dpath_mulcore_ary1_a0_c0[14] ,
         dpath_mulcore_ary1_a0_c0[13] , dpath_mulcore_ary1_a0_c0[12] ,
         dpath_mulcore_ary1_a0_c0[11] , dpath_mulcore_ary1_a0_c0[10] ,
         dpath_mulcore_ary1_a0_c0[9] , dpath_mulcore_ary1_a0_c0[8] ,
         dpath_mulcore_ary1_a0_c0[7] , dpath_mulcore_ary1_a0_c0[6] ,
         dpath_mulcore_ary1_a0_c0[5] , dpath_mulcore_ary1_a0_c0[4] ,
         dpath_mulcore_ary1_a0_c0[3] , dpath_mulcore_ary1_a0_c0[2] ,
         dpath_mulcore_ary1_a0_c0[1] , dpath_mulcore_ary1_a0_s2[3] ,
         dpath_mulcore_ary1_a0_s2[2] , dpath_mulcore_ary1_a0_s2[1] ,
         dpath_mulcore_ary1_a0_s2[0] , dpath_mulcore_ary1_a0_c2[3] ,
         dpath_mulcore_ary1_a0_c2[2] , dpath_mulcore_ary1_a0_c2[1] ,
         dpath_mulcore_ary1_a0_c1[66] , dpath_mulcore_ary1_a0_c1[65] ,
         dpath_mulcore_ary1_a0_c1[64] , dpath_mulcore_ary1_a0_c1[63] ,
         dpath_mulcore_ary1_a0_c1[62] , dpath_mulcore_ary1_a0_c1[61] ,
         dpath_mulcore_ary1_a0_c1[60] , dpath_mulcore_ary1_a0_c1[59] ,
         dpath_mulcore_ary1_a0_c1[58] , dpath_mulcore_ary1_a0_c1[57] ,
         dpath_mulcore_ary1_a0_c1[56] , dpath_mulcore_ary1_a0_c1[55] ,
         dpath_mulcore_ary1_a0_c1[54] , dpath_mulcore_ary1_a0_c1[53] ,
         dpath_mulcore_ary1_a0_c1[52] , dpath_mulcore_ary1_a0_c1[51] ,
         dpath_mulcore_ary1_a0_c1[50] , dpath_mulcore_ary1_a0_c1[49] ,
         dpath_mulcore_ary1_a0_c1[48] , dpath_mulcore_ary1_a0_c1[47] ,
         dpath_mulcore_ary1_a0_c1[46] , dpath_mulcore_ary1_a0_c1[45] ,
         dpath_mulcore_ary1_a0_c1[44] , dpath_mulcore_ary1_a0_c1[43] ,
         dpath_mulcore_ary1_a0_c1[42] , dpath_mulcore_ary1_a0_c1[41] ,
         dpath_mulcore_ary1_a0_c1[40] , dpath_mulcore_ary1_a0_c1[39] ,
         dpath_mulcore_ary1_a0_c1[38] , dpath_mulcore_ary1_a0_c1[37] ,
         dpath_mulcore_ary1_a0_c1[36] , dpath_mulcore_ary1_a0_c1[35] ,
         dpath_mulcore_ary1_a0_c1[34] , dpath_mulcore_ary1_a0_c1[33] ,
         dpath_mulcore_ary1_a0_c1[32] , dpath_mulcore_ary1_a0_c1[31] ,
         dpath_mulcore_ary1_a0_c1[30] , dpath_mulcore_ary1_a0_c1[29] ,
         dpath_mulcore_ary1_a0_c1[28] , dpath_mulcore_ary1_a0_c1[27] ,
         dpath_mulcore_ary1_a0_c1[26] , dpath_mulcore_ary1_a0_c1[25] ,
         dpath_mulcore_ary1_a0_c1[24] , dpath_mulcore_ary1_a0_c1[23] ,
         dpath_mulcore_ary1_a0_c1[22] , dpath_mulcore_ary1_a0_c1[21] ,
         dpath_mulcore_ary1_a0_c1[20] , dpath_mulcore_ary1_a0_c1[19] ,
         dpath_mulcore_ary1_a0_c1[18] , dpath_mulcore_ary1_a0_c1[17] ,
         dpath_mulcore_ary1_a0_c1[16] , dpath_mulcore_ary1_a0_c1[15] ,
         dpath_mulcore_ary1_a0_c1[14] , dpath_mulcore_ary1_a0_c1[13] ,
         dpath_mulcore_ary1_a0_c1[12] , dpath_mulcore_ary1_a0_c1[11] ,
         dpath_mulcore_ary1_a0_c1[10] , dpath_mulcore_ary1_a0_c1[9] ,
         dpath_mulcore_ary1_a0_c1[8] , dpath_mulcore_ary1_a0_c1[7] ,
         dpath_mulcore_ary1_a0_c1[6] , dpath_mulcore_ary1_a0_c1[5] ,
         dpath_mulcore_ary1_a0_c1[4] , dpath_mulcore_ary1_a0_c1[3] ,
         dpath_mulcore_ary1_a0_c1[2] , dpath_mulcore_ary1_a0_c1[1] ,
         dpath_mulcore_ary1_a0_s_1[69] , dpath_mulcore_ary1_a0_s_1[68] ,
         dpath_mulcore_ary1_a0_s_1[67] , dpath_mulcore_ary1_a0_s_1[66] ,
         dpath_mulcore_ary1_a0_s_1[65] , dpath_mulcore_ary1_a0_s_1[64] ,
         dpath_mulcore_ary1_a0_s_1[63] , dpath_mulcore_ary1_a0_s_1[62] ,
         dpath_mulcore_ary1_a0_s_1[61] , dpath_mulcore_ary1_a0_s_1[60] ,
         dpath_mulcore_ary1_a0_s_1[59] , dpath_mulcore_ary1_a0_s_1[58] ,
         dpath_mulcore_ary1_a0_s_1[57] , dpath_mulcore_ary1_a0_s_1[56] ,
         dpath_mulcore_ary1_a0_s_1[55] , dpath_mulcore_ary1_a0_s_1[54] ,
         dpath_mulcore_ary1_a0_s_1[53] , dpath_mulcore_ary1_a0_s_1[52] ,
         dpath_mulcore_ary1_a0_s_1[51] , dpath_mulcore_ary1_a0_s_1[50] ,
         dpath_mulcore_ary1_a0_s_1[49] , dpath_mulcore_ary1_a0_s_1[48] ,
         dpath_mulcore_ary1_a0_s_1[47] , dpath_mulcore_ary1_a0_s_1[46] ,
         dpath_mulcore_ary1_a0_s_1[45] , dpath_mulcore_ary1_a0_s_1[44] ,
         dpath_mulcore_ary1_a0_s_1[43] , dpath_mulcore_ary1_a0_s_1[42] ,
         dpath_mulcore_ary1_a0_s_1[41] , dpath_mulcore_ary1_a0_s_1[40] ,
         dpath_mulcore_ary1_a0_s_1[39] , dpath_mulcore_ary1_a0_s_1[38] ,
         dpath_mulcore_ary1_a0_s_1[37] , dpath_mulcore_ary1_a0_s_1[36] ,
         dpath_mulcore_ary1_a0_s_1[35] , dpath_mulcore_ary1_a0_s_1[34] ,
         dpath_mulcore_ary1_a0_s_1[33] , dpath_mulcore_ary1_a0_s_1[32] ,
         dpath_mulcore_ary1_a0_s_1[31] , dpath_mulcore_ary1_a0_s_1[30] ,
         dpath_mulcore_ary1_a0_s_1[29] , dpath_mulcore_ary1_a0_s_1[28] ,
         dpath_mulcore_ary1_a0_s_1[27] , dpath_mulcore_ary1_a0_s_1[26] ,
         dpath_mulcore_ary1_a0_s_1[25] , dpath_mulcore_ary1_a0_s_1[24] ,
         dpath_mulcore_ary1_a0_s_1[23] , dpath_mulcore_ary1_a0_s_1[22] ,
         dpath_mulcore_ary1_a0_s_1[21] , dpath_mulcore_ary1_a0_s_1[20] ,
         dpath_mulcore_ary1_a0_s_1[19] , dpath_mulcore_ary1_a0_s_1[18] ,
         dpath_mulcore_ary1_a0_s_1[17] , dpath_mulcore_ary1_a0_s_1[16] ,
         dpath_mulcore_ary1_a0_s_1[15] , dpath_mulcore_ary1_a0_s_1[14] ,
         dpath_mulcore_ary1_a0_s_1[13] , dpath_mulcore_ary1_a0_s_1[12] ,
         dpath_mulcore_ary1_a0_s_1[11] , dpath_mulcore_ary1_a0_s_1[10] ,
         dpath_mulcore_ary1_a0_s_1[9] , dpath_mulcore_ary1_a0_s_1[8] ,
         dpath_mulcore_ary1_a0_s_1[7] , dpath_mulcore_ary1_a0_s_1[6] ,
         dpath_mulcore_ary1_a0_s_1[5] , dpath_mulcore_ary1_a0_s_1[4] ,
         dpath_mulcore_ary1_a0_s1[67] , dpath_mulcore_ary1_a0_s1[66] ,
         dpath_mulcore_ary1_a0_s1[65] , dpath_mulcore_ary1_a0_s1[64] ,
         dpath_mulcore_ary1_a0_s1[63] , dpath_mulcore_ary1_a0_s1[62] ,
         dpath_mulcore_ary1_a0_s1[61] , dpath_mulcore_ary1_a0_s1[60] ,
         dpath_mulcore_ary1_a0_s1[59] , dpath_mulcore_ary1_a0_s1[58] ,
         dpath_mulcore_ary1_a0_s1[57] , dpath_mulcore_ary1_a0_s1[56] ,
         dpath_mulcore_ary1_a0_s1[55] , dpath_mulcore_ary1_a0_s1[54] ,
         dpath_mulcore_ary1_a0_s1[53] , dpath_mulcore_ary1_a0_s1[52] ,
         dpath_mulcore_ary1_a0_s1[51] , dpath_mulcore_ary1_a0_s1[50] ,
         dpath_mulcore_ary1_a0_s1[49] , dpath_mulcore_ary1_a0_s1[48] ,
         dpath_mulcore_ary1_a0_s1[47] , dpath_mulcore_ary1_a0_s1[46] ,
         dpath_mulcore_ary1_a0_s1[45] , dpath_mulcore_ary1_a0_s1[44] ,
         dpath_mulcore_ary1_a0_s1[43] , dpath_mulcore_ary1_a0_s1[42] ,
         dpath_mulcore_ary1_a0_s1[41] , dpath_mulcore_ary1_a0_s1[40] ,
         dpath_mulcore_ary1_a0_s1[39] , dpath_mulcore_ary1_a0_s1[38] ,
         dpath_mulcore_ary1_a0_s1[37] , dpath_mulcore_ary1_a0_s1[36] ,
         dpath_mulcore_ary1_a0_s1[35] , dpath_mulcore_ary1_a0_s1[34] ,
         dpath_mulcore_ary1_a0_s1[33] , dpath_mulcore_ary1_a0_s1[32] ,
         dpath_mulcore_ary1_a0_s1[31] , dpath_mulcore_ary1_a0_s1[30] ,
         dpath_mulcore_ary1_a0_s1[29] , dpath_mulcore_ary1_a0_s1[28] ,
         dpath_mulcore_ary1_a0_s1[27] , dpath_mulcore_ary1_a0_s1[26] ,
         dpath_mulcore_ary1_a0_s1[25] , dpath_mulcore_ary1_a0_s1[24] ,
         dpath_mulcore_ary1_a0_s1[23] , dpath_mulcore_ary1_a0_s1[22] ,
         dpath_mulcore_ary1_a0_s1[21] , dpath_mulcore_ary1_a0_s1[20] ,
         dpath_mulcore_ary1_a0_s1[19] , dpath_mulcore_ary1_a0_s1[18] ,
         dpath_mulcore_ary1_a0_s1[17] , dpath_mulcore_ary1_a0_s1[16] ,
         dpath_mulcore_ary1_a0_s1[15] , dpath_mulcore_ary1_a0_s1[14] ,
         dpath_mulcore_ary1_a0_s1[13] , dpath_mulcore_ary1_a0_s1[12] ,
         dpath_mulcore_ary1_a0_s1[11] , dpath_mulcore_ary1_a0_s1[10] ,
         dpath_mulcore_ary1_a0_s1[9] , dpath_mulcore_ary1_a0_s1[8] ,
         dpath_mulcore_ary1_a0_s1[7] , dpath_mulcore_ary1_a0_s1[6] ,
         dpath_mulcore_ary1_a0_s1[5] , dpath_mulcore_ary1_a0_s1[4] ,
         dpath_mulcore_ary1_a0_s1[3] , dpath_mulcore_ary1_a0_s1[2] ,
         dpath_mulcore_ary1_a0_s1[1] , dpath_mulcore_ary1_a0_s1[0] ,
         dpath_mulcore_ary1_a0_c_2[76] , dpath_mulcore_ary1_a0_c_2[75] ,
         dpath_mulcore_ary1_a0_c_2[74] , dpath_mulcore_ary1_a0_c_2[73] ,
         dpath_mulcore_ary1_a0_c_2[72] , dpath_mulcore_ary1_a0_c_2[71] ,
         dpath_mulcore_ary1_a0_c_2[70] , dpath_mulcore_ary1_a0_c_2[69] ,
         dpath_mulcore_ary1_a0_c_2[68] , dpath_mulcore_ary1_a0_c_2[67] ,
         dpath_mulcore_ary1_a0_c_2[66] , dpath_mulcore_ary1_a0_c_2[65] ,
         dpath_mulcore_ary1_a0_c_2[64] , dpath_mulcore_ary1_a0_c_2[63] ,
         dpath_mulcore_ary1_a0_c_2[62] , dpath_mulcore_ary1_a0_c_2[61] ,
         dpath_mulcore_ary1_a0_c_2[60] , dpath_mulcore_ary1_a0_c_2[59] ,
         dpath_mulcore_ary1_a0_c_2[58] , dpath_mulcore_ary1_a0_c_2[57] ,
         dpath_mulcore_ary1_a0_c_2[56] , dpath_mulcore_ary1_a0_c_2[55] ,
         dpath_mulcore_ary1_a0_c_2[54] , dpath_mulcore_ary1_a0_c_2[53] ,
         dpath_mulcore_ary1_a0_c_2[52] , dpath_mulcore_ary1_a0_c_2[51] ,
         dpath_mulcore_ary1_a0_c_2[50] , dpath_mulcore_ary1_a0_c_2[49] ,
         dpath_mulcore_ary1_a0_c_2[48] , dpath_mulcore_ary1_a0_c_2[47] ,
         dpath_mulcore_ary1_a0_c_2[46] , dpath_mulcore_ary1_a0_c_2[45] ,
         dpath_mulcore_ary1_a0_c_2[44] , dpath_mulcore_ary1_a0_c_2[43] ,
         dpath_mulcore_ary1_a0_c_2[42] , dpath_mulcore_ary1_a0_c_2[41] ,
         dpath_mulcore_ary1_a0_c_2[40] , dpath_mulcore_ary1_a0_c_2[39] ,
         dpath_mulcore_ary1_a0_c_2[38] , dpath_mulcore_ary1_a0_c_2[37] ,
         dpath_mulcore_ary1_a0_c_2[36] , dpath_mulcore_ary1_a0_c_2[35] ,
         dpath_mulcore_ary1_a0_c_2[34] , dpath_mulcore_ary1_a0_c_2[33] ,
         dpath_mulcore_ary1_a0_c_2[32] , dpath_mulcore_ary1_a0_c_2[31] ,
         dpath_mulcore_ary1_a0_c_2[30] , dpath_mulcore_ary1_a0_c_2[29] ,
         dpath_mulcore_ary1_a0_c_2[28] , dpath_mulcore_ary1_a0_c_2[27] ,
         dpath_mulcore_ary1_a0_c_2[26] , dpath_mulcore_ary1_a0_c_2[25] ,
         dpath_mulcore_ary1_a0_c_2[24] , dpath_mulcore_ary1_a0_c_2[23] ,
         dpath_mulcore_ary1_a0_c_2[22] , dpath_mulcore_ary1_a0_c_2[21] ,
         dpath_mulcore_ary1_a0_c_2[20] , dpath_mulcore_ary1_a0_c_2[19] ,
         dpath_mulcore_ary1_a0_c_2[18] , dpath_mulcore_ary1_a0_c_2[17] ,
         dpath_mulcore_ary1_a0_c_2[16] , dpath_mulcore_ary1_a0_c_2[15] ,
         dpath_mulcore_ary1_a0_c_2[14] , dpath_mulcore_ary1_a0_c_2[13] ,
         dpath_mulcore_ary1_a0_c_2[12] , dpath_mulcore_ary1_a0_c_2[11] ,
         dpath_mulcore_ary1_a0_c_2[10] , dpath_mulcore_ary1_a0_c_1[69] ,
         dpath_mulcore_ary1_a0_c_1[68] , dpath_mulcore_ary1_a0_c_1[67] ,
         dpath_mulcore_ary1_a0_c_1[66] , dpath_mulcore_ary1_a0_c_1[65] ,
         dpath_mulcore_ary1_a0_c_1[64] , dpath_mulcore_ary1_a0_c_1[63] ,
         dpath_mulcore_ary1_a0_c_1[62] , dpath_mulcore_ary1_a0_c_1[61] ,
         dpath_mulcore_ary1_a0_c_1[60] , dpath_mulcore_ary1_a0_c_1[59] ,
         dpath_mulcore_ary1_a0_c_1[58] , dpath_mulcore_ary1_a0_c_1[57] ,
         dpath_mulcore_ary1_a0_c_1[56] , dpath_mulcore_ary1_a0_c_1[55] ,
         dpath_mulcore_ary1_a0_c_1[54] , dpath_mulcore_ary1_a0_c_1[53] ,
         dpath_mulcore_ary1_a0_c_1[52] , dpath_mulcore_ary1_a0_c_1[51] ,
         dpath_mulcore_ary1_a0_c_1[50] , dpath_mulcore_ary1_a0_c_1[49] ,
         dpath_mulcore_ary1_a0_c_1[48] , dpath_mulcore_ary1_a0_c_1[47] ,
         dpath_mulcore_ary1_a0_c_1[46] , dpath_mulcore_ary1_a0_c_1[45] ,
         dpath_mulcore_ary1_a0_c_1[44] , dpath_mulcore_ary1_a0_c_1[43] ,
         dpath_mulcore_ary1_a0_c_1[42] , dpath_mulcore_ary1_a0_c_1[41] ,
         dpath_mulcore_ary1_a0_c_1[40] , dpath_mulcore_ary1_a0_c_1[39] ,
         dpath_mulcore_ary1_a0_c_1[38] , dpath_mulcore_ary1_a0_c_1[37] ,
         dpath_mulcore_ary1_a0_c_1[36] , dpath_mulcore_ary1_a0_c_1[35] ,
         dpath_mulcore_ary1_a0_c_1[34] , dpath_mulcore_ary1_a0_c_1[33] ,
         dpath_mulcore_ary1_a0_c_1[32] , dpath_mulcore_ary1_a0_c_1[31] ,
         dpath_mulcore_ary1_a0_c_1[30] , dpath_mulcore_ary1_a0_c_1[29] ,
         dpath_mulcore_ary1_a0_c_1[28] , dpath_mulcore_ary1_a0_c_1[27] ,
         dpath_mulcore_ary1_a0_c_1[26] , dpath_mulcore_ary1_a0_c_1[25] ,
         dpath_mulcore_ary1_a0_c_1[24] , dpath_mulcore_ary1_a0_c_1[23] ,
         dpath_mulcore_ary1_a0_c_1[22] , dpath_mulcore_ary1_a0_c_1[21] ,
         dpath_mulcore_ary1_a0_c_1[20] , dpath_mulcore_ary1_a0_c_1[19] ,
         dpath_mulcore_ary1_a0_c_1[18] , dpath_mulcore_ary1_a0_c_1[17] ,
         dpath_mulcore_ary1_a0_c_1[16] , dpath_mulcore_ary1_a0_c_1[15] ,
         dpath_mulcore_ary1_a0_c_1[14] , dpath_mulcore_ary1_a0_c_1[13] ,
         dpath_mulcore_ary1_a0_c_1[12] , dpath_mulcore_ary1_a0_c_1[11] ,
         dpath_mulcore_ary1_a0_c_1[10] , dpath_mulcore_ary1_a0_c_1[9] ,
         dpath_mulcore_ary1_a0_c_1[8] , dpath_mulcore_ary1_a0_c_1[7] ,
         dpath_mulcore_ary1_a0_c_1[6] , dpath_mulcore_ary1_a0_c_1[5] ,
         dpath_mulcore_ary1_a0_c_1[4] , dpath_mulcore_ary1_a0_c_1[3] ,
         dpath_mulcore_ary1_a0_c_1[2] , dpath_mulcore_ary1_a0_co[71] ,
         dpath_mulcore_ary1_a0_co[70] , dpath_mulcore_ary1_a0_co[69] ,
         dpath_mulcore_ary1_a0_co[68] , dpath_mulcore_ary1_a0_co[67] ,
         dpath_mulcore_ary1_a0_co[66] , dpath_mulcore_ary1_a0_co[65] ,
         dpath_mulcore_ary1_a0_co[64] , dpath_mulcore_ary1_a0_co[63] ,
         dpath_mulcore_ary1_a0_co[62] , dpath_mulcore_ary1_a0_co[61] ,
         dpath_mulcore_ary1_a0_co[60] , dpath_mulcore_ary1_a0_co[59] ,
         dpath_mulcore_ary1_a0_co[58] , dpath_mulcore_ary1_a0_co[57] ,
         dpath_mulcore_ary1_a0_co[56] , dpath_mulcore_ary1_a0_co[55] ,
         dpath_mulcore_ary1_a0_co[54] , dpath_mulcore_ary1_a0_co[53] ,
         dpath_mulcore_ary1_a0_co[52] , dpath_mulcore_ary1_a0_co[51] ,
         dpath_mulcore_ary1_a0_co[50] , dpath_mulcore_ary1_a0_co[49] ,
         dpath_mulcore_ary1_a0_co[48] , dpath_mulcore_ary1_a0_co[47] ,
         dpath_mulcore_ary1_a0_co[46] , dpath_mulcore_ary1_a0_co[45] ,
         dpath_mulcore_ary1_a0_co[44] , dpath_mulcore_ary1_a0_co[43] ,
         dpath_mulcore_ary1_a0_co[42] , dpath_mulcore_ary1_a0_co[41] ,
         dpath_mulcore_ary1_a0_co[40] , dpath_mulcore_ary1_a0_co[39] ,
         dpath_mulcore_ary1_a0_co[38] , dpath_mulcore_ary1_a0_co[37] ,
         dpath_mulcore_ary1_a0_co[36] , dpath_mulcore_ary1_a0_co[35] ,
         dpath_mulcore_ary1_a0_co[34] , dpath_mulcore_ary1_a0_co[33] ,
         dpath_mulcore_ary1_a0_co[32] , dpath_mulcore_ary1_a0_co[31] ,
         dpath_mulcore_ary1_a0_co[30] , dpath_mulcore_ary1_a0_co[29] ,
         dpath_mulcore_ary1_a0_co[28] , dpath_mulcore_ary1_a0_co[27] ,
         dpath_mulcore_ary1_a0_co[26] , dpath_mulcore_ary1_a0_co[25] ,
         dpath_mulcore_ary1_a0_co[24] , dpath_mulcore_ary1_a0_co[23] ,
         dpath_mulcore_ary1_a0_co[22] , dpath_mulcore_ary1_a0_co[21] ,
         dpath_mulcore_ary1_a0_co[20] , dpath_mulcore_ary1_a0_co[19] ,
         dpath_mulcore_ary1_a0_co[18] , dpath_mulcore_ary1_a0_co[17] ,
         dpath_mulcore_ary1_a0_co[16] , dpath_mulcore_ary1_a0_co[15] ,
         dpath_mulcore_ary1_a0_co[14] , dpath_mulcore_ary1_a0_co[13] ,
         dpath_mulcore_ary1_a0_co[12] , dpath_mulcore_ary1_a0_co[11] ,
         dpath_mulcore_ary1_a0_s_2[75] , dpath_mulcore_ary1_a0_s_2[74] ,
         dpath_mulcore_ary1_a0_s_2[73] , dpath_mulcore_ary1_a0_s_2[72] ,
         dpath_mulcore_ary1_a0_s_2[71] , dpath_mulcore_ary1_a0_s_2[70] ,
         dpath_mulcore_ary1_a0_s_2[69] , dpath_mulcore_ary1_a0_s_2[68] ,
         dpath_mulcore_ary1_a0_s_2[67] , dpath_mulcore_ary1_a0_s_2[66] ,
         dpath_mulcore_ary1_a0_s_2[65] , dpath_mulcore_ary1_a0_s_2[64] ,
         dpath_mulcore_ary1_a0_s_2[63] , dpath_mulcore_ary1_a0_s_2[62] ,
         dpath_mulcore_ary1_a0_s_2[61] , dpath_mulcore_ary1_a0_s_2[60] ,
         dpath_mulcore_ary1_a0_s_2[59] , dpath_mulcore_ary1_a0_s_2[58] ,
         dpath_mulcore_ary1_a0_s_2[57] , dpath_mulcore_ary1_a0_s_2[56] ,
         dpath_mulcore_ary1_a0_s_2[55] , dpath_mulcore_ary1_a0_s_2[54] ,
         dpath_mulcore_ary1_a0_s_2[53] , dpath_mulcore_ary1_a0_s_2[52] ,
         dpath_mulcore_ary1_a0_s_2[51] , dpath_mulcore_ary1_a0_s_2[50] ,
         dpath_mulcore_ary1_a0_s_2[49] , dpath_mulcore_ary1_a0_s_2[48] ,
         dpath_mulcore_ary1_a0_s_2[47] , dpath_mulcore_ary1_a0_s_2[46] ,
         dpath_mulcore_ary1_a0_s_2[45] , dpath_mulcore_ary1_a0_s_2[44] ,
         dpath_mulcore_ary1_a0_s_2[43] , dpath_mulcore_ary1_a0_s_2[42] ,
         dpath_mulcore_ary1_a0_s_2[41] , dpath_mulcore_ary1_a0_s_2[40] ,
         dpath_mulcore_ary1_a0_s_2[39] , dpath_mulcore_ary1_a0_s_2[38] ,
         dpath_mulcore_ary1_a0_s_2[37] , dpath_mulcore_ary1_a0_s_2[36] ,
         dpath_mulcore_ary1_a0_s_2[35] , dpath_mulcore_ary1_a0_s_2[34] ,
         dpath_mulcore_ary1_a0_s_2[33] , dpath_mulcore_ary1_a0_s_2[32] ,
         dpath_mulcore_ary1_a0_s_2[31] , dpath_mulcore_ary1_a0_s_2[30] ,
         dpath_mulcore_ary1_a0_s_2[29] , dpath_mulcore_ary1_a0_s_2[28] ,
         dpath_mulcore_ary1_a0_s_2[27] , dpath_mulcore_ary1_a0_s_2[26] ,
         dpath_mulcore_ary1_a0_s_2[25] , dpath_mulcore_ary1_a0_s_2[24] ,
         dpath_mulcore_ary1_a0_s_2[23] , dpath_mulcore_ary1_a0_s_2[22] ,
         dpath_mulcore_ary1_a0_s_2[21] , dpath_mulcore_ary1_a0_s_2[20] ,
         dpath_mulcore_ary1_a0_s_2[19] , dpath_mulcore_ary1_a0_s_2[18] ,
         dpath_mulcore_ary1_a0_s_2[17] , dpath_mulcore_ary1_a0_s_2[16] ,
         dpath_mulcore_ary1_a0_s_2[15] , dpath_mulcore_ary1_a0_s_2[14] ,
         dpath_mulcore_ary1_a0_s_2[13] , dpath_mulcore_ary1_a0_s_2[12] ,
         dpath_mulcore_ary1_a0_s_2[11] , dpath_mulcore_ary1_a0_s_2[10] ,
         dpath_mulcore_ary1_a0_b2n[1] , dpath_mulcore_ary1_a0_b2n[0] ,
         dpath_mulcore_ary1_a0_b5n[1] , dpath_mulcore_ary1_a0_b5n[0] ,
         dpath_mulcore_a0cot_dff_n157 , dpath_mulcore_a0cot_dff_n155 ,
         dpath_mulcore_a0cot_dff_n153 , dpath_mulcore_a0cot_dff_n151 ,
         dpath_mulcore_a0cot_dff_n149 , dpath_mulcore_a0cot_dff_n147 ,
         dpath_mulcore_a0cot_dff_n145 , dpath_mulcore_a0cot_dff_n143 ,
         dpath_mulcore_a0cot_dff_n141 , dpath_mulcore_a0cot_dff_n139 ,
         dpath_mulcore_a0cot_dff_n137 , dpath_mulcore_a0cot_dff_n135 ,
         dpath_mulcore_a0cot_dff_n133 , dpath_mulcore_a0cot_dff_n131 ,
         dpath_mulcore_a0cot_dff_n129 , dpath_mulcore_a0cot_dff_n127 ,
         dpath_mulcore_a0cot_dff_n125 , dpath_mulcore_a0cot_dff_n123 ,
         dpath_mulcore_a0cot_dff_n121 , dpath_mulcore_a0cot_dff_n119 ,
         dpath_mulcore_a0cot_dff_n117 , dpath_mulcore_a0cot_dff_n115 ,
         dpath_mulcore_a0cot_dff_n113 , dpath_mulcore_a0cot_dff_n111 ,
         dpath_mulcore_a0cot_dff_n109 , dpath_mulcore_a0cot_dff_n107 ,
         dpath_mulcore_a0cot_dff_n105 , dpath_mulcore_a0cot_dff_n103 ,
         dpath_mulcore_a0cot_dff_n101 , dpath_mulcore_a0cot_dff_n99 ,
         dpath_mulcore_a0cot_dff_n97 , dpath_mulcore_a0cot_dff_n95 ,
         dpath_mulcore_a0cot_dff_n93 , dpath_mulcore_a0cot_dff_n91 ,
         dpath_mulcore_a0cot_dff_n89 , dpath_mulcore_a0cot_dff_n87 ,
         dpath_mulcore_a0cot_dff_n85 , dpath_mulcore_a0cot_dff_n83 ,
         dpath_mulcore_a0cot_dff_n81 , dpath_mulcore_a0cot_dff_n79 ,
         dpath_mulcore_a0cot_dff_n77 , dpath_mulcore_a0cot_dff_n75 ,
         dpath_mulcore_a0cot_dff_n73 , dpath_mulcore_a0cot_dff_n71 ,
         dpath_mulcore_a0cot_dff_n69 , dpath_mulcore_a0cot_dff_n67 ,
         dpath_mulcore_a0cot_dff_n65 , dpath_mulcore_a0cot_dff_n63 ,
         dpath_mulcore_a0cot_dff_n61 , dpath_mulcore_a0cot_dff_n59 ,
         dpath_mulcore_a0cot_dff_n57 , dpath_mulcore_a0cot_dff_n55 ,
         dpath_mulcore_a0cot_dff_n53 , dpath_mulcore_a0cot_dff_n51 ,
         dpath_mulcore_a0cot_dff_n49 , dpath_mulcore_a0cot_dff_n47 ,
         dpath_mulcore_a0cot_dff_n45 , dpath_mulcore_a0cot_dff_n43 ,
         dpath_mulcore_a0cot_dff_n41 , dpath_mulcore_a0cot_dff_n39 ,
         dpath_mulcore_a0cot_dff_n37 , dpath_mulcore_a0cot_dff_n35 ,
         dpath_mulcore_a0cot_dff_n33 , dpath_mulcore_a0cot_dff_n31 ,
         dpath_mulcore_a0cot_dff_n29 , dpath_mulcore_a0cot_dff_n27 ,
         dpath_mulcore_a0cot_dff_n25 , dpath_mulcore_a0cot_dff_n23 ,
         dpath_mulcore_a0cot_dff_n21 , dpath_mulcore_a0cot_dff_n19 ,
         dpath_mulcore_a0cot_dff_n17 , dpath_mulcore_a0cot_dff_n15 ,
         dpath_mulcore_a0cot_dff_n13 , dpath_mulcore_a0cot_dff_n11 ,
         dpath_mulcore_a0cot_dff_n7 , dpath_mulcore_a0cot_dff_n3 ,
         dpath_mulcore_a0sum_dff_n165 , dpath_mulcore_a0sum_dff_n163 ,
         dpath_mulcore_a0sum_dff_n161 , dpath_mulcore_a0sum_dff_n159 ,
         dpath_mulcore_a0sum_dff_n157 , dpath_mulcore_a0sum_dff_n155 ,
         dpath_mulcore_a0sum_dff_n153 , dpath_mulcore_a0sum_dff_n151 ,
         dpath_mulcore_a0sum_dff_n149 , dpath_mulcore_a0sum_dff_n147 ,
         dpath_mulcore_a0sum_dff_n145 , dpath_mulcore_a0sum_dff_n143 ,
         dpath_mulcore_a0sum_dff_n141 , dpath_mulcore_a0sum_dff_n139 ,
         dpath_mulcore_a0sum_dff_n137 , dpath_mulcore_a0sum_dff_n135 ,
         dpath_mulcore_a0sum_dff_n133 , dpath_mulcore_a0sum_dff_n131 ,
         dpath_mulcore_a0sum_dff_n129 , dpath_mulcore_a0sum_dff_n127 ,
         dpath_mulcore_a0sum_dff_n125 , dpath_mulcore_a0sum_dff_n123 ,
         dpath_mulcore_a0sum_dff_n121 , dpath_mulcore_a0sum_dff_n119 ,
         dpath_mulcore_a0sum_dff_n117 , dpath_mulcore_a0sum_dff_n115 ,
         dpath_mulcore_a0sum_dff_n113 , dpath_mulcore_a0sum_dff_n111 ,
         dpath_mulcore_a0sum_dff_n109 , dpath_mulcore_a0sum_dff_n107 ,
         dpath_mulcore_a0sum_dff_n105 , dpath_mulcore_a0sum_dff_n103 ,
         dpath_mulcore_a0sum_dff_n101 , dpath_mulcore_a0sum_dff_n99 ,
         dpath_mulcore_a0sum_dff_n97 , dpath_mulcore_a0sum_dff_n95 ,
         dpath_mulcore_a0sum_dff_n93 , dpath_mulcore_a0sum_dff_n91 ,
         dpath_mulcore_a0sum_dff_n89 , dpath_mulcore_a0sum_dff_n87 ,
         dpath_mulcore_a0sum_dff_n85 , dpath_mulcore_a0sum_dff_n83 ,
         dpath_mulcore_a0sum_dff_n81 , dpath_mulcore_a0sum_dff_n79 ,
         dpath_mulcore_a0sum_dff_n77 , dpath_mulcore_a0sum_dff_n75 ,
         dpath_mulcore_a0sum_dff_n73 , dpath_mulcore_a0sum_dff_n71 ,
         dpath_mulcore_a0sum_dff_n69 , dpath_mulcore_a0sum_dff_n67 ,
         dpath_mulcore_a0sum_dff_n65 , dpath_mulcore_a0sum_dff_n63 ,
         dpath_mulcore_a0sum_dff_n61 , dpath_mulcore_a0sum_dff_n59 ,
         dpath_mulcore_a0sum_dff_n57 , dpath_mulcore_a0sum_dff_n55 ,
         dpath_mulcore_a0sum_dff_n53 , dpath_mulcore_a0sum_dff_n51 ,
         dpath_mulcore_a0sum_dff_n49 , dpath_mulcore_a0sum_dff_n47 ,
         dpath_mulcore_a0sum_dff_n45 , dpath_mulcore_a0sum_dff_n43 ,
         dpath_mulcore_a0sum_dff_n41 , dpath_mulcore_a0sum_dff_n39 ,
         dpath_mulcore_a0sum_dff_n37 , dpath_mulcore_a0sum_dff_n35 ,
         dpath_mulcore_a0sum_dff_n33 , dpath_mulcore_a0sum_dff_n31 ,
         dpath_mulcore_a0sum_dff_n29 , dpath_mulcore_a0sum_dff_n27 ,
         dpath_mulcore_a0sum_dff_n25 , dpath_mulcore_a0sum_dff_n23 ,
         dpath_mulcore_a0sum_dff_n21 , dpath_mulcore_a0sum_dff_n19 ,
         dpath_mulcore_a0sum_dff_n17 , dpath_mulcore_a0sum_dff_n15 ,
         dpath_mulcore_a0sum_dff_n13 , dpath_mulcore_a0sum_dff_n11 ,
         dpath_mulcore_a0sum_dff_n9 , dpath_mulcore_a0sum_dff_n3 ,
         dpath_mulcore_ary1_a1_s0[67] , dpath_mulcore_ary1_a1_s0[66] ,
         dpath_mulcore_ary1_a1_s0[65] , dpath_mulcore_ary1_a1_s0[64] ,
         dpath_mulcore_ary1_a1_s0[63] , dpath_mulcore_ary1_a1_s0[62] ,
         dpath_mulcore_ary1_a1_s0[61] , dpath_mulcore_ary1_a1_s0[60] ,
         dpath_mulcore_ary1_a1_s0[59] , dpath_mulcore_ary1_a1_s0[58] ,
         dpath_mulcore_ary1_a1_s0[57] , dpath_mulcore_ary1_a1_s0[56] ,
         dpath_mulcore_ary1_a1_s0[55] , dpath_mulcore_ary1_a1_s0[54] ,
         dpath_mulcore_ary1_a1_s0[53] , dpath_mulcore_ary1_a1_s0[52] ,
         dpath_mulcore_ary1_a1_s0[51] , dpath_mulcore_ary1_a1_s0[50] ,
         dpath_mulcore_ary1_a1_s0[49] , dpath_mulcore_ary1_a1_s0[48] ,
         dpath_mulcore_ary1_a1_s0[47] , dpath_mulcore_ary1_a1_s0[46] ,
         dpath_mulcore_ary1_a1_s0[45] , dpath_mulcore_ary1_a1_s0[44] ,
         dpath_mulcore_ary1_a1_s0[43] , dpath_mulcore_ary1_a1_s0[42] ,
         dpath_mulcore_ary1_a1_s0[41] , dpath_mulcore_ary1_a1_s0[40] ,
         dpath_mulcore_ary1_a1_s0[39] , dpath_mulcore_ary1_a1_s0[38] ,
         dpath_mulcore_ary1_a1_s0[37] , dpath_mulcore_ary1_a1_s0[36] ,
         dpath_mulcore_ary1_a1_s0[35] , dpath_mulcore_ary1_a1_s0[34] ,
         dpath_mulcore_ary1_a1_s0[33] , dpath_mulcore_ary1_a1_s0[32] ,
         dpath_mulcore_ary1_a1_s0[31] , dpath_mulcore_ary1_a1_s0[30] ,
         dpath_mulcore_ary1_a1_s0[29] , dpath_mulcore_ary1_a1_s0[28] ,
         dpath_mulcore_ary1_a1_s0[27] , dpath_mulcore_ary1_a1_s0[26] ,
         dpath_mulcore_ary1_a1_s0[25] , dpath_mulcore_ary1_a1_s0[24] ,
         dpath_mulcore_ary1_a1_s0[23] , dpath_mulcore_ary1_a1_s0[22] ,
         dpath_mulcore_ary1_a1_s0[21] , dpath_mulcore_ary1_a1_s0[20] ,
         dpath_mulcore_ary1_a1_s0[19] , dpath_mulcore_ary1_a1_s0[18] ,
         dpath_mulcore_ary1_a1_s0[17] , dpath_mulcore_ary1_a1_s0[16] ,
         dpath_mulcore_ary1_a1_s0[15] , dpath_mulcore_ary1_a1_s0[14] ,
         dpath_mulcore_ary1_a1_s0[13] , dpath_mulcore_ary1_a1_s0[12] ,
         dpath_mulcore_ary1_a1_s0[11] , dpath_mulcore_ary1_a1_s0[10] ,
         dpath_mulcore_ary1_a1_s0[9] , dpath_mulcore_ary1_a1_s0[8] ,
         dpath_mulcore_ary1_a1_s0[7] , dpath_mulcore_ary1_a1_s0[6] ,
         dpath_mulcore_ary1_a1_s0[5] , dpath_mulcore_ary1_a1_s0[4] ,
         dpath_mulcore_ary1_a1_s0[3] , dpath_mulcore_ary1_a1_s0[2] ,
         dpath_mulcore_ary1_a1_c0[66] , dpath_mulcore_ary1_a1_c0[65] ,
         dpath_mulcore_ary1_a1_c0[64] , dpath_mulcore_ary1_a1_c0[63] ,
         dpath_mulcore_ary1_a1_c0[62] , dpath_mulcore_ary1_a1_c0[61] ,
         dpath_mulcore_ary1_a1_c0[60] , dpath_mulcore_ary1_a1_c0[59] ,
         dpath_mulcore_ary1_a1_c0[58] , dpath_mulcore_ary1_a1_c0[57] ,
         dpath_mulcore_ary1_a1_c0[56] , dpath_mulcore_ary1_a1_c0[55] ,
         dpath_mulcore_ary1_a1_c0[54] , dpath_mulcore_ary1_a1_c0[53] ,
         dpath_mulcore_ary1_a1_c0[52] , dpath_mulcore_ary1_a1_c0[51] ,
         dpath_mulcore_ary1_a1_c0[50] , dpath_mulcore_ary1_a1_c0[49] ,
         dpath_mulcore_ary1_a1_c0[48] , dpath_mulcore_ary1_a1_c0[47] ,
         dpath_mulcore_ary1_a1_c0[46] , dpath_mulcore_ary1_a1_c0[45] ,
         dpath_mulcore_ary1_a1_c0[44] , dpath_mulcore_ary1_a1_c0[43] ,
         dpath_mulcore_ary1_a1_c0[42] , dpath_mulcore_ary1_a1_c0[41] ,
         dpath_mulcore_ary1_a1_c0[40] , dpath_mulcore_ary1_a1_c0[39] ,
         dpath_mulcore_ary1_a1_c0[38] , dpath_mulcore_ary1_a1_c0[37] ,
         dpath_mulcore_ary1_a1_c0[36] , dpath_mulcore_ary1_a1_c0[35] ,
         dpath_mulcore_ary1_a1_c0[34] , dpath_mulcore_ary1_a1_c0[33] ,
         dpath_mulcore_ary1_a1_c0[32] , dpath_mulcore_ary1_a1_c0[31] ,
         dpath_mulcore_ary1_a1_c0[30] , dpath_mulcore_ary1_a1_c0[29] ,
         dpath_mulcore_ary1_a1_c0[28] , dpath_mulcore_ary1_a1_c0[27] ,
         dpath_mulcore_ary1_a1_c0[26] , dpath_mulcore_ary1_a1_c0[25] ,
         dpath_mulcore_ary1_a1_c0[24] , dpath_mulcore_ary1_a1_c0[23] ,
         dpath_mulcore_ary1_a1_c0[22] , dpath_mulcore_ary1_a1_c0[21] ,
         dpath_mulcore_ary1_a1_c0[20] , dpath_mulcore_ary1_a1_c0[19] ,
         dpath_mulcore_ary1_a1_c0[18] , dpath_mulcore_ary1_a1_c0[17] ,
         dpath_mulcore_ary1_a1_c0[16] , dpath_mulcore_ary1_a1_c0[15] ,
         dpath_mulcore_ary1_a1_c0[14] , dpath_mulcore_ary1_a1_c0[13] ,
         dpath_mulcore_ary1_a1_c0[12] , dpath_mulcore_ary1_a1_c0[11] ,
         dpath_mulcore_ary1_a1_c0[10] , dpath_mulcore_ary1_a1_c0[9] ,
         dpath_mulcore_ary1_a1_c0[8] , dpath_mulcore_ary1_a1_c0[7] ,
         dpath_mulcore_ary1_a1_c0[6] , dpath_mulcore_ary1_a1_c0[5] ,
         dpath_mulcore_ary1_a1_c0[4] , dpath_mulcore_ary1_a1_c0[3] ,
         dpath_mulcore_ary1_a1_c0[2] , dpath_mulcore_ary1_a1_c0[1] ,
         dpath_mulcore_ary1_a1_s2[67] , dpath_mulcore_ary1_a1_s2[66] ,
         dpath_mulcore_ary1_a1_s2[65] , dpath_mulcore_ary1_a1_s2[64] ,
         dpath_mulcore_ary1_a1_s2[63] , dpath_mulcore_ary1_a1_s2[62] ,
         dpath_mulcore_ary1_a1_s2[61] , dpath_mulcore_ary1_a1_s2[60] ,
         dpath_mulcore_ary1_a1_s2[59] , dpath_mulcore_ary1_a1_s2[58] ,
         dpath_mulcore_ary1_a1_s2[57] , dpath_mulcore_ary1_a1_s2[56] ,
         dpath_mulcore_ary1_a1_s2[55] , dpath_mulcore_ary1_a1_s2[54] ,
         dpath_mulcore_ary1_a1_s2[53] , dpath_mulcore_ary1_a1_s2[52] ,
         dpath_mulcore_ary1_a1_s2[51] , dpath_mulcore_ary1_a1_s2[50] ,
         dpath_mulcore_ary1_a1_s2[49] , dpath_mulcore_ary1_a1_s2[48] ,
         dpath_mulcore_ary1_a1_s2[47] , dpath_mulcore_ary1_a1_s2[46] ,
         dpath_mulcore_ary1_a1_s2[45] , dpath_mulcore_ary1_a1_s2[44] ,
         dpath_mulcore_ary1_a1_s2[43] , dpath_mulcore_ary1_a1_s2[42] ,
         dpath_mulcore_ary1_a1_s2[41] , dpath_mulcore_ary1_a1_s2[40] ,
         dpath_mulcore_ary1_a1_s2[39] , dpath_mulcore_ary1_a1_s2[38] ,
         dpath_mulcore_ary1_a1_s2[37] , dpath_mulcore_ary1_a1_s2[36] ,
         dpath_mulcore_ary1_a1_s2[35] , dpath_mulcore_ary1_a1_s2[34] ,
         dpath_mulcore_ary1_a1_s2[33] , dpath_mulcore_ary1_a1_s2[32] ,
         dpath_mulcore_ary1_a1_s2[31] , dpath_mulcore_ary1_a1_s2[30] ,
         dpath_mulcore_ary1_a1_s2[29] , dpath_mulcore_ary1_a1_s2[28] ,
         dpath_mulcore_ary1_a1_s2[27] , dpath_mulcore_ary1_a1_s2[26] ,
         dpath_mulcore_ary1_a1_s2[25] , dpath_mulcore_ary1_a1_s2[24] ,
         dpath_mulcore_ary1_a1_s2[23] , dpath_mulcore_ary1_a1_s2[22] ,
         dpath_mulcore_ary1_a1_s2[21] , dpath_mulcore_ary1_a1_s2[20] ,
         dpath_mulcore_ary1_a1_s2[19] , dpath_mulcore_ary1_a1_s2[18] ,
         dpath_mulcore_ary1_a1_s2[17] , dpath_mulcore_ary1_a1_s2[16] ,
         dpath_mulcore_ary1_a1_s2[15] , dpath_mulcore_ary1_a1_s2[14] ,
         dpath_mulcore_ary1_a1_s2[13] , dpath_mulcore_ary1_a1_s2[12] ,
         dpath_mulcore_ary1_a1_s2[11] , dpath_mulcore_ary1_a1_s2[10] ,
         dpath_mulcore_ary1_a1_s2[9] , dpath_mulcore_ary1_a1_s2[8] ,
         dpath_mulcore_ary1_a1_s2[7] , dpath_mulcore_ary1_a1_s2[6] ,
         dpath_mulcore_ary1_a1_s2[5] , dpath_mulcore_ary1_a1_s2[4] ,
         dpath_mulcore_ary1_a1_s2[3] , dpath_mulcore_ary1_a1_s2[2] ,
         dpath_mulcore_ary1_a1_s2[1] , dpath_mulcore_ary1_a1_s2[0] ,
         dpath_mulcore_ary1_a1_c2[66] , dpath_mulcore_ary1_a1_c2[65] ,
         dpath_mulcore_ary1_a1_c2[64] , dpath_mulcore_ary1_a1_c2[63] ,
         dpath_mulcore_ary1_a1_c2[62] , dpath_mulcore_ary1_a1_c2[61] ,
         dpath_mulcore_ary1_a1_c2[60] , dpath_mulcore_ary1_a1_c2[59] ,
         dpath_mulcore_ary1_a1_c2[58] , dpath_mulcore_ary1_a1_c2[57] ,
         dpath_mulcore_ary1_a1_c2[56] , dpath_mulcore_ary1_a1_c2[55] ,
         dpath_mulcore_ary1_a1_c2[54] , dpath_mulcore_ary1_a1_c2[53] ,
         dpath_mulcore_ary1_a1_c2[52] , dpath_mulcore_ary1_a1_c2[51] ,
         dpath_mulcore_ary1_a1_c2[50] , dpath_mulcore_ary1_a1_c2[49] ,
         dpath_mulcore_ary1_a1_c2[48] , dpath_mulcore_ary1_a1_c2[47] ,
         dpath_mulcore_ary1_a1_c2[46] , dpath_mulcore_ary1_a1_c2[45] ,
         dpath_mulcore_ary1_a1_c2[44] , dpath_mulcore_ary1_a1_c2[43] ,
         dpath_mulcore_ary1_a1_c2[42] , dpath_mulcore_ary1_a1_c2[41] ,
         dpath_mulcore_ary1_a1_c2[40] , dpath_mulcore_ary1_a1_c2[39] ,
         dpath_mulcore_ary1_a1_c2[38] , dpath_mulcore_ary1_a1_c2[37] ,
         dpath_mulcore_ary1_a1_c2[36] , dpath_mulcore_ary1_a1_c2[35] ,
         dpath_mulcore_ary1_a1_c2[34] , dpath_mulcore_ary1_a1_c2[33] ,
         dpath_mulcore_ary1_a1_c2[32] , dpath_mulcore_ary1_a1_c2[31] ,
         dpath_mulcore_ary1_a1_c2[30] , dpath_mulcore_ary1_a1_c2[29] ,
         dpath_mulcore_ary1_a1_c2[28] , dpath_mulcore_ary1_a1_c2[27] ,
         dpath_mulcore_ary1_a1_c2[26] , dpath_mulcore_ary1_a1_c2[25] ,
         dpath_mulcore_ary1_a1_c2[24] , dpath_mulcore_ary1_a1_c2[23] ,
         dpath_mulcore_ary1_a1_c2[22] , dpath_mulcore_ary1_a1_c2[21] ,
         dpath_mulcore_ary1_a1_c2[20] , dpath_mulcore_ary1_a1_c2[19] ,
         dpath_mulcore_ary1_a1_c2[18] , dpath_mulcore_ary1_a1_c2[17] ,
         dpath_mulcore_ary1_a1_c2[16] , dpath_mulcore_ary1_a1_c2[15] ,
         dpath_mulcore_ary1_a1_c2[14] , dpath_mulcore_ary1_a1_c2[13] ,
         dpath_mulcore_ary1_a1_c2[12] , dpath_mulcore_ary1_a1_c2[11] ,
         dpath_mulcore_ary1_a1_c2[10] , dpath_mulcore_ary1_a1_c2[9] ,
         dpath_mulcore_ary1_a1_c2[8] , dpath_mulcore_ary1_a1_c2[7] ,
         dpath_mulcore_ary1_a1_c2[6] , dpath_mulcore_ary1_a1_c2[5] ,
         dpath_mulcore_ary1_a1_c2[4] , dpath_mulcore_ary1_a1_c2[3] ,
         dpath_mulcore_ary1_a1_c2[2] , dpath_mulcore_ary1_a1_c2[1] ,
         dpath_mulcore_ary1_a1_c1[66] , dpath_mulcore_ary1_a1_c1[65] ,
         dpath_mulcore_ary1_a1_c1[64] , dpath_mulcore_ary1_a1_c1[63] ,
         dpath_mulcore_ary1_a1_c1[62] , dpath_mulcore_ary1_a1_c1[61] ,
         dpath_mulcore_ary1_a1_c1[60] , dpath_mulcore_ary1_a1_c1[59] ,
         dpath_mulcore_ary1_a1_c1[58] , dpath_mulcore_ary1_a1_c1[57] ,
         dpath_mulcore_ary1_a1_c1[56] , dpath_mulcore_ary1_a1_c1[55] ,
         dpath_mulcore_ary1_a1_c1[54] , dpath_mulcore_ary1_a1_c1[53] ,
         dpath_mulcore_ary1_a1_c1[52] , dpath_mulcore_ary1_a1_c1[51] ,
         dpath_mulcore_ary1_a1_c1[50] , dpath_mulcore_ary1_a1_c1[49] ,
         dpath_mulcore_ary1_a1_c1[48] , dpath_mulcore_ary1_a1_c1[47] ,
         dpath_mulcore_ary1_a1_c1[46] , dpath_mulcore_ary1_a1_c1[45] ,
         dpath_mulcore_ary1_a1_c1[44] , dpath_mulcore_ary1_a1_c1[43] ,
         dpath_mulcore_ary1_a1_c1[42] , dpath_mulcore_ary1_a1_c1[41] ,
         dpath_mulcore_ary1_a1_c1[40] , dpath_mulcore_ary1_a1_c1[39] ,
         dpath_mulcore_ary1_a1_c1[38] , dpath_mulcore_ary1_a1_c1[37] ,
         dpath_mulcore_ary1_a1_c1[36] , dpath_mulcore_ary1_a1_c1[35] ,
         dpath_mulcore_ary1_a1_c1[34] , dpath_mulcore_ary1_a1_c1[33] ,
         dpath_mulcore_ary1_a1_c1[32] , dpath_mulcore_ary1_a1_c1[31] ,
         dpath_mulcore_ary1_a1_c1[30] , dpath_mulcore_ary1_a1_c1[29] ,
         dpath_mulcore_ary1_a1_c1[28] , dpath_mulcore_ary1_a1_c1[27] ,
         dpath_mulcore_ary1_a1_c1[26] , dpath_mulcore_ary1_a1_c1[25] ,
         dpath_mulcore_ary1_a1_c1[24] , dpath_mulcore_ary1_a1_c1[23] ,
         dpath_mulcore_ary1_a1_c1[22] , dpath_mulcore_ary1_a1_c1[21] ,
         dpath_mulcore_ary1_a1_c1[20] , dpath_mulcore_ary1_a1_c1[19] ,
         dpath_mulcore_ary1_a1_c1[18] , dpath_mulcore_ary1_a1_c1[17] ,
         dpath_mulcore_ary1_a1_c1[16] , dpath_mulcore_ary1_a1_c1[15] ,
         dpath_mulcore_ary1_a1_c1[14] , dpath_mulcore_ary1_a1_c1[13] ,
         dpath_mulcore_ary1_a1_c1[12] , dpath_mulcore_ary1_a1_c1[11] ,
         dpath_mulcore_ary1_a1_c1[10] , dpath_mulcore_ary1_a1_c1[9] ,
         dpath_mulcore_ary1_a1_c1[8] , dpath_mulcore_ary1_a1_c1[7] ,
         dpath_mulcore_ary1_a1_c1[6] , dpath_mulcore_ary1_a1_c1[5] ,
         dpath_mulcore_ary1_a1_c1[4] , dpath_mulcore_ary1_a1_c1[3] ,
         dpath_mulcore_ary1_a1_c1[2] , dpath_mulcore_ary1_a1_c1[1] ,
         dpath_mulcore_ary1_a1_s_1[69] , dpath_mulcore_ary1_a1_s_1[68] ,
         dpath_mulcore_ary1_a1_s_1[67] , dpath_mulcore_ary1_a1_s_1[66] ,
         dpath_mulcore_ary1_a1_s_1[65] , dpath_mulcore_ary1_a1_s_1[64] ,
         dpath_mulcore_ary1_a1_s_1[63] , dpath_mulcore_ary1_a1_s_1[62] ,
         dpath_mulcore_ary1_a1_s_1[61] , dpath_mulcore_ary1_a1_s_1[60] ,
         dpath_mulcore_ary1_a1_s_1[59] , dpath_mulcore_ary1_a1_s_1[58] ,
         dpath_mulcore_ary1_a1_s_1[57] , dpath_mulcore_ary1_a1_s_1[56] ,
         dpath_mulcore_ary1_a1_s_1[55] , dpath_mulcore_ary1_a1_s_1[54] ,
         dpath_mulcore_ary1_a1_s_1[53] , dpath_mulcore_ary1_a1_s_1[52] ,
         dpath_mulcore_ary1_a1_s_1[51] , dpath_mulcore_ary1_a1_s_1[50] ,
         dpath_mulcore_ary1_a1_s_1[49] , dpath_mulcore_ary1_a1_s_1[48] ,
         dpath_mulcore_ary1_a1_s_1[47] , dpath_mulcore_ary1_a1_s_1[46] ,
         dpath_mulcore_ary1_a1_s_1[45] , dpath_mulcore_ary1_a1_s_1[44] ,
         dpath_mulcore_ary1_a1_s_1[43] , dpath_mulcore_ary1_a1_s_1[42] ,
         dpath_mulcore_ary1_a1_s_1[41] , dpath_mulcore_ary1_a1_s_1[40] ,
         dpath_mulcore_ary1_a1_s_1[39] , dpath_mulcore_ary1_a1_s_1[38] ,
         dpath_mulcore_ary1_a1_s_1[37] , dpath_mulcore_ary1_a1_s_1[36] ,
         dpath_mulcore_ary1_a1_s_1[35] , dpath_mulcore_ary1_a1_s_1[34] ,
         dpath_mulcore_ary1_a1_s_1[33] , dpath_mulcore_ary1_a1_s_1[32] ,
         dpath_mulcore_ary1_a1_s_1[31] , dpath_mulcore_ary1_a1_s_1[30] ,
         dpath_mulcore_ary1_a1_s_1[29] , dpath_mulcore_ary1_a1_s_1[28] ,
         dpath_mulcore_ary1_a1_s_1[27] , dpath_mulcore_ary1_a1_s_1[26] ,
         dpath_mulcore_ary1_a1_s_1[25] , dpath_mulcore_ary1_a1_s_1[24] ,
         dpath_mulcore_ary1_a1_s_1[23] , dpath_mulcore_ary1_a1_s_1[22] ,
         dpath_mulcore_ary1_a1_s_1[21] , dpath_mulcore_ary1_a1_s_1[20] ,
         dpath_mulcore_ary1_a1_s_1[19] , dpath_mulcore_ary1_a1_s_1[18] ,
         dpath_mulcore_ary1_a1_s_1[17] , dpath_mulcore_ary1_a1_s_1[16] ,
         dpath_mulcore_ary1_a1_s_1[15] , dpath_mulcore_ary1_a1_s_1[14] ,
         dpath_mulcore_ary1_a1_s_1[13] , dpath_mulcore_ary1_a1_s_1[12] ,
         dpath_mulcore_ary1_a1_s_1[11] , dpath_mulcore_ary1_a1_s_1[10] ,
         dpath_mulcore_ary1_a1_s_1[9] , dpath_mulcore_ary1_a1_s_1[8] ,
         dpath_mulcore_ary1_a1_s_1[7] , dpath_mulcore_ary1_a1_s_1[6] ,
         dpath_mulcore_ary1_a1_s_1[5] , dpath_mulcore_ary1_a1_s_1[4] ,
         dpath_mulcore_ary1_a1_s1[67] , dpath_mulcore_ary1_a1_s1[66] ,
         dpath_mulcore_ary1_a1_s1[65] , dpath_mulcore_ary1_a1_s1[64] ,
         dpath_mulcore_ary1_a1_s1[63] , dpath_mulcore_ary1_a1_s1[62] ,
         dpath_mulcore_ary1_a1_s1[61] , dpath_mulcore_ary1_a1_s1[60] ,
         dpath_mulcore_ary1_a1_s1[59] , dpath_mulcore_ary1_a1_s1[58] ,
         dpath_mulcore_ary1_a1_s1[57] , dpath_mulcore_ary1_a1_s1[56] ,
         dpath_mulcore_ary1_a1_s1[55] , dpath_mulcore_ary1_a1_s1[54] ,
         dpath_mulcore_ary1_a1_s1[53] , dpath_mulcore_ary1_a1_s1[52] ,
         dpath_mulcore_ary1_a1_s1[51] , dpath_mulcore_ary1_a1_s1[50] ,
         dpath_mulcore_ary1_a1_s1[49] , dpath_mulcore_ary1_a1_s1[48] ,
         dpath_mulcore_ary1_a1_s1[47] , dpath_mulcore_ary1_a1_s1[46] ,
         dpath_mulcore_ary1_a1_s1[45] , dpath_mulcore_ary1_a1_s1[44] ,
         dpath_mulcore_ary1_a1_s1[43] , dpath_mulcore_ary1_a1_s1[42] ,
         dpath_mulcore_ary1_a1_s1[41] , dpath_mulcore_ary1_a1_s1[40] ,
         dpath_mulcore_ary1_a1_s1[39] , dpath_mulcore_ary1_a1_s1[38] ,
         dpath_mulcore_ary1_a1_s1[37] , dpath_mulcore_ary1_a1_s1[36] ,
         dpath_mulcore_ary1_a1_s1[35] , dpath_mulcore_ary1_a1_s1[34] ,
         dpath_mulcore_ary1_a1_s1[33] , dpath_mulcore_ary1_a1_s1[32] ,
         dpath_mulcore_ary1_a1_s1[31] , dpath_mulcore_ary1_a1_s1[30] ,
         dpath_mulcore_ary1_a1_s1[29] , dpath_mulcore_ary1_a1_s1[28] ,
         dpath_mulcore_ary1_a1_s1[27] , dpath_mulcore_ary1_a1_s1[26] ,
         dpath_mulcore_ary1_a1_s1[25] , dpath_mulcore_ary1_a1_s1[24] ,
         dpath_mulcore_ary1_a1_s1[23] , dpath_mulcore_ary1_a1_s1[22] ,
         dpath_mulcore_ary1_a1_s1[21] , dpath_mulcore_ary1_a1_s1[20] ,
         dpath_mulcore_ary1_a1_s1[19] , dpath_mulcore_ary1_a1_s1[18] ,
         dpath_mulcore_ary1_a1_s1[17] , dpath_mulcore_ary1_a1_s1[16] ,
         dpath_mulcore_ary1_a1_s1[15] , dpath_mulcore_ary1_a1_s1[14] ,
         dpath_mulcore_ary1_a1_s1[13] , dpath_mulcore_ary1_a1_s1[12] ,
         dpath_mulcore_ary1_a1_s1[11] , dpath_mulcore_ary1_a1_s1[10] ,
         dpath_mulcore_ary1_a1_s1[9] , dpath_mulcore_ary1_a1_s1[8] ,
         dpath_mulcore_ary1_a1_s1[7] , dpath_mulcore_ary1_a1_s1[6] ,
         dpath_mulcore_ary1_a1_s1[5] , dpath_mulcore_ary1_a1_s1[4] ,
         dpath_mulcore_ary1_a1_s1[3] , dpath_mulcore_ary1_a1_s1[2] ,
         dpath_mulcore_ary1_a1_s1[1] , dpath_mulcore_ary1_a1_s1[0] ,
         dpath_mulcore_ary1_a1_c_2[76] , dpath_mulcore_ary1_a1_c_2[75] ,
         dpath_mulcore_ary1_a1_c_2[74] , dpath_mulcore_ary1_a1_c_2[73] ,
         dpath_mulcore_ary1_a1_c_2[72] , dpath_mulcore_ary1_a1_c_2[71] ,
         dpath_mulcore_ary1_a1_c_2[70] , dpath_mulcore_ary1_a1_c_2[69] ,
         dpath_mulcore_ary1_a1_c_2[68] , dpath_mulcore_ary1_a1_c_2[67] ,
         dpath_mulcore_ary1_a1_c_2[66] , dpath_mulcore_ary1_a1_c_2[65] ,
         dpath_mulcore_ary1_a1_c_2[64] , dpath_mulcore_ary1_a1_c_2[63] ,
         dpath_mulcore_ary1_a1_c_2[62] , dpath_mulcore_ary1_a1_c_2[61] ,
         dpath_mulcore_ary1_a1_c_2[60] , dpath_mulcore_ary1_a1_c_2[59] ,
         dpath_mulcore_ary1_a1_c_2[58] , dpath_mulcore_ary1_a1_c_2[57] ,
         dpath_mulcore_ary1_a1_c_2[56] , dpath_mulcore_ary1_a1_c_2[55] ,
         dpath_mulcore_ary1_a1_c_2[54] , dpath_mulcore_ary1_a1_c_2[53] ,
         dpath_mulcore_ary1_a1_c_2[52] , dpath_mulcore_ary1_a1_c_2[51] ,
         dpath_mulcore_ary1_a1_c_2[50] , dpath_mulcore_ary1_a1_c_2[49] ,
         dpath_mulcore_ary1_a1_c_2[48] , dpath_mulcore_ary1_a1_c_2[47] ,
         dpath_mulcore_ary1_a1_c_2[46] , dpath_mulcore_ary1_a1_c_2[45] ,
         dpath_mulcore_ary1_a1_c_2[44] , dpath_mulcore_ary1_a1_c_2[43] ,
         dpath_mulcore_ary1_a1_c_2[42] , dpath_mulcore_ary1_a1_c_2[41] ,
         dpath_mulcore_ary1_a1_c_2[40] , dpath_mulcore_ary1_a1_c_2[39] ,
         dpath_mulcore_ary1_a1_c_2[38] , dpath_mulcore_ary1_a1_c_2[37] ,
         dpath_mulcore_ary1_a1_c_2[36] , dpath_mulcore_ary1_a1_c_2[35] ,
         dpath_mulcore_ary1_a1_c_2[34] , dpath_mulcore_ary1_a1_c_2[33] ,
         dpath_mulcore_ary1_a1_c_2[32] , dpath_mulcore_ary1_a1_c_2[31] ,
         dpath_mulcore_ary1_a1_c_2[30] , dpath_mulcore_ary1_a1_c_2[29] ,
         dpath_mulcore_ary1_a1_c_2[28] , dpath_mulcore_ary1_a1_c_2[27] ,
         dpath_mulcore_ary1_a1_c_2[26] , dpath_mulcore_ary1_a1_c_2[25] ,
         dpath_mulcore_ary1_a1_c_2[24] , dpath_mulcore_ary1_a1_c_2[23] ,
         dpath_mulcore_ary1_a1_c_2[22] , dpath_mulcore_ary1_a1_c_2[21] ,
         dpath_mulcore_ary1_a1_c_2[20] , dpath_mulcore_ary1_a1_c_2[19] ,
         dpath_mulcore_ary1_a1_c_2[18] , dpath_mulcore_ary1_a1_c_2[17] ,
         dpath_mulcore_ary1_a1_c_2[16] , dpath_mulcore_ary1_a1_c_2[15] ,
         dpath_mulcore_ary1_a1_c_2[14] , dpath_mulcore_ary1_a1_c_2[13] ,
         dpath_mulcore_ary1_a1_c_2[12] , dpath_mulcore_ary1_a1_c_2[11] ,
         dpath_mulcore_ary1_a1_c_2[10] , dpath_mulcore_ary1_a1_c_1[69] ,
         dpath_mulcore_ary1_a1_c_1[68] , dpath_mulcore_ary1_a1_c_1[67] ,
         dpath_mulcore_ary1_a1_c_1[66] , dpath_mulcore_ary1_a1_c_1[65] ,
         dpath_mulcore_ary1_a1_c_1[64] , dpath_mulcore_ary1_a1_c_1[63] ,
         dpath_mulcore_ary1_a1_c_1[62] , dpath_mulcore_ary1_a1_c_1[61] ,
         dpath_mulcore_ary1_a1_c_1[60] , dpath_mulcore_ary1_a1_c_1[59] ,
         dpath_mulcore_ary1_a1_c_1[58] , dpath_mulcore_ary1_a1_c_1[57] ,
         dpath_mulcore_ary1_a1_c_1[56] , dpath_mulcore_ary1_a1_c_1[55] ,
         dpath_mulcore_ary1_a1_c_1[54] , dpath_mulcore_ary1_a1_c_1[53] ,
         dpath_mulcore_ary1_a1_c_1[52] , dpath_mulcore_ary1_a1_c_1[51] ,
         dpath_mulcore_ary1_a1_c_1[50] , dpath_mulcore_ary1_a1_c_1[49] ,
         dpath_mulcore_ary1_a1_c_1[48] , dpath_mulcore_ary1_a1_c_1[47] ,
         dpath_mulcore_ary1_a1_c_1[46] , dpath_mulcore_ary1_a1_c_1[45] ,
         dpath_mulcore_ary1_a1_c_1[44] , dpath_mulcore_ary1_a1_c_1[43] ,
         dpath_mulcore_ary1_a1_c_1[42] , dpath_mulcore_ary1_a1_c_1[41] ,
         dpath_mulcore_ary1_a1_c_1[40] , dpath_mulcore_ary1_a1_c_1[39] ,
         dpath_mulcore_ary1_a1_c_1[38] , dpath_mulcore_ary1_a1_c_1[37] ,
         dpath_mulcore_ary1_a1_c_1[36] , dpath_mulcore_ary1_a1_c_1[35] ,
         dpath_mulcore_ary1_a1_c_1[34] , dpath_mulcore_ary1_a1_c_1[33] ,
         dpath_mulcore_ary1_a1_c_1[32] , dpath_mulcore_ary1_a1_c_1[31] ,
         dpath_mulcore_ary1_a1_c_1[30] , dpath_mulcore_ary1_a1_c_1[29] ,
         dpath_mulcore_ary1_a1_c_1[28] , dpath_mulcore_ary1_a1_c_1[27] ,
         dpath_mulcore_ary1_a1_c_1[26] , dpath_mulcore_ary1_a1_c_1[25] ,
         dpath_mulcore_ary1_a1_c_1[24] , dpath_mulcore_ary1_a1_c_1[23] ,
         dpath_mulcore_ary1_a1_c_1[22] , dpath_mulcore_ary1_a1_c_1[21] ,
         dpath_mulcore_ary1_a1_c_1[20] , dpath_mulcore_ary1_a1_c_1[19] ,
         dpath_mulcore_ary1_a1_c_1[18] , dpath_mulcore_ary1_a1_c_1[17] ,
         dpath_mulcore_ary1_a1_c_1[16] , dpath_mulcore_ary1_a1_c_1[15] ,
         dpath_mulcore_ary1_a1_c_1[14] , dpath_mulcore_ary1_a1_c_1[13] ,
         dpath_mulcore_ary1_a1_c_1[12] , dpath_mulcore_ary1_a1_c_1[11] ,
         dpath_mulcore_ary1_a1_c_1[10] , dpath_mulcore_ary1_a1_c_1[9] ,
         dpath_mulcore_ary1_a1_c_1[8] , dpath_mulcore_ary1_a1_c_1[7] ,
         dpath_mulcore_ary1_a1_c_1[6] , dpath_mulcore_ary1_a1_c_1[5] ,
         dpath_mulcore_ary1_a1_c_1[4] , dpath_mulcore_ary1_a1_c_1[3] ,
         dpath_mulcore_ary1_a1_c_1[2] , dpath_mulcore_ary1_a1_co[71] ,
         dpath_mulcore_ary1_a1_co[70] , dpath_mulcore_ary1_a1_co[69] ,
         dpath_mulcore_ary1_a1_co[68] , dpath_mulcore_ary1_a1_co[67] ,
         dpath_mulcore_ary1_a1_co[66] , dpath_mulcore_ary1_a1_co[65] ,
         dpath_mulcore_ary1_a1_co[64] , dpath_mulcore_ary1_a1_co[63] ,
         dpath_mulcore_ary1_a1_co[62] , dpath_mulcore_ary1_a1_co[61] ,
         dpath_mulcore_ary1_a1_co[60] , dpath_mulcore_ary1_a1_co[59] ,
         dpath_mulcore_ary1_a1_co[58] , dpath_mulcore_ary1_a1_co[57] ,
         dpath_mulcore_ary1_a1_co[56] , dpath_mulcore_ary1_a1_co[55] ,
         dpath_mulcore_ary1_a1_co[54] , dpath_mulcore_ary1_a1_co[53] ,
         dpath_mulcore_ary1_a1_co[52] , dpath_mulcore_ary1_a1_co[51] ,
         dpath_mulcore_ary1_a1_co[50] , dpath_mulcore_ary1_a1_co[49] ,
         dpath_mulcore_ary1_a1_co[48] , dpath_mulcore_ary1_a1_co[47] ,
         dpath_mulcore_ary1_a1_co[46] , dpath_mulcore_ary1_a1_co[45] ,
         dpath_mulcore_ary1_a1_co[44] , dpath_mulcore_ary1_a1_co[43] ,
         dpath_mulcore_ary1_a1_co[42] , dpath_mulcore_ary1_a1_co[41] ,
         dpath_mulcore_ary1_a1_co[40] , dpath_mulcore_ary1_a1_co[39] ,
         dpath_mulcore_ary1_a1_co[38] , dpath_mulcore_ary1_a1_co[37] ,
         dpath_mulcore_ary1_a1_co[36] , dpath_mulcore_ary1_a1_co[35] ,
         dpath_mulcore_ary1_a1_co[34] , dpath_mulcore_ary1_a1_co[33] ,
         dpath_mulcore_ary1_a1_co[32] , dpath_mulcore_ary1_a1_co[31] ,
         dpath_mulcore_ary1_a1_co[30] , dpath_mulcore_ary1_a1_co[29] ,
         dpath_mulcore_ary1_a1_co[28] , dpath_mulcore_ary1_a1_co[27] ,
         dpath_mulcore_ary1_a1_co[26] , dpath_mulcore_ary1_a1_co[25] ,
         dpath_mulcore_ary1_a1_co[24] , dpath_mulcore_ary1_a1_co[23] ,
         dpath_mulcore_ary1_a1_co[22] , dpath_mulcore_ary1_a1_co[21] ,
         dpath_mulcore_ary1_a1_co[20] , dpath_mulcore_ary1_a1_co[19] ,
         dpath_mulcore_ary1_a1_co[18] , dpath_mulcore_ary1_a1_co[17] ,
         dpath_mulcore_ary1_a1_co[16] , dpath_mulcore_ary1_a1_co[15] ,
         dpath_mulcore_ary1_a1_co[14] , dpath_mulcore_ary1_a1_co[13] ,
         dpath_mulcore_ary1_a1_co[12] , dpath_mulcore_ary1_a1_co[11] ,
         dpath_mulcore_ary1_a1_s_2[75] , dpath_mulcore_ary1_a1_s_2[74] ,
         dpath_mulcore_ary1_a1_s_2[73] , dpath_mulcore_ary1_a1_s_2[72] ,
         dpath_mulcore_ary1_a1_s_2[71] , dpath_mulcore_ary1_a1_s_2[70] ,
         dpath_mulcore_ary1_a1_s_2[69] , dpath_mulcore_ary1_a1_s_2[68] ,
         dpath_mulcore_ary1_a1_s_2[67] , dpath_mulcore_ary1_a1_s_2[66] ,
         dpath_mulcore_ary1_a1_s_2[65] , dpath_mulcore_ary1_a1_s_2[64] ,
         dpath_mulcore_ary1_a1_s_2[63] , dpath_mulcore_ary1_a1_s_2[62] ,
         dpath_mulcore_ary1_a1_s_2[61] , dpath_mulcore_ary1_a1_s_2[60] ,
         dpath_mulcore_ary1_a1_s_2[59] , dpath_mulcore_ary1_a1_s_2[58] ,
         dpath_mulcore_ary1_a1_s_2[57] , dpath_mulcore_ary1_a1_s_2[56] ,
         dpath_mulcore_ary1_a1_s_2[55] , dpath_mulcore_ary1_a1_s_2[54] ,
         dpath_mulcore_ary1_a1_s_2[53] , dpath_mulcore_ary1_a1_s_2[52] ,
         dpath_mulcore_ary1_a1_s_2[51] , dpath_mulcore_ary1_a1_s_2[50] ,
         dpath_mulcore_ary1_a1_s_2[49] , dpath_mulcore_ary1_a1_s_2[48] ,
         dpath_mulcore_ary1_a1_s_2[47] , dpath_mulcore_ary1_a1_s_2[46] ,
         dpath_mulcore_ary1_a1_s_2[45] , dpath_mulcore_ary1_a1_s_2[44] ,
         dpath_mulcore_ary1_a1_s_2[43] , dpath_mulcore_ary1_a1_s_2[42] ,
         dpath_mulcore_ary1_a1_s_2[41] , dpath_mulcore_ary1_a1_s_2[40] ,
         dpath_mulcore_ary1_a1_s_2[39] , dpath_mulcore_ary1_a1_s_2[38] ,
         dpath_mulcore_ary1_a1_s_2[37] , dpath_mulcore_ary1_a1_s_2[36] ,
         dpath_mulcore_ary1_a1_s_2[35] , dpath_mulcore_ary1_a1_s_2[34] ,
         dpath_mulcore_ary1_a1_s_2[33] , dpath_mulcore_ary1_a1_s_2[32] ,
         dpath_mulcore_ary1_a1_s_2[31] , dpath_mulcore_ary1_a1_s_2[30] ,
         dpath_mulcore_ary1_a1_s_2[29] , dpath_mulcore_ary1_a1_s_2[28] ,
         dpath_mulcore_ary1_a1_s_2[27] , dpath_mulcore_ary1_a1_s_2[26] ,
         dpath_mulcore_ary1_a1_s_2[25] , dpath_mulcore_ary1_a1_s_2[24] ,
         dpath_mulcore_ary1_a1_s_2[23] , dpath_mulcore_ary1_a1_s_2[22] ,
         dpath_mulcore_ary1_a1_s_2[21] , dpath_mulcore_ary1_a1_s_2[20] ,
         dpath_mulcore_ary1_a1_s_2[19] , dpath_mulcore_ary1_a1_s_2[18] ,
         dpath_mulcore_ary1_a1_s_2[17] , dpath_mulcore_ary1_a1_s_2[16] ,
         dpath_mulcore_ary1_a1_s_2[15] , dpath_mulcore_ary1_a1_s_2[14] ,
         dpath_mulcore_ary1_a1_s_2[13] , dpath_mulcore_ary1_a1_s_2[12] ,
         dpath_mulcore_ary1_a1_s_2[11] , dpath_mulcore_ary1_a1_s_2[10] ,
         dpath_mulcore_ary1_a1_b2n[1] , dpath_mulcore_ary1_a1_b2n[0] ,
         dpath_mulcore_ary1_a1_b5n[1] , dpath_mulcore_ary1_a1_b5n[0] ,
         dpath_mulcore_array2_c1x2 , dpath_mulcore_array2_s1x2 ,
         dpath_mulcore_array2_c1[82] , dpath_mulcore_array2_c1[81] ,
         dpath_mulcore_array2_c1[80] , dpath_mulcore_array2_c1[79] ,
         dpath_mulcore_array2_c1[78] , dpath_mulcore_array2_c1[77] ,
         dpath_mulcore_array2_c1[76] , dpath_mulcore_array2_c1[75] ,
         dpath_mulcore_array2_c1[74] , dpath_mulcore_array2_c1[73] ,
         dpath_mulcore_array2_c1[72] , dpath_mulcore_array2_c1[71] ,
         dpath_mulcore_array2_c1[70] , dpath_mulcore_array2_c1[69] ,
         dpath_mulcore_array2_c1[68] , dpath_mulcore_array2_c1[67] ,
         dpath_mulcore_array2_c1[66] , dpath_mulcore_array2_c1[65] ,
         dpath_mulcore_array2_c1[64] , dpath_mulcore_array2_c1[63] ,
         dpath_mulcore_array2_c1[62] , dpath_mulcore_array2_c1[61] ,
         dpath_mulcore_array2_c1[60] , dpath_mulcore_array2_c1[59] ,
         dpath_mulcore_array2_c1[58] , dpath_mulcore_array2_c1[57] ,
         dpath_mulcore_array2_c1[56] , dpath_mulcore_array2_c1[55] ,
         dpath_mulcore_array2_c1[54] , dpath_mulcore_array2_c1[53] ,
         dpath_mulcore_array2_c1[52] , dpath_mulcore_array2_c1[51] ,
         dpath_mulcore_array2_c1[50] , dpath_mulcore_array2_c1[49] ,
         dpath_mulcore_array2_c1[48] , dpath_mulcore_array2_c1[47] ,
         dpath_mulcore_array2_c1[46] , dpath_mulcore_array2_c1[45] ,
         dpath_mulcore_array2_c1[44] , dpath_mulcore_array2_c1[43] ,
         dpath_mulcore_array2_c1[42] , dpath_mulcore_array2_c1[41] ,
         dpath_mulcore_array2_c1[40] , dpath_mulcore_array2_c1[39] ,
         dpath_mulcore_array2_c1[38] , dpath_mulcore_array2_c1[37] ,
         dpath_mulcore_array2_c1[36] , dpath_mulcore_array2_c1[35] ,
         dpath_mulcore_array2_c1[34] , dpath_mulcore_array2_c1[33] ,
         dpath_mulcore_array2_c1[32] , dpath_mulcore_array2_c1[31] ,
         dpath_mulcore_array2_c1[30] , dpath_mulcore_array2_c1[29] ,
         dpath_mulcore_array2_c1[28] , dpath_mulcore_array2_c1[27] ,
         dpath_mulcore_array2_c1[26] , dpath_mulcore_array2_c1[25] ,
         dpath_mulcore_array2_c1[24] , dpath_mulcore_array2_c1[23] ,
         dpath_mulcore_array2_c1[22] , dpath_mulcore_array2_c1[21] ,
         dpath_mulcore_array2_c1[20] , dpath_mulcore_array2_c1[19] ,
         dpath_mulcore_array2_c1[18] , dpath_mulcore_array2_c1[17] ,
         dpath_mulcore_array2_c1[16] , dpath_mulcore_array2_c1[14] ,
         dpath_mulcore_array2_c1[13] , dpath_mulcore_array2_c1[12] ,
         dpath_mulcore_array2_c1[11] , dpath_mulcore_array2_c1[10] ,
         dpath_mulcore_array2_c1[9] , dpath_mulcore_array2_c1[8] ,
         dpath_mulcore_array2_c1[7] , dpath_mulcore_array2_c1[6] ,
         dpath_mulcore_array2_c1[5] , dpath_mulcore_array2_c1[4] ,
         dpath_mulcore_array2_c1[3] , dpath_mulcore_array2_c1[2] ,
         dpath_mulcore_array2_c1[1] , dpath_mulcore_array2_c1[0] ,
         dpath_mulcore_array2_s1[82] , dpath_mulcore_array2_s1[81] ,
         dpath_mulcore_array2_s1[80] , dpath_mulcore_array2_s1[79] ,
         dpath_mulcore_array2_s1[78] , dpath_mulcore_array2_s1[77] ,
         dpath_mulcore_array2_s1[76] , dpath_mulcore_array2_s1[75] ,
         dpath_mulcore_array2_s1[74] , dpath_mulcore_array2_s1[73] ,
         dpath_mulcore_array2_s1[72] , dpath_mulcore_array2_s1[71] ,
         dpath_mulcore_array2_s1[70] , dpath_mulcore_array2_s1[69] ,
         dpath_mulcore_array2_s1[68] , dpath_mulcore_array2_s1[67] ,
         dpath_mulcore_array2_s1[66] , dpath_mulcore_array2_s1[65] ,
         dpath_mulcore_array2_s1[64] , dpath_mulcore_array2_s1[63] ,
         dpath_mulcore_array2_s1[62] , dpath_mulcore_array2_s1[61] ,
         dpath_mulcore_array2_s1[60] , dpath_mulcore_array2_s1[59] ,
         dpath_mulcore_array2_s1[58] , dpath_mulcore_array2_s1[57] ,
         dpath_mulcore_array2_s1[56] , dpath_mulcore_array2_s1[55] ,
         dpath_mulcore_array2_s1[54] , dpath_mulcore_array2_s1[53] ,
         dpath_mulcore_array2_s1[52] , dpath_mulcore_array2_s1[51] ,
         dpath_mulcore_array2_s1[50] , dpath_mulcore_array2_s1[49] ,
         dpath_mulcore_array2_s1[48] , dpath_mulcore_array2_s1[47] ,
         dpath_mulcore_array2_s1[46] , dpath_mulcore_array2_s1[45] ,
         dpath_mulcore_array2_s1[44] , dpath_mulcore_array2_s1[43] ,
         dpath_mulcore_array2_s1[42] , dpath_mulcore_array2_s1[41] ,
         dpath_mulcore_array2_s1[40] , dpath_mulcore_array2_s1[39] ,
         dpath_mulcore_array2_s1[38] , dpath_mulcore_array2_s1[37] ,
         dpath_mulcore_array2_s1[36] , dpath_mulcore_array2_s1[35] ,
         dpath_mulcore_array2_s1[34] , dpath_mulcore_array2_s1[33] ,
         dpath_mulcore_array2_s1[32] , dpath_mulcore_array2_s1[31] ,
         dpath_mulcore_array2_s1[30] , dpath_mulcore_array2_s1[29] ,
         dpath_mulcore_array2_s1[28] , dpath_mulcore_array2_s1[27] ,
         dpath_mulcore_array2_s1[26] , dpath_mulcore_array2_s1[25] ,
         dpath_mulcore_array2_s1[24] , dpath_mulcore_array2_s1[23] ,
         dpath_mulcore_array2_s1[22] , dpath_mulcore_array2_s1[21] ,
         dpath_mulcore_array2_s1[20] , dpath_mulcore_array2_s1[19] ,
         dpath_mulcore_array2_s1[18] , dpath_mulcore_array2_s1[17] ,
         dpath_mulcore_array2_s1[16] , dpath_mulcore_array2_s1[14] ,
         dpath_mulcore_array2_s1[13] , dpath_mulcore_array2_s1[12] ,
         dpath_mulcore_array2_s1[11] , dpath_mulcore_array2_s1[10] ,
         dpath_mulcore_array2_s1[9] , dpath_mulcore_array2_s1[8] ,
         dpath_mulcore_array2_s1[7] , dpath_mulcore_array2_s1[6] ,
         dpath_mulcore_array2_s1[5] , dpath_mulcore_array2_s1[4] ,
         dpath_mulcore_array2_s1[3] , dpath_mulcore_array2_s1[2] ,
         dpath_mulcore_array2_s1[1] , dpath_mulcore_array2_s1[0] ,
         dpath_mulcore_array2_s3[81] , dpath_mulcore_array2_s3[80] ,
         dpath_mulcore_array2_s3[79] , dpath_mulcore_array2_s3[78] ,
         dpath_mulcore_array2_s3[77] , dpath_mulcore_array2_s3[76] ,
         dpath_mulcore_array2_s3[75] , dpath_mulcore_array2_s3[74] ,
         dpath_mulcore_array2_s3[73] , dpath_mulcore_array2_s3[72] ,
         dpath_mulcore_array2_s3[71] , dpath_mulcore_array2_s3[70] ,
         dpath_mulcore_array2_s3[69] , dpath_mulcore_array2_s3[68] ,
         dpath_mulcore_array2_s3[67] , dpath_mulcore_array2_s3[66] ,
         dpath_mulcore_array2_s3[65] , dpath_mulcore_array2_s3[64] ,
         dpath_mulcore_array2_s3[63] , dpath_mulcore_array2_s3[62] ,
         dpath_mulcore_array2_s3[61] , dpath_mulcore_array2_s3[60] ,
         dpath_mulcore_array2_s3[59] , dpath_mulcore_array2_s3[58] ,
         dpath_mulcore_array2_s3[57] , dpath_mulcore_array2_s3[56] ,
         dpath_mulcore_array2_s3[55] , dpath_mulcore_array2_s3[54] ,
         dpath_mulcore_array2_s3[53] , dpath_mulcore_array2_s3[52] ,
         dpath_mulcore_array2_s3[51] , dpath_mulcore_array2_s3[50] ,
         dpath_mulcore_array2_s3[49] , dpath_mulcore_array2_s3[48] ,
         dpath_mulcore_array2_s3[47] , dpath_mulcore_array2_s3[46] ,
         dpath_mulcore_array2_s3[45] , dpath_mulcore_array2_s3[44] ,
         dpath_mulcore_array2_s3[43] , dpath_mulcore_array2_s3[42] ,
         dpath_mulcore_array2_s3[41] , dpath_mulcore_array2_s3[40] ,
         dpath_mulcore_array2_s3[39] , dpath_mulcore_array2_s3[38] ,
         dpath_mulcore_array2_s3[37] , dpath_mulcore_array2_s3[36] ,
         dpath_mulcore_array2_s3[35] , dpath_mulcore_array2_s3[34] ,
         dpath_mulcore_array2_s3[33] , dpath_mulcore_array2_s3[32] ,
         dpath_mulcore_array2_s3[31] , dpath_mulcore_array2_s3[30] ,
         dpath_mulcore_array2_s3[29] , dpath_mulcore_array2_s3[28] ,
         dpath_mulcore_array2_s3[27] , dpath_mulcore_array2_s3[26] ,
         dpath_mulcore_array2_s3[25] , dpath_mulcore_array2_s3[24] ,
         dpath_mulcore_array2_s3[23] , dpath_mulcore_array2_s3[22] ,
         dpath_mulcore_array2_s3[21] , dpath_mulcore_array2_s3[19] ,
         dpath_mulcore_array2_s3[18] , dpath_mulcore_array2_s3[17] ,
         dpath_mulcore_array2_s3[16] , dpath_mulcore_array2_s3[15] ,
         dpath_mulcore_array2_s2[96] , dpath_mulcore_array2_s2[95] ,
         dpath_mulcore_array2_s2[94] , dpath_mulcore_array2_s2[93] ,
         dpath_mulcore_array2_s2[92] , dpath_mulcore_array2_s2[91] ,
         dpath_mulcore_array2_s2[90] , dpath_mulcore_array2_s2[89] ,
         dpath_mulcore_array2_s2[88] , dpath_mulcore_array2_s2[87] ,
         dpath_mulcore_array2_s2[86] , dpath_mulcore_array2_s2[85] ,
         dpath_mulcore_array2_s2[84] , dpath_mulcore_array2_s2[83] ,
         dpath_mulcore_array2_s2[82] , dpath_mulcore_array2_s2[81] ,
         dpath_mulcore_array2_s2[80] , dpath_mulcore_array2_s2[79] ,
         dpath_mulcore_array2_s2[78] , dpath_mulcore_array2_s2[77] ,
         dpath_mulcore_array2_s2[76] , dpath_mulcore_array2_s2[75] ,
         dpath_mulcore_array2_s2[74] , dpath_mulcore_array2_s2[73] ,
         dpath_mulcore_array2_s2[72] , dpath_mulcore_array2_s2[71] ,
         dpath_mulcore_array2_s2[70] , dpath_mulcore_array2_s2[69] ,
         dpath_mulcore_array2_s2[68] , dpath_mulcore_array2_s2[67] ,
         dpath_mulcore_array2_s2[66] , dpath_mulcore_array2_s2[65] ,
         dpath_mulcore_array2_s2[64] , dpath_mulcore_array2_s2[63] ,
         dpath_mulcore_array2_s2[62] , dpath_mulcore_array2_s2[61] ,
         dpath_mulcore_array2_s2[60] , dpath_mulcore_array2_s2[59] ,
         dpath_mulcore_array2_s2[58] , dpath_mulcore_array2_s2[57] ,
         dpath_mulcore_array2_s2[56] , dpath_mulcore_array2_s2[55] ,
         dpath_mulcore_array2_s2[54] , dpath_mulcore_array2_s2[53] ,
         dpath_mulcore_array2_s2[52] , dpath_mulcore_array2_s2[51] ,
         dpath_mulcore_array2_s2[50] , dpath_mulcore_array2_s2[49] ,
         dpath_mulcore_array2_s2[48] , dpath_mulcore_array2_s2[47] ,
         dpath_mulcore_array2_s2[46] , dpath_mulcore_array2_s2[45] ,
         dpath_mulcore_array2_s2[44] , dpath_mulcore_array2_s2[43] ,
         dpath_mulcore_array2_s2[42] , dpath_mulcore_array2_s2[41] ,
         dpath_mulcore_array2_s2[40] , dpath_mulcore_array2_s2[39] ,
         dpath_mulcore_array2_s2[38] , dpath_mulcore_array2_s2[37] ,
         dpath_mulcore_array2_s2[36] , dpath_mulcore_array2_s2[35] ,
         dpath_mulcore_array2_s2[34] , dpath_mulcore_array2_s2[33] ,
         dpath_mulcore_array2_s2[32] , dpath_mulcore_array2_s2[31] ,
         dpath_mulcore_array2_s2[30] , dpath_mulcore_array2_s2[29] ,
         dpath_mulcore_array2_s2[28] , dpath_mulcore_array2_s2[27] ,
         dpath_mulcore_array2_s2[26] , dpath_mulcore_array2_s2[25] ,
         dpath_mulcore_array2_s2[24] , dpath_mulcore_array2_s2[23] ,
         dpath_mulcore_array2_s2[22] , dpath_mulcore_array2_s2[21] ,
         dpath_mulcore_array2_s2[20] , dpath_mulcore_array2_s2[19] ,
         dpath_mulcore_array2_s2[18] , dpath_mulcore_array2_s2[17] ,
         dpath_mulcore_array2_s2[16] , dpath_mulcore_array2_s2[15] ,
         dpath_mulcore_array2_s2[14] , dpath_mulcore_array2_s2[13] ,
         dpath_mulcore_array2_s2[12] , dpath_mulcore_array2_s2[11] ,
         dpath_mulcore_array2_s2[10] , dpath_mulcore_array2_s2[9] ,
         dpath_mulcore_array2_s2[8] , dpath_mulcore_array2_s2[7] ,
         dpath_mulcore_array2_s2[6] , dpath_mulcore_array2_s2[5] ,
         dpath_mulcore_array2_s2[4] , dpath_mulcore_array2_s2[3] ,
         dpath_mulcore_array2_s2[2] , dpath_mulcore_array2_s2[1] ,
         dpath_mulcore_array2_s2[0] , dpath_mulcore_array2_c2[96] ,
         dpath_mulcore_array2_c2[95] , dpath_mulcore_array2_c2[94] ,
         dpath_mulcore_array2_c2[93] , dpath_mulcore_array2_c2[92] ,
         dpath_mulcore_array2_c2[91] , dpath_mulcore_array2_c2[90] ,
         dpath_mulcore_array2_c2[89] , dpath_mulcore_array2_c2[88] ,
         dpath_mulcore_array2_c2[87] , dpath_mulcore_array2_c2[86] ,
         dpath_mulcore_array2_c2[85] , dpath_mulcore_array2_c2[84] ,
         dpath_mulcore_array2_c2[83] , dpath_mulcore_array2_c2[82] ,
         dpath_mulcore_array2_c2[81] , dpath_mulcore_array2_c2[80] ,
         dpath_mulcore_array2_c2[79] , dpath_mulcore_array2_c2[78] ,
         dpath_mulcore_array2_c2[77] , dpath_mulcore_array2_c2[76] ,
         dpath_mulcore_array2_c2[75] , dpath_mulcore_array2_c2[74] ,
         dpath_mulcore_array2_c2[73] , dpath_mulcore_array2_c2[72] ,
         dpath_mulcore_array2_c2[71] , dpath_mulcore_array2_c2[70] ,
         dpath_mulcore_array2_c2[69] , dpath_mulcore_array2_c2[68] ,
         dpath_mulcore_array2_c2[67] , dpath_mulcore_array2_c2[66] ,
         dpath_mulcore_array2_c2[65] , dpath_mulcore_array2_c2[64] ,
         dpath_mulcore_array2_c2[63] , dpath_mulcore_array2_c2[62] ,
         dpath_mulcore_array2_c2[61] , dpath_mulcore_array2_c2[60] ,
         dpath_mulcore_array2_c2[59] , dpath_mulcore_array2_c2[58] ,
         dpath_mulcore_array2_c2[57] , dpath_mulcore_array2_c2[56] ,
         dpath_mulcore_array2_c2[55] , dpath_mulcore_array2_c2[54] ,
         dpath_mulcore_array2_c2[53] , dpath_mulcore_array2_c2[52] ,
         dpath_mulcore_array2_c2[51] , dpath_mulcore_array2_c2[50] ,
         dpath_mulcore_array2_c2[49] , dpath_mulcore_array2_c2[48] ,
         dpath_mulcore_array2_c2[47] , dpath_mulcore_array2_c2[46] ,
         dpath_mulcore_array2_c2[45] , dpath_mulcore_array2_c2[44] ,
         dpath_mulcore_array2_c2[43] , dpath_mulcore_array2_c2[42] ,
         dpath_mulcore_array2_c2[41] , dpath_mulcore_array2_c2[40] ,
         dpath_mulcore_array2_c2[39] , dpath_mulcore_array2_c2[38] ,
         dpath_mulcore_array2_c2[37] , dpath_mulcore_array2_c2[36] ,
         dpath_mulcore_array2_c2[35] , dpath_mulcore_array2_c2[34] ,
         dpath_mulcore_array2_c2[33] , dpath_mulcore_array2_c2[32] ,
         dpath_mulcore_array2_c2[31] , dpath_mulcore_array2_c2[30] ,
         dpath_mulcore_array2_c2[29] , dpath_mulcore_array2_c2[28] ,
         dpath_mulcore_array2_c2[27] , dpath_mulcore_array2_c2[26] ,
         dpath_mulcore_array2_c2[25] , dpath_mulcore_array2_c2[24] ,
         dpath_mulcore_array2_c2[23] , dpath_mulcore_array2_c2[22] ,
         dpath_mulcore_array2_c2[21] , dpath_mulcore_array2_c2[19] ,
         dpath_mulcore_array2_c2[18] , dpath_mulcore_array2_c2[17] ,
         dpath_mulcore_array2_c2[16] , dpath_mulcore_array2_c2[15] ,
         dpath_mulcore_array2_c2[14] , dpath_mulcore_array2_c2[13] ,
         dpath_mulcore_array2_c2[12] , dpath_mulcore_array2_c2[11] ,
         dpath_mulcore_array2_c2[10] , dpath_mulcore_array2_c2[9] ,
         dpath_mulcore_array2_c2[8] , dpath_mulcore_array2_c2[7] ,
         dpath_mulcore_array2_c2[6] , dpath_mulcore_array2_c2[5] ,
         dpath_mulcore_array2_c2[4] , dpath_mulcore_array2_c2[3] ,
         dpath_mulcore_array2_c2[2] , dpath_mulcore_array2_c2[1] ,
         dpath_mulcore_array2_c2[0] , dpath_mulcore_array2_c3[81] ,
         dpath_mulcore_array2_c3[80] , dpath_mulcore_array2_c3[79] ,
         dpath_mulcore_array2_c3[78] , dpath_mulcore_array2_c3[77] ,
         dpath_mulcore_array2_c3[76] , dpath_mulcore_array2_c3[75] ,
         dpath_mulcore_array2_c3[74] , dpath_mulcore_array2_c3[73] ,
         dpath_mulcore_array2_c3[72] , dpath_mulcore_array2_c3[71] ,
         dpath_mulcore_array2_c3[70] , dpath_mulcore_array2_c3[69] ,
         dpath_mulcore_array2_c3[68] , dpath_mulcore_array2_c3[67] ,
         dpath_mulcore_array2_c3[66] , dpath_mulcore_array2_c3[65] ,
         dpath_mulcore_array2_c3[64] , dpath_mulcore_array2_c3[63] ,
         dpath_mulcore_array2_c3[62] , dpath_mulcore_array2_c3[61] ,
         dpath_mulcore_array2_c3[60] , dpath_mulcore_array2_c3[59] ,
         dpath_mulcore_array2_c3[58] , dpath_mulcore_array2_c3[57] ,
         dpath_mulcore_array2_c3[56] , dpath_mulcore_array2_c3[55] ,
         dpath_mulcore_array2_c3[54] , dpath_mulcore_array2_c3[53] ,
         dpath_mulcore_array2_c3[52] , dpath_mulcore_array2_c3[51] ,
         dpath_mulcore_array2_c3[50] , dpath_mulcore_array2_c3[49] ,
         dpath_mulcore_array2_c3[48] , dpath_mulcore_array2_c3[47] ,
         dpath_mulcore_array2_c3[46] , dpath_mulcore_array2_c3[45] ,
         dpath_mulcore_array2_c3[44] , dpath_mulcore_array2_c3[43] ,
         dpath_mulcore_array2_c3[42] , dpath_mulcore_array2_c3[41] ,
         dpath_mulcore_array2_c3[40] , dpath_mulcore_array2_c3[39] ,
         dpath_mulcore_array2_c3[38] , dpath_mulcore_array2_c3[37] ,
         dpath_mulcore_array2_c3[36] , dpath_mulcore_array2_c3[35] ,
         dpath_mulcore_array2_c3[34] , dpath_mulcore_array2_c3[33] ,
         dpath_mulcore_array2_c3[32] , dpath_mulcore_array2_c3[31] ,
         dpath_mulcore_array2_c3[30] , dpath_mulcore_array2_c3[29] ,
         dpath_mulcore_array2_c3[28] , dpath_mulcore_array2_c3[27] ,
         dpath_mulcore_array2_c3[26] , dpath_mulcore_array2_c3[25] ,
         dpath_mulcore_array2_c3[24] , dpath_mulcore_array2_c3[23] ,
         dpath_mulcore_array2_c3[22] , dpath_mulcore_array2_c3[21] ,
         dpath_mulcore_array2_c3[19] , dpath_mulcore_array2_c3[18] ,
         dpath_mulcore_array2_c3[17] , dpath_mulcore_array2_c3[16] ,
         dpath_mulcore_array2_c3[15] , dpath_mulcore_array2_co[66] ,
         dpath_mulcore_array2_co[65] , dpath_mulcore_array2_co[64] ,
         dpath_mulcore_array2_co[63] , dpath_mulcore_array2_co[62] ,
         dpath_mulcore_array2_co[61] , dpath_mulcore_array2_co[60] ,
         dpath_mulcore_array2_co[59] , dpath_mulcore_array2_co[58] ,
         dpath_mulcore_array2_co[57] , dpath_mulcore_array2_co[56] ,
         dpath_mulcore_array2_co[55] , dpath_mulcore_array2_co[54] ,
         dpath_mulcore_array2_co[53] , dpath_mulcore_array2_co[52] ,
         dpath_mulcore_array2_co[51] , dpath_mulcore_array2_co[50] ,
         dpath_mulcore_array2_co[49] , dpath_mulcore_array2_co[48] ,
         dpath_mulcore_array2_co[47] , dpath_mulcore_array2_co[46] ,
         dpath_mulcore_array2_co[45] , dpath_mulcore_array2_co[44] ,
         dpath_mulcore_array2_co[43] , dpath_mulcore_array2_co[42] ,
         dpath_mulcore_array2_co[41] , dpath_mulcore_array2_co[40] ,
         dpath_mulcore_array2_co[39] , dpath_mulcore_array2_co[38] ,
         dpath_mulcore_array2_co[37] , dpath_mulcore_array2_co[36] ,
         dpath_mulcore_array2_co[35] , dpath_mulcore_array2_co[34] ,
         dpath_mulcore_array2_co[33] , dpath_mulcore_array2_co[32] ,
         dpath_mulcore_array2_co[31] , dpath_mulcore_array2_co[30] ,
         dpath_mulcore_array2_co[29] , dpath_mulcore_array2_co[28] ,
         dpath_mulcore_array2_co[27] , dpath_mulcore_array2_co[26] ,
         dpath_mulcore_array2_co[25] , dpath_mulcore_array2_co[24] ,
         dpath_mulcore_array2_co[23] , dpath_mulcore_array2_co[22] ,
         dpath_mulcore_array2_co[21] , dpath_mulcore_array2_co[20] ,
         dpath_mulcore_array2_ain[95] , dpath_mulcore_array2_ain[94] ,
         dpath_mulcore_array2_ain[93] , dpath_mulcore_array2_ain[92] ,
         dpath_mulcore_array2_ain[91] , dpath_mulcore_array2_ain[90] ,
         dpath_mulcore_array2_ain[89] , dpath_mulcore_array2_ain[88] ,
         dpath_mulcore_array2_ain[87] , dpath_mulcore_array2_ain[86] ,
         dpath_mulcore_array2_ain[85] , dpath_mulcore_array2_ain[84] ,
         dpath_mulcore_array2_ain[83] , dpath_mulcore_array2_ain[82] ,
         dpath_mulcore_array2_ain[81] , dpath_mulcore_array2_ain[80] ,
         dpath_mulcore_array2_ain[79] , dpath_mulcore_array2_ain[78] ,
         dpath_mulcore_array2_ain[77] , dpath_mulcore_array2_ain[76] ,
         dpath_mulcore_array2_ain[75] , dpath_mulcore_array2_ain[74] ,
         dpath_mulcore_array2_ain[73] , dpath_mulcore_array2_ain[72] ,
         dpath_mulcore_array2_ain[71] , dpath_mulcore_array2_ain[70] ,
         dpath_mulcore_array2_ain[69] , dpath_mulcore_array2_ain[68] ,
         dpath_mulcore_array2_ain[67] , dpath_mulcore_array2_ain[66] ,
         dpath_mulcore_array2_ain[65] , dpath_mulcore_array2_ain[64] ,
         dpath_mulcore_array2_ain[63] , dpath_mulcore_array2_ain[62] ,
         dpath_mulcore_array2_ain[61] , dpath_mulcore_array2_ain[60] ,
         dpath_mulcore_array2_ain[59] , dpath_mulcore_array2_ain[58] ,
         dpath_mulcore_array2_ain[57] , dpath_mulcore_array2_ain[56] ,
         dpath_mulcore_array2_ain[55] , dpath_mulcore_array2_ain[54] ,
         dpath_mulcore_array2_ain[53] , dpath_mulcore_array2_ain[52] ,
         dpath_mulcore_array2_ain[51] , dpath_mulcore_array2_ain[50] ,
         dpath_mulcore_array2_ain[49] , dpath_mulcore_array2_ain[48] ,
         dpath_mulcore_array2_ain[47] , dpath_mulcore_array2_ain[46] ,
         dpath_mulcore_array2_ain[45] , dpath_mulcore_array2_ain[44] ,
         dpath_mulcore_array2_ain[43] , dpath_mulcore_array2_ain[42] ,
         dpath_mulcore_array2_ain[41] , dpath_mulcore_array2_ain[40] ,
         dpath_mulcore_array2_ain[39] , dpath_mulcore_array2_ain[38] ,
         dpath_mulcore_array2_ain[37] , dpath_mulcore_array2_ain[36] ,
         dpath_mulcore_array2_ain[35] , dpath_mulcore_array2_ain[34] ,
         dpath_mulcore_array2_ain[33] , dpath_mulcore_array2_ain[32] ,
         dpath_mulcore_array2_ain[31] , dpath_mulcore_array2_ain[30] ,
         dpath_mulcore_array2_ain[29] , dpath_mulcore_array2_ain[28] ,
         dpath_mulcore_array2_ain[27] , dpath_mulcore_array2_ain[26] ,
         dpath_mulcore_array2_ain[25] , dpath_mulcore_array2_ain[24] ,
         dpath_mulcore_array2_ain[23] , dpath_mulcore_array2_ain[22] ,
         dpath_mulcore_array2_ain[21] , dpath_mulcore_array2_ain[20] ,
         dpath_mulcore_array2_ain[19] , dpath_mulcore_array2_ain[18] ,
         dpath_mulcore_array2_ain[17] , dpath_mulcore_array2_ain[16] ,
         dpath_mulcore_array2_ain[15] , dpath_mulcore_array2_ain[14] ,
         dpath_mulcore_array2_ain[13] , dpath_mulcore_array2_ain[12] ,
         dpath_mulcore_array2_ain[11] , dpath_mulcore_array2_ain[10] ,
         dpath_mulcore_array2_ain[9] , dpath_mulcore_array2_ain[8] ,
         dpath_mulcore_array2_ain[7] , dpath_mulcore_array2_ain[6] ,
         dpath_mulcore_array2_ain[5] , dpath_mulcore_array2_ain[4] ,
         dpath_mulcore_array2_ain[3] , dpath_mulcore_array2_ain[2] ,
         dpath_mulcore_array2_ain[1] , dpath_mulcore_array2_ain[0] ,
         dpath_mulcore_ary2_cmux_n195 , dpath_mulcore_ary2_cmux_n194 ,
         dpath_mulcore_ary2_cmux_n193 , dpath_mulcore_ary2_cmux_n192 ,
         dpath_mulcore_ary2_cmux_n191 , dpath_mulcore_ary2_cmux_n190 ,
         dpath_mulcore_ary2_cmux_n189 , dpath_mulcore_ary2_cmux_n188 ,
         dpath_mulcore_ary2_cmux_n187 , dpath_mulcore_ary2_cmux_n186 ,
         dpath_mulcore_ary2_cmux_n185 , dpath_mulcore_ary2_cmux_n184 ,
         dpath_mulcore_ary2_cmux_n183 , dpath_mulcore_ary2_cmux_n182 ,
         dpath_mulcore_ary2_cmux_n181 , dpath_mulcore_ary2_cmux_n180 ,
         dpath_mulcore_ary2_cmux_n179 , dpath_mulcore_ary2_cmux_n178 ,
         dpath_mulcore_ary2_cmux_n177 , dpath_mulcore_ary2_cmux_n176 ,
         dpath_mulcore_ary2_cmux_n175 , dpath_mulcore_ary2_cmux_n174 ,
         dpath_mulcore_ary2_cmux_n173 , dpath_mulcore_ary2_cmux_n172 ,
         dpath_mulcore_ary2_cmux_n171 , dpath_mulcore_ary2_cmux_n170 ,
         dpath_mulcore_ary2_cmux_n169 , dpath_mulcore_ary2_cmux_n168 ,
         dpath_mulcore_ary2_cmux_n167 , dpath_mulcore_ary2_cmux_n166 ,
         dpath_mulcore_ary2_cmux_n165 , dpath_mulcore_ary2_cmux_n164 ,
         dpath_mulcore_ary2_cmux_n163 , dpath_mulcore_ary2_cmux_n162 ,
         dpath_mulcore_ary2_cmux_n161 , dpath_mulcore_ary2_cmux_n160 ,
         dpath_mulcore_ary2_cmux_n159 , dpath_mulcore_ary2_cmux_n158 ,
         dpath_mulcore_ary2_cmux_n157 , dpath_mulcore_ary2_cmux_n156 ,
         dpath_mulcore_ary2_cmux_n155 , dpath_mulcore_ary2_cmux_n154 ,
         dpath_mulcore_ary2_cmux_n153 , dpath_mulcore_ary2_cmux_n152 ,
         dpath_mulcore_ary2_cmux_n151 , dpath_mulcore_ary2_cmux_n150 ,
         dpath_mulcore_ary2_cmux_n149 , dpath_mulcore_ary2_cmux_n148 ,
         dpath_mulcore_ary2_cmux_n147 , dpath_mulcore_ary2_cmux_n146 ,
         dpath_mulcore_ary2_cmux_n145 , dpath_mulcore_ary2_cmux_n144 ,
         dpath_mulcore_ary2_cmux_n143 , dpath_mulcore_ary2_cmux_n142 ,
         dpath_mulcore_ary2_cmux_n141 , dpath_mulcore_ary2_cmux_n140 ,
         dpath_mulcore_ary2_cmux_n139 , dpath_mulcore_ary2_cmux_n138 ,
         dpath_mulcore_ary2_cmux_n137 , dpath_mulcore_ary2_cmux_n136 ,
         dpath_mulcore_ary2_cmux_n135 , dpath_mulcore_ary2_cmux_n134 ,
         dpath_mulcore_ary2_cmux_n133 , dpath_mulcore_ary2_cmux_n132 ,
         dpath_mulcore_ary2_cmux_n131 , dpath_mulcore_ary2_cmux_n130 ,
         dpath_mulcore_ary2_cmux_n129 , dpath_mulcore_ary2_cmux_n128 ,
         dpath_mulcore_ary2_cmux_n127 , dpath_mulcore_ary2_cmux_n126 ,
         dpath_mulcore_ary2_cmux_n125 , dpath_mulcore_ary2_cmux_n124 ,
         dpath_mulcore_ary2_cmux_n123 , dpath_mulcore_ary2_cmux_n122 ,
         dpath_mulcore_ary2_cmux_n121 , dpath_mulcore_ary2_cmux_n120 ,
         dpath_mulcore_ary2_cmux_n119 , dpath_mulcore_ary2_cmux_n118 ,
         dpath_mulcore_ary2_cmux_n117 , dpath_mulcore_ary2_cmux_n116 ,
         dpath_mulcore_ary2_cmux_n115 , dpath_mulcore_ary2_cmux_n114 ,
         dpath_mulcore_ary2_cmux_n113 , dpath_mulcore_ary2_cmux_n112 ,
         dpath_mulcore_ary2_cmux_n111 , dpath_mulcore_ary2_cmux_n110 ,
         dpath_mulcore_ary2_cmux_n109 , dpath_mulcore_ary2_cmux_n108 ,
         dpath_mulcore_ary2_cmux_n107 , dpath_mulcore_ary2_cmux_n106 ,
         dpath_mulcore_ary2_cmux_n105 , dpath_mulcore_ary2_cmux_n104 ,
         dpath_mulcore_ary2_cmux_n103 , dpath_mulcore_ary2_cmux_n102 ,
         dpath_mulcore_ary2_cmux_n101 , dpath_mulcore_ary2_cmux_n100 ,
         dpath_mulcore_ary2_cmux_n99 , dpath_mulcore_ary2_cmux_n98 ,
         dpath_mulcore_ary2_cmux_n97 , dpath_mulcore_ary2_cmux_n96 ,
         dpath_mulcore_ary2_cmux_n95 , dpath_mulcore_ary2_cmux_n94 ,
         dpath_mulcore_ary2_cmux_n93 , dpath_mulcore_ary2_cmux_n92 ,
         dpath_mulcore_ary2_cmux_n91 , dpath_mulcore_ary2_cmux_n90 ,
         dpath_mulcore_ary2_cmux_n89 , dpath_mulcore_ary2_cmux_n88 ,
         dpath_mulcore_ary2_cmux_n87 , dpath_mulcore_ary2_cmux_n86 ,
         dpath_mulcore_ary2_cmux_n85 , dpath_mulcore_ary2_cmux_n84 ,
         dpath_mulcore_ary2_cmux_n83 , dpath_mulcore_ary2_cmux_n82 ,
         dpath_mulcore_ary2_cmux_n81 , dpath_mulcore_ary2_cmux_n80 ,
         dpath_mulcore_ary2_cmux_n79 , dpath_mulcore_ary2_cmux_n78 ,
         dpath_mulcore_ary2_cmux_n77 , dpath_mulcore_ary2_cmux_n76 ,
         dpath_mulcore_ary2_cmux_n75 , dpath_mulcore_ary2_cmux_n74 ,
         dpath_mulcore_ary2_cmux_n73 , dpath_mulcore_ary2_cmux_n72 ,
         dpath_mulcore_ary2_cmux_n71 , dpath_mulcore_ary2_cmux_n70 ,
         dpath_mulcore_ary2_cmux_n69 , dpath_mulcore_ary2_cmux_n68 ,
         dpath_mulcore_ary2_cmux_n67 , dpath_mulcore_ary2_cmux_n66 ,
         dpath_mulcore_ary2_cmux_n65 , dpath_mulcore_ary2_cmux_n64 ,
         dpath_mulcore_ary2_cmux_n63 , dpath_mulcore_ary2_cmux_n62 ,
         dpath_mulcore_ary2_cmux_n61 , dpath_mulcore_ary2_cmux_n60 ,
         dpath_mulcore_ary2_cmux_n59 , dpath_mulcore_ary2_cmux_n58 ,
         dpath_mulcore_ary2_cmux_n57 , dpath_mulcore_ary2_cmux_n56 ,
         dpath_mulcore_ary2_cmux_n55 , dpath_mulcore_ary2_cmux_n54 ,
         dpath_mulcore_ary2_cmux_n53 , dpath_mulcore_ary2_cmux_n52 ,
         dpath_mulcore_ary2_cmux_n51 , dpath_mulcore_ary2_cmux_n50 ,
         dpath_mulcore_ary2_cmux_n49 , dpath_mulcore_ary2_cmux_n48 ,
         dpath_mulcore_ary2_cmux_n47 , dpath_mulcore_ary2_cmux_n46 ,
         dpath_mulcore_ary2_cmux_n45 , dpath_mulcore_ary2_cmux_n44 ,
         dpath_mulcore_ary2_cmux_n43 , dpath_mulcore_ary2_cmux_n42 ,
         dpath_mulcore_ary2_cmux_n41 , dpath_mulcore_ary2_cmux_n40 ,
         dpath_mulcore_ary2_cmux_n39 , dpath_mulcore_ary2_cmux_n38 ,
         dpath_mulcore_ary2_cmux_n37 , dpath_mulcore_ary2_cmux_n36 ,
         dpath_mulcore_ary2_cmux_n35 , dpath_mulcore_ary2_cmux_n34 ,
         dpath_mulcore_ary2_cmux_n33 , dpath_mulcore_ary2_cmux_n32 ,
         dpath_mulcore_ary2_cmux_n31 , dpath_mulcore_ary2_cmux_n30 ,
         dpath_mulcore_ary2_cmux_n29 , dpath_mulcore_ary2_cmux_n28 ,
         dpath_mulcore_ary2_cmux_n27 , dpath_mulcore_ary2_cmux_n26 ,
         dpath_mulcore_ary2_cmux_n25 , dpath_mulcore_ary2_cmux_n24 ,
         dpath_mulcore_ary2_cmux_n23 , dpath_mulcore_ary2_cmux_n22 ,
         dpath_mulcore_ary2_cmux_n21 , dpath_mulcore_ary2_cmux_n20 ,
         dpath_mulcore_ary2_cmux_n19 , dpath_mulcore_ary2_cmux_n18 ,
         dpath_mulcore_ary2_cmux_n17 , dpath_mulcore_ary2_cmux_n16 ,
         dpath_mulcore_ary2_cmux_n15 , dpath_mulcore_ary2_cmux_n14 ,
         dpath_mulcore_ary2_cmux_n13 , dpath_mulcore_ary2_cmux_n12 ,
         dpath_mulcore_ary2_cmux_n11 , dpath_mulcore_ary2_cmux_n10 ,
         dpath_mulcore_ary2_cmux_n9 , dpath_mulcore_ary2_cmux_n8 ,
         dpath_mulcore_ary2_cmux_n7 , dpath_mulcore_ary2_cmux_n6 ,
         dpath_mulcore_ary2_cmux_n5 , dpath_mulcore_ary2_cmux_n4 ,
         dpath_mulcore_ary2_cmux_n3 , dpath_mulcore_ary2_cmux_n2 ,
         dpath_mulcore_a2cot_dff_n195 , dpath_mulcore_a2cot_dff_n193 ,
         dpath_mulcore_a2cot_dff_n191 , dpath_mulcore_a2cot_dff_n189 ,
         dpath_mulcore_a2cot_dff_n187 , dpath_mulcore_a2cot_dff_n185 ,
         dpath_mulcore_a2cot_dff_n183 , dpath_mulcore_a2cot_dff_n181 ,
         dpath_mulcore_a2cot_dff_n179 , dpath_mulcore_a2cot_dff_n177 ,
         dpath_mulcore_a2cot_dff_n175 , dpath_mulcore_a2cot_dff_n173 ,
         dpath_mulcore_a2cot_dff_n171 , dpath_mulcore_a2cot_dff_n169 ,
         dpath_mulcore_a2cot_dff_n167 , dpath_mulcore_a2cot_dff_n165 ,
         dpath_mulcore_a2cot_dff_n163 , dpath_mulcore_a2cot_dff_n161 ,
         dpath_mulcore_a2cot_dff_n159 , dpath_mulcore_a2cot_dff_n157 ,
         dpath_mulcore_a2cot_dff_n155 , dpath_mulcore_a2cot_dff_n153 ,
         dpath_mulcore_a2cot_dff_n151 , dpath_mulcore_a2cot_dff_n149 ,
         dpath_mulcore_a2cot_dff_n147 , dpath_mulcore_a2cot_dff_n145 ,
         dpath_mulcore_a2cot_dff_n143 , dpath_mulcore_a2cot_dff_n141 ,
         dpath_mulcore_a2cot_dff_n139 , dpath_mulcore_a2cot_dff_n137 ,
         dpath_mulcore_a2cot_dff_n135 , dpath_mulcore_a2cot_dff_n133 ,
         dpath_mulcore_a2cot_dff_n131 , dpath_mulcore_a2cot_dff_n129 ,
         dpath_mulcore_a2cot_dff_n127 , dpath_mulcore_a2cot_dff_n125 ,
         dpath_mulcore_a2cot_dff_n123 , dpath_mulcore_a2cot_dff_n121 ,
         dpath_mulcore_a2cot_dff_n119 , dpath_mulcore_a2cot_dff_n117 ,
         dpath_mulcore_a2cot_dff_n115 , dpath_mulcore_a2cot_dff_n113 ,
         dpath_mulcore_a2cot_dff_n111 , dpath_mulcore_a2cot_dff_n109 ,
         dpath_mulcore_a2cot_dff_n107 , dpath_mulcore_a2cot_dff_n105 ,
         dpath_mulcore_a2cot_dff_n103 , dpath_mulcore_a2cot_dff_n101 ,
         dpath_mulcore_a2cot_dff_n99 , dpath_mulcore_a2cot_dff_n97 ,
         dpath_mulcore_a2cot_dff_n95 , dpath_mulcore_a2cot_dff_n93 ,
         dpath_mulcore_a2cot_dff_n91 , dpath_mulcore_a2cot_dff_n89 ,
         dpath_mulcore_a2cot_dff_n87 , dpath_mulcore_a2cot_dff_n85 ,
         dpath_mulcore_a2cot_dff_n83 , dpath_mulcore_a2cot_dff_n81 ,
         dpath_mulcore_a2cot_dff_n79 , dpath_mulcore_a2cot_dff_n77 ,
         dpath_mulcore_a2cot_dff_n75 , dpath_mulcore_a2cot_dff_n73 ,
         dpath_mulcore_a2cot_dff_n71 , dpath_mulcore_a2cot_dff_n69 ,
         dpath_mulcore_a2cot_dff_n67 , dpath_mulcore_a2cot_dff_n65 ,
         dpath_mulcore_a2cot_dff_n63 , dpath_mulcore_a2cot_dff_n61 ,
         dpath_mulcore_a2cot_dff_n59 , dpath_mulcore_a2cot_dff_n57 ,
         dpath_mulcore_a2cot_dff_n55 , dpath_mulcore_a2cot_dff_n53 ,
         dpath_mulcore_a2cot_dff_n51 , dpath_mulcore_a2cot_dff_n49 ,
         dpath_mulcore_a2cot_dff_n47 , dpath_mulcore_a2cot_dff_n45 ,
         dpath_mulcore_a2cot_dff_n43 , dpath_mulcore_a2cot_dff_n41 ,
         dpath_mulcore_a2cot_dff_n39 , dpath_mulcore_a2cot_dff_n37 ,
         dpath_mulcore_a2cot_dff_n35 , dpath_mulcore_a2cot_dff_n33 ,
         dpath_mulcore_a2cot_dff_n31 , dpath_mulcore_a2cot_dff_n29 ,
         dpath_mulcore_a2cot_dff_n27 , dpath_mulcore_a2cot_dff_n25 ,
         dpath_mulcore_a2cot_dff_n23 , dpath_mulcore_a2cot_dff_n21 ,
         dpath_mulcore_a2cot_dff_n19 , dpath_mulcore_a2cot_dff_n17 ,
         dpath_mulcore_a2cot_dff_n15 , dpath_mulcore_a2cot_dff_n13 ,
         dpath_mulcore_a2cot_dff_n11 , dpath_mulcore_a2cot_dff_n9 ,
         dpath_mulcore_a2cot_dff_n7 , dpath_mulcore_a2cot_dff_n5 ,
         dpath_mulcore_a2cot_dff_n3 , dpath_mulcore_ary2_smux_n197 ,
         dpath_mulcore_ary2_smux_n196 , dpath_mulcore_ary2_smux_n195 ,
         dpath_mulcore_ary2_smux_n194 , dpath_mulcore_ary2_smux_n193 ,
         dpath_mulcore_ary2_smux_n192 , dpath_mulcore_ary2_smux_n191 ,
         dpath_mulcore_ary2_smux_n190 , dpath_mulcore_ary2_smux_n189 ,
         dpath_mulcore_ary2_smux_n188 , dpath_mulcore_ary2_smux_n187 ,
         dpath_mulcore_ary2_smux_n186 , dpath_mulcore_ary2_smux_n185 ,
         dpath_mulcore_ary2_smux_n184 , dpath_mulcore_ary2_smux_n183 ,
         dpath_mulcore_ary2_smux_n182 , dpath_mulcore_ary2_smux_n181 ,
         dpath_mulcore_ary2_smux_n180 , dpath_mulcore_ary2_smux_n179 ,
         dpath_mulcore_ary2_smux_n178 , dpath_mulcore_ary2_smux_n177 ,
         dpath_mulcore_ary2_smux_n176 , dpath_mulcore_ary2_smux_n175 ,
         dpath_mulcore_ary2_smux_n174 , dpath_mulcore_ary2_smux_n173 ,
         dpath_mulcore_ary2_smux_n172 , dpath_mulcore_ary2_smux_n171 ,
         dpath_mulcore_ary2_smux_n170 , dpath_mulcore_ary2_smux_n169 ,
         dpath_mulcore_ary2_smux_n168 , dpath_mulcore_ary2_smux_n167 ,
         dpath_mulcore_ary2_smux_n166 , dpath_mulcore_ary2_smux_n165 ,
         dpath_mulcore_ary2_smux_n164 , dpath_mulcore_ary2_smux_n163 ,
         dpath_mulcore_ary2_smux_n162 , dpath_mulcore_ary2_smux_n161 ,
         dpath_mulcore_ary2_smux_n160 , dpath_mulcore_ary2_smux_n159 ,
         dpath_mulcore_ary2_smux_n158 , dpath_mulcore_ary2_smux_n157 ,
         dpath_mulcore_ary2_smux_n156 , dpath_mulcore_ary2_smux_n155 ,
         dpath_mulcore_ary2_smux_n154 , dpath_mulcore_ary2_smux_n153 ,
         dpath_mulcore_ary2_smux_n152 , dpath_mulcore_ary2_smux_n151 ,
         dpath_mulcore_ary2_smux_n150 , dpath_mulcore_ary2_smux_n149 ,
         dpath_mulcore_ary2_smux_n148 , dpath_mulcore_ary2_smux_n147 ,
         dpath_mulcore_ary2_smux_n146 , dpath_mulcore_ary2_smux_n145 ,
         dpath_mulcore_ary2_smux_n144 , dpath_mulcore_ary2_smux_n143 ,
         dpath_mulcore_ary2_smux_n142 , dpath_mulcore_ary2_smux_n141 ,
         dpath_mulcore_ary2_smux_n140 , dpath_mulcore_ary2_smux_n139 ,
         dpath_mulcore_ary2_smux_n138 , dpath_mulcore_ary2_smux_n137 ,
         dpath_mulcore_ary2_smux_n136 , dpath_mulcore_ary2_smux_n135 ,
         dpath_mulcore_ary2_smux_n134 , dpath_mulcore_ary2_smux_n133 ,
         dpath_mulcore_ary2_smux_n132 , dpath_mulcore_ary2_smux_n131 ,
         dpath_mulcore_ary2_smux_n130 , dpath_mulcore_ary2_smux_n129 ,
         dpath_mulcore_ary2_smux_n128 , dpath_mulcore_ary2_smux_n127 ,
         dpath_mulcore_ary2_smux_n126 , dpath_mulcore_ary2_smux_n125 ,
         dpath_mulcore_ary2_smux_n124 , dpath_mulcore_ary2_smux_n123 ,
         dpath_mulcore_ary2_smux_n122 , dpath_mulcore_ary2_smux_n121 ,
         dpath_mulcore_ary2_smux_n120 , dpath_mulcore_ary2_smux_n119 ,
         dpath_mulcore_ary2_smux_n118 , dpath_mulcore_ary2_smux_n117 ,
         dpath_mulcore_ary2_smux_n116 , dpath_mulcore_ary2_smux_n115 ,
         dpath_mulcore_ary2_smux_n114 , dpath_mulcore_ary2_smux_n113 ,
         dpath_mulcore_ary2_smux_n112 , dpath_mulcore_ary2_smux_n111 ,
         dpath_mulcore_ary2_smux_n110 , dpath_mulcore_ary2_smux_n109 ,
         dpath_mulcore_ary2_smux_n108 , dpath_mulcore_ary2_smux_n107 ,
         dpath_mulcore_ary2_smux_n106 , dpath_mulcore_ary2_smux_n105 ,
         dpath_mulcore_ary2_smux_n104 , dpath_mulcore_ary2_smux_n103 ,
         dpath_mulcore_ary2_smux_n102 , dpath_mulcore_ary2_smux_n101 ,
         dpath_mulcore_ary2_smux_n100 , dpath_mulcore_ary2_smux_n99 ,
         dpath_mulcore_ary2_smux_n98 , dpath_mulcore_ary2_smux_n97 ,
         dpath_mulcore_ary2_smux_n96 , dpath_mulcore_ary2_smux_n95 ,
         dpath_mulcore_ary2_smux_n94 , dpath_mulcore_ary2_smux_n93 ,
         dpath_mulcore_ary2_smux_n92 , dpath_mulcore_ary2_smux_n91 ,
         dpath_mulcore_ary2_smux_n90 , dpath_mulcore_ary2_smux_n89 ,
         dpath_mulcore_ary2_smux_n88 , dpath_mulcore_ary2_smux_n87 ,
         dpath_mulcore_ary2_smux_n86 , dpath_mulcore_ary2_smux_n85 ,
         dpath_mulcore_ary2_smux_n84 , dpath_mulcore_ary2_smux_n83 ,
         dpath_mulcore_ary2_smux_n82 , dpath_mulcore_ary2_smux_n81 ,
         dpath_mulcore_ary2_smux_n80 , dpath_mulcore_ary2_smux_n79 ,
         dpath_mulcore_ary2_smux_n78 , dpath_mulcore_ary2_smux_n77 ,
         dpath_mulcore_ary2_smux_n76 , dpath_mulcore_ary2_smux_n75 ,
         dpath_mulcore_ary2_smux_n74 , dpath_mulcore_ary2_smux_n73 ,
         dpath_mulcore_ary2_smux_n72 , dpath_mulcore_ary2_smux_n71 ,
         dpath_mulcore_ary2_smux_n70 , dpath_mulcore_ary2_smux_n69 ,
         dpath_mulcore_ary2_smux_n68 , dpath_mulcore_ary2_smux_n67 ,
         dpath_mulcore_ary2_smux_n66 , dpath_mulcore_ary2_smux_n65 ,
         dpath_mulcore_ary2_smux_n64 , dpath_mulcore_ary2_smux_n63 ,
         dpath_mulcore_ary2_smux_n62 , dpath_mulcore_ary2_smux_n61 ,
         dpath_mulcore_ary2_smux_n60 , dpath_mulcore_ary2_smux_n59 ,
         dpath_mulcore_ary2_smux_n58 , dpath_mulcore_ary2_smux_n57 ,
         dpath_mulcore_ary2_smux_n56 , dpath_mulcore_ary2_smux_n55 ,
         dpath_mulcore_ary2_smux_n54 , dpath_mulcore_ary2_smux_n53 ,
         dpath_mulcore_ary2_smux_n52 , dpath_mulcore_ary2_smux_n51 ,
         dpath_mulcore_ary2_smux_n50 , dpath_mulcore_ary2_smux_n49 ,
         dpath_mulcore_ary2_smux_n48 , dpath_mulcore_ary2_smux_n47 ,
         dpath_mulcore_ary2_smux_n46 , dpath_mulcore_ary2_smux_n45 ,
         dpath_mulcore_ary2_smux_n44 , dpath_mulcore_ary2_smux_n43 ,
         dpath_mulcore_ary2_smux_n42 , dpath_mulcore_ary2_smux_n41 ,
         dpath_mulcore_ary2_smux_n40 , dpath_mulcore_ary2_smux_n39 ,
         dpath_mulcore_ary2_smux_n38 , dpath_mulcore_ary2_smux_n37 ,
         dpath_mulcore_ary2_smux_n36 , dpath_mulcore_ary2_smux_n35 ,
         dpath_mulcore_ary2_smux_n34 , dpath_mulcore_ary2_smux_n33 ,
         dpath_mulcore_ary2_smux_n32 , dpath_mulcore_ary2_smux_n31 ,
         dpath_mulcore_ary2_smux_n30 , dpath_mulcore_ary2_smux_n29 ,
         dpath_mulcore_ary2_smux_n28 , dpath_mulcore_ary2_smux_n27 ,
         dpath_mulcore_ary2_smux_n26 , dpath_mulcore_ary2_smux_n25 ,
         dpath_mulcore_ary2_smux_n24 , dpath_mulcore_ary2_smux_n23 ,
         dpath_mulcore_ary2_smux_n22 , dpath_mulcore_ary2_smux_n21 ,
         dpath_mulcore_ary2_smux_n20 , dpath_mulcore_ary2_smux_n19 ,
         dpath_mulcore_ary2_smux_n18 , dpath_mulcore_ary2_smux_n17 ,
         dpath_mulcore_ary2_smux_n16 , dpath_mulcore_ary2_smux_n15 ,
         dpath_mulcore_ary2_smux_n14 , dpath_mulcore_ary2_smux_n13 ,
         dpath_mulcore_ary2_smux_n12 , dpath_mulcore_ary2_smux_n11 ,
         dpath_mulcore_ary2_smux_n10 , dpath_mulcore_ary2_smux_n9 ,
         dpath_mulcore_ary2_smux_n8 , dpath_mulcore_ary2_smux_n7 ,
         dpath_mulcore_ary2_smux_n6 , dpath_mulcore_ary2_smux_n5 ,
         dpath_mulcore_ary2_smux_n4 , dpath_mulcore_ary2_smux_n3 ,
         dpath_mulcore_ary2_smux_n2 , dpath_mulcore_a2sum_dff_n197 ,
         dpath_mulcore_a2sum_dff_n195 , dpath_mulcore_a2sum_dff_n193 ,
         dpath_mulcore_a2sum_dff_n191 , dpath_mulcore_a2sum_dff_n189 ,
         dpath_mulcore_a2sum_dff_n187 , dpath_mulcore_a2sum_dff_n185 ,
         dpath_mulcore_a2sum_dff_n183 , dpath_mulcore_a2sum_dff_n181 ,
         dpath_mulcore_a2sum_dff_n179 , dpath_mulcore_a2sum_dff_n177 ,
         dpath_mulcore_a2sum_dff_n175 , dpath_mulcore_a2sum_dff_n173 ,
         dpath_mulcore_a2sum_dff_n171 , dpath_mulcore_a2sum_dff_n169 ,
         dpath_mulcore_a2sum_dff_n167 , dpath_mulcore_a2sum_dff_n165 ,
         dpath_mulcore_a2sum_dff_n163 , dpath_mulcore_a2sum_dff_n161 ,
         dpath_mulcore_a2sum_dff_n159 , dpath_mulcore_a2sum_dff_n157 ,
         dpath_mulcore_a2sum_dff_n155 , dpath_mulcore_a2sum_dff_n153 ,
         dpath_mulcore_a2sum_dff_n151 , dpath_mulcore_a2sum_dff_n149 ,
         dpath_mulcore_a2sum_dff_n147 , dpath_mulcore_a2sum_dff_n145 ,
         dpath_mulcore_a2sum_dff_n143 , dpath_mulcore_a2sum_dff_n141 ,
         dpath_mulcore_a2sum_dff_n139 , dpath_mulcore_a2sum_dff_n137 ,
         dpath_mulcore_a2sum_dff_n135 , dpath_mulcore_a2sum_dff_n133 ,
         dpath_mulcore_a2sum_dff_n131 , dpath_mulcore_a2sum_dff_n129 ,
         dpath_mulcore_a2sum_dff_n127 , dpath_mulcore_a2sum_dff_n125 ,
         dpath_mulcore_a2sum_dff_n123 , dpath_mulcore_a2sum_dff_n121 ,
         dpath_mulcore_a2sum_dff_n119 , dpath_mulcore_a2sum_dff_n117 ,
         dpath_mulcore_a2sum_dff_n115 , dpath_mulcore_a2sum_dff_n113 ,
         dpath_mulcore_a2sum_dff_n111 , dpath_mulcore_a2sum_dff_n109 ,
         dpath_mulcore_a2sum_dff_n107 , dpath_mulcore_a2sum_dff_n105 ,
         dpath_mulcore_a2sum_dff_n103 , dpath_mulcore_a2sum_dff_n101 ,
         dpath_mulcore_a2sum_dff_n99 , dpath_mulcore_a2sum_dff_n97 ,
         dpath_mulcore_a2sum_dff_n95 , dpath_mulcore_a2sum_dff_n93 ,
         dpath_mulcore_a2sum_dff_n91 , dpath_mulcore_a2sum_dff_n89 ,
         dpath_mulcore_a2sum_dff_n87 , dpath_mulcore_a2sum_dff_n85 ,
         dpath_mulcore_a2sum_dff_n83 , dpath_mulcore_a2sum_dff_n81 ,
         dpath_mulcore_a2sum_dff_n79 , dpath_mulcore_a2sum_dff_n77 ,
         dpath_mulcore_a2sum_dff_n75 , dpath_mulcore_a2sum_dff_n73 ,
         dpath_mulcore_a2sum_dff_n71 , dpath_mulcore_a2sum_dff_n69 ,
         dpath_mulcore_a2sum_dff_n67 , dpath_mulcore_a2sum_dff_n65 ,
         dpath_mulcore_a2sum_dff_n63 , dpath_mulcore_a2sum_dff_n61 ,
         dpath_mulcore_a2sum_dff_n59 , dpath_mulcore_a2sum_dff_n57 ,
         dpath_mulcore_a2sum_dff_n55 , dpath_mulcore_a2sum_dff_n53 ,
         dpath_mulcore_a2sum_dff_n51 , dpath_mulcore_a2sum_dff_n49 ,
         dpath_mulcore_a2sum_dff_n47 , dpath_mulcore_a2sum_dff_n45 ,
         dpath_mulcore_a2sum_dff_n43 , dpath_mulcore_a2sum_dff_n41 ,
         dpath_mulcore_a2sum_dff_n39 , dpath_mulcore_a2sum_dff_n37 ,
         dpath_mulcore_a2sum_dff_n35 , dpath_mulcore_a2sum_dff_n33 ,
         dpath_mulcore_a2sum_dff_n31 , dpath_mulcore_a2sum_dff_n29 ,
         dpath_mulcore_a2sum_dff_n27 , dpath_mulcore_a2sum_dff_n25 ,
         dpath_mulcore_a2sum_dff_n23 , dpath_mulcore_a2sum_dff_n21 ,
         dpath_mulcore_a2sum_dff_n19 , dpath_mulcore_a2sum_dff_n17 ,
         dpath_mulcore_a2sum_dff_n15 , dpath_mulcore_a2sum_dff_n13 ,
         dpath_mulcore_a2sum_dff_n11 , dpath_mulcore_a2sum_dff_n9 ,
         dpath_mulcore_a2sum_dff_n7 , dpath_mulcore_a2sum_dff_n5 ,
         dpath_mulcore_a2sum_dff_n3 , dpath_mulcore_psum_dff_n137 ,
         dpath_mulcore_psum_dff_n135 , dpath_mulcore_psum_dff_n133 ,
         dpath_mulcore_psum_dff_n131 , dpath_mulcore_psum_dff_n129 ,
         dpath_mulcore_psum_dff_n127 , dpath_mulcore_psum_dff_n125 ,
         dpath_mulcore_psum_dff_n123 , dpath_mulcore_psum_dff_n121 ,
         dpath_mulcore_psum_dff_n119 , dpath_mulcore_psum_dff_n117 ,
         dpath_mulcore_psum_dff_n115 , dpath_mulcore_psum_dff_n113 ,
         dpath_mulcore_psum_dff_n111 , dpath_mulcore_psum_dff_n109 ,
         dpath_mulcore_psum_dff_n107 , dpath_mulcore_psum_dff_n105 ,
         dpath_mulcore_psum_dff_n103 , dpath_mulcore_psum_dff_n101 ,
         dpath_mulcore_psum_dff_n99 , dpath_mulcore_psum_dff_n97 ,
         dpath_mulcore_psum_dff_n95 , dpath_mulcore_psum_dff_n93 ,
         dpath_mulcore_psum_dff_n91 , dpath_mulcore_psum_dff_n89 ,
         dpath_mulcore_psum_dff_n87 , dpath_mulcore_psum_dff_n85 ,
         dpath_mulcore_psum_dff_n83 , dpath_mulcore_psum_dff_n81 ,
         dpath_mulcore_psum_dff_n79 , dpath_mulcore_psum_dff_n77 ,
         dpath_mulcore_psum_dff_n75 , dpath_mulcore_psum_dff_n73 ,
         dpath_mulcore_psum_dff_n71 , dpath_mulcore_psum_dff_n69 ,
         dpath_mulcore_psum_dff_n67 , dpath_mulcore_psum_dff_n65 ,
         dpath_mulcore_psum_dff_n63 , dpath_mulcore_psum_dff_n61 ,
         dpath_mulcore_psum_dff_n59 , dpath_mulcore_psum_dff_n57 ,
         dpath_mulcore_psum_dff_n55 , dpath_mulcore_psum_dff_n53 ,
         dpath_mulcore_psum_dff_n51 , dpath_mulcore_psum_dff_n49 ,
         dpath_mulcore_psum_dff_n47 , dpath_mulcore_psum_dff_n45 ,
         dpath_mulcore_psum_dff_n43 , dpath_mulcore_psum_dff_n41 ,
         dpath_mulcore_psum_dff_n39 , dpath_mulcore_psum_dff_n37 ,
         dpath_mulcore_psum_dff_n35 , dpath_mulcore_psum_dff_n33 ,
         dpath_mulcore_psum_dff_n31 , dpath_mulcore_psum_dff_n29 ,
         dpath_mulcore_psum_dff_n27 , dpath_mulcore_psum_dff_n25 ,
         dpath_mulcore_psum_dff_n23 , dpath_mulcore_psum_dff_n21 ,
         dpath_mulcore_psum_dff_n19 , dpath_mulcore_psum_dff_n17 ,
         dpath_mulcore_psum_dff_n15 , dpath_mulcore_psum_dff_n13 ,
         dpath_mulcore_psum_dff_n11 , dpath_mulcore_psum_dff_n9 ,
         dpath_mulcore_psum_dff_n7 , dpath_mulcore_psum_dff_n5 ,
         dpath_mulcore_psum_dff_n3 , dpath_mulcore_pcout_dff_n139 ,
         dpath_mulcore_pcout_dff_n137 , dpath_mulcore_pcout_dff_n135 ,
         dpath_mulcore_pcout_dff_n133 , dpath_mulcore_pcout_dff_n131 ,
         dpath_mulcore_pcout_dff_n129 , dpath_mulcore_pcout_dff_n127 ,
         dpath_mulcore_pcout_dff_n125 , dpath_mulcore_pcout_dff_n123 ,
         dpath_mulcore_pcout_dff_n121 , dpath_mulcore_pcout_dff_n119 ,
         dpath_mulcore_pcout_dff_n117 , dpath_mulcore_pcout_dff_n115 ,
         dpath_mulcore_pcout_dff_n113 , dpath_mulcore_pcout_dff_n111 ,
         dpath_mulcore_pcout_dff_n109 , dpath_mulcore_pcout_dff_n107 ,
         dpath_mulcore_pcout_dff_n105 , dpath_mulcore_pcout_dff_n103 ,
         dpath_mulcore_pcout_dff_n101 , dpath_mulcore_pcout_dff_n99 ,
         dpath_mulcore_pcout_dff_n97 , dpath_mulcore_pcout_dff_n95 ,
         dpath_mulcore_pcout_dff_n93 , dpath_mulcore_pcout_dff_n91 ,
         dpath_mulcore_pcout_dff_n89 , dpath_mulcore_pcout_dff_n87 ,
         dpath_mulcore_pcout_dff_n85 , dpath_mulcore_pcout_dff_n83 ,
         dpath_mulcore_pcout_dff_n81 , dpath_mulcore_pcout_dff_n79 ,
         dpath_mulcore_pcout_dff_n77 , dpath_mulcore_pcout_dff_n75 ,
         dpath_mulcore_pcout_dff_n73 , dpath_mulcore_pcout_dff_n71 ,
         dpath_mulcore_pcout_dff_n69 , dpath_mulcore_pcout_dff_n67 ,
         dpath_mulcore_pcout_dff_n65 , dpath_mulcore_pcout_dff_n63 ,
         dpath_mulcore_pcout_dff_n61 , dpath_mulcore_pcout_dff_n59 ,
         dpath_mulcore_pcout_dff_n57 , dpath_mulcore_pcout_dff_n55 ,
         dpath_mulcore_pcout_dff_n53 , dpath_mulcore_pcout_dff_n51 ,
         dpath_mulcore_pcout_dff_n49 , dpath_mulcore_pcout_dff_n47 ,
         dpath_mulcore_pcout_dff_n45 , dpath_mulcore_pcout_dff_n43 ,
         dpath_mulcore_pcout_dff_n41 , dpath_mulcore_pcout_dff_n39 ,
         dpath_mulcore_pcout_dff_n37 , dpath_mulcore_pcout_dff_n35 ,
         dpath_mulcore_pcout_dff_n33 , dpath_mulcore_pcout_dff_n31 ,
         dpath_mulcore_pcout_dff_n29 , dpath_mulcore_pcout_dff_n27 ,
         dpath_mulcore_pcout_dff_n25 , dpath_mulcore_pcout_dff_n23 ,
         dpath_mulcore_pcout_dff_n21 , dpath_mulcore_pcout_dff_n19 ,
         dpath_mulcore_pcout_dff_n17 , dpath_mulcore_pcout_dff_n15 ,
         dpath_mulcore_pcout_dff_n13 , dpath_mulcore_pcout_dff_n11 ,
         dpath_mulcore_pcout_dff_n9 , dpath_mulcore_pcout_dff_n5 ,
         dpath_mulcore_pcout_dff_n3 , dpath_mulcore_out_dff_n209 ,
         dpath_mulcore_out_dff_n207 , dpath_mulcore_out_dff_n205 ,
         dpath_mulcore_out_dff_n203 , dpath_mulcore_out_dff_n201 ,
         dpath_mulcore_out_dff_n199 , dpath_mulcore_out_dff_n197 ,
         dpath_mulcore_out_dff_n195 , dpath_mulcore_out_dff_n193 ,
         dpath_mulcore_out_dff_n191 , dpath_mulcore_out_dff_n189 ,
         dpath_mulcore_out_dff_n187 , dpath_mulcore_out_dff_n185 ,
         dpath_mulcore_out_dff_n183 , dpath_mulcore_out_dff_n181 ,
         dpath_mulcore_out_dff_n179 , dpath_mulcore_out_dff_n177 ,
         dpath_mulcore_out_dff_n175 , dpath_mulcore_out_dff_n173 ,
         dpath_mulcore_out_dff_n171 , dpath_mulcore_out_dff_n169 ,
         dpath_mulcore_out_dff_n167 , dpath_mulcore_out_dff_n165 ,
         dpath_mulcore_out_dff_n163 , dpath_mulcore_out_dff_n161 ,
         dpath_mulcore_out_dff_n159 , dpath_mulcore_out_dff_n157 ,
         dpath_mulcore_out_dff_n155 , dpath_mulcore_out_dff_n153 ,
         dpath_mulcore_out_dff_n151 , dpath_mulcore_out_dff_n149 ,
         dpath_mulcore_out_dff_n147 , dpath_mulcore_out_dff_n145 ,
         dpath_mulcore_out_dff_n143 , dpath_mulcore_out_dff_n141 ,
         dpath_mulcore_out_dff_n139 , dpath_mulcore_out_dff_n137 ,
         dpath_mulcore_out_dff_n135 , dpath_mulcore_out_dff_n133 ,
         dpath_mulcore_out_dff_n131 , dpath_mulcore_out_dff_n129 ,
         dpath_mulcore_out_dff_n127 , dpath_mulcore_out_dff_n125 ,
         dpath_mulcore_out_dff_n123 , dpath_mulcore_out_dff_n121 ,
         dpath_mulcore_out_dff_n119 , dpath_mulcore_out_dff_n117 ,
         dpath_mulcore_out_dff_n115 , dpath_mulcore_out_dff_n113 ,
         dpath_mulcore_out_dff_n111 , dpath_mulcore_out_dff_n109 ,
         dpath_mulcore_out_dff_n107 , dpath_mulcore_out_dff_n105 ,
         dpath_mulcore_out_dff_n103 , dpath_mulcore_out_dff_n101 ,
         dpath_mulcore_out_dff_n99 , dpath_mulcore_out_dff_n97 ,
         dpath_mulcore_out_dff_n95 , dpath_mulcore_out_dff_n93 ,
         dpath_mulcore_out_dff_n91 , dpath_mulcore_out_dff_n89 ,
         dpath_mulcore_out_dff_n87 , dpath_mulcore_out_dff_n85 ,
         dpath_mulcore_out_dff_n83 , dpath_mulcore_out_dff_n81 ,
         dpath_mulcore_out_dff_n79 , dpath_mulcore_out_dff_n77 ,
         dpath_mulcore_out_dff_n75 , dpath_mulcore_out_dff_n73 ,
         dpath_mulcore_out_dff_n71 , dpath_mulcore_out_dff_n69 ,
         dpath_mulcore_out_dff_n67 , dpath_mulcore_out_dff_n65 ,
         dpath_mulcore_out_dff_n63 , dpath_mulcore_out_dff_n61 ,
         dpath_mulcore_out_dff_n59 , dpath_mulcore_out_dff_n57 ,
         dpath_mulcore_out_dff_n55 , dpath_mulcore_out_dff_n53 ,
         dpath_mulcore_out_dff_n51 , dpath_mulcore_out_dff_n49 ,
         dpath_mulcore_out_dff_n47 , dpath_mulcore_out_dff_n45 ,
         dpath_mulcore_out_dff_n43 , dpath_mulcore_out_dff_n41 ,
         dpath_mulcore_out_dff_n39 , dpath_mulcore_out_dff_n37 ,
         dpath_mulcore_out_dff_n35 , dpath_mulcore_out_dff_n33 ,
         dpath_mulcore_out_dff_n31 , dpath_mulcore_out_dff_n29 ,
         dpath_mulcore_out_dff_n27 , dpath_mulcore_out_dff_n25 ,
         dpath_mulcore_out_dff_n23 , dpath_mulcore_out_dff_n21 ,
         dpath_mulcore_out_dff_n19 , dpath_mulcore_out_dff_n17 ,
         dpath_mulcore_out_dff_n15 , dpath_mulcore_out_dff_n13 ,
         dpath_mulcore_out_dff_n11 , dpath_mulcore_out_dff_n9 ,
         dpath_mulcore_out_dff_n7 , dpath_mulcore_out_dff_n5 ,
         dpath_mulcore_out_dff_n3 , dpath_mulcore_pip_dff_n65 ,
         dpath_mulcore_pip_dff_n63 , dpath_mulcore_pip_dff_n61 ,
         dpath_mulcore_pip_dff_n59 , dpath_mulcore_pip_dff_n57 ,
         dpath_mulcore_pip_dff_n55 , dpath_mulcore_pip_dff_n53 ,
         dpath_mulcore_pip_dff_n51 , dpath_mulcore_pip_dff_n49 ,
         dpath_mulcore_pip_dff_n47 , dpath_mulcore_pip_dff_n45 ,
         dpath_mulcore_pip_dff_n43 , dpath_mulcore_pip_dff_n41 ,
         dpath_mulcore_pip_dff_n39 , dpath_mulcore_pip_dff_n37 ,
         dpath_mulcore_pip_dff_n35 , dpath_mulcore_pip_dff_n33 ,
         dpath_mulcore_pip_dff_n31 , dpath_mulcore_pip_dff_n29 ,
         dpath_mulcore_pip_dff_n27 , dpath_mulcore_pip_dff_n25 ,
         dpath_mulcore_pip_dff_n23 , dpath_mulcore_pip_dff_n21 ,
         dpath_mulcore_pip_dff_n19 , dpath_mulcore_pip_dff_n17 ,
         dpath_mulcore_pip_dff_n15 , dpath_mulcore_pip_dff_n13 ,
         dpath_mulcore_pip_dff_n11 , dpath_mulcore_pip_dff_n9 ,
         dpath_mulcore_pip_dff_n7 , dpath_mulcore_pip_dff_n5 ,
         dpath_mulcore_pip_dff_n3 , dpath_mulcore_booth_encode0_a_n75 ,
         dpath_mulcore_booth_encode0_a_n74 ,
         dpath_mulcore_booth_encode0_a_n73 ,
         dpath_mulcore_booth_encode0_a_n72 ,
         dpath_mulcore_booth_encode0_a_n71 ,
         dpath_mulcore_booth_encode0_a_n70 ,
         dpath_mulcore_booth_encode0_a_n69 ,
         dpath_mulcore_booth_encode0_a_n68 ,
         dpath_mulcore_booth_encode0_a_n67 ,
         dpath_mulcore_booth_encode0_a_n66 ,
         dpath_mulcore_booth_encode0_a_n65 ,
         dpath_mulcore_booth_encode0_a_n64 ,
         dpath_mulcore_booth_encode0_a_n63 ,
         dpath_mulcore_booth_encode0_a_n62 ,
         dpath_mulcore_booth_encode0_a_n61 ,
         dpath_mulcore_booth_encode0_a_n60 ,
         dpath_mulcore_booth_encode0_a_n59 ,
         dpath_mulcore_booth_encode0_a_n58 ,
         dpath_mulcore_booth_encode0_a_n57 ,
         dpath_mulcore_booth_encode0_a_n56 ,
         dpath_mulcore_booth_encode0_a_n55 ,
         dpath_mulcore_booth_encode0_a_n54 ,
         dpath_mulcore_booth_encode0_a_n53 ,
         dpath_mulcore_booth_encode0_a_n52 ,
         dpath_mulcore_booth_encode0_a_n51 ,
         dpath_mulcore_booth_encode0_a_n50 ,
         dpath_mulcore_booth_encode0_a_n49 ,
         dpath_mulcore_booth_encode0_a_n48 ,
         dpath_mulcore_booth_encode0_a_n47 ,
         dpath_mulcore_booth_encode0_a_n46 ,
         dpath_mulcore_booth_encode0_a_n45 ,
         dpath_mulcore_booth_encode0_a_n44 ,
         dpath_mulcore_booth_encode0_a_n43 ,
         dpath_mulcore_booth_encode0_a_n42 ,
         dpath_mulcore_booth_encode0_a_n41 ,
         dpath_mulcore_booth_encode0_a_n40 ,
         dpath_mulcore_booth_encode0_a_n39 ,
         dpath_mulcore_booth_encode0_a_n38 ,
         dpath_mulcore_booth_encode0_a_n37 ,
         dpath_mulcore_booth_encode0_a_n36 ,
         dpath_mulcore_booth_encode0_a_n35 ,
         dpath_mulcore_booth_encode0_a_n34 ,
         dpath_mulcore_booth_encode0_a_n33 ,
         dpath_mulcore_booth_encode0_a_n32 ,
         dpath_mulcore_booth_encode0_a_n31 ,
         dpath_mulcore_booth_encode0_a_n30 ,
         dpath_mulcore_booth_encode0_a_n29 ,
         dpath_mulcore_booth_encode0_a_n28 ,
         dpath_mulcore_booth_encode0_a_n27 ,
         dpath_mulcore_booth_encode0_a_n26 ,
         dpath_mulcore_booth_encode0_a_n25 ,
         dpath_mulcore_booth_encode0_a_n24 ,
         dpath_mulcore_booth_encode0_a_n23 ,
         dpath_mulcore_booth_encode0_a_n22 ,
         dpath_mulcore_booth_encode0_a_n21 ,
         dpath_mulcore_booth_encode0_a_n20 ,
         dpath_mulcore_booth_encode0_a_n19 ,
         dpath_mulcore_booth_encode0_a_n17 ,
         dpath_mulcore_booth_out_mux0_n7 , dpath_mulcore_booth_out_mux0_n6 ,
         dpath_mulcore_booth_out_mux0_n5 , dpath_mulcore_booth_out_mux0_n4 ,
         dpath_mulcore_booth_out_mux0_n3 , dpath_mulcore_booth_out_mux0_n2 ,
         dpath_mulcore_booth_out_mux16_n2 , dpath_mulcore_booth_out_dff0_n7 ,
         dpath_mulcore_booth_out_dff0_n5 , dpath_mulcore_booth_out_dff0_n3 ,
         dpath_mulcore_ary1_a0_p1n_n5 , dpath_mulcore_ary1_a0_p1n_n4 ,
         dpath_mulcore_ary1_a0_sc3_71__n8 ,
         dpath_mulcore_ary1_a0_sc3_71__n7 ,
         dpath_mulcore_ary1_a0_sc3_71__n6 ,
         dpath_mulcore_ary1_a0_sc3_71__n5 ,
         dpath_mulcore_ary1_a0_sc3_71__n4 ,
         dpath_mulcore_ary1_a0_sc3_71__n3 ,
         dpath_mulcore_ary1_a0_sc3_71__n2 , dpath_mulcore_ary1_a0_sc3_71__z ,
         dpath_mulcore_ary1_a0_sc2_2_70__n3 ,
         dpath_mulcore_ary1_a0_sc2_2_70__n2 ,
         dpath_mulcore_ary1_a0_sc2_2_70__n1 ,
         dpath_mulcore_ary1_a0_I2_p0_l[63] ,
         dpath_mulcore_ary1_a0_I2_p0_l[62] ,
         dpath_mulcore_ary1_a0_I2_p0_l[61] ,
         dpath_mulcore_ary1_a0_I2_p0_l[60] ,
         dpath_mulcore_ary1_a0_I2_p0_l[59] ,
         dpath_mulcore_ary1_a0_I2_p0_l[58] ,
         dpath_mulcore_ary1_a0_I2_p0_l[57] ,
         dpath_mulcore_ary1_a0_I2_p0_l[56] ,
         dpath_mulcore_ary1_a0_I2_p0_l[55] ,
         dpath_mulcore_ary1_a0_I2_p0_l[54] ,
         dpath_mulcore_ary1_a0_I2_p0_l[53] ,
         dpath_mulcore_ary1_a0_I2_p0_l[52] ,
         dpath_mulcore_ary1_a0_I2_p0_l[51] ,
         dpath_mulcore_ary1_a0_I2_p0_l[50] ,
         dpath_mulcore_ary1_a0_I2_p0_l[49] ,
         dpath_mulcore_ary1_a0_I2_p0_l[48] ,
         dpath_mulcore_ary1_a0_I2_p0_l[47] ,
         dpath_mulcore_ary1_a0_I2_p0_l[46] ,
         dpath_mulcore_ary1_a0_I2_p0_l[45] ,
         dpath_mulcore_ary1_a0_I2_p0_l[44] ,
         dpath_mulcore_ary1_a0_I2_p0_l[43] ,
         dpath_mulcore_ary1_a0_I2_p0_l[42] ,
         dpath_mulcore_ary1_a0_I2_p0_l[41] ,
         dpath_mulcore_ary1_a0_I2_p0_l[40] ,
         dpath_mulcore_ary1_a0_I2_p0_l[39] ,
         dpath_mulcore_ary1_a0_I2_p0_l[38] ,
         dpath_mulcore_ary1_a0_I2_p0_l[37] ,
         dpath_mulcore_ary1_a0_I2_p0_l[36] ,
         dpath_mulcore_ary1_a0_I2_p0_l[35] ,
         dpath_mulcore_ary1_a0_I2_p0_l[34] ,
         dpath_mulcore_ary1_a0_I2_p0_l[33] ,
         dpath_mulcore_ary1_a0_I2_p0_l[32] ,
         dpath_mulcore_ary1_a0_I2_p0_l[31] ,
         dpath_mulcore_ary1_a0_I2_p0_l[30] ,
         dpath_mulcore_ary1_a0_I2_p0_l[29] ,
         dpath_mulcore_ary1_a0_I2_p0_l[28] ,
         dpath_mulcore_ary1_a0_I2_p0_l[27] ,
         dpath_mulcore_ary1_a0_I2_p0_l[26] ,
         dpath_mulcore_ary1_a0_I2_p0_l[25] ,
         dpath_mulcore_ary1_a0_I2_p0_l[24] ,
         dpath_mulcore_ary1_a0_I2_p0_l[23] ,
         dpath_mulcore_ary1_a0_I2_p0_l[22] ,
         dpath_mulcore_ary1_a0_I2_p0_l[21] ,
         dpath_mulcore_ary1_a0_I2_p0_l[20] ,
         dpath_mulcore_ary1_a0_I2_p0_l[19] ,
         dpath_mulcore_ary1_a0_I2_p0_l[18] ,
         dpath_mulcore_ary1_a0_I2_p0_l[17] ,
         dpath_mulcore_ary1_a0_I2_p0_l[16] ,
         dpath_mulcore_ary1_a0_I2_p0_l[15] ,
         dpath_mulcore_ary1_a0_I2_p0_l[14] ,
         dpath_mulcore_ary1_a0_I2_p0_l[13] ,
         dpath_mulcore_ary1_a0_I2_p0_l[12] ,
         dpath_mulcore_ary1_a0_I2_p0_l[11] ,
         dpath_mulcore_ary1_a0_I2_p0_l[10] ,
         dpath_mulcore_ary1_a0_I2_p0_l[9] ,
         dpath_mulcore_ary1_a0_I2_p0_l[8] ,
         dpath_mulcore_ary1_a0_I2_p0_l[7] ,
         dpath_mulcore_ary1_a0_I2_p0_l[6] ,
         dpath_mulcore_ary1_a0_I2_p0_l[5] ,
         dpath_mulcore_ary1_a0_I2_p0_l[4] ,
         dpath_mulcore_ary1_a0_I2_p0_l[3] ,
         dpath_mulcore_ary1_a0_I2_p1_l[63] ,
         dpath_mulcore_ary1_a0_I2_p1_l[62] ,
         dpath_mulcore_ary1_a0_I2_p1_l[61] ,
         dpath_mulcore_ary1_a0_I2_p1_l[60] ,
         dpath_mulcore_ary1_a0_I2_p1_l[59] ,
         dpath_mulcore_ary1_a0_I2_p1_l[58] ,
         dpath_mulcore_ary1_a0_I2_p1_l[57] ,
         dpath_mulcore_ary1_a0_I2_p1_l[56] ,
         dpath_mulcore_ary1_a0_I2_p1_l[55] ,
         dpath_mulcore_ary1_a0_I2_p1_l[54] ,
         dpath_mulcore_ary1_a0_I2_p1_l[53] ,
         dpath_mulcore_ary1_a0_I2_p1_l[52] ,
         dpath_mulcore_ary1_a0_I2_p1_l[51] ,
         dpath_mulcore_ary1_a0_I2_p1_l[50] ,
         dpath_mulcore_ary1_a0_I2_p1_l[49] ,
         dpath_mulcore_ary1_a0_I2_p1_l[48] ,
         dpath_mulcore_ary1_a0_I2_p1_l[47] ,
         dpath_mulcore_ary1_a0_I2_p1_l[46] ,
         dpath_mulcore_ary1_a0_I2_p1_l[45] ,
         dpath_mulcore_ary1_a0_I2_p1_l[44] ,
         dpath_mulcore_ary1_a0_I2_p1_l[43] ,
         dpath_mulcore_ary1_a0_I2_p1_l[42] ,
         dpath_mulcore_ary1_a0_I2_p1_l[41] ,
         dpath_mulcore_ary1_a0_I2_p1_l[40] ,
         dpath_mulcore_ary1_a0_I2_p1_l[39] ,
         dpath_mulcore_ary1_a0_I2_p1_l[38] ,
         dpath_mulcore_ary1_a0_I2_p1_l[37] ,
         dpath_mulcore_ary1_a0_I2_p1_l[36] ,
         dpath_mulcore_ary1_a0_I2_p1_l[35] ,
         dpath_mulcore_ary1_a0_I2_p1_l[34] ,
         dpath_mulcore_ary1_a0_I2_p1_l[33] ,
         dpath_mulcore_ary1_a0_I2_p1_l[32] ,
         dpath_mulcore_ary1_a0_I2_p1_l[31] ,
         dpath_mulcore_ary1_a0_I2_p1_l[30] ,
         dpath_mulcore_ary1_a0_I2_p1_l[29] ,
         dpath_mulcore_ary1_a0_I2_p1_l[28] ,
         dpath_mulcore_ary1_a0_I2_p1_l[27] ,
         dpath_mulcore_ary1_a0_I2_p1_l[26] ,
         dpath_mulcore_ary1_a0_I2_p1_l[25] ,
         dpath_mulcore_ary1_a0_I2_p1_l[24] ,
         dpath_mulcore_ary1_a0_I2_p1_l[23] ,
         dpath_mulcore_ary1_a0_I2_p1_l[22] ,
         dpath_mulcore_ary1_a0_I2_p1_l[21] ,
         dpath_mulcore_ary1_a0_I2_p1_l[20] ,
         dpath_mulcore_ary1_a0_I2_p1_l[19] ,
         dpath_mulcore_ary1_a0_I2_p1_l[18] ,
         dpath_mulcore_ary1_a0_I2_p1_l[17] ,
         dpath_mulcore_ary1_a0_I2_p1_l[16] ,
         dpath_mulcore_ary1_a0_I2_p1_l[15] ,
         dpath_mulcore_ary1_a0_I2_p1_l[14] ,
         dpath_mulcore_ary1_a0_I2_p1_l[13] ,
         dpath_mulcore_ary1_a0_I2_p1_l[12] ,
         dpath_mulcore_ary1_a0_I2_p1_l[11] ,
         dpath_mulcore_ary1_a0_I2_p1_l[10] ,
         dpath_mulcore_ary1_a0_I2_p1_l[9] ,
         dpath_mulcore_ary1_a0_I2_p1_l[8] ,
         dpath_mulcore_ary1_a0_I2_p1_l[7] ,
         dpath_mulcore_ary1_a0_I2_p1_l[6] ,
         dpath_mulcore_ary1_a0_I2_p1_l[5] ,
         dpath_mulcore_ary1_a0_I2_p1_l[4] ,
         dpath_mulcore_ary1_a0_I2_p1_l[3] ,
         dpath_mulcore_ary1_a0_I1_p0_l[63] ,
         dpath_mulcore_ary1_a0_I1_p0_l[62] ,
         dpath_mulcore_ary1_a0_I1_p0_l[61] ,
         dpath_mulcore_ary1_a0_I1_p0_l[60] ,
         dpath_mulcore_ary1_a0_I1_p0_l[59] ,
         dpath_mulcore_ary1_a0_I1_p0_l[58] ,
         dpath_mulcore_ary1_a0_I1_p0_l[57] ,
         dpath_mulcore_ary1_a0_I1_p0_l[56] ,
         dpath_mulcore_ary1_a0_I1_p0_l[55] ,
         dpath_mulcore_ary1_a0_I1_p0_l[54] ,
         dpath_mulcore_ary1_a0_I1_p0_l[53] ,
         dpath_mulcore_ary1_a0_I1_p0_l[52] ,
         dpath_mulcore_ary1_a0_I1_p0_l[51] ,
         dpath_mulcore_ary1_a0_I1_p0_l[50] ,
         dpath_mulcore_ary1_a0_I1_p0_l[49] ,
         dpath_mulcore_ary1_a0_I1_p0_l[48] ,
         dpath_mulcore_ary1_a0_I1_p0_l[47] ,
         dpath_mulcore_ary1_a0_I1_p0_l[46] ,
         dpath_mulcore_ary1_a0_I1_p0_l[45] ,
         dpath_mulcore_ary1_a0_I1_p0_l[44] ,
         dpath_mulcore_ary1_a0_I1_p0_l[43] ,
         dpath_mulcore_ary1_a0_I1_p0_l[42] ,
         dpath_mulcore_ary1_a0_I1_p0_l[41] ,
         dpath_mulcore_ary1_a0_I1_p0_l[40] ,
         dpath_mulcore_ary1_a0_I1_p0_l[39] ,
         dpath_mulcore_ary1_a0_I1_p0_l[38] ,
         dpath_mulcore_ary1_a0_I1_p0_l[37] ,
         dpath_mulcore_ary1_a0_I1_p0_l[36] ,
         dpath_mulcore_ary1_a0_I1_p0_l[35] ,
         dpath_mulcore_ary1_a0_I1_p0_l[34] ,
         dpath_mulcore_ary1_a0_I1_p0_l[33] ,
         dpath_mulcore_ary1_a0_I1_p0_l[32] ,
         dpath_mulcore_ary1_a0_I1_p0_l[31] ,
         dpath_mulcore_ary1_a0_I1_p0_l[30] ,
         dpath_mulcore_ary1_a0_I1_p0_l[29] ,
         dpath_mulcore_ary1_a0_I1_p0_l[28] ,
         dpath_mulcore_ary1_a0_I1_p0_l[27] ,
         dpath_mulcore_ary1_a0_I1_p0_l[26] ,
         dpath_mulcore_ary1_a0_I1_p0_l[25] ,
         dpath_mulcore_ary1_a0_I1_p0_l[24] ,
         dpath_mulcore_ary1_a0_I1_p0_l[23] ,
         dpath_mulcore_ary1_a0_I1_p0_l[22] ,
         dpath_mulcore_ary1_a0_I1_p0_l[21] ,
         dpath_mulcore_ary1_a0_I1_p0_l[20] ,
         dpath_mulcore_ary1_a0_I1_p0_l[19] ,
         dpath_mulcore_ary1_a0_I1_p0_l[18] ,
         dpath_mulcore_ary1_a0_I1_p0_l[17] ,
         dpath_mulcore_ary1_a0_I1_p0_l[16] ,
         dpath_mulcore_ary1_a0_I1_p0_l[15] ,
         dpath_mulcore_ary1_a0_I1_p0_l[14] ,
         dpath_mulcore_ary1_a0_I1_p0_l[13] ,
         dpath_mulcore_ary1_a0_I1_p0_l[12] ,
         dpath_mulcore_ary1_a0_I1_p0_l[11] ,
         dpath_mulcore_ary1_a0_I1_p0_l[10] ,
         dpath_mulcore_ary1_a0_I1_p0_l[9] ,
         dpath_mulcore_ary1_a0_I1_p0_l[8] ,
         dpath_mulcore_ary1_a0_I1_p0_l[7] ,
         dpath_mulcore_ary1_a0_I1_p0_l[6] ,
         dpath_mulcore_ary1_a0_I1_p0_l[5] ,
         dpath_mulcore_ary1_a0_I1_p0_l[4] ,
         dpath_mulcore_ary1_a0_I1_p0_l[3] ,
         dpath_mulcore_ary1_a0_I1_p1_l[63] ,
         dpath_mulcore_ary1_a0_I1_p1_l[62] ,
         dpath_mulcore_ary1_a0_I1_p1_l[61] ,
         dpath_mulcore_ary1_a0_I1_p1_l[60] ,
         dpath_mulcore_ary1_a0_I1_p1_l[59] ,
         dpath_mulcore_ary1_a0_I1_p1_l[58] ,
         dpath_mulcore_ary1_a0_I1_p1_l[57] ,
         dpath_mulcore_ary1_a0_I1_p1_l[56] ,
         dpath_mulcore_ary1_a0_I1_p1_l[55] ,
         dpath_mulcore_ary1_a0_I1_p1_l[54] ,
         dpath_mulcore_ary1_a0_I1_p1_l[53] ,
         dpath_mulcore_ary1_a0_I1_p1_l[52] ,
         dpath_mulcore_ary1_a0_I1_p1_l[51] ,
         dpath_mulcore_ary1_a0_I1_p1_l[50] ,
         dpath_mulcore_ary1_a0_I1_p1_l[49] ,
         dpath_mulcore_ary1_a0_I1_p1_l[48] ,
         dpath_mulcore_ary1_a0_I1_p1_l[47] ,
         dpath_mulcore_ary1_a0_I1_p1_l[46] ,
         dpath_mulcore_ary1_a0_I1_p1_l[45] ,
         dpath_mulcore_ary1_a0_I1_p1_l[44] ,
         dpath_mulcore_ary1_a0_I1_p1_l[43] ,
         dpath_mulcore_ary1_a0_I1_p1_l[42] ,
         dpath_mulcore_ary1_a0_I1_p1_l[41] ,
         dpath_mulcore_ary1_a0_I1_p1_l[40] ,
         dpath_mulcore_ary1_a0_I1_p1_l[39] ,
         dpath_mulcore_ary1_a0_I1_p1_l[38] ,
         dpath_mulcore_ary1_a0_I1_p1_l[37] ,
         dpath_mulcore_ary1_a0_I1_p1_l[36] ,
         dpath_mulcore_ary1_a0_I1_p1_l[35] ,
         dpath_mulcore_ary1_a0_I1_p1_l[34] ,
         dpath_mulcore_ary1_a0_I1_p1_l[33] ,
         dpath_mulcore_ary1_a0_I1_p1_l[32] ,
         dpath_mulcore_ary1_a0_I1_p1_l[31] ,
         dpath_mulcore_ary1_a0_I1_p1_l[30] ,
         dpath_mulcore_ary1_a0_I1_p1_l[29] ,
         dpath_mulcore_ary1_a0_I1_p1_l[28] ,
         dpath_mulcore_ary1_a0_I1_p1_l[27] ,
         dpath_mulcore_ary1_a0_I1_p1_l[26] ,
         dpath_mulcore_ary1_a0_I1_p1_l[25] ,
         dpath_mulcore_ary1_a0_I1_p1_l[24] ,
         dpath_mulcore_ary1_a0_I1_p1_l[23] ,
         dpath_mulcore_ary1_a0_I1_p1_l[22] ,
         dpath_mulcore_ary1_a0_I1_p1_l[21] ,
         dpath_mulcore_ary1_a0_I1_p1_l[20] ,
         dpath_mulcore_ary1_a0_I1_p1_l[19] ,
         dpath_mulcore_ary1_a0_I1_p1_l[18] ,
         dpath_mulcore_ary1_a0_I1_p1_l[17] ,
         dpath_mulcore_ary1_a0_I1_p1_l[16] ,
         dpath_mulcore_ary1_a0_I1_p1_l[15] ,
         dpath_mulcore_ary1_a0_I1_p1_l[14] ,
         dpath_mulcore_ary1_a0_I1_p1_l[13] ,
         dpath_mulcore_ary1_a0_I1_p1_l[12] ,
         dpath_mulcore_ary1_a0_I1_p1_l[11] ,
         dpath_mulcore_ary1_a0_I1_p1_l[10] ,
         dpath_mulcore_ary1_a0_I1_p1_l[9] ,
         dpath_mulcore_ary1_a0_I1_p1_l[8] ,
         dpath_mulcore_ary1_a0_I1_p1_l[7] ,
         dpath_mulcore_ary1_a0_I1_p1_l[6] ,
         dpath_mulcore_ary1_a0_I1_p1_l[5] ,
         dpath_mulcore_ary1_a0_I1_p1_l[4] ,
         dpath_mulcore_ary1_a0_I1_p1_l[3] ,
         dpath_mulcore_ary1_a0_I1_p2_l[63] ,
         dpath_mulcore_ary1_a0_I1_p2_l[62] ,
         dpath_mulcore_ary1_a0_I1_p2_l[61] ,
         dpath_mulcore_ary1_a0_I1_p2_l[60] ,
         dpath_mulcore_ary1_a0_I1_p2_l[59] ,
         dpath_mulcore_ary1_a0_I1_p2_l[58] ,
         dpath_mulcore_ary1_a0_I1_p2_l[57] ,
         dpath_mulcore_ary1_a0_I1_p2_l[56] ,
         dpath_mulcore_ary1_a0_I1_p2_l[55] ,
         dpath_mulcore_ary1_a0_I1_p2_l[54] ,
         dpath_mulcore_ary1_a0_I1_p2_l[53] ,
         dpath_mulcore_ary1_a0_I1_p2_l[52] ,
         dpath_mulcore_ary1_a0_I1_p2_l[51] ,
         dpath_mulcore_ary1_a0_I1_p2_l[50] ,
         dpath_mulcore_ary1_a0_I1_p2_l[49] ,
         dpath_mulcore_ary1_a0_I1_p2_l[48] ,
         dpath_mulcore_ary1_a0_I1_p2_l[47] ,
         dpath_mulcore_ary1_a0_I1_p2_l[46] ,
         dpath_mulcore_ary1_a0_I1_p2_l[45] ,
         dpath_mulcore_ary1_a0_I1_p2_l[44] ,
         dpath_mulcore_ary1_a0_I1_p2_l[43] ,
         dpath_mulcore_ary1_a0_I1_p2_l[42] ,
         dpath_mulcore_ary1_a0_I1_p2_l[41] ,
         dpath_mulcore_ary1_a0_I1_p2_l[40] ,
         dpath_mulcore_ary1_a0_I1_p2_l[39] ,
         dpath_mulcore_ary1_a0_I1_p2_l[38] ,
         dpath_mulcore_ary1_a0_I1_p2_l[37] ,
         dpath_mulcore_ary1_a0_I1_p2_l[36] ,
         dpath_mulcore_ary1_a0_I1_p2_l[35] ,
         dpath_mulcore_ary1_a0_I1_p2_l[34] ,
         dpath_mulcore_ary1_a0_I1_p2_l[33] ,
         dpath_mulcore_ary1_a0_I1_p2_l[32] ,
         dpath_mulcore_ary1_a0_I1_p2_l[31] ,
         dpath_mulcore_ary1_a0_I1_p2_l[30] ,
         dpath_mulcore_ary1_a0_I1_p2_l[29] ,
         dpath_mulcore_ary1_a0_I1_p2_l[28] ,
         dpath_mulcore_ary1_a0_I1_p2_l[27] ,
         dpath_mulcore_ary1_a0_I1_p2_l[26] ,
         dpath_mulcore_ary1_a0_I1_p2_l[25] ,
         dpath_mulcore_ary1_a0_I1_p2_l[24] ,
         dpath_mulcore_ary1_a0_I1_p2_l[23] ,
         dpath_mulcore_ary1_a0_I1_p2_l[22] ,
         dpath_mulcore_ary1_a0_I1_p2_l[21] ,
         dpath_mulcore_ary1_a0_I1_p2_l[20] ,
         dpath_mulcore_ary1_a0_I1_p2_l[19] ,
         dpath_mulcore_ary1_a0_I1_p2_l[18] ,
         dpath_mulcore_ary1_a0_I1_p2_l[17] ,
         dpath_mulcore_ary1_a0_I1_p2_l[16] ,
         dpath_mulcore_ary1_a0_I1_p2_l[15] ,
         dpath_mulcore_ary1_a0_I1_p2_l[14] ,
         dpath_mulcore_ary1_a0_I1_p2_l[13] ,
         dpath_mulcore_ary1_a0_I1_p2_l[12] ,
         dpath_mulcore_ary1_a0_I1_p2_l[11] ,
         dpath_mulcore_ary1_a0_I1_p2_l[10] ,
         dpath_mulcore_ary1_a0_I1_p2_l[9] ,
         dpath_mulcore_ary1_a0_I1_p2_l[8] ,
         dpath_mulcore_ary1_a0_I1_p2_l[7] ,
         dpath_mulcore_ary1_a0_I1_p2_l[6] ,
         dpath_mulcore_ary1_a0_I1_p2_l[5] ,
         dpath_mulcore_ary1_a0_I1_p2_l[4] , dpath_mulcore_array2_sh_82__n3 ,
         dpath_mulcore_array2_sh_82__n2 , dpath_mulcore_ary1_a0_I2_I2_net48 ,
         dpath_mulcore_ary1_a0_I2_I2_net43 ,
         dpath_mulcore_ary1_a0_I2_I2_p1_l_64 ,
         dpath_mulcore_ary1_a0_I2_I2_net0118 ,
         dpath_mulcore_ary1_a0_I2_I2_net38 ,
         dpath_mulcore_ary1_a0_I2_I2_p1_l_65 ,
         dpath_mulcore_ary1_a0_I2_I2_net47 ,
         dpath_mulcore_ary1_a0_I2_I2_net088 ,
         dpath_mulcore_ary1_a0_I2_I1_63__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_63__net046 ,
         dpath_mulcore_ary1_a0_I2_I0_n1 ,
         dpath_mulcore_ary1_a0_I2_I0_p0_l_0 ,
         dpath_mulcore_ary1_a0_I2_I0_p0_l_1 ,
         dpath_mulcore_ary1_a0_I2_I0_p1_l_2 ,
         dpath_mulcore_ary1_a0_I2_I0_p0_l_2 ,
         dpath_mulcore_ary1_a0_I2_I0_p0_1 ,
         dpath_mulcore_ary1_a0_I2_I0_p1_3 ,
         dpath_mulcore_ary1_a0_I2_I0_p0_3 ,
         dpath_mulcore_ary1_a0_I2_I0_p0_2 ,
         dpath_mulcore_ary1_a0_I2_I0_b1n_0 ,
         dpath_mulcore_ary1_a0_I2_I0_b1n_1 ,
         dpath_mulcore_ary1_a0_I2_I0_b0n ,
         dpath_mulcore_ary1_a0_I2_I0_b0n_0 ,
         dpath_mulcore_ary1_a0_I2_I0_b0n_1 ,
         dpath_mulcore_ary1_a0_I1_I2_net35 ,
         dpath_mulcore_ary1_a0_I1_I2_net48 ,
         dpath_mulcore_ary1_a0_I1_I2_net43 ,
         dpath_mulcore_ary1_a0_I1_I2_p1_l_64 ,
         dpath_mulcore_ary1_a0_I1_I2_net15 ,
         dpath_mulcore_ary1_a0_I1_I2_p2_l_64 ,
         dpath_mulcore_ary1_a0_I1_I2_net8 ,
         dpath_mulcore_ary1_a0_I1_I2_p2_l_65 ,
         dpath_mulcore_ary1_a0_I1_I2_net078 ,
         dpath_mulcore_ary1_a0_I1_I2_p2_l_66 ,
         dpath_mulcore_ary1_a0_I1_I2_net0118 ,
         dpath_mulcore_ary1_a0_I1_I2_net38 ,
         dpath_mulcore_ary1_a0_I1_I2_p1_l_65 ,
         dpath_mulcore_ary1_a0_I1_I2_net073 ,
         dpath_mulcore_ary1_a0_I1_I2_p2_l_67 ,
         dpath_mulcore_ary1_a0_I1_I2_net47 ,
         dpath_mulcore_ary1_a0_I1_I2_net088 ,
         dpath_mulcore_ary1_a0_I1_I2_net075 ,
         dpath_mulcore_ary1_a0_I2_I2_p0_64__n3 ,
         dpath_mulcore_ary1_a0_I2_I2_p0_64__n2 ,
         dpath_mulcore_booth_ckbuf_1_clken , dpath_mulcore_booth_ckbuf_1_N1 ,
         dpath_mulcore_ckbuf_1_clken , dpath_mulcore_array2_sc3_20__z ,
         dpath_mulcore_array2_sc3_21__z , dpath_mulcore_array2_sc3_22__z ,
         dpath_mulcore_array2_sc3_23__z , dpath_mulcore_array2_sc3_24__z ,
         dpath_mulcore_array2_sc3_25__z , dpath_mulcore_array2_sc3_26__z ,
         dpath_mulcore_array2_sc3_27__z , dpath_mulcore_array2_sc3_28__z ,
         dpath_mulcore_array2_sc3_29__z , dpath_mulcore_array2_sc3_30__z ,
         dpath_mulcore_array2_sc3_31__z , dpath_mulcore_array2_sc3_32__z ,
         dpath_mulcore_array2_sc3_33__z , dpath_mulcore_array2_sc3_34__z ,
         dpath_mulcore_array2_sc3_35__z , dpath_mulcore_array2_sc3_36__z ,
         dpath_mulcore_array2_sc3_37__z , dpath_mulcore_array2_sc3_38__z ,
         dpath_mulcore_array2_sc3_39__z , dpath_mulcore_array2_sc3_40__z ,
         dpath_mulcore_array2_sc3_41__z , dpath_mulcore_array2_sc3_42__z ,
         dpath_mulcore_array2_sc3_43__z , dpath_mulcore_array2_sc3_44__z ,
         dpath_mulcore_array2_sc3_45__z , dpath_mulcore_array2_sc3_46__z ,
         dpath_mulcore_array2_sc3_47__z , dpath_mulcore_array2_sc3_48__z ,
         dpath_mulcore_array2_sc3_49__z , dpath_mulcore_array2_sc3_50__z ,
         dpath_mulcore_array2_sc3_51__z , dpath_mulcore_array2_sc3_52__z ,
         dpath_mulcore_array2_sc3_53__z , dpath_mulcore_array2_sc3_54__z ,
         dpath_mulcore_array2_sc3_55__z , dpath_mulcore_array2_sc3_56__z ,
         dpath_mulcore_array2_sc3_57__z , dpath_mulcore_array2_sc3_58__z ,
         dpath_mulcore_array2_sc3_59__z , dpath_mulcore_array2_sc3_60__z ,
         dpath_mulcore_array2_sc3_61__z , dpath_mulcore_array2_sc3_62__z ,
         dpath_mulcore_array2_sc3_63__z , dpath_mulcore_array2_sc3_64__z ,
         dpath_mulcore_array2_sc3_65__z , dpath_mulcore_array2_sc3_66__z ,
         dpath_mulcore_array2_sc3_67__z , dpath_mulcore_array2_sc3_68__z ,
         dpath_mulcore_ary1_a1_sc3_11__z , dpath_mulcore_ary1_a1_sc3_12__z ,
         dpath_mulcore_ary1_a1_sc3_13__z , dpath_mulcore_ary1_a1_sc3_14__z ,
         dpath_mulcore_ary1_a1_sc3_15__z , dpath_mulcore_ary1_a1_sc3_16__z ,
         dpath_mulcore_ary1_a1_sc3_17__z , dpath_mulcore_ary1_a1_sc3_18__z ,
         dpath_mulcore_ary1_a1_sc3_19__z , dpath_mulcore_ary1_a1_sc3_20__z ,
         dpath_mulcore_ary1_a1_sc3_21__z , dpath_mulcore_ary1_a1_sc3_22__z ,
         dpath_mulcore_ary1_a1_sc3_23__z , dpath_mulcore_ary1_a1_sc3_24__z ,
         dpath_mulcore_ary1_a1_sc3_25__z , dpath_mulcore_ary1_a1_sc3_26__z ,
         dpath_mulcore_ary1_a1_sc3_27__z , dpath_mulcore_ary1_a1_sc3_28__z ,
         dpath_mulcore_ary1_a1_sc3_29__z , dpath_mulcore_ary1_a1_sc3_30__z ,
         dpath_mulcore_ary1_a1_sc3_31__z , dpath_mulcore_ary1_a1_sc3_32__z ,
         dpath_mulcore_ary1_a1_sc3_33__z , dpath_mulcore_ary1_a1_sc3_34__z ,
         dpath_mulcore_ary1_a1_sc3_35__z , dpath_mulcore_ary1_a1_sc3_36__z ,
         dpath_mulcore_ary1_a1_sc3_37__z , dpath_mulcore_ary1_a1_sc3_38__z ,
         dpath_mulcore_ary1_a1_sc3_39__z , dpath_mulcore_ary1_a1_sc3_40__z ,
         dpath_mulcore_ary1_a1_sc3_41__z , dpath_mulcore_ary1_a1_sc3_42__z ,
         dpath_mulcore_ary1_a1_sc3_43__z , dpath_mulcore_ary1_a1_sc3_44__z ,
         dpath_mulcore_ary1_a1_sc3_45__z , dpath_mulcore_ary1_a1_sc3_46__z ,
         dpath_mulcore_ary1_a1_sc3_47__z , dpath_mulcore_ary1_a1_sc3_48__z ,
         dpath_mulcore_ary1_a1_sc3_49__z , dpath_mulcore_ary1_a1_sc3_50__z ,
         dpath_mulcore_ary1_a1_sc3_51__z , dpath_mulcore_ary1_a1_sc3_52__z ,
         dpath_mulcore_ary1_a1_sc3_53__z , dpath_mulcore_ary1_a1_sc3_54__z ,
         dpath_mulcore_ary1_a1_sc3_55__z , dpath_mulcore_ary1_a1_sc3_56__z ,
         dpath_mulcore_ary1_a1_sc3_57__z , dpath_mulcore_ary1_a1_sc3_58__z ,
         dpath_mulcore_ary1_a1_sc3_59__z , dpath_mulcore_ary1_a1_sc3_60__z ,
         dpath_mulcore_ary1_a1_sc3_61__z , dpath_mulcore_ary1_a1_sc3_62__z ,
         dpath_mulcore_ary1_a1_sc3_63__z , dpath_mulcore_ary1_a1_sc3_64__z ,
         dpath_mulcore_ary1_a1_sc3_65__z , dpath_mulcore_ary1_a1_sc3_66__z ,
         dpath_mulcore_ary1_a1_sc3_67__z , dpath_mulcore_ary1_a1_sc3_68__z ,
         dpath_mulcore_ary1_a1_sc3_69__z , dpath_mulcore_ary1_a1_sc3_70__z ,
         dpath_mulcore_ary1_a1_sc3_76__z , dpath_mulcore_ary1_a1_sc3_72__z ,
         dpath_mulcore_ary1_a1_sc3_73__z , dpath_mulcore_ary1_a1_sc3_74__z ,
         dpath_mulcore_ary1_a1_sc3_75__z , dpath_mulcore_ary1_a1_sc3_71__z ,
         dpath_mulcore_ary1_a0_sc3_11__z , dpath_mulcore_ary1_a0_sc3_12__z ,
         dpath_mulcore_ary1_a0_sc3_13__z , dpath_mulcore_ary1_a0_sc3_14__z ,
         dpath_mulcore_ary1_a0_sc3_15__z , dpath_mulcore_ary1_a0_sc3_16__z ,
         dpath_mulcore_ary1_a0_sc3_17__z , dpath_mulcore_ary1_a0_sc3_18__z ,
         dpath_mulcore_ary1_a0_sc3_19__z , dpath_mulcore_ary1_a0_sc3_20__z ,
         dpath_mulcore_ary1_a0_sc3_21__z , dpath_mulcore_ary1_a0_sc3_22__z ,
         dpath_mulcore_ary1_a0_sc3_23__z , dpath_mulcore_ary1_a0_sc3_24__z ,
         dpath_mulcore_ary1_a0_sc3_25__z , dpath_mulcore_ary1_a0_sc3_26__z ,
         dpath_mulcore_ary1_a0_sc3_27__z , dpath_mulcore_ary1_a0_sc3_28__z ,
         dpath_mulcore_ary1_a0_sc3_29__z , dpath_mulcore_ary1_a0_sc3_30__z ,
         dpath_mulcore_ary1_a0_sc3_31__z , dpath_mulcore_ary1_a0_sc3_32__z ,
         dpath_mulcore_ary1_a0_sc3_33__z , dpath_mulcore_ary1_a0_sc3_34__z ,
         dpath_mulcore_ary1_a0_sc3_35__z , dpath_mulcore_ary1_a0_sc3_36__z ,
         dpath_mulcore_ary1_a0_sc3_37__z , dpath_mulcore_ary1_a0_sc3_38__z ,
         dpath_mulcore_ary1_a0_sc3_39__z , dpath_mulcore_ary1_a0_sc3_40__z ,
         dpath_mulcore_ary1_a0_sc3_41__z , dpath_mulcore_ary1_a0_sc3_42__z ,
         dpath_mulcore_ary1_a0_sc3_43__z , dpath_mulcore_ary1_a0_sc3_44__z ,
         dpath_mulcore_ary1_a0_sc3_45__z , dpath_mulcore_ary1_a0_sc3_46__z ,
         dpath_mulcore_ary1_a0_sc3_47__z , dpath_mulcore_ary1_a0_sc3_48__z ,
         dpath_mulcore_ary1_a0_sc3_49__z , dpath_mulcore_ary1_a0_sc3_50__z ,
         dpath_mulcore_ary1_a0_sc3_51__z , dpath_mulcore_ary1_a0_sc3_52__z ,
         dpath_mulcore_ary1_a0_sc3_53__z , dpath_mulcore_ary1_a0_sc3_54__z ,
         dpath_mulcore_ary1_a0_sc3_55__z , dpath_mulcore_ary1_a0_sc3_56__z ,
         dpath_mulcore_ary1_a0_sc3_57__z , dpath_mulcore_ary1_a0_sc3_58__z ,
         dpath_mulcore_ary1_a0_sc3_59__z , dpath_mulcore_ary1_a0_sc3_60__z ,
         dpath_mulcore_ary1_a0_sc3_61__z , dpath_mulcore_ary1_a0_sc3_62__z ,
         dpath_mulcore_ary1_a0_sc3_63__z , dpath_mulcore_ary1_a0_sc3_64__z ,
         dpath_mulcore_ary1_a0_sc3_65__z , dpath_mulcore_ary1_a0_sc3_66__z ,
         dpath_mulcore_ary1_a0_sc3_67__z , dpath_mulcore_ary1_a0_sc3_68__z ,
         dpath_mulcore_ary1_a0_sc3_69__z , dpath_mulcore_ary1_a0_sc3_70__z ,
         dpath_mulcore_ary1_a0_sc3_76__z , dpath_mulcore_ary1_a0_sc3_72__z ,
         dpath_mulcore_ary1_a0_sc3_73__z , dpath_mulcore_ary1_a0_sc3_74__z ,
         dpath_mulcore_ary1_a0_sc3_75__z ,
         dpath_mulcore_ary1_a1_I0_p0_l[63] ,
         dpath_mulcore_ary1_a1_I0_p0_l[62] ,
         dpath_mulcore_ary1_a1_I0_p0_l[61] ,
         dpath_mulcore_ary1_a1_I0_p0_l[60] ,
         dpath_mulcore_ary1_a1_I0_p0_l[59] ,
         dpath_mulcore_ary1_a1_I0_p0_l[58] ,
         dpath_mulcore_ary1_a1_I0_p0_l[57] ,
         dpath_mulcore_ary1_a1_I0_p0_l[56] ,
         dpath_mulcore_ary1_a1_I0_p0_l[55] ,
         dpath_mulcore_ary1_a1_I0_p0_l[54] ,
         dpath_mulcore_ary1_a1_I0_p0_l[53] ,
         dpath_mulcore_ary1_a1_I0_p0_l[52] ,
         dpath_mulcore_ary1_a1_I0_p0_l[51] ,
         dpath_mulcore_ary1_a1_I0_p0_l[50] ,
         dpath_mulcore_ary1_a1_I0_p0_l[49] ,
         dpath_mulcore_ary1_a1_I0_p0_l[48] ,
         dpath_mulcore_ary1_a1_I0_p0_l[47] ,
         dpath_mulcore_ary1_a1_I0_p0_l[46] ,
         dpath_mulcore_ary1_a1_I0_p0_l[45] ,
         dpath_mulcore_ary1_a1_I0_p0_l[44] ,
         dpath_mulcore_ary1_a1_I0_p0_l[43] ,
         dpath_mulcore_ary1_a1_I0_p0_l[42] ,
         dpath_mulcore_ary1_a1_I0_p0_l[41] ,
         dpath_mulcore_ary1_a1_I0_p0_l[40] ,
         dpath_mulcore_ary1_a1_I0_p0_l[39] ,
         dpath_mulcore_ary1_a1_I0_p0_l[38] ,
         dpath_mulcore_ary1_a1_I0_p0_l[37] ,
         dpath_mulcore_ary1_a1_I0_p0_l[36] ,
         dpath_mulcore_ary1_a1_I0_p0_l[35] ,
         dpath_mulcore_ary1_a1_I0_p0_l[34] ,
         dpath_mulcore_ary1_a1_I0_p0_l[33] ,
         dpath_mulcore_ary1_a1_I0_p0_l[32] ,
         dpath_mulcore_ary1_a1_I0_p0_l[31] ,
         dpath_mulcore_ary1_a1_I0_p0_l[30] ,
         dpath_mulcore_ary1_a1_I0_p0_l[29] ,
         dpath_mulcore_ary1_a1_I0_p0_l[28] ,
         dpath_mulcore_ary1_a1_I0_p0_l[27] ,
         dpath_mulcore_ary1_a1_I0_p0_l[26] ,
         dpath_mulcore_ary1_a1_I0_p0_l[25] ,
         dpath_mulcore_ary1_a1_I0_p0_l[24] ,
         dpath_mulcore_ary1_a1_I0_p0_l[23] ,
         dpath_mulcore_ary1_a1_I0_p0_l[22] ,
         dpath_mulcore_ary1_a1_I0_p0_l[21] ,
         dpath_mulcore_ary1_a1_I0_p0_l[20] ,
         dpath_mulcore_ary1_a1_I0_p0_l[19] ,
         dpath_mulcore_ary1_a1_I0_p0_l[18] ,
         dpath_mulcore_ary1_a1_I0_p0_l[17] ,
         dpath_mulcore_ary1_a1_I0_p0_l[16] ,
         dpath_mulcore_ary1_a1_I0_p0_l[15] ,
         dpath_mulcore_ary1_a1_I0_p0_l[14] ,
         dpath_mulcore_ary1_a1_I0_p0_l[13] ,
         dpath_mulcore_ary1_a1_I0_p0_l[12] ,
         dpath_mulcore_ary1_a1_I0_p0_l[11] ,
         dpath_mulcore_ary1_a1_I0_p0_l[10] ,
         dpath_mulcore_ary1_a1_I0_p0_l[9] ,
         dpath_mulcore_ary1_a1_I0_p0_l[8] ,
         dpath_mulcore_ary1_a1_I0_p0_l[7] ,
         dpath_mulcore_ary1_a1_I0_p0_l[6] ,
         dpath_mulcore_ary1_a1_I0_p0_l[5] ,
         dpath_mulcore_ary1_a1_I0_p0_l[4] ,
         dpath_mulcore_ary1_a1_I0_p0_l[3] ,
         dpath_mulcore_ary1_a1_I0_p1_l[63] ,
         dpath_mulcore_ary1_a1_I0_p1_l[62] ,
         dpath_mulcore_ary1_a1_I0_p1_l[61] ,
         dpath_mulcore_ary1_a1_I0_p1_l[60] ,
         dpath_mulcore_ary1_a1_I0_p1_l[59] ,
         dpath_mulcore_ary1_a1_I0_p1_l[58] ,
         dpath_mulcore_ary1_a1_I0_p1_l[57] ,
         dpath_mulcore_ary1_a1_I0_p1_l[56] ,
         dpath_mulcore_ary1_a1_I0_p1_l[55] ,
         dpath_mulcore_ary1_a1_I0_p1_l[54] ,
         dpath_mulcore_ary1_a1_I0_p1_l[53] ,
         dpath_mulcore_ary1_a1_I0_p1_l[52] ,
         dpath_mulcore_ary1_a1_I0_p1_l[51] ,
         dpath_mulcore_ary1_a1_I0_p1_l[50] ,
         dpath_mulcore_ary1_a1_I0_p1_l[49] ,
         dpath_mulcore_ary1_a1_I0_p1_l[48] ,
         dpath_mulcore_ary1_a1_I0_p1_l[47] ,
         dpath_mulcore_ary1_a1_I0_p1_l[46] ,
         dpath_mulcore_ary1_a1_I0_p1_l[45] ,
         dpath_mulcore_ary1_a1_I0_p1_l[44] ,
         dpath_mulcore_ary1_a1_I0_p1_l[43] ,
         dpath_mulcore_ary1_a1_I0_p1_l[42] ,
         dpath_mulcore_ary1_a1_I0_p1_l[41] ,
         dpath_mulcore_ary1_a1_I0_p1_l[40] ,
         dpath_mulcore_ary1_a1_I0_p1_l[39] ,
         dpath_mulcore_ary1_a1_I0_p1_l[38] ,
         dpath_mulcore_ary1_a1_I0_p1_l[37] ,
         dpath_mulcore_ary1_a1_I0_p1_l[36] ,
         dpath_mulcore_ary1_a1_I0_p1_l[35] ,
         dpath_mulcore_ary1_a1_I0_p1_l[34] ,
         dpath_mulcore_ary1_a1_I0_p1_l[33] ,
         dpath_mulcore_ary1_a1_I0_p1_l[32] ,
         dpath_mulcore_ary1_a1_I0_p1_l[31] ,
         dpath_mulcore_ary1_a1_I0_p1_l[30] ,
         dpath_mulcore_ary1_a1_I0_p1_l[29] ,
         dpath_mulcore_ary1_a1_I0_p1_l[28] ,
         dpath_mulcore_ary1_a1_I0_p1_l[27] ,
         dpath_mulcore_ary1_a1_I0_p1_l[26] ,
         dpath_mulcore_ary1_a1_I0_p1_l[25] ,
         dpath_mulcore_ary1_a1_I0_p1_l[24] ,
         dpath_mulcore_ary1_a1_I0_p1_l[23] ,
         dpath_mulcore_ary1_a1_I0_p1_l[22] ,
         dpath_mulcore_ary1_a1_I0_p1_l[21] ,
         dpath_mulcore_ary1_a1_I0_p1_l[20] ,
         dpath_mulcore_ary1_a1_I0_p1_l[19] ,
         dpath_mulcore_ary1_a1_I0_p1_l[18] ,
         dpath_mulcore_ary1_a1_I0_p1_l[17] ,
         dpath_mulcore_ary1_a1_I0_p1_l[16] ,
         dpath_mulcore_ary1_a1_I0_p1_l[15] ,
         dpath_mulcore_ary1_a1_I0_p1_l[14] ,
         dpath_mulcore_ary1_a1_I0_p1_l[13] ,
         dpath_mulcore_ary1_a1_I0_p1_l[12] ,
         dpath_mulcore_ary1_a1_I0_p1_l[11] ,
         dpath_mulcore_ary1_a1_I0_p1_l[10] ,
         dpath_mulcore_ary1_a1_I0_p1_l[9] ,
         dpath_mulcore_ary1_a1_I0_p1_l[8] ,
         dpath_mulcore_ary1_a1_I0_p1_l[7] ,
         dpath_mulcore_ary1_a1_I0_p1_l[6] ,
         dpath_mulcore_ary1_a1_I0_p1_l[5] ,
         dpath_mulcore_ary1_a1_I0_p1_l[4] ,
         dpath_mulcore_ary1_a1_I0_p1_l[3] ,
         dpath_mulcore_ary1_a1_I0_p2_l[63] ,
         dpath_mulcore_ary1_a1_I0_p2_l[62] ,
         dpath_mulcore_ary1_a1_I0_p2_l[61] ,
         dpath_mulcore_ary1_a1_I0_p2_l[60] ,
         dpath_mulcore_ary1_a1_I0_p2_l[59] ,
         dpath_mulcore_ary1_a1_I0_p2_l[58] ,
         dpath_mulcore_ary1_a1_I0_p2_l[57] ,
         dpath_mulcore_ary1_a1_I0_p2_l[56] ,
         dpath_mulcore_ary1_a1_I0_p2_l[55] ,
         dpath_mulcore_ary1_a1_I0_p2_l[54] ,
         dpath_mulcore_ary1_a1_I0_p2_l[53] ,
         dpath_mulcore_ary1_a1_I0_p2_l[52] ,
         dpath_mulcore_ary1_a1_I0_p2_l[51] ,
         dpath_mulcore_ary1_a1_I0_p2_l[50] ,
         dpath_mulcore_ary1_a1_I0_p2_l[49] ,
         dpath_mulcore_ary1_a1_I0_p2_l[48] ,
         dpath_mulcore_ary1_a1_I0_p2_l[47] ,
         dpath_mulcore_ary1_a1_I0_p2_l[46] ,
         dpath_mulcore_ary1_a1_I0_p2_l[45] ,
         dpath_mulcore_ary1_a1_I0_p2_l[44] ,
         dpath_mulcore_ary1_a1_I0_p2_l[43] ,
         dpath_mulcore_ary1_a1_I0_p2_l[42] ,
         dpath_mulcore_ary1_a1_I0_p2_l[41] ,
         dpath_mulcore_ary1_a1_I0_p2_l[40] ,
         dpath_mulcore_ary1_a1_I0_p2_l[39] ,
         dpath_mulcore_ary1_a1_I0_p2_l[38] ,
         dpath_mulcore_ary1_a1_I0_p2_l[37] ,
         dpath_mulcore_ary1_a1_I0_p2_l[36] ,
         dpath_mulcore_ary1_a1_I0_p2_l[35] ,
         dpath_mulcore_ary1_a1_I0_p2_l[34] ,
         dpath_mulcore_ary1_a1_I0_p2_l[33] ,
         dpath_mulcore_ary1_a1_I0_p2_l[32] ,
         dpath_mulcore_ary1_a1_I0_p2_l[31] ,
         dpath_mulcore_ary1_a1_I0_p2_l[30] ,
         dpath_mulcore_ary1_a1_I0_p2_l[29] ,
         dpath_mulcore_ary1_a1_I0_p2_l[28] ,
         dpath_mulcore_ary1_a1_I0_p2_l[27] ,
         dpath_mulcore_ary1_a1_I0_p2_l[26] ,
         dpath_mulcore_ary1_a1_I0_p2_l[25] ,
         dpath_mulcore_ary1_a1_I0_p2_l[24] ,
         dpath_mulcore_ary1_a1_I0_p2_l[23] ,
         dpath_mulcore_ary1_a1_I0_p2_l[22] ,
         dpath_mulcore_ary1_a1_I0_p2_l[21] ,
         dpath_mulcore_ary1_a1_I0_p2_l[20] ,
         dpath_mulcore_ary1_a1_I0_p2_l[19] ,
         dpath_mulcore_ary1_a1_I0_p2_l[18] ,
         dpath_mulcore_ary1_a1_I0_p2_l[17] ,
         dpath_mulcore_ary1_a1_I0_p2_l[16] ,
         dpath_mulcore_ary1_a1_I0_p2_l[15] ,
         dpath_mulcore_ary1_a1_I0_p2_l[14] ,
         dpath_mulcore_ary1_a1_I0_p2_l[13] ,
         dpath_mulcore_ary1_a1_I0_p2_l[12] ,
         dpath_mulcore_ary1_a1_I0_p2_l[11] ,
         dpath_mulcore_ary1_a1_I0_p2_l[10] ,
         dpath_mulcore_ary1_a1_I0_p2_l[9] ,
         dpath_mulcore_ary1_a1_I0_p2_l[8] ,
         dpath_mulcore_ary1_a1_I0_p2_l[7] ,
         dpath_mulcore_ary1_a1_I0_p2_l[6] ,
         dpath_mulcore_ary1_a1_I0_p2_l[5] ,
         dpath_mulcore_ary1_a1_I0_p2_l[4] ,
         dpath_mulcore_ary1_a1_I1_p0_l[63] ,
         dpath_mulcore_ary1_a1_I1_p0_l[62] ,
         dpath_mulcore_ary1_a1_I1_p0_l[61] ,
         dpath_mulcore_ary1_a1_I1_p0_l[60] ,
         dpath_mulcore_ary1_a1_I1_p0_l[59] ,
         dpath_mulcore_ary1_a1_I1_p0_l[58] ,
         dpath_mulcore_ary1_a1_I1_p0_l[57] ,
         dpath_mulcore_ary1_a1_I1_p0_l[56] ,
         dpath_mulcore_ary1_a1_I1_p0_l[55] ,
         dpath_mulcore_ary1_a1_I1_p0_l[54] ,
         dpath_mulcore_ary1_a1_I1_p0_l[53] ,
         dpath_mulcore_ary1_a1_I1_p0_l[52] ,
         dpath_mulcore_ary1_a1_I1_p0_l[51] ,
         dpath_mulcore_ary1_a1_I1_p0_l[50] ,
         dpath_mulcore_ary1_a1_I1_p0_l[49] ,
         dpath_mulcore_ary1_a1_I1_p0_l[48] ,
         dpath_mulcore_ary1_a1_I1_p0_l[47] ,
         dpath_mulcore_ary1_a1_I1_p0_l[46] ,
         dpath_mulcore_ary1_a1_I1_p0_l[45] ,
         dpath_mulcore_ary1_a1_I1_p0_l[44] ,
         dpath_mulcore_ary1_a1_I1_p0_l[43] ,
         dpath_mulcore_ary1_a1_I1_p0_l[42] ,
         dpath_mulcore_ary1_a1_I1_p0_l[41] ,
         dpath_mulcore_ary1_a1_I1_p0_l[40] ,
         dpath_mulcore_ary1_a1_I1_p0_l[39] ,
         dpath_mulcore_ary1_a1_I1_p0_l[38] ,
         dpath_mulcore_ary1_a1_I1_p0_l[37] ,
         dpath_mulcore_ary1_a1_I1_p0_l[36] ,
         dpath_mulcore_ary1_a1_I1_p0_l[35] ,
         dpath_mulcore_ary1_a1_I1_p0_l[34] ,
         dpath_mulcore_ary1_a1_I1_p0_l[33] ,
         dpath_mulcore_ary1_a1_I1_p0_l[32] ,
         dpath_mulcore_ary1_a1_I1_p0_l[31] ,
         dpath_mulcore_ary1_a1_I1_p0_l[30] ,
         dpath_mulcore_ary1_a1_I1_p0_l[29] ,
         dpath_mulcore_ary1_a1_I1_p0_l[28] ,
         dpath_mulcore_ary1_a1_I1_p0_l[27] ,
         dpath_mulcore_ary1_a1_I1_p0_l[26] ,
         dpath_mulcore_ary1_a1_I1_p0_l[25] ,
         dpath_mulcore_ary1_a1_I1_p0_l[24] ,
         dpath_mulcore_ary1_a1_I1_p0_l[23] ,
         dpath_mulcore_ary1_a1_I1_p0_l[22] ,
         dpath_mulcore_ary1_a1_I1_p0_l[21] ,
         dpath_mulcore_ary1_a1_I1_p0_l[20] ,
         dpath_mulcore_ary1_a1_I1_p0_l[19] ,
         dpath_mulcore_ary1_a1_I1_p0_l[18] ,
         dpath_mulcore_ary1_a1_I1_p0_l[17] ,
         dpath_mulcore_ary1_a1_I1_p0_l[16] ,
         dpath_mulcore_ary1_a1_I1_p0_l[15] ,
         dpath_mulcore_ary1_a1_I1_p0_l[14] ,
         dpath_mulcore_ary1_a1_I1_p0_l[13] ,
         dpath_mulcore_ary1_a1_I1_p0_l[12] ,
         dpath_mulcore_ary1_a1_I1_p0_l[11] ,
         dpath_mulcore_ary1_a1_I1_p0_l[10] ,
         dpath_mulcore_ary1_a1_I1_p0_l[9] ,
         dpath_mulcore_ary1_a1_I1_p0_l[8] ,
         dpath_mulcore_ary1_a1_I1_p0_l[7] ,
         dpath_mulcore_ary1_a1_I1_p0_l[6] ,
         dpath_mulcore_ary1_a1_I1_p0_l[5] ,
         dpath_mulcore_ary1_a1_I1_p0_l[4] ,
         dpath_mulcore_ary1_a1_I1_p0_l[3] ,
         dpath_mulcore_ary1_a1_I1_p1_l[63] ,
         dpath_mulcore_ary1_a1_I1_p1_l[62] ,
         dpath_mulcore_ary1_a1_I1_p1_l[61] ,
         dpath_mulcore_ary1_a1_I1_p1_l[60] ,
         dpath_mulcore_ary1_a1_I1_p1_l[59] ,
         dpath_mulcore_ary1_a1_I1_p1_l[58] ,
         dpath_mulcore_ary1_a1_I1_p1_l[57] ,
         dpath_mulcore_ary1_a1_I1_p1_l[56] ,
         dpath_mulcore_ary1_a1_I1_p1_l[55] ,
         dpath_mulcore_ary1_a1_I1_p1_l[54] ,
         dpath_mulcore_ary1_a1_I1_p1_l[53] ,
         dpath_mulcore_ary1_a1_I1_p1_l[52] ,
         dpath_mulcore_ary1_a1_I1_p1_l[51] ,
         dpath_mulcore_ary1_a1_I1_p1_l[50] ,
         dpath_mulcore_ary1_a1_I1_p1_l[49] ,
         dpath_mulcore_ary1_a1_I1_p1_l[48] ,
         dpath_mulcore_ary1_a1_I1_p1_l[47] ,
         dpath_mulcore_ary1_a1_I1_p1_l[46] ,
         dpath_mulcore_ary1_a1_I1_p1_l[45] ,
         dpath_mulcore_ary1_a1_I1_p1_l[44] ,
         dpath_mulcore_ary1_a1_I1_p1_l[43] ,
         dpath_mulcore_ary1_a1_I1_p1_l[42] ,
         dpath_mulcore_ary1_a1_I1_p1_l[41] ,
         dpath_mulcore_ary1_a1_I1_p1_l[40] ,
         dpath_mulcore_ary1_a1_I1_p1_l[39] ,
         dpath_mulcore_ary1_a1_I1_p1_l[38] ,
         dpath_mulcore_ary1_a1_I1_p1_l[37] ,
         dpath_mulcore_ary1_a1_I1_p1_l[36] ,
         dpath_mulcore_ary1_a1_I1_p1_l[35] ,
         dpath_mulcore_ary1_a1_I1_p1_l[34] ,
         dpath_mulcore_ary1_a1_I1_p1_l[33] ,
         dpath_mulcore_ary1_a1_I1_p1_l[32] ,
         dpath_mulcore_ary1_a1_I1_p1_l[31] ,
         dpath_mulcore_ary1_a1_I1_p1_l[30] ,
         dpath_mulcore_ary1_a1_I1_p1_l[29] ,
         dpath_mulcore_ary1_a1_I1_p1_l[28] ,
         dpath_mulcore_ary1_a1_I1_p1_l[27] ,
         dpath_mulcore_ary1_a1_I1_p1_l[26] ,
         dpath_mulcore_ary1_a1_I1_p1_l[25] ,
         dpath_mulcore_ary1_a1_I1_p1_l[24] ,
         dpath_mulcore_ary1_a1_I1_p1_l[23] ,
         dpath_mulcore_ary1_a1_I1_p1_l[22] ,
         dpath_mulcore_ary1_a1_I1_p1_l[21] ,
         dpath_mulcore_ary1_a1_I1_p1_l[20] ,
         dpath_mulcore_ary1_a1_I1_p1_l[19] ,
         dpath_mulcore_ary1_a1_I1_p1_l[18] ,
         dpath_mulcore_ary1_a1_I1_p1_l[17] ,
         dpath_mulcore_ary1_a1_I1_p1_l[16] ,
         dpath_mulcore_ary1_a1_I1_p1_l[15] ,
         dpath_mulcore_ary1_a1_I1_p1_l[14] ,
         dpath_mulcore_ary1_a1_I1_p1_l[13] ,
         dpath_mulcore_ary1_a1_I1_p1_l[12] ,
         dpath_mulcore_ary1_a1_I1_p1_l[11] ,
         dpath_mulcore_ary1_a1_I1_p1_l[10] ,
         dpath_mulcore_ary1_a1_I1_p1_l[9] ,
         dpath_mulcore_ary1_a1_I1_p1_l[8] ,
         dpath_mulcore_ary1_a1_I1_p1_l[7] ,
         dpath_mulcore_ary1_a1_I1_p1_l[6] ,
         dpath_mulcore_ary1_a1_I1_p1_l[5] ,
         dpath_mulcore_ary1_a1_I1_p1_l[4] ,
         dpath_mulcore_ary1_a1_I1_p1_l[3] ,
         dpath_mulcore_ary1_a1_I1_p2_l[63] ,
         dpath_mulcore_ary1_a1_I1_p2_l[62] ,
         dpath_mulcore_ary1_a1_I1_p2_l[61] ,
         dpath_mulcore_ary1_a1_I1_p2_l[60] ,
         dpath_mulcore_ary1_a1_I1_p2_l[59] ,
         dpath_mulcore_ary1_a1_I1_p2_l[58] ,
         dpath_mulcore_ary1_a1_I1_p2_l[57] ,
         dpath_mulcore_ary1_a1_I1_p2_l[56] ,
         dpath_mulcore_ary1_a1_I1_p2_l[55] ,
         dpath_mulcore_ary1_a1_I1_p2_l[54] ,
         dpath_mulcore_ary1_a1_I1_p2_l[53] ,
         dpath_mulcore_ary1_a1_I1_p2_l[52] ,
         dpath_mulcore_ary1_a1_I1_p2_l[51] ,
         dpath_mulcore_ary1_a1_I1_p2_l[50] ,
         dpath_mulcore_ary1_a1_I1_p2_l[49] ,
         dpath_mulcore_ary1_a1_I1_p2_l[48] ,
         dpath_mulcore_ary1_a1_I1_p2_l[47] ,
         dpath_mulcore_ary1_a1_I1_p2_l[46] ,
         dpath_mulcore_ary1_a1_I1_p2_l[45] ,
         dpath_mulcore_ary1_a1_I1_p2_l[44] ,
         dpath_mulcore_ary1_a1_I1_p2_l[43] ,
         dpath_mulcore_ary1_a1_I1_p2_l[42] ,
         dpath_mulcore_ary1_a1_I1_p2_l[41] ,
         dpath_mulcore_ary1_a1_I1_p2_l[40] ,
         dpath_mulcore_ary1_a1_I1_p2_l[39] ,
         dpath_mulcore_ary1_a1_I1_p2_l[38] ,
         dpath_mulcore_ary1_a1_I1_p2_l[37] ,
         dpath_mulcore_ary1_a1_I1_p2_l[36] ,
         dpath_mulcore_ary1_a1_I1_p2_l[35] ,
         dpath_mulcore_ary1_a1_I1_p2_l[34] ,
         dpath_mulcore_ary1_a1_I1_p2_l[33] ,
         dpath_mulcore_ary1_a1_I1_p2_l[32] ,
         dpath_mulcore_ary1_a1_I1_p2_l[31] ,
         dpath_mulcore_ary1_a1_I1_p2_l[30] ,
         dpath_mulcore_ary1_a1_I1_p2_l[29] ,
         dpath_mulcore_ary1_a1_I1_p2_l[28] ,
         dpath_mulcore_ary1_a1_I1_p2_l[27] ,
         dpath_mulcore_ary1_a1_I1_p2_l[26] ,
         dpath_mulcore_ary1_a1_I1_p2_l[25] ,
         dpath_mulcore_ary1_a1_I1_p2_l[24] ,
         dpath_mulcore_ary1_a1_I1_p2_l[23] ,
         dpath_mulcore_ary1_a1_I1_p2_l[22] ,
         dpath_mulcore_ary1_a1_I1_p2_l[21] ,
         dpath_mulcore_ary1_a1_I1_p2_l[20] ,
         dpath_mulcore_ary1_a1_I1_p2_l[19] ,
         dpath_mulcore_ary1_a1_I1_p2_l[18] ,
         dpath_mulcore_ary1_a1_I1_p2_l[17] ,
         dpath_mulcore_ary1_a1_I1_p2_l[16] ,
         dpath_mulcore_ary1_a1_I1_p2_l[15] ,
         dpath_mulcore_ary1_a1_I1_p2_l[14] ,
         dpath_mulcore_ary1_a1_I1_p2_l[13] ,
         dpath_mulcore_ary1_a1_I1_p2_l[12] ,
         dpath_mulcore_ary1_a1_I1_p2_l[11] ,
         dpath_mulcore_ary1_a1_I1_p2_l[10] ,
         dpath_mulcore_ary1_a1_I1_p2_l[9] ,
         dpath_mulcore_ary1_a1_I1_p2_l[8] ,
         dpath_mulcore_ary1_a1_I1_p2_l[7] ,
         dpath_mulcore_ary1_a1_I1_p2_l[6] ,
         dpath_mulcore_ary1_a1_I1_p2_l[5] ,
         dpath_mulcore_ary1_a1_I1_p2_l[4] ,
         dpath_mulcore_ary1_a1_I2_p0_l[63] ,
         dpath_mulcore_ary1_a1_I2_p0_l[62] ,
         dpath_mulcore_ary1_a1_I2_p0_l[61] ,
         dpath_mulcore_ary1_a1_I2_p0_l[60] ,
         dpath_mulcore_ary1_a1_I2_p0_l[59] ,
         dpath_mulcore_ary1_a1_I2_p0_l[58] ,
         dpath_mulcore_ary1_a1_I2_p0_l[57] ,
         dpath_mulcore_ary1_a1_I2_p0_l[56] ,
         dpath_mulcore_ary1_a1_I2_p0_l[55] ,
         dpath_mulcore_ary1_a1_I2_p0_l[54] ,
         dpath_mulcore_ary1_a1_I2_p0_l[53] ,
         dpath_mulcore_ary1_a1_I2_p0_l[52] ,
         dpath_mulcore_ary1_a1_I2_p0_l[51] ,
         dpath_mulcore_ary1_a1_I2_p0_l[50] ,
         dpath_mulcore_ary1_a1_I2_p0_l[49] ,
         dpath_mulcore_ary1_a1_I2_p0_l[48] ,
         dpath_mulcore_ary1_a1_I2_p0_l[47] ,
         dpath_mulcore_ary1_a1_I2_p0_l[46] ,
         dpath_mulcore_ary1_a1_I2_p0_l[45] ,
         dpath_mulcore_ary1_a1_I2_p0_l[44] ,
         dpath_mulcore_ary1_a1_I2_p0_l[43] ,
         dpath_mulcore_ary1_a1_I2_p0_l[42] ,
         dpath_mulcore_ary1_a1_I2_p0_l[41] ,
         dpath_mulcore_ary1_a1_I2_p0_l[40] ,
         dpath_mulcore_ary1_a1_I2_p0_l[39] ,
         dpath_mulcore_ary1_a1_I2_p0_l[38] ,
         dpath_mulcore_ary1_a1_I2_p0_l[37] ,
         dpath_mulcore_ary1_a1_I2_p0_l[36] ,
         dpath_mulcore_ary1_a1_I2_p0_l[35] ,
         dpath_mulcore_ary1_a1_I2_p0_l[34] ,
         dpath_mulcore_ary1_a1_I2_p0_l[33] ,
         dpath_mulcore_ary1_a1_I2_p0_l[32] ,
         dpath_mulcore_ary1_a1_I2_p0_l[31] ,
         dpath_mulcore_ary1_a1_I2_p0_l[30] ,
         dpath_mulcore_ary1_a1_I2_p0_l[29] ,
         dpath_mulcore_ary1_a1_I2_p0_l[28] ,
         dpath_mulcore_ary1_a1_I2_p0_l[27] ,
         dpath_mulcore_ary1_a1_I2_p0_l[26] ,
         dpath_mulcore_ary1_a1_I2_p0_l[25] ,
         dpath_mulcore_ary1_a1_I2_p0_l[24] ,
         dpath_mulcore_ary1_a1_I2_p0_l[23] ,
         dpath_mulcore_ary1_a1_I2_p0_l[22] ,
         dpath_mulcore_ary1_a1_I2_p0_l[21] ,
         dpath_mulcore_ary1_a1_I2_p0_l[20] ,
         dpath_mulcore_ary1_a1_I2_p0_l[19] ,
         dpath_mulcore_ary1_a1_I2_p0_l[18] ,
         dpath_mulcore_ary1_a1_I2_p0_l[17] ,
         dpath_mulcore_ary1_a1_I2_p0_l[16] ,
         dpath_mulcore_ary1_a1_I2_p0_l[15] ,
         dpath_mulcore_ary1_a1_I2_p0_l[14] ,
         dpath_mulcore_ary1_a1_I2_p0_l[13] ,
         dpath_mulcore_ary1_a1_I2_p0_l[12] ,
         dpath_mulcore_ary1_a1_I2_p0_l[11] ,
         dpath_mulcore_ary1_a1_I2_p0_l[10] ,
         dpath_mulcore_ary1_a1_I2_p0_l[9] ,
         dpath_mulcore_ary1_a1_I2_p0_l[8] ,
         dpath_mulcore_ary1_a1_I2_p0_l[7] ,
         dpath_mulcore_ary1_a1_I2_p0_l[6] ,
         dpath_mulcore_ary1_a1_I2_p0_l[5] ,
         dpath_mulcore_ary1_a1_I2_p0_l[4] ,
         dpath_mulcore_ary1_a1_I2_p0_l[3] ,
         dpath_mulcore_ary1_a1_I2_p1_l[63] ,
         dpath_mulcore_ary1_a1_I2_p1_l[62] ,
         dpath_mulcore_ary1_a1_I2_p1_l[61] ,
         dpath_mulcore_ary1_a1_I2_p1_l[60] ,
         dpath_mulcore_ary1_a1_I2_p1_l[59] ,
         dpath_mulcore_ary1_a1_I2_p1_l[58] ,
         dpath_mulcore_ary1_a1_I2_p1_l[57] ,
         dpath_mulcore_ary1_a1_I2_p1_l[56] ,
         dpath_mulcore_ary1_a1_I2_p1_l[55] ,
         dpath_mulcore_ary1_a1_I2_p1_l[54] ,
         dpath_mulcore_ary1_a1_I2_p1_l[53] ,
         dpath_mulcore_ary1_a1_I2_p1_l[52] ,
         dpath_mulcore_ary1_a1_I2_p1_l[51] ,
         dpath_mulcore_ary1_a1_I2_p1_l[50] ,
         dpath_mulcore_ary1_a1_I2_p1_l[49] ,
         dpath_mulcore_ary1_a1_I2_p1_l[48] ,
         dpath_mulcore_ary1_a1_I2_p1_l[47] ,
         dpath_mulcore_ary1_a1_I2_p1_l[46] ,
         dpath_mulcore_ary1_a1_I2_p1_l[45] ,
         dpath_mulcore_ary1_a1_I2_p1_l[44] ,
         dpath_mulcore_ary1_a1_I2_p1_l[43] ,
         dpath_mulcore_ary1_a1_I2_p1_l[42] ,
         dpath_mulcore_ary1_a1_I2_p1_l[41] ,
         dpath_mulcore_ary1_a1_I2_p1_l[40] ,
         dpath_mulcore_ary1_a1_I2_p1_l[39] ,
         dpath_mulcore_ary1_a1_I2_p1_l[38] ,
         dpath_mulcore_ary1_a1_I2_p1_l[37] ,
         dpath_mulcore_ary1_a1_I2_p1_l[36] ,
         dpath_mulcore_ary1_a1_I2_p1_l[35] ,
         dpath_mulcore_ary1_a1_I2_p1_l[34] ,
         dpath_mulcore_ary1_a1_I2_p1_l[33] ,
         dpath_mulcore_ary1_a1_I2_p1_l[32] ,
         dpath_mulcore_ary1_a1_I2_p1_l[31] ,
         dpath_mulcore_ary1_a1_I2_p1_l[30] ,
         dpath_mulcore_ary1_a1_I2_p1_l[29] ,
         dpath_mulcore_ary1_a1_I2_p1_l[28] ,
         dpath_mulcore_ary1_a1_I2_p1_l[27] ,
         dpath_mulcore_ary1_a1_I2_p1_l[26] ,
         dpath_mulcore_ary1_a1_I2_p1_l[25] ,
         dpath_mulcore_ary1_a1_I2_p1_l[24] ,
         dpath_mulcore_ary1_a1_I2_p1_l[23] ,
         dpath_mulcore_ary1_a1_I2_p1_l[22] ,
         dpath_mulcore_ary1_a1_I2_p1_l[21] ,
         dpath_mulcore_ary1_a1_I2_p1_l[20] ,
         dpath_mulcore_ary1_a1_I2_p1_l[19] ,
         dpath_mulcore_ary1_a1_I2_p1_l[18] ,
         dpath_mulcore_ary1_a1_I2_p1_l[17] ,
         dpath_mulcore_ary1_a1_I2_p1_l[16] ,
         dpath_mulcore_ary1_a1_I2_p1_l[15] ,
         dpath_mulcore_ary1_a1_I2_p1_l[14] ,
         dpath_mulcore_ary1_a1_I2_p1_l[13] ,
         dpath_mulcore_ary1_a1_I2_p1_l[12] ,
         dpath_mulcore_ary1_a1_I2_p1_l[11] ,
         dpath_mulcore_ary1_a1_I2_p1_l[10] ,
         dpath_mulcore_ary1_a1_I2_p1_l[9] ,
         dpath_mulcore_ary1_a1_I2_p1_l[8] ,
         dpath_mulcore_ary1_a1_I2_p1_l[7] ,
         dpath_mulcore_ary1_a1_I2_p1_l[6] ,
         dpath_mulcore_ary1_a1_I2_p1_l[5] ,
         dpath_mulcore_ary1_a1_I2_p1_l[4] ,
         dpath_mulcore_ary1_a1_I2_p1_l[3] ,
         dpath_mulcore_ary1_a1_I2_p2_l[63] ,
         dpath_mulcore_ary1_a1_I2_p2_l[62] ,
         dpath_mulcore_ary1_a1_I2_p2_l[61] ,
         dpath_mulcore_ary1_a1_I2_p2_l[60] ,
         dpath_mulcore_ary1_a1_I2_p2_l[59] ,
         dpath_mulcore_ary1_a1_I2_p2_l[58] ,
         dpath_mulcore_ary1_a1_I2_p2_l[57] ,
         dpath_mulcore_ary1_a1_I2_p2_l[56] ,
         dpath_mulcore_ary1_a1_I2_p2_l[55] ,
         dpath_mulcore_ary1_a1_I2_p2_l[54] ,
         dpath_mulcore_ary1_a1_I2_p2_l[53] ,
         dpath_mulcore_ary1_a1_I2_p2_l[52] ,
         dpath_mulcore_ary1_a1_I2_p2_l[51] ,
         dpath_mulcore_ary1_a1_I2_p2_l[50] ,
         dpath_mulcore_ary1_a1_I2_p2_l[49] ,
         dpath_mulcore_ary1_a1_I2_p2_l[48] ,
         dpath_mulcore_ary1_a1_I2_p2_l[47] ,
         dpath_mulcore_ary1_a1_I2_p2_l[46] ,
         dpath_mulcore_ary1_a1_I2_p2_l[45] ,
         dpath_mulcore_ary1_a1_I2_p2_l[44] ,
         dpath_mulcore_ary1_a1_I2_p2_l[43] ,
         dpath_mulcore_ary1_a1_I2_p2_l[42] ,
         dpath_mulcore_ary1_a1_I2_p2_l[41] ,
         dpath_mulcore_ary1_a1_I2_p2_l[40] ,
         dpath_mulcore_ary1_a1_I2_p2_l[39] ,
         dpath_mulcore_ary1_a1_I2_p2_l[38] ,
         dpath_mulcore_ary1_a1_I2_p2_l[37] ,
         dpath_mulcore_ary1_a1_I2_p2_l[36] ,
         dpath_mulcore_ary1_a1_I2_p2_l[35] ,
         dpath_mulcore_ary1_a1_I2_p2_l[34] ,
         dpath_mulcore_ary1_a1_I2_p2_l[33] ,
         dpath_mulcore_ary1_a1_I2_p2_l[32] ,
         dpath_mulcore_ary1_a1_I2_p2_l[31] ,
         dpath_mulcore_ary1_a1_I2_p2_l[30] ,
         dpath_mulcore_ary1_a1_I2_p2_l[29] ,
         dpath_mulcore_ary1_a1_I2_p2_l[28] ,
         dpath_mulcore_ary1_a1_I2_p2_l[27] ,
         dpath_mulcore_ary1_a1_I2_p2_l[26] ,
         dpath_mulcore_ary1_a1_I2_p2_l[25] ,
         dpath_mulcore_ary1_a1_I2_p2_l[24] ,
         dpath_mulcore_ary1_a1_I2_p2_l[23] ,
         dpath_mulcore_ary1_a1_I2_p2_l[22] ,
         dpath_mulcore_ary1_a1_I2_p2_l[21] ,
         dpath_mulcore_ary1_a1_I2_p2_l[20] ,
         dpath_mulcore_ary1_a1_I2_p2_l[19] ,
         dpath_mulcore_ary1_a1_I2_p2_l[18] ,
         dpath_mulcore_ary1_a1_I2_p2_l[17] ,
         dpath_mulcore_ary1_a1_I2_p2_l[16] ,
         dpath_mulcore_ary1_a1_I2_p2_l[15] ,
         dpath_mulcore_ary1_a1_I2_p2_l[14] ,
         dpath_mulcore_ary1_a1_I2_p2_l[13] ,
         dpath_mulcore_ary1_a1_I2_p2_l[12] ,
         dpath_mulcore_ary1_a1_I2_p2_l[11] ,
         dpath_mulcore_ary1_a1_I2_p2_l[10] ,
         dpath_mulcore_ary1_a1_I2_p2_l[9] ,
         dpath_mulcore_ary1_a1_I2_p2_l[8] ,
         dpath_mulcore_ary1_a1_I2_p2_l[7] ,
         dpath_mulcore_ary1_a1_I2_p2_l[6] ,
         dpath_mulcore_ary1_a1_I2_p2_l[5] ,
         dpath_mulcore_ary1_a1_I2_p2_l[4] ,
         dpath_mulcore_ary1_a0_I0_p0_l[63] ,
         dpath_mulcore_ary1_a0_I0_p0_l[62] ,
         dpath_mulcore_ary1_a0_I0_p0_l[61] ,
         dpath_mulcore_ary1_a0_I0_p0_l[60] ,
         dpath_mulcore_ary1_a0_I0_p0_l[59] ,
         dpath_mulcore_ary1_a0_I0_p0_l[58] ,
         dpath_mulcore_ary1_a0_I0_p0_l[57] ,
         dpath_mulcore_ary1_a0_I0_p0_l[56] ,
         dpath_mulcore_ary1_a0_I0_p0_l[55] ,
         dpath_mulcore_ary1_a0_I0_p0_l[54] ,
         dpath_mulcore_ary1_a0_I0_p0_l[53] ,
         dpath_mulcore_ary1_a0_I0_p0_l[52] ,
         dpath_mulcore_ary1_a0_I0_p0_l[51] ,
         dpath_mulcore_ary1_a0_I0_p0_l[50] ,
         dpath_mulcore_ary1_a0_I0_p0_l[49] ,
         dpath_mulcore_ary1_a0_I0_p0_l[48] ,
         dpath_mulcore_ary1_a0_I0_p0_l[47] ,
         dpath_mulcore_ary1_a0_I0_p0_l[46] ,
         dpath_mulcore_ary1_a0_I0_p0_l[45] ,
         dpath_mulcore_ary1_a0_I0_p0_l[44] ,
         dpath_mulcore_ary1_a0_I0_p0_l[43] ,
         dpath_mulcore_ary1_a0_I0_p0_l[42] ,
         dpath_mulcore_ary1_a0_I0_p0_l[41] ,
         dpath_mulcore_ary1_a0_I0_p0_l[40] ,
         dpath_mulcore_ary1_a0_I0_p0_l[39] ,
         dpath_mulcore_ary1_a0_I0_p0_l[38] ,
         dpath_mulcore_ary1_a0_I0_p0_l[37] ,
         dpath_mulcore_ary1_a0_I0_p0_l[36] ,
         dpath_mulcore_ary1_a0_I0_p0_l[35] ,
         dpath_mulcore_ary1_a0_I0_p0_l[34] ,
         dpath_mulcore_ary1_a0_I0_p0_l[33] ,
         dpath_mulcore_ary1_a0_I0_p0_l[32] ,
         dpath_mulcore_ary1_a0_I0_p0_l[31] ,
         dpath_mulcore_ary1_a0_I0_p0_l[30] ,
         dpath_mulcore_ary1_a0_I0_p0_l[29] ,
         dpath_mulcore_ary1_a0_I0_p0_l[28] ,
         dpath_mulcore_ary1_a0_I0_p0_l[27] ,
         dpath_mulcore_ary1_a0_I0_p0_l[26] ,
         dpath_mulcore_ary1_a0_I0_p0_l[25] ,
         dpath_mulcore_ary1_a0_I0_p0_l[24] ,
         dpath_mulcore_ary1_a0_I0_p0_l[23] ,
         dpath_mulcore_ary1_a0_I0_p0_l[22] ,
         dpath_mulcore_ary1_a0_I0_p0_l[21] ,
         dpath_mulcore_ary1_a0_I0_p0_l[20] ,
         dpath_mulcore_ary1_a0_I0_p0_l[19] ,
         dpath_mulcore_ary1_a0_I0_p0_l[18] ,
         dpath_mulcore_ary1_a0_I0_p0_l[17] ,
         dpath_mulcore_ary1_a0_I0_p0_l[16] ,
         dpath_mulcore_ary1_a0_I0_p0_l[15] ,
         dpath_mulcore_ary1_a0_I0_p0_l[14] ,
         dpath_mulcore_ary1_a0_I0_p0_l[13] ,
         dpath_mulcore_ary1_a0_I0_p0_l[12] ,
         dpath_mulcore_ary1_a0_I0_p0_l[11] ,
         dpath_mulcore_ary1_a0_I0_p0_l[10] ,
         dpath_mulcore_ary1_a0_I0_p0_l[9] ,
         dpath_mulcore_ary1_a0_I0_p0_l[8] ,
         dpath_mulcore_ary1_a0_I0_p0_l[7] ,
         dpath_mulcore_ary1_a0_I0_p0_l[6] ,
         dpath_mulcore_ary1_a0_I0_p0_l[5] ,
         dpath_mulcore_ary1_a0_I0_p0_l[4] ,
         dpath_mulcore_ary1_a0_I0_p0_l[3] ,
         dpath_mulcore_ary1_a0_I0_p1_l[63] ,
         dpath_mulcore_ary1_a0_I0_p1_l[62] ,
         dpath_mulcore_ary1_a0_I0_p1_l[61] ,
         dpath_mulcore_ary1_a0_I0_p1_l[60] ,
         dpath_mulcore_ary1_a0_I0_p1_l[59] ,
         dpath_mulcore_ary1_a0_I0_p1_l[58] ,
         dpath_mulcore_ary1_a0_I0_p1_l[57] ,
         dpath_mulcore_ary1_a0_I0_p1_l[56] ,
         dpath_mulcore_ary1_a0_I0_p1_l[55] ,
         dpath_mulcore_ary1_a0_I0_p1_l[54] ,
         dpath_mulcore_ary1_a0_I0_p1_l[53] ,
         dpath_mulcore_ary1_a0_I0_p1_l[52] ,
         dpath_mulcore_ary1_a0_I0_p1_l[51] ,
         dpath_mulcore_ary1_a0_I0_p1_l[50] ,
         dpath_mulcore_ary1_a0_I0_p1_l[49] ,
         dpath_mulcore_ary1_a0_I0_p1_l[48] ,
         dpath_mulcore_ary1_a0_I0_p1_l[47] ,
         dpath_mulcore_ary1_a0_I0_p1_l[46] ,
         dpath_mulcore_ary1_a0_I0_p1_l[45] ,
         dpath_mulcore_ary1_a0_I0_p1_l[44] ,
         dpath_mulcore_ary1_a0_I0_p1_l[43] ,
         dpath_mulcore_ary1_a0_I0_p1_l[42] ,
         dpath_mulcore_ary1_a0_I0_p1_l[41] ,
         dpath_mulcore_ary1_a0_I0_p1_l[40] ,
         dpath_mulcore_ary1_a0_I0_p1_l[39] ,
         dpath_mulcore_ary1_a0_I0_p1_l[38] ,
         dpath_mulcore_ary1_a0_I0_p1_l[37] ,
         dpath_mulcore_ary1_a0_I0_p1_l[36] ,
         dpath_mulcore_ary1_a0_I0_p1_l[35] ,
         dpath_mulcore_ary1_a0_I0_p1_l[34] ,
         dpath_mulcore_ary1_a0_I0_p1_l[33] ,
         dpath_mulcore_ary1_a0_I0_p1_l[32] ,
         dpath_mulcore_ary1_a0_I0_p1_l[31] ,
         dpath_mulcore_ary1_a0_I0_p1_l[30] ,
         dpath_mulcore_ary1_a0_I0_p1_l[29] ,
         dpath_mulcore_ary1_a0_I0_p1_l[28] ,
         dpath_mulcore_ary1_a0_I0_p1_l[27] ,
         dpath_mulcore_ary1_a0_I0_p1_l[26] ,
         dpath_mulcore_ary1_a0_I0_p1_l[25] ,
         dpath_mulcore_ary1_a0_I0_p1_l[24] ,
         dpath_mulcore_ary1_a0_I0_p1_l[23] ,
         dpath_mulcore_ary1_a0_I0_p1_l[22] ,
         dpath_mulcore_ary1_a0_I0_p1_l[21] ,
         dpath_mulcore_ary1_a0_I0_p1_l[20] ,
         dpath_mulcore_ary1_a0_I0_p1_l[19] ,
         dpath_mulcore_ary1_a0_I0_p1_l[18] ,
         dpath_mulcore_ary1_a0_I0_p1_l[17] ,
         dpath_mulcore_ary1_a0_I0_p1_l[16] ,
         dpath_mulcore_ary1_a0_I0_p1_l[15] ,
         dpath_mulcore_ary1_a0_I0_p1_l[14] ,
         dpath_mulcore_ary1_a0_I0_p1_l[13] ,
         dpath_mulcore_ary1_a0_I0_p1_l[12] ,
         dpath_mulcore_ary1_a0_I0_p1_l[11] ,
         dpath_mulcore_ary1_a0_I0_p1_l[10] ,
         dpath_mulcore_ary1_a0_I0_p1_l[9] ,
         dpath_mulcore_ary1_a0_I0_p1_l[8] ,
         dpath_mulcore_ary1_a0_I0_p1_l[7] ,
         dpath_mulcore_ary1_a0_I0_p1_l[6] ,
         dpath_mulcore_ary1_a0_I0_p1_l[5] ,
         dpath_mulcore_ary1_a0_I0_p1_l[4] ,
         dpath_mulcore_ary1_a0_I0_p1_l[3] ,
         dpath_mulcore_ary1_a0_I0_p2_l[63] ,
         dpath_mulcore_ary1_a0_I0_p2_l[62] ,
         dpath_mulcore_ary1_a0_I0_p2_l[61] ,
         dpath_mulcore_ary1_a0_I0_p2_l[60] ,
         dpath_mulcore_ary1_a0_I0_p2_l[59] ,
         dpath_mulcore_ary1_a0_I0_p2_l[58] ,
         dpath_mulcore_ary1_a0_I0_p2_l[57] ,
         dpath_mulcore_ary1_a0_I0_p2_l[56] ,
         dpath_mulcore_ary1_a0_I0_p2_l[55] ,
         dpath_mulcore_ary1_a0_I0_p2_l[54] ,
         dpath_mulcore_ary1_a0_I0_p2_l[53] ,
         dpath_mulcore_ary1_a0_I0_p2_l[52] ,
         dpath_mulcore_ary1_a0_I0_p2_l[51] ,
         dpath_mulcore_ary1_a0_I0_p2_l[50] ,
         dpath_mulcore_ary1_a0_I0_p2_l[49] ,
         dpath_mulcore_ary1_a0_I0_p2_l[48] ,
         dpath_mulcore_ary1_a0_I0_p2_l[47] ,
         dpath_mulcore_ary1_a0_I0_p2_l[46] ,
         dpath_mulcore_ary1_a0_I0_p2_l[45] ,
         dpath_mulcore_ary1_a0_I0_p2_l[44] ,
         dpath_mulcore_ary1_a0_I0_p2_l[43] ,
         dpath_mulcore_ary1_a0_I0_p2_l[42] ,
         dpath_mulcore_ary1_a0_I0_p2_l[41] ,
         dpath_mulcore_ary1_a0_I0_p2_l[40] ,
         dpath_mulcore_ary1_a0_I0_p2_l[39] ,
         dpath_mulcore_ary1_a0_I0_p2_l[38] ,
         dpath_mulcore_ary1_a0_I0_p2_l[37] ,
         dpath_mulcore_ary1_a0_I0_p2_l[36] ,
         dpath_mulcore_ary1_a0_I0_p2_l[35] ,
         dpath_mulcore_ary1_a0_I0_p2_l[34] ,
         dpath_mulcore_ary1_a0_I0_p2_l[33] ,
         dpath_mulcore_ary1_a0_I0_p2_l[32] ,
         dpath_mulcore_ary1_a0_I0_p2_l[31] ,
         dpath_mulcore_ary1_a0_I0_p2_l[30] ,
         dpath_mulcore_ary1_a0_I0_p2_l[29] ,
         dpath_mulcore_ary1_a0_I0_p2_l[28] ,
         dpath_mulcore_ary1_a0_I0_p2_l[27] ,
         dpath_mulcore_ary1_a0_I0_p2_l[26] ,
         dpath_mulcore_ary1_a0_I0_p2_l[25] ,
         dpath_mulcore_ary1_a0_I0_p2_l[24] ,
         dpath_mulcore_ary1_a0_I0_p2_l[23] ,
         dpath_mulcore_ary1_a0_I0_p2_l[22] ,
         dpath_mulcore_ary1_a0_I0_p2_l[21] ,
         dpath_mulcore_ary1_a0_I0_p2_l[20] ,
         dpath_mulcore_ary1_a0_I0_p2_l[19] ,
         dpath_mulcore_ary1_a0_I0_p2_l[18] ,
         dpath_mulcore_ary1_a0_I0_p2_l[17] ,
         dpath_mulcore_ary1_a0_I0_p2_l[16] ,
         dpath_mulcore_ary1_a0_I0_p2_l[15] ,
         dpath_mulcore_ary1_a0_I0_p2_l[14] ,
         dpath_mulcore_ary1_a0_I0_p2_l[13] ,
         dpath_mulcore_ary1_a0_I0_p2_l[12] ,
         dpath_mulcore_ary1_a0_I0_p2_l[11] ,
         dpath_mulcore_ary1_a0_I0_p2_l[10] ,
         dpath_mulcore_ary1_a0_I0_p2_l[9] ,
         dpath_mulcore_ary1_a0_I0_p2_l[8] ,
         dpath_mulcore_ary1_a0_I0_p2_l[7] ,
         dpath_mulcore_ary1_a0_I0_p2_l[6] ,
         dpath_mulcore_ary1_a0_I0_p2_l[5] ,
         dpath_mulcore_ary1_a0_I0_p2_l[4] ,
         dpath_mulcore_ary1_a1_I0_I2_net35 ,
         dpath_mulcore_ary1_a1_I0_I2_net48 ,
         dpath_mulcore_ary1_a1_I0_I2_net43 ,
         dpath_mulcore_ary1_a1_I0_I2_p1_l_64 ,
         dpath_mulcore_ary1_a1_I0_I2_net15 ,
         dpath_mulcore_ary1_a1_I0_I2_p2_l_64 ,
         dpath_mulcore_ary1_a1_I0_I2_net8 ,
         dpath_mulcore_ary1_a1_I0_I2_p2_l_65 ,
         dpath_mulcore_ary1_a1_I0_I2_net078 ,
         dpath_mulcore_ary1_a1_I0_I2_p2_l_66 ,
         dpath_mulcore_ary1_a1_I0_I2_net0118 ,
         dpath_mulcore_ary1_a1_I0_I2_net38 ,
         dpath_mulcore_ary1_a1_I0_I2_p1_l_65 ,
         dpath_mulcore_ary1_a1_I0_I2_net073 ,
         dpath_mulcore_ary1_a1_I0_I2_p2_l_67 ,
         dpath_mulcore_ary1_a1_I0_I2_net47 ,
         dpath_mulcore_ary1_a1_I0_I2_net088 ,
         dpath_mulcore_ary1_a1_I0_I2_net075 ,
         dpath_mulcore_ary1_a1_I1_I2_net35 ,
         dpath_mulcore_ary1_a1_I1_I2_net48 ,
         dpath_mulcore_ary1_a1_I1_I2_net43 ,
         dpath_mulcore_ary1_a1_I1_I2_p1_l_64 ,
         dpath_mulcore_ary1_a1_I1_I2_net15 ,
         dpath_mulcore_ary1_a1_I1_I2_p2_l_64 ,
         dpath_mulcore_ary1_a1_I1_I2_net8 ,
         dpath_mulcore_ary1_a1_I1_I2_p2_l_65 ,
         dpath_mulcore_ary1_a1_I1_I2_net078 ,
         dpath_mulcore_ary1_a1_I1_I2_p2_l_66 ,
         dpath_mulcore_ary1_a1_I1_I2_net0118 ,
         dpath_mulcore_ary1_a1_I1_I2_net38 ,
         dpath_mulcore_ary1_a1_I1_I2_p1_l_65 ,
         dpath_mulcore_ary1_a1_I1_I2_net073 ,
         dpath_mulcore_ary1_a1_I1_I2_p2_l_67 ,
         dpath_mulcore_ary1_a1_I1_I2_net47 ,
         dpath_mulcore_ary1_a1_I1_I2_net088 ,
         dpath_mulcore_ary1_a1_I1_I2_net075 ,
         dpath_mulcore_ary1_a1_I2_I2_net48 ,
         dpath_mulcore_ary1_a1_I2_I2_net43 ,
         dpath_mulcore_ary1_a1_I2_I2_p1_l_64 ,
         dpath_mulcore_ary1_a1_I2_I2_p2_l_64 ,
         dpath_mulcore_ary1_a1_I2_I2_p2_l_65 ,
         dpath_mulcore_ary1_a1_I2_I2_p2_l_66 ,
         dpath_mulcore_ary1_a1_I2_I2_net0118 ,
         dpath_mulcore_ary1_a1_I2_I2_net38 ,
         dpath_mulcore_ary1_a1_I2_I2_p1_l_65 ,
         dpath_mulcore_ary1_a1_I2_I2_p2_l_67 ,
         dpath_mulcore_ary1_a1_I2_I2_net47 ,
         dpath_mulcore_ary1_a1_I2_I2_net088 ,
         dpath_mulcore_ary1_a0_I0_I2_sc1_66__b ,
         dpath_mulcore_ary1_a0_I0_I2_net35 ,
         dpath_mulcore_ary1_a0_I0_I2_net48 ,
         dpath_mulcore_ary1_a0_I0_I2_net43 ,
         dpath_mulcore_ary1_a0_I0_I2_p1_l_64 ,
         dpath_mulcore_ary1_a0_I0_I2_net15 ,
         dpath_mulcore_ary1_a0_I0_I2_p2_l_64 ,
         dpath_mulcore_ary1_a0_I0_I2_net8 ,
         dpath_mulcore_ary1_a0_I0_I2_p2_l_65 ,
         dpath_mulcore_ary1_a0_I0_I2_net078 ,
         dpath_mulcore_ary1_a0_I0_I2_p2_l_66 ,
         dpath_mulcore_ary1_a0_I0_I2_net0118 ,
         dpath_mulcore_ary1_a0_I0_I2_net38 ,
         dpath_mulcore_ary1_a0_I0_I2_p1_l_65 ,
         dpath_mulcore_ary1_a0_I0_I2_net073 ,
         dpath_mulcore_ary1_a0_I0_I2_p2_l_67 ,
         dpath_mulcore_ary1_a0_I0_I2_net47 ,
         dpath_mulcore_ary1_a0_I0_I2_net42 ,
         dpath_mulcore_ary1_a0_I0_I2_net088 ,
         dpath_mulcore_ary1_a0_I0_I2_net075 ,
         dpath_mulcore_ary1_a1_I0_I1_4__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_4__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_5__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_5__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_5__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_6__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_6__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_6__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_7__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_7__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_7__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_8__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_8__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_8__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_9__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_9__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_9__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_10__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_10__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_10__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_11__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_11__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_11__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_12__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_12__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_12__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_13__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_13__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_13__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_14__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_14__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_14__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_15__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_15__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_15__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_16__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_16__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_16__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_17__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_17__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_17__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_18__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_18__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_18__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_19__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_19__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_19__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_20__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_20__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_20__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_21__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_21__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_21__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_22__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_22__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_22__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_23__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_23__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_23__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_24__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_24__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_24__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_25__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_25__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_25__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_26__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_26__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_26__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_27__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_27__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_27__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_28__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_28__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_28__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_29__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_29__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_29__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_30__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_30__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_30__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_31__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_31__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_31__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_32__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_32__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_32__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_33__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_33__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_33__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_34__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_34__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_34__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_35__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_35__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_35__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_36__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_36__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_36__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_37__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_37__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_37__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_38__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_38__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_38__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_39__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_39__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_39__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_40__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_40__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_40__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_41__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_41__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_41__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_42__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_42__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_42__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_43__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_43__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_43__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_44__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_44__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_44__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_45__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_45__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_45__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_46__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_46__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_46__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_47__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_47__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_47__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_48__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_48__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_48__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_49__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_49__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_49__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_50__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_50__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_50__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_51__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_51__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_51__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_52__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_52__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_52__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_53__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_53__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_53__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_54__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_54__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_54__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_55__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_55__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_55__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_56__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_56__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_56__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_57__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_57__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_57__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_58__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_58__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_58__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_59__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_59__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_59__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_60__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_60__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_60__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_61__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_61__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_61__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_62__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_62__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_62__net046 ,
         dpath_mulcore_ary1_a1_I0_I1_63__net043 ,
         dpath_mulcore_ary1_a1_I0_I1_63__net32 ,
         dpath_mulcore_ary1_a1_I0_I1_63__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_4__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_4__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_5__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_5__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_5__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_6__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_6__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_6__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_7__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_7__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_7__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_8__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_8__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_8__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_9__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_9__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_9__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_10__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_10__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_10__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_11__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_11__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_11__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_12__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_12__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_12__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_13__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_13__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_13__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_14__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_14__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_14__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_15__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_15__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_15__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_16__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_16__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_16__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_17__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_17__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_17__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_18__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_18__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_18__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_19__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_19__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_19__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_20__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_20__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_20__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_21__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_21__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_21__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_22__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_22__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_22__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_23__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_23__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_23__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_24__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_24__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_24__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_25__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_25__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_25__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_26__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_26__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_26__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_27__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_27__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_27__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_28__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_28__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_28__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_29__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_29__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_29__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_30__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_30__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_30__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_31__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_31__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_31__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_32__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_32__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_32__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_33__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_33__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_33__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_34__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_34__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_34__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_35__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_35__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_35__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_36__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_36__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_36__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_37__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_37__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_37__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_38__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_38__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_38__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_39__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_39__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_39__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_40__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_40__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_40__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_41__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_41__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_41__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_42__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_42__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_42__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_43__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_43__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_43__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_44__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_44__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_44__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_45__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_45__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_45__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_46__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_46__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_46__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_47__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_47__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_47__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_48__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_48__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_48__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_49__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_49__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_49__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_50__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_50__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_50__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_51__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_51__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_51__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_52__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_52__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_52__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_53__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_53__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_53__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_54__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_54__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_54__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_55__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_55__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_55__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_56__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_56__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_56__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_57__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_57__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_57__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_58__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_58__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_58__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_59__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_59__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_59__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_60__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_60__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_60__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_61__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_61__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_61__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_62__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_62__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_62__net046 ,
         dpath_mulcore_ary1_a1_I1_I1_63__net043 ,
         dpath_mulcore_ary1_a1_I1_I1_63__net32 ,
         dpath_mulcore_ary1_a1_I1_I1_63__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_4__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_4__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_5__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_5__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_6__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_6__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_7__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_7__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_8__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_8__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_9__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_9__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_10__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_10__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_11__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_11__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_12__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_12__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_13__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_13__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_14__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_14__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_15__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_15__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_16__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_16__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_17__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_17__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_18__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_18__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_19__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_19__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_20__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_20__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_21__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_21__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_22__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_22__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_23__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_23__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_24__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_24__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_25__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_25__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_26__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_26__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_27__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_27__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_28__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_28__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_29__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_29__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_30__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_30__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_31__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_31__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_32__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_32__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_33__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_33__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_34__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_34__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_35__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_35__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_36__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_36__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_37__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_37__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_38__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_38__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_39__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_39__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_40__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_40__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_41__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_41__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_42__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_42__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_43__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_43__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_44__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_44__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_45__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_45__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_46__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_46__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_47__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_47__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_48__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_48__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_49__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_49__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_50__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_50__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_51__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_51__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_52__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_52__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_53__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_53__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_54__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_54__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_55__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_55__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_56__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_56__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_57__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_57__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_58__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_58__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_59__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_59__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_60__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_60__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_61__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_61__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_62__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_62__net046 ,
         dpath_mulcore_ary1_a1_I2_I1_63__net32 ,
         dpath_mulcore_ary1_a1_I2_I1_63__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_4__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_4__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_5__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_5__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_5__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_6__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_6__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_6__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_7__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_7__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_7__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_8__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_8__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_8__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_9__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_9__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_9__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_10__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_10__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_10__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_11__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_11__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_11__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_12__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_12__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_12__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_13__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_13__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_13__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_14__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_14__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_14__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_15__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_15__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_15__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_16__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_16__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_16__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_17__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_17__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_17__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_18__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_18__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_18__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_19__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_19__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_19__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_20__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_20__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_20__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_21__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_21__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_21__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_22__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_22__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_22__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_23__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_23__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_23__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_24__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_24__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_24__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_25__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_25__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_25__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_26__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_26__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_26__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_27__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_27__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_27__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_28__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_28__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_28__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_29__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_29__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_29__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_30__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_30__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_30__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_31__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_31__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_31__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_32__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_32__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_32__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_33__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_33__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_33__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_34__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_34__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_34__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_35__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_35__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_35__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_36__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_36__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_36__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_37__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_37__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_37__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_38__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_38__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_38__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_39__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_39__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_39__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_40__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_40__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_40__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_41__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_41__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_41__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_42__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_42__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_42__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_43__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_43__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_43__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_44__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_44__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_44__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_45__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_45__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_45__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_46__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_46__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_46__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_47__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_47__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_47__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_48__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_48__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_48__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_49__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_49__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_49__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_50__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_50__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_50__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_51__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_51__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_51__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_52__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_52__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_52__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_53__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_53__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_53__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_54__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_54__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_54__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_55__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_55__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_55__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_56__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_56__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_56__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_57__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_57__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_57__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_58__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_58__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_58__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_59__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_59__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_59__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_60__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_60__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_60__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_61__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_61__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_61__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_62__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_62__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_62__net046 ,
         dpath_mulcore_ary1_a0_I0_I1_63__net043 ,
         dpath_mulcore_ary1_a0_I0_I1_63__net32 ,
         dpath_mulcore_ary1_a0_I0_I1_63__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_4__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_4__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_5__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_5__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_5__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_6__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_6__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_6__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_7__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_7__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_7__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_8__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_8__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_8__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_9__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_9__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_9__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_10__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_10__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_10__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_11__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_11__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_11__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_12__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_12__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_12__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_13__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_13__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_13__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_14__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_14__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_14__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_15__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_15__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_15__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_16__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_16__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_16__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_17__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_17__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_17__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_18__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_18__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_18__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_19__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_19__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_19__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_20__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_20__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_20__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_21__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_21__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_21__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_22__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_22__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_22__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_23__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_23__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_23__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_24__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_24__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_24__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_25__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_25__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_25__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_26__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_26__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_26__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_27__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_27__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_27__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_28__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_28__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_28__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_29__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_29__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_29__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_30__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_30__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_30__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_31__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_31__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_31__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_32__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_32__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_32__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_33__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_33__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_33__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_34__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_34__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_34__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_35__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_35__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_35__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_36__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_36__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_36__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_37__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_37__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_37__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_38__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_38__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_38__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_39__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_39__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_39__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_40__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_40__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_40__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_41__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_41__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_41__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_42__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_42__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_42__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_43__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_43__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_43__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_44__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_44__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_44__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_45__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_45__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_45__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_46__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_46__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_46__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_47__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_47__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_47__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_48__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_48__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_48__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_49__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_49__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_49__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_50__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_50__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_50__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_51__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_51__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_51__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_52__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_52__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_52__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_53__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_53__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_53__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_54__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_54__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_54__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_55__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_55__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_55__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_56__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_56__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_56__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_57__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_57__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_57__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_58__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_58__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_58__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_59__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_59__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_59__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_60__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_60__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_60__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_61__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_61__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_61__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_62__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_62__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_62__net046 ,
         dpath_mulcore_ary1_a0_I1_I1_63__net043 ,
         dpath_mulcore_ary1_a0_I1_I1_63__net32 ,
         dpath_mulcore_ary1_a0_I1_I1_63__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_4__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_4__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_5__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_5__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_6__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_6__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_7__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_7__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_8__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_8__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_9__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_9__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_10__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_10__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_11__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_11__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_12__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_12__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_13__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_13__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_14__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_14__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_15__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_15__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_16__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_16__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_17__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_17__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_18__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_18__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_19__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_19__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_20__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_20__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_21__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_21__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_22__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_22__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_23__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_23__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_24__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_24__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_25__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_25__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_26__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_26__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_27__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_27__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_28__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_28__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_29__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_29__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_30__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_30__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_31__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_31__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_32__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_32__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_33__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_33__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_34__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_34__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_35__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_35__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_36__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_36__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_37__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_37__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_38__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_38__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_39__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_39__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_40__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_40__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_41__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_41__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_42__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_42__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_43__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_43__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_44__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_44__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_45__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_45__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_46__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_46__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_47__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_47__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_48__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_48__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_49__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_49__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_50__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_50__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_51__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_51__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_52__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_52__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_53__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_53__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_54__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_54__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_55__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_55__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_56__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_56__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_57__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_57__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_58__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_58__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_59__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_59__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_60__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_60__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_61__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_61__net046 ,
         dpath_mulcore_ary1_a0_I2_I1_62__net32 ,
         dpath_mulcore_ary1_a0_I2_I1_62__net046 ,
         dpath_mulcore_ary1_a1_I0_I0_p0_l_0 ,
         dpath_mulcore_ary1_a1_I0_I0_p0_l_1 ,
         dpath_mulcore_ary1_a1_I0_I0_p1_l_2 ,
         dpath_mulcore_ary1_a1_I0_I0_p0_l_2 ,
         dpath_mulcore_ary1_a1_I0_I0_p0_1 ,
         dpath_mulcore_ary1_a1_I0_I0_p1_3 ,
         dpath_mulcore_ary1_a1_I0_I0_p0_3 ,
         dpath_mulcore_ary1_a1_I0_I0_p0_2 ,
         dpath_mulcore_ary1_a1_I0_I0_b1n_0 ,
         dpath_mulcore_ary1_a1_I0_I0_b1n_1 ,
         dpath_mulcore_ary1_a1_I0_I0_b0n ,
         dpath_mulcore_ary1_a1_I0_I0_b0n_0 ,
         dpath_mulcore_ary1_a1_I0_I0_b0n_1 ,
         dpath_mulcore_ary1_a1_I1_I0_p0_l_0 ,
         dpath_mulcore_ary1_a1_I1_I0_p0_l_1 ,
         dpath_mulcore_ary1_a1_I1_I0_p1_l_2 ,
         dpath_mulcore_ary1_a1_I1_I0_p0_l_2 ,
         dpath_mulcore_ary1_a1_I1_I0_p0_1 ,
         dpath_mulcore_ary1_a1_I1_I0_p1_3 ,
         dpath_mulcore_ary1_a1_I1_I0_p0_3 ,
         dpath_mulcore_ary1_a1_I1_I0_p0_2 ,
         dpath_mulcore_ary1_a1_I1_I0_b1n_0 ,
         dpath_mulcore_ary1_a1_I1_I0_b1n_1 ,
         dpath_mulcore_ary1_a1_I1_I0_b0n ,
         dpath_mulcore_ary1_a1_I1_I0_b0n_0 ,
         dpath_mulcore_ary1_a1_I1_I0_b0n_1 ,
         dpath_mulcore_ary1_a1_I2_I0_p0_l_0 ,
         dpath_mulcore_ary1_a1_I2_I0_p0_l_1 ,
         dpath_mulcore_ary1_a1_I2_I0_p1_l_2 ,
         dpath_mulcore_ary1_a1_I2_I0_p0_l_2 ,
         dpath_mulcore_ary1_a1_I2_I0_p0_1 ,
         dpath_mulcore_ary1_a1_I2_I0_p1_3 ,
         dpath_mulcore_ary1_a1_I2_I0_p0_3 ,
         dpath_mulcore_ary1_a1_I2_I0_p0_2 ,
         dpath_mulcore_ary1_a1_I2_I0_b1n_0 ,
         dpath_mulcore_ary1_a1_I2_I0_b1n_1 ,
         dpath_mulcore_ary1_a1_I2_I0_b0n ,
         dpath_mulcore_ary1_a1_I2_I0_b0n_0 ,
         dpath_mulcore_ary1_a1_I2_I0_b0n_1 ,
         dpath_mulcore_ary1_a0_I0_I0_p0_l_0 ,
         dpath_mulcore_ary1_a0_I0_I0_p0_l_1 ,
         dpath_mulcore_ary1_a0_I0_I0_p1_l_2 ,
         dpath_mulcore_ary1_a0_I0_I0_p0_l_2 ,
         dpath_mulcore_ary1_a0_I0_I0_p0_1 ,
         dpath_mulcore_ary1_a0_I0_I0_p1_3 ,
         dpath_mulcore_ary1_a0_I0_I0_p0_3 ,
         dpath_mulcore_ary1_a0_I0_I0_p0_2 ,
         dpath_mulcore_ary1_a0_I0_I0_b1n_0 ,
         dpath_mulcore_ary1_a0_I0_I0_b1n_1 ,
         dpath_mulcore_ary1_a0_I0_I0_b0n ,
         dpath_mulcore_ary1_a0_I0_I0_b0n_0 ,
         dpath_mulcore_ary1_a0_I0_I0_b0n_1 ,
         dpath_mulcore_ary1_a0_I1_I0_p0_l_0 ,
         dpath_mulcore_ary1_a0_I1_I0_p0_l_1 ,
         dpath_mulcore_ary1_a0_I1_I0_p1_l_2 ,
         dpath_mulcore_ary1_a0_I1_I0_p0_l_2 ,
         dpath_mulcore_ary1_a0_I1_I0_p0_1 ,
         dpath_mulcore_ary1_a0_I1_I0_p1_3 ,
         dpath_mulcore_ary1_a0_I1_I0_p0_3 ,
         dpath_mulcore_ary1_a0_I1_I0_p0_2 ,
         dpath_mulcore_ary1_a0_I1_I0_b1n_0 ,
         dpath_mulcore_ary1_a0_I1_I0_b1n_1 ,
         dpath_mulcore_ary1_a0_I1_I0_b0n ,
         dpath_mulcore_ary1_a0_I1_I0_b0n_0 ,
         dpath_mulcore_ary1_a0_I1_I0_b0n_1 , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337;
  assign dpath_mulcore_clk_enb0  = rclk;
DFFSR rstff_q_reg[0] ( .D(rstff_n4 ), .CLK(dpath_mulcore_clk_enb0 ), .R(arst_l), .S(1'b1), .Q(rst_l) );
DFFPOSX1 control_acc_reg_rst_reg(.D(spu_mul_areg_rst), .CLK(dpath_mulcore_clk_enb0), .Q(acc_reg_rst));
DFFPOSX1 control_acc_reg_shf_reg(.D(n3087), .CLK(dpath_mulcore_clk_enb0), .Q(acc_reg_shf));
DFFPOSX1 control_acc_actc5_reg(.D(control_N11), .CLK(dpath_mulcore_clk_enb0), .Q(byp_imm));
DFFPOSX1 control_acc_actc1_reg(.D(control_N6), .CLK(dpath_mulcore_clk_enb0), .Q(control_acc_actc1));
DFFPOSX1 control_mul_spu_ack_d_reg(.D(mul_spu_ack), .CLK(dpath_mulcore_clk_enb0), .Q(control_mul_spu_ack_d));
DFFPOSX1 control_c3_act_reg(.D(control_N4), .CLK(dpath_mulcore_clk_enb0), .Q(control_c3_act));
DFFPOSX1 control_c2_act_reg(.D(control_N3), .CLK(dpath_mulcore_clk_enb0), .Q(control_c2_act));
DFFPOSX1 control_c1_act_reg(.D(control_N2), .CLK(dpath_mulcore_clk_enb0), .Q(control_c1_act));
DFFPOSX1 control_favor_e_reg(.D(control_N5), .CLK(dpath_mulcore_clk_enb0), .Q(control_favor_e));
DFFPOSX1 control_mul_ecl_ack_d_reg(.D(mul_exu_ack), .CLK(dpath_mulcore_clk_enb0), .Q(control_mul_ecl_ack_d));
DFFPOSX1 control_acc_actc4_reg(.D(control_N9), .CLK(dpath_mulcore_clk_enb0), .Q(control_acc_actc4));
DFFPOSX1 control_acc_actc3_reg(.D(control_N8), .CLK(dpath_mulcore_clk_enb0), .Q(acc_actc3));
DFFPOSX1 control_acc_actc2_reg(.D(control_N7), .CLK(dpath_mulcore_clk_enb0), .Q(acc_actc2));
NAND2X1 mul_dpath_U947(.A(n5756), .B(n5135), .Y(mul_data_out[0]));
NAND2X1 mul_dpath_U944(.A(n5755), .B(n5134), .Y(mul_data_out[10]));
NAND2X1 mul_dpath_U941(.A(n5754), .B(n5133), .Y(mul_data_out[11]));
NAND2X1 mul_dpath_U938(.A(n5753), .B(n5132), .Y(mul_data_out[12]));
NAND2X1 mul_dpath_U935(.A(n5752), .B(n5131), .Y(mul_data_out[13]));
NAND2X1 mul_dpath_U932(.A(n5751), .B(n5130), .Y(mul_data_out[14]));
NAND2X1 mul_dpath_U929(.A(n5750), .B(n5129), .Y(mul_data_out[15]));
NAND2X1 mul_dpath_U926(.A(n5749), .B(n5128), .Y(mul_data_out[16]));
NAND2X1 mul_dpath_U923(.A(n5748), .B(n5127), .Y(mul_data_out[17]));
NAND2X1 mul_dpath_U920(.A(n5747), .B(n5126), .Y(mul_data_out[18]));
NAND2X1 mul_dpath_U917(.A(n5746), .B(n5125), .Y(mul_data_out[19]));
NAND2X1 mul_dpath_U914(.A(n5745), .B(n5124), .Y(mul_data_out[1]));
NAND2X1 mul_dpath_U911(.A(n5744), .B(n5123), .Y(mul_data_out[20]));
NAND2X1 mul_dpath_U908(.A(n5743), .B(n5122), .Y(mul_data_out[21]));
NAND2X1 mul_dpath_U905(.A(n5742), .B(n5121), .Y(mul_data_out[22]));
NAND2X1 mul_dpath_U902(.A(n5741), .B(n5120), .Y(mul_data_out[23]));
NAND2X1 mul_dpath_U899(.A(n5740), .B(n5119), .Y(mul_data_out[24]));
NAND2X1 mul_dpath_U896(.A(n5739), .B(n5118), .Y(mul_data_out[25]));
NAND2X1 mul_dpath_U893(.A(n5738), .B(n5117), .Y(mul_data_out[26]));
NAND2X1 mul_dpath_U890(.A(n5737), .B(n5116), .Y(mul_data_out[27]));
NAND2X1 mul_dpath_U887(.A(n5736), .B(n5115), .Y(mul_data_out[28]));
NAND2X1 mul_dpath_U884(.A(n5735), .B(n5114), .Y(mul_data_out[29]));
NAND2X1 mul_dpath_U881(.A(n5734), .B(n5113), .Y(mul_data_out[2]));
NAND2X1 mul_dpath_U878(.A(n5733), .B(n5112), .Y(mul_data_out[30]));
NAND2X1 mul_dpath_U875(.A(n5732), .B(n5111), .Y(mul_data_out[31]));
NAND2X1 mul_dpath_U872(.A(n5731), .B(n5110), .Y(mul_data_out[32]));
NAND2X1 mul_dpath_U869(.A(n5730), .B(n5109), .Y(mul_data_out[33]));
NAND2X1 mul_dpath_U866(.A(n5729), .B(n5108), .Y(mul_data_out[34]));
NAND2X1 mul_dpath_U863(.A(n5728), .B(n5107), .Y(mul_data_out[35]));
NAND2X1 mul_dpath_U860(.A(n5727), .B(n5106), .Y(mul_data_out[36]));
NAND2X1 mul_dpath_U857(.A(n5726), .B(n5105), .Y(mul_data_out[37]));
NAND2X1 mul_dpath_U854(.A(n5725), .B(n5104), .Y(mul_data_out[38]));
NAND2X1 mul_dpath_U851(.A(n5724), .B(n5103), .Y(mul_data_out[39]));
NAND2X1 mul_dpath_U848(.A(n5723), .B(n5102), .Y(mul_data_out[3]));
NAND2X1 mul_dpath_U845(.A(n5722), .B(n5101), .Y(mul_data_out[40]));
NAND2X1 mul_dpath_U842(.A(n5721), .B(n5100), .Y(mul_data_out[41]));
NAND2X1 mul_dpath_U839(.A(n5720), .B(n5099), .Y(mul_data_out[42]));
NAND2X1 mul_dpath_U836(.A(n5719), .B(n5098), .Y(mul_data_out[43]));
NAND2X1 mul_dpath_U833(.A(n5718), .B(n5097), .Y(mul_data_out[44]));
NAND2X1 mul_dpath_U830(.A(n5717), .B(n5096), .Y(mul_data_out[45]));
NAND2X1 mul_dpath_U827(.A(n5716), .B(n5095), .Y(mul_data_out[46]));
NAND2X1 mul_dpath_U824(.A(n5715), .B(n5094), .Y(mul_data_out[47]));
NAND2X1 mul_dpath_U821(.A(n5714), .B(n5093), .Y(mul_data_out[48]));
NAND2X1 mul_dpath_U818(.A(n5713), .B(n5092), .Y(mul_data_out[49]));
NAND2X1 mul_dpath_U815(.A(n5712), .B(n5091), .Y(mul_data_out[4]));
NAND2X1 mul_dpath_U812(.A(n5711), .B(n5090), .Y(mul_data_out[50]));
NAND2X1 mul_dpath_U809(.A(n5710), .B(n5089), .Y(mul_data_out[51]));
NAND2X1 mul_dpath_U806(.A(n5709), .B(n5088), .Y(mul_data_out[52]));
NAND2X1 mul_dpath_U803(.A(n5708), .B(n5087), .Y(mul_data_out[53]));
NAND2X1 mul_dpath_U800(.A(n5707), .B(n5086), .Y(mul_data_out[54]));
NAND2X1 mul_dpath_U797(.A(n5706), .B(n5085), .Y(mul_data_out[55]));
NAND2X1 mul_dpath_U794(.A(n5705), .B(n5084), .Y(mul_data_out[56]));
NAND2X1 mul_dpath_U791(.A(n5704), .B(n5083), .Y(mul_data_out[57]));
NAND2X1 mul_dpath_U788(.A(n5703), .B(n5082), .Y(mul_data_out[58]));
NAND2X1 mul_dpath_U785(.A(n5702), .B(n5081), .Y(mul_data_out[59]));
NAND2X1 mul_dpath_U782(.A(n5701), .B(n5080), .Y(mul_data_out[5]));
NAND2X1 mul_dpath_U779(.A(n5700), .B(n5079), .Y(mul_data_out[60]));
NAND2X1 mul_dpath_U776(.A(n5699), .B(n5078), .Y(mul_data_out[61]));
NAND2X1 mul_dpath_U773(.A(n5698), .B(n5077), .Y(mul_data_out[62]));
NAND2X1 mul_dpath_U770(.A(n5697), .B(n5076), .Y(mul_data_out[63]));
NAND2X1 mul_dpath_U767(.A(n5696), .B(n5075), .Y(mul_data_out[6]));
NAND2X1 mul_dpath_U764(.A(n5695), .B(n5074), .Y(mul_data_out[7]));
NAND2X1 mul_dpath_U761(.A(n5694), .B(n5073), .Y(mul_data_out[8]));
NAND2X1 mul_dpath_U758(.A(n5693), .B(n5072), .Y(mul_data_out[9]));
DFFPOSX1 dpath_dffshf_q_reg[0](.D(dpath_dffshf_n3), .CLK(dpath_mulcore_clk_enb0), .Q(dpath_acc_reg_shf2));
DFFPOSX1 dpath_accum_q_reg[0](.D(dpath_accum_n273), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[0]));
DFFPOSX1 dpath_accum_q_reg[1](.D(dpath_accum_n271), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[1]));
DFFPOSX1 dpath_accum_q_reg[2](.D(dpath_accum_n269), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[2]));
DFFPOSX1 dpath_accum_q_reg[3](.D(dpath_accum_n267), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[3]));
DFFPOSX1 dpath_accum_q_reg[4](.D(dpath_accum_n265), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[4]));
DFFPOSX1 dpath_accum_q_reg[5](.D(dpath_accum_n263), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[5]));
DFFPOSX1 dpath_accum_q_reg[6](.D(dpath_accum_n261), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[6]));
DFFPOSX1 dpath_accum_q_reg[7](.D(dpath_accum_n259), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[7]));
DFFPOSX1 dpath_accum_q_reg[8](.D(dpath_accum_n257), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[8]));
DFFPOSX1 dpath_accum_q_reg[9](.D(dpath_accum_n255), .CLK(n9757), .Q(dpath_acc_reg[9]));
DFFPOSX1 dpath_accum_q_reg[10](.D(dpath_accum_n253), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[10]));
DFFPOSX1 dpath_accum_q_reg[11](.D(dpath_accum_n251), .CLK(n9756), .Q(dpath_acc_reg[11]));
DFFPOSX1 dpath_accum_q_reg[12](.D(dpath_accum_n249), .CLK(n9758), .Q(dpath_acc_reg[12]));
DFFPOSX1 dpath_accum_q_reg[13](.D(dpath_accum_n247), .CLK(n9759), .Q(dpath_acc_reg[13]));
DFFPOSX1 dpath_accum_q_reg[14](.D(dpath_accum_n245), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[14]));
DFFPOSX1 dpath_accum_q_reg[15](.D(dpath_accum_n243), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[15]));
DFFPOSX1 dpath_accum_q_reg[16](.D(dpath_accum_n241), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[16]));
DFFPOSX1 dpath_accum_q_reg[17](.D(dpath_accum_n239), .CLK(n9757), .Q(dpath_acc_reg[17]));
DFFPOSX1 dpath_accum_q_reg[18](.D(dpath_accum_n237), .CLK(n9755), .Q(dpath_acc_reg[18]));
DFFPOSX1 dpath_accum_q_reg[19](.D(dpath_accum_n235), .CLK(n9758), .Q(dpath_acc_reg[19]));
DFFPOSX1 dpath_accum_q_reg[20](.D(dpath_accum_n233), .CLK(n9755), .Q(dpath_acc_reg[20]));
DFFPOSX1 dpath_accum_q_reg[21](.D(dpath_accum_n231), .CLK(n9757), .Q(dpath_acc_reg[21]));
DFFPOSX1 dpath_accum_q_reg[22](.D(dpath_accum_n229), .CLK(n9759), .Q(dpath_acc_reg[22]));
DFFPOSX1 dpath_accum_q_reg[23](.D(dpath_accum_n227), .CLK(n9756), .Q(dpath_acc_reg[23]));
DFFPOSX1 dpath_accum_q_reg[24](.D(dpath_accum_n225), .CLK(n9755), .Q(dpath_acc_reg[24]));
DFFPOSX1 dpath_accum_q_reg[25](.D(dpath_accum_n223), .CLK(n9756), .Q(dpath_acc_reg[25]));
DFFPOSX1 dpath_accum_q_reg[26](.D(dpath_accum_n221), .CLK(n9758), .Q(dpath_acc_reg[26]));
DFFPOSX1 dpath_accum_q_reg[27](.D(dpath_accum_n219), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[27]));
DFFPOSX1 dpath_accum_q_reg[28](.D(dpath_accum_n217), .CLK(n9756), .Q(dpath_acc_reg[28]));
DFFPOSX1 dpath_accum_q_reg[29](.D(dpath_accum_n215), .CLK(n9759), .Q(dpath_acc_reg[29]));
DFFPOSX1 dpath_accum_q_reg[30](.D(dpath_accum_n213), .CLK(n9758), .Q(dpath_acc_reg[30]));
DFFPOSX1 dpath_accum_q_reg[31](.D(dpath_accum_n211), .CLK(n9755), .Q(dpath_acc_reg[31]));
DFFPOSX1 dpath_accum_q_reg[32](.D(dpath_accum_n209), .CLK(n9757), .Q(dpath_acc_reg[32]));
DFFPOSX1 dpath_accum_q_reg[33](.D(dpath_accum_n207), .CLK(n9759), .Q(dpath_acc_reg[33]));
DFFPOSX1 dpath_accum_q_reg[34](.D(dpath_accum_n205), .CLK(n9755), .Q(dpath_acc_reg[34]));
DFFPOSX1 dpath_accum_q_reg[35](.D(dpath_accum_n203), .CLK(n9755), .Q(dpath_acc_reg[35]));
DFFPOSX1 dpath_accum_q_reg[36](.D(dpath_accum_n201), .CLK(n9756), .Q(dpath_acc_reg[36]));
DFFPOSX1 dpath_accum_q_reg[37](.D(dpath_accum_n199), .CLK(n9758), .Q(dpath_acc_reg[37]));
DFFPOSX1 dpath_accum_q_reg[38](.D(dpath_accum_n197), .CLK(n9757), .Q(dpath_acc_reg[38]));
DFFPOSX1 dpath_accum_q_reg[39](.D(dpath_accum_n195), .CLK(n9759), .Q(dpath_acc_reg[39]));
DFFPOSX1 dpath_accum_q_reg[40](.D(dpath_accum_n193), .CLK(n9757), .Q(dpath_acc_reg[40]));
DFFPOSX1 dpath_accum_q_reg[41](.D(dpath_accum_n191), .CLK(n9755), .Q(dpath_acc_reg[41]));
DFFPOSX1 dpath_accum_q_reg[42](.D(dpath_accum_n189), .CLK(n9758), .Q(dpath_acc_reg[42]));
DFFPOSX1 dpath_accum_q_reg[43](.D(dpath_accum_n187), .CLK(n9757), .Q(dpath_acc_reg[43]));
DFFPOSX1 dpath_accum_q_reg[44](.D(dpath_accum_n185), .CLK(n9756), .Q(dpath_acc_reg[44]));
DFFPOSX1 dpath_accum_q_reg[45](.D(dpath_accum_n183), .CLK(n9757), .Q(dpath_acc_reg[45]));
DFFPOSX1 dpath_accum_q_reg[46](.D(dpath_accum_n181), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[46]));
DFFPOSX1 dpath_accum_q_reg[47](.D(dpath_accum_n179), .CLK(n9759), .Q(dpath_acc_reg[47]));
DFFPOSX1 dpath_accum_q_reg[48](.D(dpath_accum_n177), .CLK(n9755), .Q(dpath_acc_reg[48]));
DFFPOSX1 dpath_accum_q_reg[49](.D(dpath_accum_n175), .CLK(n9756), .Q(dpath_acc_reg[49]));
DFFPOSX1 dpath_accum_q_reg[50](.D(dpath_accum_n173), .CLK(n9758), .Q(dpath_acc_reg[50]));
DFFPOSX1 dpath_accum_q_reg[51](.D(dpath_accum_n171), .CLK(n9756), .Q(dpath_acc_reg[51]));
DFFPOSX1 dpath_accum_q_reg[52](.D(dpath_accum_n169), .CLK(n9759), .Q(dpath_acc_reg[52]));
DFFPOSX1 dpath_accum_q_reg[53](.D(dpath_accum_n167), .CLK(n9759), .Q(dpath_acc_reg[53]));
DFFPOSX1 dpath_accum_q_reg[54](.D(dpath_accum_n165), .CLK(n9757), .Q(dpath_acc_reg[54]));
DFFPOSX1 dpath_accum_q_reg[55](.D(dpath_accum_n163), .CLK(dpath_clk_enb1), .Q(dpath_acc_reg[55]));
DFFPOSX1 dpath_accum_q_reg[56](.D(dpath_accum_n161), .CLK(n9758), .Q(dpath_acc_reg[56]));
DFFPOSX1 dpath_accum_q_reg[57](.D(dpath_accum_n159), .CLK(n9759), .Q(dpath_acc_reg[57]));
DFFPOSX1 dpath_accum_q_reg[58](.D(dpath_accum_n157), .CLK(n9759), .Q(dpath_acc_reg[58]));
DFFPOSX1 dpath_accum_q_reg[59](.D(dpath_accum_n155), .CLK(n9759), .Q(dpath_acc_reg[59]));
DFFPOSX1 dpath_accum_q_reg[60](.D(dpath_accum_n153), .CLK(n9759), .Q(dpath_acc_reg[60]));
DFFPOSX1 dpath_accum_q_reg[61](.D(dpath_accum_n151), .CLK(n9759), .Q(dpath_acc_reg[61]));
DFFPOSX1 dpath_accum_q_reg[62](.D(dpath_accum_n149), .CLK(n9759), .Q(dpath_acc_reg[62]));
DFFPOSX1 dpath_accum_q_reg[63](.D(dpath_accum_n147), .CLK(n9759), .Q(dpath_acc_reg[63]));
DFFPOSX1 dpath_accum_q_reg[64](.D(dpath_accum_n145), .CLK(n9759), .Q(dpath_acc_reg[64]));
DFFPOSX1 dpath_accum_q_reg[65](.D(dpath_accum_n143), .CLK(n9759), .Q(dpath_acc_reg[65]));
DFFPOSX1 dpath_accum_q_reg[66](.D(dpath_accum_n141), .CLK(n9759), .Q(dpath_acc_reg[66]));
DFFPOSX1 dpath_accum_q_reg[67](.D(dpath_accum_n139), .CLK(n9759), .Q(dpath_acc_reg[67]));
DFFPOSX1 dpath_accum_q_reg[68](.D(dpath_accum_n137), .CLK(n9759), .Q(dpath_acc_reg[68]));
DFFPOSX1 dpath_accum_q_reg[69](.D(dpath_accum_n135), .CLK(n9759), .Q(dpath_acc_reg[69]));
DFFPOSX1 dpath_accum_q_reg[70](.D(dpath_accum_n133), .CLK(n9759), .Q(dpath_acc_reg[70]));
DFFPOSX1 dpath_accum_q_reg[71](.D(dpath_accum_n131), .CLK(n9758), .Q(dpath_acc_reg[71]));
DFFPOSX1 dpath_accum_q_reg[72](.D(dpath_accum_n129), .CLK(n9758), .Q(dpath_acc_reg[72]));
DFFPOSX1 dpath_accum_q_reg[73](.D(dpath_accum_n127), .CLK(n9758), .Q(dpath_acc_reg[73]));
DFFPOSX1 dpath_accum_q_reg[74](.D(dpath_accum_n125), .CLK(n9758), .Q(dpath_acc_reg[74]));
DFFPOSX1 dpath_accum_q_reg[75](.D(dpath_accum_n123), .CLK(n9758), .Q(dpath_acc_reg[75]));
DFFPOSX1 dpath_accum_q_reg[76](.D(dpath_accum_n121), .CLK(n9758), .Q(dpath_acc_reg[76]));
DFFPOSX1 dpath_accum_q_reg[77](.D(dpath_accum_n119), .CLK(n9758), .Q(dpath_acc_reg[77]));
DFFPOSX1 dpath_accum_q_reg[78](.D(dpath_accum_n117), .CLK(n9758), .Q(dpath_acc_reg[78]));
DFFPOSX1 dpath_accum_q_reg[79](.D(dpath_accum_n115), .CLK(n9758), .Q(dpath_acc_reg[79]));
DFFPOSX1 dpath_accum_q_reg[80](.D(dpath_accum_n113), .CLK(n9758), .Q(dpath_acc_reg[80]));
DFFPOSX1 dpath_accum_q_reg[81](.D(dpath_accum_n111), .CLK(n9758), .Q(dpath_acc_reg[81]));
DFFPOSX1 dpath_accum_q_reg[82](.D(dpath_accum_n109), .CLK(n9758), .Q(dpath_acc_reg[82]));
DFFPOSX1 dpath_accum_q_reg[83](.D(dpath_accum_n107), .CLK(n9758), .Q(dpath_acc_reg[83]));
DFFPOSX1 dpath_accum_q_reg[84](.D(dpath_accum_n105), .CLK(n9757), .Q(dpath_acc_reg[84]));
DFFPOSX1 dpath_accum_q_reg[85](.D(dpath_accum_n103), .CLK(n9757), .Q(dpath_acc_reg[85]));
DFFPOSX1 dpath_accum_q_reg[86](.D(dpath_accum_n101), .CLK(n9757), .Q(dpath_acc_reg[86]));
DFFPOSX1 dpath_accum_q_reg[87](.D(dpath_accum_n99), .CLK(n9757), .Q(dpath_acc_reg[87]));
DFFPOSX1 dpath_accum_q_reg[88](.D(dpath_accum_n97), .CLK(n9757), .Q(dpath_acc_reg[88]));
DFFPOSX1 dpath_accum_q_reg[89](.D(dpath_accum_n95), .CLK(n9757), .Q(dpath_acc_reg[89]));
DFFPOSX1 dpath_accum_q_reg[90](.D(dpath_accum_n93), .CLK(n9757), .Q(dpath_acc_reg[90]));
DFFPOSX1 dpath_accum_q_reg[91](.D(dpath_accum_n91), .CLK(n9757), .Q(dpath_acc_reg[91]));
DFFPOSX1 dpath_accum_q_reg[92](.D(dpath_accum_n89), .CLK(n9757), .Q(dpath_acc_reg[92]));
DFFPOSX1 dpath_accum_q_reg[93](.D(dpath_accum_n87), .CLK(n9757), .Q(dpath_acc_reg[93]));
DFFPOSX1 dpath_accum_q_reg[94](.D(dpath_accum_n85), .CLK(n9757), .Q(dpath_acc_reg[94]));
DFFPOSX1 dpath_accum_q_reg[95](.D(dpath_accum_n83), .CLK(n9757), .Q(dpath_acc_reg[95]));
DFFPOSX1 dpath_accum_q_reg[96](.D(dpath_accum_n81), .CLK(n9757), .Q(dpath_acc_reg[96]));
DFFPOSX1 dpath_accum_q_reg[97](.D(dpath_accum_n79), .CLK(n9756), .Q(dpath_acc_reg[97]));
DFFPOSX1 dpath_accum_q_reg[98](.D(dpath_accum_n77), .CLK(n9756), .Q(dpath_acc_reg[98]));
DFFPOSX1 dpath_accum_q_reg[99](.D(dpath_accum_n75), .CLK(n9756), .Q(dpath_acc_reg[99]));
DFFPOSX1 dpath_accum_q_reg[100](.D(dpath_accum_n73), .CLK(n9756), .Q(dpath_acc_reg[100]));
DFFPOSX1 dpath_accum_q_reg[101](.D(dpath_accum_n71), .CLK(n9756), .Q(dpath_acc_reg[101]));
DFFPOSX1 dpath_accum_q_reg[102](.D(dpath_accum_n69), .CLK(n9756), .Q(dpath_acc_reg[102]));
DFFPOSX1 dpath_accum_q_reg[103](.D(dpath_accum_n67), .CLK(n9756), .Q(dpath_acc_reg[103]));
DFFPOSX1 dpath_accum_q_reg[104](.D(dpath_accum_n65), .CLK(n9756), .Q(dpath_acc_reg[104]));
DFFPOSX1 dpath_accum_q_reg[105](.D(dpath_accum_n63), .CLK(n9756), .Q(dpath_acc_reg[105]));
DFFPOSX1 dpath_accum_q_reg[106](.D(dpath_accum_n61), .CLK(n9756), .Q(dpath_acc_reg[106]));
DFFPOSX1 dpath_accum_q_reg[107](.D(dpath_accum_n59), .CLK(n9756), .Q(dpath_acc_reg[107]));
DFFPOSX1 dpath_accum_q_reg[108](.D(dpath_accum_n57), .CLK(n9756), .Q(dpath_acc_reg[108]));
DFFPOSX1 dpath_accum_q_reg[109](.D(dpath_accum_n55), .CLK(n9756), .Q(dpath_acc_reg[109]));
DFFPOSX1 dpath_accum_q_reg[110](.D(dpath_accum_n53), .CLK(n9757), .Q(dpath_acc_reg[110]));
DFFPOSX1 dpath_accum_q_reg[111](.D(dpath_accum_n51), .CLK(n9759), .Q(dpath_acc_reg[111]));
DFFPOSX1 dpath_accum_q_reg[112](.D(dpath_accum_n49), .CLK(n9756), .Q(dpath_acc_reg[112]));
DFFPOSX1 dpath_accum_q_reg[113](.D(dpath_accum_n47), .CLK(n9758), .Q(dpath_acc_reg[113]));
DFFPOSX1 dpath_accum_q_reg[114](.D(dpath_accum_n45), .CLK(n9755), .Q(dpath_acc_reg[114]));
DFFPOSX1 dpath_accum_q_reg[115](.D(dpath_accum_n43), .CLK(n9756), .Q(dpath_acc_reg[115]));
DFFPOSX1 dpath_accum_q_reg[116](.D(dpath_accum_n41), .CLK(n9758), .Q(dpath_acc_reg[116]));
DFFPOSX1 dpath_accum_q_reg[117](.D(dpath_accum_n39), .CLK(n9755), .Q(dpath_acc_reg[117]));
DFFPOSX1 dpath_accum_q_reg[118](.D(dpath_accum_n37), .CLK(n9757), .Q(dpath_acc_reg[118]));
DFFPOSX1 dpath_accum_q_reg[119](.D(dpath_accum_n35), .CLK(n9759), .Q(dpath_acc_reg[119]));
DFFPOSX1 dpath_accum_q_reg[120](.D(dpath_accum_n33), .CLK(n9756), .Q(dpath_acc_reg[120]));
DFFPOSX1 dpath_accum_q_reg[121](.D(dpath_accum_n31), .CLK(n9758), .Q(dpath_acc_reg[121]));
DFFPOSX1 dpath_accum_q_reg[122](.D(dpath_accum_n29), .CLK(n9755), .Q(dpath_acc_reg[122]));
DFFPOSX1 dpath_accum_q_reg[123](.D(dpath_accum_n27), .CLK(n9755), .Q(dpath_acc_reg[123]));
DFFPOSX1 dpath_accum_q_reg[124](.D(dpath_accum_n25), .CLK(n9755), .Q(dpath_acc_reg[124]));
DFFPOSX1 dpath_accum_q_reg[125](.D(dpath_accum_n23), .CLK(n9755), .Q(dpath_acc_reg[125]));
DFFPOSX1 dpath_accum_q_reg[126](.D(dpath_accum_n21), .CLK(n9755), .Q(dpath_acc_reg[126]));
DFFPOSX1 dpath_accum_q_reg[127](.D(dpath_accum_n19), .CLK(n9755), .Q(dpath_acc_reg[127]));
DFFPOSX1 dpath_accum_q_reg[128](.D(dpath_accum_n17), .CLK(n9755), .Q(dpath_acc_reg[128]));
DFFPOSX1 dpath_accum_q_reg[129](.D(dpath_accum_n15), .CLK(n9755), .Q(dpath_acc_reg[129]));
DFFPOSX1 dpath_accum_q_reg[130](.D(dpath_accum_n13), .CLK(n9755), .Q(dpath_acc_reg[130]));
DFFPOSX1 dpath_accum_q_reg[131](.D(dpath_accum_n11), .CLK(n9755), .Q(dpath_acc_reg[131]));
DFFPOSX1 dpath_accum_q_reg[132](.D(dpath_accum_n9), .CLK(n9755), .Q(dpath_acc_reg[132]));
DFFPOSX1 dpath_accum_q_reg[133](.D(dpath_accum_n7), .CLK(n9755), .Q(dpath_acc_reg[133]));
DFFPOSX1 dpath_accum_q_reg[134](.D(dpath_accum_n5), .CLK(n9755), .Q(dpath_acc_reg[134]));
DFFPOSX1 dpath_accum_q_reg[135](.D(dpath_accum_n2), .CLK(n9755), .Q(dpath_acc_reg[135]));
LATCH dpath_ckbuf_1_clken_reg(.D(n9785), .CLK(n4), .Q(dpath_ckbuf_1_clken));
DFFPOSX1 dpath_mulcore_cyc1_dff_q_reg[0](.D(dpath_mulcore_cyc1_dff_n2), .CLK(dpath_mulcore_clk_enb0), .Q(dpath_mulcore_cyc1));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[0](.D(dpath_mulcore_ffrs1_n89), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[0]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[1](.D(dpath_mulcore_ffrs1_n67), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[1]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[2](.D(dpath_mulcore_ffrs1_n45), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[2]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[3](.D(dpath_mulcore_ffrs1_n23), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[3]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[4](.D(dpath_mulcore_ffrs1_n7), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[4]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[5](.D(dpath_mulcore_ffrs1_n5), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[5]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[6](.D(dpath_mulcore_ffrs1_n3), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[6]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[7](.D(dpath_mulcore_ffrs1_n129), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[7]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[8](.D(dpath_mulcore_ffrs1_n127), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[8]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[9](.D(dpath_mulcore_ffrs1_n125), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[9]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[10](.D(dpath_mulcore_ffrs1_n123), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[10]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[11](.D(dpath_mulcore_ffrs1_n121), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[11]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[12](.D(dpath_mulcore_ffrs1_n119), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[12]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[13](.D(dpath_mulcore_ffrs1_n117), .CLK(n9718), .Q(dpath_mulcore_op1_l[13]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[14](.D(dpath_mulcore_ffrs1_n115), .CLK(n9719), .Q(dpath_mulcore_op1_l[14]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[15](.D(dpath_mulcore_ffrs1_n113), .CLK(n9719), .Q(dpath_mulcore_op1_l[15]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[16](.D(dpath_mulcore_ffrs1_n111), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[16]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[17](.D(dpath_mulcore_ffrs1_n109), .CLK(n9718), .Q(dpath_mulcore_op1_l[17]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[18](.D(dpath_mulcore_ffrs1_n107), .CLK(n9719), .Q(dpath_mulcore_op1_l[18]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[19](.D(dpath_mulcore_ffrs1_n105), .CLK(n9718), .Q(dpath_mulcore_op1_l[19]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[20](.D(dpath_mulcore_ffrs1_n103), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[20]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[21](.D(dpath_mulcore_ffrs1_n101), .CLK(n9718), .Q(dpath_mulcore_op1_l[21]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[22](.D(dpath_mulcore_ffrs1_n99), .CLK(n9719), .Q(dpath_mulcore_op1_l[22]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[23](.D(dpath_mulcore_ffrs1_n97), .CLK(n9719), .Q(dpath_mulcore_op1_l[23]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[24](.D(dpath_mulcore_ffrs1_n95), .CLK(dpath_mulcore_clk_enb1), .Q(dpath_mulcore_op1_l[24]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[25](.D(dpath_mulcore_ffrs1_n93), .CLK(n9718), .Q(dpath_mulcore_op1_l[25]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[26](.D(dpath_mulcore_ffrs1_n91), .CLK(n9719), .Q(dpath_mulcore_op1_l[26]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[27](.D(dpath_mulcore_ffrs1_n87), .CLK(n9718), .Q(dpath_mulcore_op1_l[27]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[28](.D(dpath_mulcore_ffrs1_n85), .CLK(n9719), .Q(dpath_mulcore_op1_l[28]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[29](.D(dpath_mulcore_ffrs1_n83), .CLK(n9718), .Q(dpath_mulcore_op1_l[29]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[30](.D(dpath_mulcore_ffrs1_n81), .CLK(n9719), .Q(dpath_mulcore_op1_l[30]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[31](.D(dpath_mulcore_ffrs1_n79), .CLK(n9718), .Q(dpath_mulcore_op1_l[31]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[32](.D(dpath_mulcore_ffrs1_n77), .CLK(n9719), .Q(dpath_mulcore_op1_l[32]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[33](.D(dpath_mulcore_ffrs1_n75), .CLK(n9718), .Q(dpath_mulcore_op1_l[33]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[34](.D(dpath_mulcore_ffrs1_n73), .CLK(n9719), .Q(dpath_mulcore_op1_l[34]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[35](.D(dpath_mulcore_ffrs1_n71), .CLK(n9718), .Q(dpath_mulcore_op1_l[35]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[36](.D(dpath_mulcore_ffrs1_n69), .CLK(n9719), .Q(dpath_mulcore_op1_l[36]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[37](.D(dpath_mulcore_ffrs1_n65), .CLK(n9718), .Q(dpath_mulcore_op1_l[37]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[38](.D(dpath_mulcore_ffrs1_n63), .CLK(n9719), .Q(dpath_mulcore_op1_l[38]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[39](.D(dpath_mulcore_ffrs1_n61), .CLK(n9719), .Q(dpath_mulcore_op1_l[39]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[40](.D(dpath_mulcore_ffrs1_n59), .CLK(n9719), .Q(dpath_mulcore_op1_l[40]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[41](.D(dpath_mulcore_ffrs1_n57), .CLK(n9719), .Q(dpath_mulcore_op1_l[41]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[42](.D(dpath_mulcore_ffrs1_n55), .CLK(n9719), .Q(dpath_mulcore_op1_l[42]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[43](.D(dpath_mulcore_ffrs1_n53), .CLK(n9719), .Q(dpath_mulcore_op1_l[43]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[44](.D(dpath_mulcore_ffrs1_n51), .CLK(n9719), .Q(dpath_mulcore_op1_l[44]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[45](.D(dpath_mulcore_ffrs1_n49), .CLK(n9719), .Q(dpath_mulcore_op1_l[45]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[46](.D(dpath_mulcore_ffrs1_n47), .CLK(n9719), .Q(dpath_mulcore_op1_l[46]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[47](.D(dpath_mulcore_ffrs1_n43), .CLK(n9719), .Q(dpath_mulcore_op1_l[47]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[48](.D(dpath_mulcore_ffrs1_n41), .CLK(n9719), .Q(dpath_mulcore_op1_l[48]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[49](.D(dpath_mulcore_ffrs1_n39), .CLK(n9719), .Q(dpath_mulcore_op1_l[49]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[50](.D(dpath_mulcore_ffrs1_n37), .CLK(n9719), .Q(dpath_mulcore_op1_l[50]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[51](.D(dpath_mulcore_ffrs1_n35), .CLK(n9718), .Q(dpath_mulcore_op1_l[51]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[52](.D(dpath_mulcore_ffrs1_n33), .CLK(n9718), .Q(dpath_mulcore_op1_l[52]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[53](.D(dpath_mulcore_ffrs1_n31), .CLK(n9718), .Q(dpath_mulcore_op1_l[53]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[54](.D(dpath_mulcore_ffrs1_n29), .CLK(n9718), .Q(dpath_mulcore_op1_l[54]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[55](.D(dpath_mulcore_ffrs1_n27), .CLK(n9718), .Q(dpath_mulcore_op1_l[55]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[56](.D(dpath_mulcore_ffrs1_n25), .CLK(n9718), .Q(dpath_mulcore_op1_l[56]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[57](.D(dpath_mulcore_ffrs1_n21), .CLK(n9718), .Q(dpath_mulcore_op1_l[57]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[58](.D(dpath_mulcore_ffrs1_n19), .CLK(n9718), .Q(dpath_mulcore_op1_l[58]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[59](.D(dpath_mulcore_ffrs1_n17), .CLK(n9718), .Q(dpath_mulcore_op1_l[59]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[60](.D(dpath_mulcore_ffrs1_n15), .CLK(n9718), .Q(dpath_mulcore_op1_l[60]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[61](.D(dpath_mulcore_ffrs1_n13), .CLK(n9718), .Q(dpath_mulcore_op1_l[61]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[62](.D(dpath_mulcore_ffrs1_n11), .CLK(n9718), .Q(dpath_mulcore_op1_l[62]));
DFFPOSX1 dpath_mulcore_ffrs1_q_reg[63](.D(dpath_mulcore_ffrs1_n9), .CLK(n9718), .Q(dpath_mulcore_op1_l[63]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[0](.D(dpath_mulcore_a0cot_dff_n117), .CLK(dpath_mulcore_clk_enb0), .Q(dpath_mulcore_a0c[4]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[1](.D(dpath_mulcore_a0cot_dff_n95), .CLK(n9658), .Q(dpath_mulcore_a0c[5]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[2](.D(dpath_mulcore_a0cot_dff_n73), .CLK(n9658), .Q(dpath_mulcore_a0c[6]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[3](.D(dpath_mulcore_a0cot_dff_n51), .CLK(n9658), .Q(dpath_mulcore_a0c[7]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[4](.D(dpath_mulcore_a0cot_dff_n29), .CLK(n9658), .Q(dpath_mulcore_a0c[8]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[5](.D(dpath_mulcore_a0cot_dff_n7), .CLK(n9658), .Q(dpath_mulcore_a0c[9]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[6](.D(dpath_mulcore_a0cot_dff_n3), .CLK(n9658), .Q(dpath_mulcore_a0c[10]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[7](.D(dpath_mulcore_a0cot_dff_n157), .CLK(n9658), .Q(dpath_mulcore_a0c[11]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[8](.D(dpath_mulcore_a0cot_dff_n155), .CLK(n9658), .Q(dpath_mulcore_a0c[12]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[9](.D(dpath_mulcore_a0cot_dff_n153), .CLK(n9658), .Q(dpath_mulcore_a0c[13]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[10](.D(dpath_mulcore_a0cot_dff_n151), .CLK(n9658), .Q(dpath_mulcore_a0c[14]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[11](.D(dpath_mulcore_a0cot_dff_n149), .CLK(n9658), .Q(dpath_mulcore_a0c[15]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[12](.D(dpath_mulcore_a0cot_dff_n147), .CLK(n9658), .Q(dpath_mulcore_a0c[16]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[13](.D(dpath_mulcore_a0cot_dff_n145), .CLK(n9658), .Q(dpath_mulcore_a0c[17]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[14](.D(dpath_mulcore_a0cot_dff_n143), .CLK(n9657), .Q(dpath_mulcore_a0c[18]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[15](.D(dpath_mulcore_a0cot_dff_n141), .CLK(n9657), .Q(dpath_mulcore_a0c[19]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[16](.D(dpath_mulcore_a0cot_dff_n139), .CLK(n9657), .Q(dpath_mulcore_a0c[20]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[17](.D(dpath_mulcore_a0cot_dff_n137), .CLK(n9657), .Q(dpath_mulcore_a0c[21]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[18](.D(dpath_mulcore_a0cot_dff_n135), .CLK(n9657), .Q(dpath_mulcore_a0c[22]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[19](.D(dpath_mulcore_a0cot_dff_n133), .CLK(n9657), .Q(dpath_mulcore_a0c[23]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[20](.D(dpath_mulcore_a0cot_dff_n131), .CLK(n9657), .Q(dpath_mulcore_a0c[24]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[21](.D(dpath_mulcore_a0cot_dff_n129), .CLK(n9657), .Q(dpath_mulcore_a0c[25]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[22](.D(dpath_mulcore_a0cot_dff_n127), .CLK(n9657), .Q(dpath_mulcore_a0c[26]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[23](.D(dpath_mulcore_a0cot_dff_n125), .CLK(n9657), .Q(dpath_mulcore_a0c[27]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[24](.D(dpath_mulcore_a0cot_dff_n123), .CLK(n9657), .Q(dpath_mulcore_a0c[28]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[25](.D(dpath_mulcore_a0cot_dff_n121), .CLK(n9657), .Q(dpath_mulcore_a0c[29]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[26](.D(dpath_mulcore_a0cot_dff_n119), .CLK(n9657), .Q(dpath_mulcore_a0c[30]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[27](.D(dpath_mulcore_a0cot_dff_n115), .CLK(n9656), .Q(dpath_mulcore_a0c[31]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[28](.D(dpath_mulcore_a0cot_dff_n113), .CLK(n9656), .Q(dpath_mulcore_a0c[32]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[29](.D(dpath_mulcore_a0cot_dff_n111), .CLK(n9656), .Q(dpath_mulcore_a0c[33]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[30](.D(dpath_mulcore_a0cot_dff_n109), .CLK(n9656), .Q(dpath_mulcore_a0c[34]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[31](.D(dpath_mulcore_a0cot_dff_n107), .CLK(n9656), .Q(dpath_mulcore_a0c[35]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[32](.D(dpath_mulcore_a0cot_dff_n105), .CLK(n9656), .Q(dpath_mulcore_a0c[36]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[33](.D(dpath_mulcore_a0cot_dff_n103), .CLK(n9656), .Q(dpath_mulcore_a0c[37]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[34](.D(dpath_mulcore_a0cot_dff_n101), .CLK(n9656), .Q(dpath_mulcore_a0c[38]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[35](.D(dpath_mulcore_a0cot_dff_n99), .CLK(n9656), .Q(dpath_mulcore_a0c[39]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[36](.D(dpath_mulcore_a0cot_dff_n97), .CLK(n9656), .Q(dpath_mulcore_a0c[40]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[37](.D(dpath_mulcore_a0cot_dff_n93), .CLK(n9656), .Q(dpath_mulcore_a0c[41]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[38](.D(dpath_mulcore_a0cot_dff_n91), .CLK(n9656), .Q(dpath_mulcore_a0c[42]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[39](.D(dpath_mulcore_a0cot_dff_n89), .CLK(n9656), .Q(dpath_mulcore_a0c[43]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[40](.D(dpath_mulcore_a0cot_dff_n87), .CLK(n9655), .Q(dpath_mulcore_a0c[44]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[41](.D(dpath_mulcore_a0cot_dff_n85), .CLK(n9655), .Q(dpath_mulcore_a0c[45]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[42](.D(dpath_mulcore_a0cot_dff_n83), .CLK(n9655), .Q(dpath_mulcore_a0c[46]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[43](.D(dpath_mulcore_a0cot_dff_n81), .CLK(n9655), .Q(dpath_mulcore_a0c[47]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[44](.D(dpath_mulcore_a0cot_dff_n79), .CLK(n9655), .Q(dpath_mulcore_a0c[48]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[45](.D(dpath_mulcore_a0cot_dff_n77), .CLK(n9655), .Q(dpath_mulcore_a0c[49]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[46](.D(dpath_mulcore_a0cot_dff_n75), .CLK(n9655), .Q(dpath_mulcore_a0c[50]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[47](.D(dpath_mulcore_a0cot_dff_n71), .CLK(n9655), .Q(dpath_mulcore_a0c[51]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[48](.D(dpath_mulcore_a0cot_dff_n69), .CLK(n9655), .Q(dpath_mulcore_a0c[52]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[49](.D(dpath_mulcore_a0cot_dff_n67), .CLK(n9655), .Q(dpath_mulcore_a0c[53]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[50](.D(dpath_mulcore_a0cot_dff_n65), .CLK(n9655), .Q(dpath_mulcore_a0c[54]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[51](.D(dpath_mulcore_a0cot_dff_n63), .CLK(n9655), .Q(dpath_mulcore_a0c[55]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[52](.D(dpath_mulcore_a0cot_dff_n61), .CLK(n9655), .Q(dpath_mulcore_a0c[56]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[53](.D(dpath_mulcore_a0cot_dff_n59), .CLK(n9654), .Q(dpath_mulcore_a0c[57]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[54](.D(dpath_mulcore_a0cot_dff_n57), .CLK(n9654), .Q(dpath_mulcore_a0c[58]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[55](.D(dpath_mulcore_a0cot_dff_n55), .CLK(n9654), .Q(dpath_mulcore_a0c[59]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[56](.D(dpath_mulcore_a0cot_dff_n53), .CLK(n9654), .Q(dpath_mulcore_a0c[60]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[57](.D(dpath_mulcore_a0cot_dff_n49), .CLK(n9654), .Q(dpath_mulcore_a0c[61]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[58](.D(dpath_mulcore_a0cot_dff_n47), .CLK(n9654), .Q(dpath_mulcore_a0c[62]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[59](.D(dpath_mulcore_a0cot_dff_n45), .CLK(n9654), .Q(dpath_mulcore_a0c[63]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[60](.D(dpath_mulcore_a0cot_dff_n43), .CLK(n9654), .Q(dpath_mulcore_a0c[64]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[61](.D(dpath_mulcore_a0cot_dff_n41), .CLK(n9654), .Q(dpath_mulcore_a0c[65]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[62](.D(dpath_mulcore_a0cot_dff_n39), .CLK(n9654), .Q(dpath_mulcore_a0c[66]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[63](.D(dpath_mulcore_a0cot_dff_n37), .CLK(n9654), .Q(dpath_mulcore_a0c[67]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[64](.D(dpath_mulcore_a0cot_dff_n35), .CLK(n9654), .Q(dpath_mulcore_a0c[68]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[65](.D(dpath_mulcore_a0cot_dff_n33), .CLK(n9654), .Q(dpath_mulcore_a0c[69]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[66](.D(dpath_mulcore_a0cot_dff_n31), .CLK(n9653), .Q(dpath_mulcore_a0c[70]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[67](.D(dpath_mulcore_a0cot_dff_n27), .CLK(n9653), .Q(dpath_mulcore_a0c[71]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[68](.D(dpath_mulcore_a0cot_dff_n25), .CLK(n9653), .Q(dpath_mulcore_a0c[72]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[69](.D(dpath_mulcore_a0cot_dff_n23), .CLK(n9653), .Q(dpath_mulcore_a0c[73]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[70](.D(dpath_mulcore_a0cot_dff_n21), .CLK(n9653), .Q(dpath_mulcore_a0c[74]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[71](.D(dpath_mulcore_a0cot_dff_n19), .CLK(n9653), .Q(dpath_mulcore_a0c[75]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[72](.D(dpath_mulcore_a0cot_dff_n17), .CLK(n9653), .Q(dpath_mulcore_a0c[76]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[73](.D(dpath_mulcore_a0cot_dff_n15), .CLK(n9653), .Q(dpath_mulcore_a0c[77]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[74](.D(dpath_mulcore_a0cot_dff_n13), .CLK(n9653), .Q(dpath_mulcore_a0c[78]));
DFFPOSX1 dpath_mulcore_a0cot_dff_q_reg[75](.D(dpath_mulcore_a0cot_dff_n11), .CLK(n9653), .Q(dpath_mulcore_a0c[79]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[0](.D(dpath_mulcore_a0sum_dff_n125), .CLK(n9653), .Q(dpath_mulcore_a0s[0]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[1](.D(dpath_mulcore_a0sum_dff_n103), .CLK(n9652), .Q(dpath_mulcore_a0s[1]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[2](.D(dpath_mulcore_a0sum_dff_n81), .CLK(n9652), .Q(dpath_mulcore_a0s[2]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[3](.D(dpath_mulcore_a0sum_dff_n59), .CLK(n9652), .Q(dpath_mulcore_a0s[3]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[4](.D(dpath_mulcore_a0sum_dff_n37), .CLK(n9652), .Q(dpath_mulcore_a0s[4]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[5](.D(dpath_mulcore_a0sum_dff_n15), .CLK(n9652), .Q(dpath_mulcore_a0s[5]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[6](.D(dpath_mulcore_a0sum_dff_n3), .CLK(n9652), .Q(dpath_mulcore_a0s[6]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[7](.D(dpath_mulcore_a0sum_dff_n165), .CLK(n9652), .Q(dpath_mulcore_a0s[7]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[8](.D(dpath_mulcore_a0sum_dff_n163), .CLK(n9652), .Q(dpath_mulcore_a0s[8]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[9](.D(dpath_mulcore_a0sum_dff_n161), .CLK(n9652), .Q(dpath_mulcore_a0s[9]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[10](.D(dpath_mulcore_a0sum_dff_n159), .CLK(n9652), .Q(dpath_mulcore_a0s[10]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[11](.D(dpath_mulcore_a0sum_dff_n157), .CLK(n9652), .Q(dpath_mulcore_a0s[11]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[12](.D(dpath_mulcore_a0sum_dff_n155), .CLK(n9652), .Q(dpath_mulcore_a0s[12]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[13](.D(dpath_mulcore_a0sum_dff_n153), .CLK(n9652), .Q(dpath_mulcore_a0s[13]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[14](.D(dpath_mulcore_a0sum_dff_n151), .CLK(n9651), .Q(dpath_mulcore_a0s[14]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[15](.D(dpath_mulcore_a0sum_dff_n149), .CLK(n9651), .Q(dpath_mulcore_a0s[15]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[16](.D(dpath_mulcore_a0sum_dff_n147), .CLK(n9651), .Q(dpath_mulcore_a0s[16]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[17](.D(dpath_mulcore_a0sum_dff_n145), .CLK(n9651), .Q(dpath_mulcore_a0s[17]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[18](.D(dpath_mulcore_a0sum_dff_n143), .CLK(n9651), .Q(dpath_mulcore_a0s[18]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[19](.D(dpath_mulcore_a0sum_dff_n141), .CLK(n9651), .Q(dpath_mulcore_a0s[19]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[20](.D(dpath_mulcore_a0sum_dff_n139), .CLK(n9651), .Q(dpath_mulcore_a0s[20]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[21](.D(dpath_mulcore_a0sum_dff_n137), .CLK(n9651), .Q(dpath_mulcore_a0s[21]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[22](.D(dpath_mulcore_a0sum_dff_n135), .CLK(n9651), .Q(dpath_mulcore_a0s[22]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[23](.D(dpath_mulcore_a0sum_dff_n133), .CLK(n9651), .Q(dpath_mulcore_a0s[23]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[24](.D(dpath_mulcore_a0sum_dff_n131), .CLK(n9651), .Q(dpath_mulcore_a0s[24]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[25](.D(dpath_mulcore_a0sum_dff_n129), .CLK(n9651), .Q(dpath_mulcore_a0s[25]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[26](.D(dpath_mulcore_a0sum_dff_n127), .CLK(n9651), .Q(dpath_mulcore_a0s[26]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[27](.D(dpath_mulcore_a0sum_dff_n123), .CLK(n9650), .Q(dpath_mulcore_a0s[27]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[28](.D(dpath_mulcore_a0sum_dff_n121), .CLK(n9650), .Q(dpath_mulcore_a0s[28]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[29](.D(dpath_mulcore_a0sum_dff_n119), .CLK(n9650), .Q(dpath_mulcore_a0s[29]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[30](.D(dpath_mulcore_a0sum_dff_n117), .CLK(n9650), .Q(dpath_mulcore_a0s[30]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[31](.D(dpath_mulcore_a0sum_dff_n115), .CLK(n9650), .Q(dpath_mulcore_a0s[31]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[32](.D(dpath_mulcore_a0sum_dff_n113), .CLK(n9650), .Q(dpath_mulcore_a0s[32]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[33](.D(dpath_mulcore_a0sum_dff_n111), .CLK(n9650), .Q(dpath_mulcore_a0s[33]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[34](.D(dpath_mulcore_a0sum_dff_n109), .CLK(n9650), .Q(dpath_mulcore_a0s[34]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[35](.D(dpath_mulcore_a0sum_dff_n107), .CLK(n9650), .Q(dpath_mulcore_a0s[35]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[36](.D(dpath_mulcore_a0sum_dff_n105), .CLK(n9650), .Q(dpath_mulcore_a0s[36]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[37](.D(dpath_mulcore_a0sum_dff_n101), .CLK(n9650), .Q(dpath_mulcore_a0s[37]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[38](.D(dpath_mulcore_a0sum_dff_n99), .CLK(n9650), .Q(dpath_mulcore_a0s[38]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[39](.D(dpath_mulcore_a0sum_dff_n97), .CLK(n9650), .Q(dpath_mulcore_a0s[39]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[40](.D(dpath_mulcore_a0sum_dff_n95), .CLK(n9649), .Q(dpath_mulcore_a0s[40]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[41](.D(dpath_mulcore_a0sum_dff_n93), .CLK(n9649), .Q(dpath_mulcore_a0s[41]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[42](.D(dpath_mulcore_a0sum_dff_n91), .CLK(n9649), .Q(dpath_mulcore_a0s[42]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[43](.D(dpath_mulcore_a0sum_dff_n89), .CLK(n9649), .Q(dpath_mulcore_a0s[43]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[44](.D(dpath_mulcore_a0sum_dff_n87), .CLK(n9649), .Q(dpath_mulcore_a0s[44]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[45](.D(dpath_mulcore_a0sum_dff_n85), .CLK(n9649), .Q(dpath_mulcore_a0s[45]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[46](.D(dpath_mulcore_a0sum_dff_n83), .CLK(n9649), .Q(dpath_mulcore_a0s[46]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[47](.D(dpath_mulcore_a0sum_dff_n79), .CLK(n9649), .Q(dpath_mulcore_a0s[47]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[48](.D(dpath_mulcore_a0sum_dff_n77), .CLK(n9649), .Q(dpath_mulcore_a0s[48]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[49](.D(dpath_mulcore_a0sum_dff_n75), .CLK(n9649), .Q(dpath_mulcore_a0s[49]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[50](.D(dpath_mulcore_a0sum_dff_n73), .CLK(n9649), .Q(dpath_mulcore_a0s[50]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[51](.D(dpath_mulcore_a0sum_dff_n71), .CLK(n9649), .Q(dpath_mulcore_a0s[51]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[52](.D(dpath_mulcore_a0sum_dff_n69), .CLK(n9649), .Q(dpath_mulcore_a0s[52]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[53](.D(dpath_mulcore_a0sum_dff_n67), .CLK(n9648), .Q(dpath_mulcore_a0s[53]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[54](.D(dpath_mulcore_a0sum_dff_n65), .CLK(n9648), .Q(dpath_mulcore_a0s[54]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[55](.D(dpath_mulcore_a0sum_dff_n63), .CLK(n9648), .Q(dpath_mulcore_a0s[55]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[56](.D(dpath_mulcore_a0sum_dff_n61), .CLK(n9648), .Q(dpath_mulcore_a0s[56]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[57](.D(dpath_mulcore_a0sum_dff_n57), .CLK(n9648), .Q(dpath_mulcore_a0s[57]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[58](.D(dpath_mulcore_a0sum_dff_n55), .CLK(n9648), .Q(dpath_mulcore_a0s[58]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[59](.D(dpath_mulcore_a0sum_dff_n53), .CLK(n9648), .Q(dpath_mulcore_a0s[59]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[60](.D(dpath_mulcore_a0sum_dff_n51), .CLK(n9648), .Q(dpath_mulcore_a0s[60]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[61](.D(dpath_mulcore_a0sum_dff_n49), .CLK(n9648), .Q(dpath_mulcore_a0s[61]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[62](.D(dpath_mulcore_a0sum_dff_n47), .CLK(n9648), .Q(dpath_mulcore_a0s[62]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[63](.D(dpath_mulcore_a0sum_dff_n45), .CLK(n9648), .Q(dpath_mulcore_a0s[63]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[64](.D(dpath_mulcore_a0sum_dff_n43), .CLK(n9648), .Q(dpath_mulcore_a0s[64]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[65](.D(dpath_mulcore_a0sum_dff_n41), .CLK(n9648), .Q(dpath_mulcore_a0s[65]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[66](.D(dpath_mulcore_a0sum_dff_n39), .CLK(n9647), .Q(dpath_mulcore_a0s[66]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[67](.D(dpath_mulcore_a0sum_dff_n35), .CLK(n9647), .Q(dpath_mulcore_a0s[67]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[68](.D(dpath_mulcore_a0sum_dff_n33), .CLK(n9647), .Q(dpath_mulcore_a0s[68]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[69](.D(dpath_mulcore_a0sum_dff_n31), .CLK(n9647), .Q(dpath_mulcore_a0s[69]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[70](.D(dpath_mulcore_a0sum_dff_n29), .CLK(n9647), .Q(dpath_mulcore_a0s[70]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[71](.D(dpath_mulcore_a0sum_dff_n27), .CLK(n9647), .Q(dpath_mulcore_a0s[71]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[72](.D(dpath_mulcore_a0sum_dff_n25), .CLK(n9647), .Q(dpath_mulcore_a0s[72]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[73](.D(dpath_mulcore_a0sum_dff_n23), .CLK(n9647), .Q(dpath_mulcore_a0s[73]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[74](.D(dpath_mulcore_a0sum_dff_n21), .CLK(n9647), .Q(dpath_mulcore_a0s[74]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[75](.D(dpath_mulcore_a0sum_dff_n19), .CLK(n9647), .Q(dpath_mulcore_a0s[75]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[76](.D(dpath_mulcore_a0sum_dff_n17), .CLK(n9647), .Q(dpath_mulcore_a0s[76]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[77](.D(dpath_mulcore_a0sum_dff_n13), .CLK(n9647), .Q(dpath_mulcore_a0s[77]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[78](.D(dpath_mulcore_a0sum_dff_n11), .CLK(n9647), .Q(dpath_mulcore_a0s[78]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[79](.D(dpath_mulcore_a0sum_dff_n9), .CLK(n9646), .Q(dpath_mulcore_a0s[79]));
DFFPOSX1 dpath_mulcore_a0sum_dff_q_reg[80](.D(n9550), .CLK(n9646), .Q(dpath_mulcore_a0s[80]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[0](.D(dpath_mulcore_a2cot_dff_n155), .CLK(n9646), .Q(dpath_mulcore_addin_cout[0]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[1](.D(dpath_mulcore_a2cot_dff_n133), .CLK(n9646), .Q(dpath_mulcore_addin_cout[1]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[2](.D(dpath_mulcore_a2cot_dff_n111), .CLK(n9646), .Q(dpath_mulcore_addin_cout[2]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[3](.D(dpath_mulcore_a2cot_dff_n89), .CLK(n9646), .Q(dpath_mulcore_addin_cout[3]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[4](.D(dpath_mulcore_a2cot_dff_n67), .CLK(n9646), .Q(dpath_mulcore_addin_cout[4]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[5](.D(dpath_mulcore_a2cot_dff_n45), .CLK(n9646), .Q(dpath_mulcore_addin_cout[5]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[6](.D(dpath_mulcore_a2cot_dff_n23), .CLK(n9646), .Q(dpath_mulcore_addin_cout[6]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[7](.D(dpath_mulcore_a2cot_dff_n195), .CLK(n9646), .Q(dpath_mulcore_addin_cout[7]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[8](.D(dpath_mulcore_a2cot_dff_n193), .CLK(n9646), .Q(dpath_mulcore_addin_cout[8]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[9](.D(dpath_mulcore_a2cot_dff_n191), .CLK(n9646), .Q(dpath_mulcore_addin_cout[9]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[10](.D(dpath_mulcore_a2cot_dff_n189), .CLK(n9645), .Q(dpath_mulcore_addin_cout[10]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[11](.D(dpath_mulcore_a2cot_dff_n187), .CLK(n9645), .Q(dpath_mulcore_addin_cout[11]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[12](.D(dpath_mulcore_a2cot_dff_n185), .CLK(n9645), .Q(dpath_mulcore_addin_cout[12]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[13](.D(dpath_mulcore_a2cot_dff_n183), .CLK(n9645), .Q(dpath_mulcore_addin_cout[13]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[14](.D(dpath_mulcore_a2cot_dff_n181), .CLK(n9645), .Q(dpath_mulcore_addin_cout[14]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[15](.D(dpath_mulcore_a2cot_dff_n179), .CLK(n9645), .Q(dpath_mulcore_addin_cout[15]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[16](.D(dpath_mulcore_a2cot_dff_n177), .CLK(n9645), .Q(dpath_mulcore_addin_cout[16]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[17](.D(dpath_mulcore_a2cot_dff_n175), .CLK(n9645), .Q(dpath_mulcore_addin_cout[17]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[18](.D(dpath_mulcore_a2cot_dff_n173), .CLK(n9645), .Q(dpath_mulcore_addin_cout[18]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[19](.D(dpath_mulcore_a2cot_dff_n171), .CLK(n9645), .Q(dpath_mulcore_addin_cout[19]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[20](.D(dpath_mulcore_a2cot_dff_n169), .CLK(n9645), .Q(dpath_mulcore_addin_cout[20]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[21](.D(dpath_mulcore_a2cot_dff_n167), .CLK(n9645), .Q(dpath_mulcore_addin_cout[21]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[22](.D(dpath_mulcore_a2cot_dff_n165), .CLK(n9645), .Q(dpath_mulcore_addin_cout[22]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[23](.D(dpath_mulcore_a2cot_dff_n163), .CLK(n9644), .Q(dpath_mulcore_addin_cout[23]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[24](.D(dpath_mulcore_a2cot_dff_n161), .CLK(n9644), .Q(dpath_mulcore_addin_cout[24]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[25](.D(dpath_mulcore_a2cot_dff_n159), .CLK(n9644), .Q(dpath_mulcore_addin_cout[25]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[26](.D(dpath_mulcore_a2cot_dff_n157), .CLK(n9644), .Q(dpath_mulcore_addin_cout[26]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[27](.D(dpath_mulcore_a2cot_dff_n153), .CLK(n9644), .Q(dpath_mulcore_addin_cout[27]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[28](.D(dpath_mulcore_a2cot_dff_n151), .CLK(n9644), .Q(dpath_mulcore_addin_cout[28]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[29](.D(dpath_mulcore_a2cot_dff_n149), .CLK(n9644), .Q(dpath_mulcore_addin_cout[29]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[30](.D(dpath_mulcore_a2cot_dff_n147), .CLK(n9644), .Q(dpath_mulcore_addin_cout[30]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[31](.D(dpath_mulcore_a2cot_dff_n145), .CLK(n9644), .Q(dpath_mulcore_addin_cout[31]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[32](.D(dpath_mulcore_a2cot_dff_n143), .CLK(n9644), .Q(dpath_mulcore_addin_cout[32]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[33](.D(dpath_mulcore_a2cot_dff_n141), .CLK(n9644), .Q(dpath_mulcore_addin_cout[33]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[34](.D(dpath_mulcore_a2cot_dff_n139), .CLK(n9644), .Q(dpath_mulcore_addin_cout[34]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[35](.D(dpath_mulcore_a2cot_dff_n137), .CLK(n9644), .Q(dpath_mulcore_addin_cout[35]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[36](.D(dpath_mulcore_a2cot_dff_n135), .CLK(n9643), .Q(dpath_mulcore_addin_cout[36]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[37](.D(dpath_mulcore_a2cot_dff_n131), .CLK(n9643), .Q(dpath_mulcore_addin_cout[37]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[38](.D(dpath_mulcore_a2cot_dff_n129), .CLK(n9643), .Q(dpath_mulcore_addin_cout[38]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[39](.D(dpath_mulcore_a2cot_dff_n127), .CLK(n9643), .Q(dpath_mulcore_addin_cout[39]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[40](.D(dpath_mulcore_a2cot_dff_n125), .CLK(n9643), .Q(dpath_mulcore_addin_cout[40]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[41](.D(dpath_mulcore_a2cot_dff_n123), .CLK(n9643), .Q(dpath_mulcore_addin_cout[41]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[42](.D(dpath_mulcore_a2cot_dff_n121), .CLK(n9643), .Q(dpath_mulcore_addin_cout[42]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[43](.D(dpath_mulcore_a2cot_dff_n119), .CLK(n9643), .Q(dpath_mulcore_addin_cout[43]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[44](.D(dpath_mulcore_a2cot_dff_n117), .CLK(n9643), .Q(dpath_mulcore_addin_cout[44]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[45](.D(dpath_mulcore_a2cot_dff_n115), .CLK(n9643), .Q(dpath_mulcore_addin_cout[45]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[46](.D(dpath_mulcore_a2cot_dff_n113), .CLK(n9643), .Q(dpath_mulcore_addin_cout[46]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[47](.D(dpath_mulcore_a2cot_dff_n109), .CLK(n9643), .Q(dpath_mulcore_addin_cout[47]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[48](.D(dpath_mulcore_a2cot_dff_n107), .CLK(n9643), .Q(dpath_mulcore_addin_cout[48]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[49](.D(dpath_mulcore_a2cot_dff_n105), .CLK(n9642), .Q(dpath_mulcore_addin_cout[49]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[50](.D(dpath_mulcore_a2cot_dff_n103), .CLK(n9642), .Q(dpath_mulcore_addin_cout[50]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[51](.D(dpath_mulcore_a2cot_dff_n101), .CLK(n9642), .Q(dpath_mulcore_addin_cout[51]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[52](.D(dpath_mulcore_a2cot_dff_n99), .CLK(n9642), .Q(dpath_mulcore_addin_cout[52]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[53](.D(dpath_mulcore_a2cot_dff_n97), .CLK(n9642), .Q(dpath_mulcore_addin_cout[53]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[54](.D(dpath_mulcore_a2cot_dff_n95), .CLK(n9642), .Q(dpath_mulcore_addin_cout[54]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[55](.D(dpath_mulcore_a2cot_dff_n93), .CLK(n9642), .Q(dpath_mulcore_addin_cout[55]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[56](.D(dpath_mulcore_a2cot_dff_n91), .CLK(n9642), .Q(dpath_mulcore_addin_cout[56]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[57](.D(dpath_mulcore_a2cot_dff_n87), .CLK(n9642), .Q(dpath_mulcore_addin_cout[57]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[58](.D(dpath_mulcore_a2cot_dff_n85), .CLK(n9642), .Q(dpath_mulcore_addin_cout[58]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[59](.D(dpath_mulcore_a2cot_dff_n83), .CLK(n9642), .Q(dpath_mulcore_addin_cout[59]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[60](.D(dpath_mulcore_a2cot_dff_n81), .CLK(n9642), .Q(dpath_mulcore_addin_cout[60]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[61](.D(dpath_mulcore_a2cot_dff_n79), .CLK(n9642), .Q(dpath_mulcore_addin_cout[61]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[62](.D(dpath_mulcore_a2cot_dff_n77), .CLK(n9641), .Q(dpath_mulcore_addin_cout[62]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[63](.D(dpath_mulcore_a2cot_dff_n75), .CLK(n9641), .Q(dpath_mulcore_addin_cout[63]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[64](.D(dpath_mulcore_a2cot_dff_n73), .CLK(n9641), .Q(dpath_mulcore_addin_cout[64]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[65](.D(dpath_mulcore_a2cot_dff_n71), .CLK(n9641), .Q(dpath_mulcore_addin_cout[65]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[66](.D(dpath_mulcore_a2cot_dff_n69), .CLK(n9641), .Q(dpath_mulcore_addin_cout[66]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[67](.D(dpath_mulcore_a2cot_dff_n65), .CLK(n9641), .Q(dpath_mulcore_addin_cout[67]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[68](.D(dpath_mulcore_a2cot_dff_n63), .CLK(n9641), .Q(dpath_mulcore_addin_cout[68]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[69](.D(dpath_mulcore_a2cot_dff_n61), .CLK(n9641), .Q(dpath_mulcore_addin_cout[69]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[70](.D(dpath_mulcore_a2cot_dff_n59), .CLK(n9641), .Q(dpath_mulcore_addin_cout[70]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[71](.D(dpath_mulcore_a2cot_dff_n57), .CLK(n9641), .Q(dpath_mulcore_addin_cout[71]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[72](.D(dpath_mulcore_a2cot_dff_n55), .CLK(n9641), .Q(dpath_mulcore_addin_cout[72]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[73](.D(dpath_mulcore_a2cot_dff_n53), .CLK(n9641), .Q(dpath_mulcore_addin_cout[73]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[74](.D(dpath_mulcore_a2cot_dff_n51), .CLK(n9641), .Q(dpath_mulcore_addin_cout[74]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[75](.D(dpath_mulcore_a2cot_dff_n49), .CLK(n9640), .Q(dpath_mulcore_addin_cout[75]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[76](.D(dpath_mulcore_a2cot_dff_n47), .CLK(n9640), .Q(dpath_mulcore_addin_cout[76]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[77](.D(dpath_mulcore_a2cot_dff_n43), .CLK(n9640), .Q(dpath_mulcore_addin_cout[77]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[78](.D(dpath_mulcore_a2cot_dff_n41), .CLK(n9640), .Q(dpath_mulcore_addin_cout[78]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[79](.D(dpath_mulcore_a2cot_dff_n39), .CLK(n9640), .Q(dpath_mulcore_addin_cout[79]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[80](.D(dpath_mulcore_a2cot_dff_n37), .CLK(n9640), .Q(dpath_mulcore_addin_cout[80]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[81](.D(dpath_mulcore_a2cot_dff_n35), .CLK(n9640), .Q(dpath_mulcore_addin_cout[81]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[82](.D(dpath_mulcore_a2cot_dff_n33), .CLK(n9640), .Q(dpath_mulcore_addin_cout[82]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[83](.D(dpath_mulcore_a2cot_dff_n31), .CLK(n9640), .Q(dpath_mulcore_addin_cout[83]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[84](.D(dpath_mulcore_a2cot_dff_n29), .CLK(n9640), .Q(dpath_mulcore_addin_cout[84]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[85](.D(dpath_mulcore_a2cot_dff_n27), .CLK(n9640), .Q(dpath_mulcore_addin_cout[85]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[86](.D(dpath_mulcore_a2cot_dff_n25), .CLK(n9640), .Q(dpath_mulcore_addin_cout[86]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[87](.D(dpath_mulcore_a2cot_dff_n21), .CLK(n9640), .Q(dpath_mulcore_addin_cout[87]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[88](.D(dpath_mulcore_a2cot_dff_n19), .CLK(n9639), .Q(dpath_mulcore_addin_cout[88]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[89](.D(dpath_mulcore_a2cot_dff_n17), .CLK(n9639), .Q(dpath_mulcore_addin_cout[89]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[90](.D(dpath_mulcore_a2cot_dff_n15), .CLK(n9639), .Q(dpath_mulcore_addin_cout[90]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[91](.D(dpath_mulcore_a2cot_dff_n13), .CLK(n9639), .Q(dpath_mulcore_addin_cout[91]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[92](.D(dpath_mulcore_a2cot_dff_n11), .CLK(n9639), .Q(dpath_mulcore_addin_cout[92]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[93](.D(dpath_mulcore_a2cot_dff_n9), .CLK(n9639), .Q(dpath_mulcore_addin_cout[93]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[94](.D(dpath_mulcore_a2cot_dff_n7), .CLK(n9639), .Q(dpath_mulcore_addin_cout[94]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[95](.D(dpath_mulcore_a2cot_dff_n5), .CLK(n9639), .Q(dpath_mulcore_addin_cout[95]));
DFFPOSX1 dpath_mulcore_a2cot_dff_q_reg[96](.D(dpath_mulcore_a2cot_dff_n3), .CLK(n9639), .Q(dpath_mulcore_addin_cout[96]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[0](.D(dpath_mulcore_a2sum_dff_n155), .CLK(n9639), .Q(dpath_mulcore_addin_sum[0]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[1](.D(dpath_mulcore_a2sum_dff_n133), .CLK(n9639), .Q(dpath_mulcore_addin_sum[1]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[2](.D(dpath_mulcore_a2sum_dff_n111), .CLK(n9639), .Q(dpath_mulcore_addin_sum[2]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[3](.D(dpath_mulcore_a2sum_dff_n89), .CLK(n9639), .Q(dpath_mulcore_addin_sum[3]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[4](.D(dpath_mulcore_a2sum_dff_n67), .CLK(n9638), .Q(dpath_mulcore_addin_sum[4]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[5](.D(dpath_mulcore_a2sum_dff_n45), .CLK(n9638), .Q(dpath_mulcore_addin_sum[5]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[6](.D(dpath_mulcore_a2sum_dff_n23), .CLK(n9638), .Q(dpath_mulcore_addin_sum[6]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[7](.D(dpath_mulcore_a2sum_dff_n197), .CLK(n9638), .Q(dpath_mulcore_addin_sum[7]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[8](.D(dpath_mulcore_a2sum_dff_n193), .CLK(n9638), .Q(dpath_mulcore_addin_sum[8]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[9](.D(dpath_mulcore_a2sum_dff_n191), .CLK(n9638), .Q(dpath_mulcore_addin_sum[9]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[10](.D(dpath_mulcore_a2sum_dff_n189), .CLK(n9638), .Q(dpath_mulcore_addin_sum[10]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[11](.D(dpath_mulcore_a2sum_dff_n187), .CLK(n9638), .Q(dpath_mulcore_addin_sum[11]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[12](.D(dpath_mulcore_a2sum_dff_n185), .CLK(n9638), .Q(dpath_mulcore_addin_sum[12]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[13](.D(dpath_mulcore_a2sum_dff_n183), .CLK(n9638), .Q(dpath_mulcore_addin_sum[13]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[14](.D(dpath_mulcore_a2sum_dff_n181), .CLK(n9638), .Q(dpath_mulcore_addin_sum[14]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[15](.D(dpath_mulcore_a2sum_dff_n179), .CLK(n9638), .Q(dpath_mulcore_addin_sum[15]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[16](.D(dpath_mulcore_a2sum_dff_n177), .CLK(n9638), .Q(dpath_mulcore_addin_sum[16]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[17](.D(dpath_mulcore_a2sum_dff_n175), .CLK(n9637), .Q(dpath_mulcore_addin_sum[17]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[18](.D(dpath_mulcore_a2sum_dff_n173), .CLK(n9637), .Q(dpath_mulcore_addin_sum[18]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[19](.D(dpath_mulcore_a2sum_dff_n171), .CLK(n9637), .Q(dpath_mulcore_addin_sum[19]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[20](.D(dpath_mulcore_a2sum_dff_n169), .CLK(n9637), .Q(dpath_mulcore_addin_sum[20]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[21](.D(dpath_mulcore_a2sum_dff_n167), .CLK(n9637), .Q(dpath_mulcore_addin_sum[21]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[22](.D(dpath_mulcore_a2sum_dff_n165), .CLK(n9637), .Q(dpath_mulcore_addin_sum[22]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[23](.D(dpath_mulcore_a2sum_dff_n163), .CLK(n9637), .Q(dpath_mulcore_addin_sum[23]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[24](.D(dpath_mulcore_a2sum_dff_n161), .CLK(n9637), .Q(dpath_mulcore_addin_sum[24]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[25](.D(dpath_mulcore_a2sum_dff_n159), .CLK(n9637), .Q(dpath_mulcore_addin_sum[25]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[26](.D(dpath_mulcore_a2sum_dff_n157), .CLK(n9637), .Q(dpath_mulcore_addin_sum[26]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[27](.D(dpath_mulcore_a2sum_dff_n153), .CLK(n9637), .Q(dpath_mulcore_addin_sum[27]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[28](.D(dpath_mulcore_a2sum_dff_n151), .CLK(n9637), .Q(dpath_mulcore_addin_sum[28]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[29](.D(dpath_mulcore_a2sum_dff_n149), .CLK(n9637), .Q(dpath_mulcore_addin_sum[29]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[30](.D(dpath_mulcore_a2sum_dff_n147), .CLK(n9636), .Q(dpath_mulcore_addin_sum[30]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[31](.D(dpath_mulcore_a2sum_dff_n145), .CLK(n9636), .Q(dpath_mulcore_addin_sum[31]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[32](.D(dpath_mulcore_a2sum_dff_n143), .CLK(n9636), .Q(dpath_mulcore_addin_sum[32]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[33](.D(dpath_mulcore_a2sum_dff_n141), .CLK(n9636), .Q(dpath_mulcore_addin_sum[33]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[34](.D(dpath_mulcore_a2sum_dff_n139), .CLK(n9636), .Q(dpath_mulcore_addin_sum[34]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[35](.D(dpath_mulcore_a2sum_dff_n137), .CLK(n9636), .Q(dpath_mulcore_addin_sum[35]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[36](.D(dpath_mulcore_a2sum_dff_n135), .CLK(n9636), .Q(dpath_mulcore_addin_sum[36]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[37](.D(dpath_mulcore_a2sum_dff_n131), .CLK(n9636), .Q(dpath_mulcore_addin_sum[37]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[38](.D(dpath_mulcore_a2sum_dff_n129), .CLK(n9636), .Q(dpath_mulcore_addin_sum[38]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[39](.D(dpath_mulcore_a2sum_dff_n127), .CLK(n9636), .Q(dpath_mulcore_addin_sum[39]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[40](.D(dpath_mulcore_a2sum_dff_n125), .CLK(n9636), .Q(dpath_mulcore_addin_sum[40]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[41](.D(dpath_mulcore_a2sum_dff_n123), .CLK(n9636), .Q(dpath_mulcore_addin_sum[41]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[42](.D(dpath_mulcore_a2sum_dff_n121), .CLK(n9636), .Q(dpath_mulcore_addin_sum[42]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[43](.D(dpath_mulcore_a2sum_dff_n119), .CLK(n9635), .Q(dpath_mulcore_addin_sum[43]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[44](.D(dpath_mulcore_a2sum_dff_n117), .CLK(n9635), .Q(dpath_mulcore_addin_sum[44]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[45](.D(dpath_mulcore_a2sum_dff_n115), .CLK(n9635), .Q(dpath_mulcore_addin_sum[45]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[46](.D(dpath_mulcore_a2sum_dff_n113), .CLK(n9635), .Q(dpath_mulcore_addin_sum[46]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[47](.D(dpath_mulcore_a2sum_dff_n109), .CLK(n9635), .Q(dpath_mulcore_addin_sum[47]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[48](.D(dpath_mulcore_a2sum_dff_n107), .CLK(n9635), .Q(dpath_mulcore_addin_sum[48]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[49](.D(dpath_mulcore_a2sum_dff_n105), .CLK(n9635), .Q(dpath_mulcore_addin_sum[49]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[50](.D(dpath_mulcore_a2sum_dff_n103), .CLK(n9635), .Q(dpath_mulcore_addin_sum[50]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[51](.D(dpath_mulcore_a2sum_dff_n101), .CLK(n9635), .Q(dpath_mulcore_addin_sum[51]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[52](.D(dpath_mulcore_a2sum_dff_n99), .CLK(n9635), .Q(dpath_mulcore_addin_sum[52]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[53](.D(dpath_mulcore_a2sum_dff_n97), .CLK(n9635), .Q(dpath_mulcore_addin_sum[53]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[54](.D(dpath_mulcore_a2sum_dff_n95), .CLK(n9635), .Q(dpath_mulcore_addin_sum[54]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[55](.D(dpath_mulcore_a2sum_dff_n93), .CLK(n9635), .Q(dpath_mulcore_addin_sum[55]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[56](.D(dpath_mulcore_a2sum_dff_n91), .CLK(n9634), .Q(dpath_mulcore_addin_sum[56]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[57](.D(dpath_mulcore_a2sum_dff_n87), .CLK(n9634), .Q(dpath_mulcore_addin_sum[57]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[58](.D(dpath_mulcore_a2sum_dff_n85), .CLK(n9634), .Q(dpath_mulcore_addin_sum[58]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[59](.D(dpath_mulcore_a2sum_dff_n83), .CLK(n9634), .Q(dpath_mulcore_addin_sum[59]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[60](.D(dpath_mulcore_a2sum_dff_n81), .CLK(n9634), .Q(dpath_mulcore_addin_sum[60]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[61](.D(dpath_mulcore_a2sum_dff_n79), .CLK(n9634), .Q(dpath_mulcore_addin_sum[61]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[62](.D(dpath_mulcore_a2sum_dff_n77), .CLK(n9634), .Q(dpath_mulcore_addin_sum[62]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[63](.D(dpath_mulcore_a2sum_dff_n75), .CLK(n9634), .Q(dpath_mulcore_addin_sum[63]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[64](.D(dpath_mulcore_a2sum_dff_n73), .CLK(n9634), .Q(dpath_mulcore_addin_sum[64]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[65](.D(dpath_mulcore_a2sum_dff_n71), .CLK(n9634), .Q(dpath_mulcore_addin_sum[65]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[66](.D(dpath_mulcore_a2sum_dff_n69), .CLK(n9634), .Q(dpath_mulcore_addin_sum[66]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[67](.D(dpath_mulcore_a2sum_dff_n65), .CLK(n9634), .Q(dpath_mulcore_addin_sum[67]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[68](.D(dpath_mulcore_a2sum_dff_n63), .CLK(n9634), .Q(dpath_mulcore_addin_sum[68]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[69](.D(dpath_mulcore_a2sum_dff_n61), .CLK(n9633), .Q(dpath_mulcore_addin_sum[69]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[70](.D(dpath_mulcore_a2sum_dff_n59), .CLK(n9633), .Q(dpath_mulcore_addin_sum[70]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[71](.D(dpath_mulcore_a2sum_dff_n57), .CLK(n9633), .Q(dpath_mulcore_addin_sum[71]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[72](.D(dpath_mulcore_a2sum_dff_n55), .CLK(n9633), .Q(dpath_mulcore_addin_sum[72]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[73](.D(dpath_mulcore_a2sum_dff_n53), .CLK(n9633), .Q(dpath_mulcore_addin_sum[73]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[74](.D(dpath_mulcore_a2sum_dff_n51), .CLK(n9633), .Q(dpath_mulcore_addin_sum[74]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[75](.D(dpath_mulcore_a2sum_dff_n49), .CLK(n9633), .Q(dpath_mulcore_addin_sum[75]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[76](.D(dpath_mulcore_a2sum_dff_n47), .CLK(n9633), .Q(dpath_mulcore_addin_sum[76]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[77](.D(dpath_mulcore_a2sum_dff_n43), .CLK(n9633), .Q(dpath_mulcore_addin_sum[77]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[78](.D(dpath_mulcore_a2sum_dff_n41), .CLK(n9633), .Q(dpath_mulcore_addin_sum[78]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[79](.D(dpath_mulcore_a2sum_dff_n39), .CLK(n9633), .Q(dpath_mulcore_addin_sum[79]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[80](.D(dpath_mulcore_a2sum_dff_n37), .CLK(n9633), .Q(dpath_mulcore_addin_sum[80]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[81](.D(dpath_mulcore_a2sum_dff_n35), .CLK(n9633), .Q(dpath_mulcore_addin_sum[81]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[82](.D(dpath_mulcore_a2sum_dff_n33), .CLK(n9632), .Q(dpath_mulcore_addin_sum[82]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[83](.D(dpath_mulcore_a2sum_dff_n31), .CLK(n9632), .Q(dpath_mulcore_addin_sum[83]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[84](.D(dpath_mulcore_a2sum_dff_n29), .CLK(n9632), .Q(dpath_mulcore_addin_sum[84]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[85](.D(dpath_mulcore_a2sum_dff_n27), .CLK(n9632), .Q(dpath_mulcore_addin_sum[85]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[86](.D(dpath_mulcore_a2sum_dff_n25), .CLK(n9632), .Q(dpath_mulcore_addin_sum[86]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[87](.D(dpath_mulcore_a2sum_dff_n21), .CLK(n9632), .Q(dpath_mulcore_addin_sum[87]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[88](.D(dpath_mulcore_a2sum_dff_n19), .CLK(n9632), .Q(dpath_mulcore_addin_sum[88]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[89](.D(dpath_mulcore_a2sum_dff_n17), .CLK(n9632), .Q(dpath_mulcore_addin_sum[89]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[90](.D(dpath_mulcore_a2sum_dff_n15), .CLK(n9632), .Q(dpath_mulcore_addin_sum[90]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[91](.D(dpath_mulcore_a2sum_dff_n13), .CLK(n9632), .Q(dpath_mulcore_addin_sum[91]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[92](.D(dpath_mulcore_a2sum_dff_n11), .CLK(n9632), .Q(dpath_mulcore_addin_sum[92]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[93](.D(dpath_mulcore_a2sum_dff_n9), .CLK(n9632), .Q(dpath_mulcore_addin_sum[93]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[94](.D(dpath_mulcore_a2sum_dff_n7), .CLK(n9632), .Q(dpath_mulcore_addin_sum[94]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[95](.D(dpath_mulcore_a2sum_dff_n5), .CLK(n9631), .Q(dpath_mulcore_addin_sum[95]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[96](.D(dpath_mulcore_a2sum_dff_n3), .CLK(n9631), .Q(dpath_mulcore_addin_sum[96]));
DFFPOSX1 dpath_mulcore_a2sum_dff_q_reg[97](.D(dpath_mulcore_a2sum_dff_n195), .CLK(n9631), .Q(dpath_mulcore_addin_sum[97]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[0](.D(dpath_mulcore_psum_dff_n97), .CLK(n9631), .Q(dpath_mulcore_ps[31]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[1](.D(dpath_mulcore_psum_dff_n75), .CLK(n9631), .Q(dpath_mulcore_ps[32]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[2](.D(dpath_mulcore_psum_dff_n53), .CLK(n9631), .Q(dpath_mulcore_ps[33]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[3](.D(dpath_mulcore_psum_dff_n31), .CLK(n9631), .Q(dpath_mulcore_ps[34]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[4](.D(dpath_mulcore_psum_dff_n9), .CLK(n9631), .Q(dpath_mulcore_ps[35]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[5](.D(dpath_mulcore_psum_dff_n5), .CLK(n9631), .Q(dpath_mulcore_ps[36]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[6](.D(dpath_mulcore_psum_dff_n3), .CLK(n9631), .Q(dpath_mulcore_ps[37]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[7](.D(dpath_mulcore_psum_dff_n137), .CLK(n9631), .Q(dpath_mulcore_ps[38]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[8](.D(dpath_mulcore_psum_dff_n135), .CLK(n9631), .Q(dpath_mulcore_ps[39]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[9](.D(dpath_mulcore_psum_dff_n133), .CLK(n9631), .Q(dpath_mulcore_ps[40]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[10](.D(dpath_mulcore_psum_dff_n131), .CLK(n9630), .Q(dpath_mulcore_ps[41]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[11](.D(dpath_mulcore_psum_dff_n129), .CLK(n9630), .Q(dpath_mulcore_ps[42]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[12](.D(dpath_mulcore_psum_dff_n127), .CLK(n9630), .Q(dpath_mulcore_ps[43]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[13](.D(dpath_mulcore_psum_dff_n125), .CLK(n9630), .Q(dpath_mulcore_ps[44]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[14](.D(dpath_mulcore_psum_dff_n123), .CLK(n9630), .Q(dpath_mulcore_ps[45]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[15](.D(dpath_mulcore_psum_dff_n121), .CLK(n9630), .Q(dpath_mulcore_ps[46]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[16](.D(dpath_mulcore_psum_dff_n119), .CLK(n9630), .Q(dpath_mulcore_ps[47]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[17](.D(dpath_mulcore_psum_dff_n117), .CLK(n9630), .Q(dpath_mulcore_ps[48]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[18](.D(dpath_mulcore_psum_dff_n115), .CLK(n9630), .Q(dpath_mulcore_ps[49]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[19](.D(dpath_mulcore_psum_dff_n113), .CLK(n9630), .Q(dpath_mulcore_ps[50]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[20](.D(dpath_mulcore_psum_dff_n111), .CLK(n9630), .Q(dpath_mulcore_ps[51]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[21](.D(dpath_mulcore_psum_dff_n109), .CLK(n9630), .Q(dpath_mulcore_ps[52]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[22](.D(dpath_mulcore_psum_dff_n107), .CLK(n9630), .Q(dpath_mulcore_ps[53]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[23](.D(dpath_mulcore_psum_dff_n105), .CLK(n9629), .Q(dpath_mulcore_ps[54]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[24](.D(dpath_mulcore_psum_dff_n103), .CLK(n9629), .Q(dpath_mulcore_ps[55]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[25](.D(dpath_mulcore_psum_dff_n101), .CLK(n9629), .Q(dpath_mulcore_ps[56]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[26](.D(dpath_mulcore_psum_dff_n99), .CLK(n9629), .Q(dpath_mulcore_ps[57]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[27](.D(dpath_mulcore_psum_dff_n95), .CLK(n9629), .Q(dpath_mulcore_ps[58]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[28](.D(dpath_mulcore_psum_dff_n93), .CLK(n9629), .Q(dpath_mulcore_ps[59]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[29](.D(dpath_mulcore_psum_dff_n91), .CLK(n9629), .Q(dpath_mulcore_ps[60]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[30](.D(dpath_mulcore_psum_dff_n89), .CLK(n9629), .Q(dpath_mulcore_ps[61]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[31](.D(dpath_mulcore_psum_dff_n87), .CLK(n9629), .Q(dpath_mulcore_ps[62]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[32](.D(dpath_mulcore_psum_dff_n85), .CLK(n9629), .Q(dpath_mulcore_ps[63]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[33](.D(dpath_mulcore_psum_dff_n83), .CLK(n9629), .Q(dpath_mulcore_ps[64]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[34](.D(dpath_mulcore_psum_dff_n81), .CLK(n9629), .Q(dpath_mulcore_ps[65]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[35](.D(dpath_mulcore_psum_dff_n79), .CLK(n9629), .Q(dpath_mulcore_ps[66]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[36](.D(dpath_mulcore_psum_dff_n77), .CLK(n9628), .Q(dpath_mulcore_ps[67]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[37](.D(dpath_mulcore_psum_dff_n73), .CLK(n9628), .Q(dpath_mulcore_ps[68]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[38](.D(dpath_mulcore_psum_dff_n71), .CLK(n9628), .Q(dpath_mulcore_ps[69]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[39](.D(dpath_mulcore_psum_dff_n69), .CLK(n9628), .Q(dpath_mulcore_ps[70]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[40](.D(dpath_mulcore_psum_dff_n67), .CLK(n9628), .Q(dpath_mulcore_ps[71]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[41](.D(dpath_mulcore_psum_dff_n65), .CLK(n9628), .Q(dpath_mulcore_ps[72]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[42](.D(dpath_mulcore_psum_dff_n63), .CLK(n9628), .Q(dpath_mulcore_ps[73]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[43](.D(dpath_mulcore_psum_dff_n61), .CLK(n9628), .Q(dpath_mulcore_ps[74]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[44](.D(dpath_mulcore_psum_dff_n59), .CLK(n9628), .Q(dpath_mulcore_ps[75]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[45](.D(dpath_mulcore_psum_dff_n57), .CLK(n9628), .Q(dpath_mulcore_ps[76]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[46](.D(dpath_mulcore_psum_dff_n55), .CLK(n9628), .Q(dpath_mulcore_ps[77]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[47](.D(dpath_mulcore_psum_dff_n51), .CLK(n9628), .Q(dpath_mulcore_ps[78]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[48](.D(dpath_mulcore_psum_dff_n49), .CLK(n9628), .Q(dpath_mulcore_ps[79]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[49](.D(dpath_mulcore_psum_dff_n47), .CLK(n9627), .Q(dpath_mulcore_ps[80]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[50](.D(dpath_mulcore_psum_dff_n45), .CLK(n9627), .Q(dpath_mulcore_ps[81]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[51](.D(dpath_mulcore_psum_dff_n43), .CLK(n9627), .Q(dpath_mulcore_ps[82]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[52](.D(dpath_mulcore_psum_dff_n41), .CLK(n9627), .Q(dpath_mulcore_ps[83]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[53](.D(dpath_mulcore_psum_dff_n39), .CLK(n9627), .Q(dpath_mulcore_ps[84]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[54](.D(dpath_mulcore_psum_dff_n37), .CLK(n9627), .Q(dpath_mulcore_ps[85]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[55](.D(dpath_mulcore_psum_dff_n35), .CLK(n9627), .Q(dpath_mulcore_ps[86]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[56](.D(dpath_mulcore_psum_dff_n33), .CLK(n9627), .Q(dpath_mulcore_ps[87]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[57](.D(dpath_mulcore_psum_dff_n29), .CLK(n9627), .Q(dpath_mulcore_ps[88]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[58](.D(dpath_mulcore_psum_dff_n27), .CLK(n9627), .Q(dpath_mulcore_ps[89]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[59](.D(dpath_mulcore_psum_dff_n25), .CLK(n9627), .Q(dpath_mulcore_ps[90]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[60](.D(dpath_mulcore_psum_dff_n23), .CLK(n9627), .Q(dpath_mulcore_ps[91]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[61](.D(dpath_mulcore_psum_dff_n21), .CLK(n9627), .Q(dpath_mulcore_ps[92]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[62](.D(dpath_mulcore_psum_dff_n19), .CLK(n9626), .Q(dpath_mulcore_ps[93]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[63](.D(dpath_mulcore_psum_dff_n17), .CLK(n9626), .Q(dpath_mulcore_ps[94]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[64](.D(dpath_mulcore_psum_dff_n15), .CLK(n9626), .Q(dpath_mulcore_ps[95]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[65](.D(dpath_mulcore_psum_dff_n13), .CLK(n9626), .Q(dpath_mulcore_ps[96]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[66](.D(dpath_mulcore_psum_dff_n11), .CLK(n9626), .Q(dpath_mulcore_ps[97]));
DFFPOSX1 dpath_mulcore_psum_dff_q_reg[67](.D(dpath_mulcore_psum_dff_n7), .CLK(n9626), .Q(dpath_mulcore_ps[98]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[0](.D(dpath_mulcore_pcout_dff_n99), .CLK(n9626), .Q(dpath_mulcore_pc[30]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[1](.D(dpath_mulcore_pcout_dff_n77), .CLK(n9626), .Q(dpath_mulcore_pc[31]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[2](.D(dpath_mulcore_pcout_dff_n55), .CLK(n9626), .Q(dpath_mulcore_pc[32]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[3](.D(dpath_mulcore_pcout_dff_n33), .CLK(n9626), .Q(dpath_mulcore_pc[33]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[4](.D(dpath_mulcore_pcout_dff_n11), .CLK(n9626), .Q(dpath_mulcore_pc[34]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[5](.D(dpath_mulcore_pcout_dff_n5), .CLK(n9626), .Q(dpath_mulcore_pc[35]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[6](.D(dpath_mulcore_pcout_dff_n3), .CLK(n9626), .Q(dpath_mulcore_pc[36]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[7](.D(dpath_mulcore_pcout_dff_n139), .CLK(n9625), .Q(dpath_mulcore_pc[37]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[8](.D(dpath_mulcore_pcout_dff_n137), .CLK(n9625), .Q(dpath_mulcore_pc[38]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[9](.D(dpath_mulcore_pcout_dff_n135), .CLK(n9625), .Q(dpath_mulcore_pc[39]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[10](.D(dpath_mulcore_pcout_dff_n133), .CLK(n9625), .Q(dpath_mulcore_pc[40]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[11](.D(dpath_mulcore_pcout_dff_n131), .CLK(n9625), .Q(dpath_mulcore_pc[41]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[12](.D(dpath_mulcore_pcout_dff_n129), .CLK(n9625), .Q(dpath_mulcore_pc[42]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[13](.D(dpath_mulcore_pcout_dff_n127), .CLK(n9625), .Q(dpath_mulcore_pc[43]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[14](.D(dpath_mulcore_pcout_dff_n125), .CLK(n9625), .Q(dpath_mulcore_pc[44]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[15](.D(dpath_mulcore_pcout_dff_n123), .CLK(n9625), .Q(dpath_mulcore_pc[45]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[16](.D(dpath_mulcore_pcout_dff_n121), .CLK(n9625), .Q(dpath_mulcore_pc[46]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[17](.D(dpath_mulcore_pcout_dff_n119), .CLK(n9625), .Q(dpath_mulcore_pc[47]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[18](.D(dpath_mulcore_pcout_dff_n117), .CLK(n9625), .Q(dpath_mulcore_pc[48]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[19](.D(dpath_mulcore_pcout_dff_n115), .CLK(n9625), .Q(dpath_mulcore_pc[49]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[20](.D(dpath_mulcore_pcout_dff_n113), .CLK(n9624), .Q(dpath_mulcore_pc[50]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[21](.D(dpath_mulcore_pcout_dff_n111), .CLK(n9624), .Q(dpath_mulcore_pc[51]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[22](.D(dpath_mulcore_pcout_dff_n109), .CLK(n9624), .Q(dpath_mulcore_pc[52]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[23](.D(dpath_mulcore_pcout_dff_n107), .CLK(n9624), .Q(dpath_mulcore_pc[53]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[24](.D(dpath_mulcore_pcout_dff_n105), .CLK(n9624), .Q(dpath_mulcore_pc[54]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[25](.D(dpath_mulcore_pcout_dff_n103), .CLK(n9624), .Q(dpath_mulcore_pc[55]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[26](.D(dpath_mulcore_pcout_dff_n101), .CLK(n9624), .Q(dpath_mulcore_pc[56]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[27](.D(dpath_mulcore_pcout_dff_n97), .CLK(n9624), .Q(dpath_mulcore_pc[57]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[28](.D(dpath_mulcore_pcout_dff_n95), .CLK(n9624), .Q(dpath_mulcore_pc[58]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[29](.D(dpath_mulcore_pcout_dff_n93), .CLK(n9624), .Q(dpath_mulcore_pc[59]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[30](.D(dpath_mulcore_pcout_dff_n91), .CLK(n9624), .Q(dpath_mulcore_pc[60]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[31](.D(dpath_mulcore_pcout_dff_n89), .CLK(n9624), .Q(dpath_mulcore_pc[61]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[32](.D(dpath_mulcore_pcout_dff_n87), .CLK(n9624), .Q(dpath_mulcore_pc[62]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[33](.D(dpath_mulcore_pcout_dff_n85), .CLK(n9623), .Q(dpath_mulcore_pc[63]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[34](.D(dpath_mulcore_pcout_dff_n83), .CLK(n9623), .Q(dpath_mulcore_pc[64]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[35](.D(dpath_mulcore_pcout_dff_n81), .CLK(n9623), .Q(dpath_mulcore_pc[65]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[36](.D(dpath_mulcore_pcout_dff_n79), .CLK(n9623), .Q(dpath_mulcore_pc[66]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[37](.D(dpath_mulcore_pcout_dff_n75), .CLK(n9623), .Q(dpath_mulcore_pc[67]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[38](.D(dpath_mulcore_pcout_dff_n73), .CLK(n9623), .Q(dpath_mulcore_pc[68]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[39](.D(dpath_mulcore_pcout_dff_n71), .CLK(n9623), .Q(dpath_mulcore_pc[69]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[40](.D(dpath_mulcore_pcout_dff_n69), .CLK(n9623), .Q(dpath_mulcore_pc[70]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[41](.D(dpath_mulcore_pcout_dff_n67), .CLK(n9623), .Q(dpath_mulcore_pc[71]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[42](.D(dpath_mulcore_pcout_dff_n65), .CLK(n9623), .Q(dpath_mulcore_pc[72]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[43](.D(dpath_mulcore_pcout_dff_n63), .CLK(n9623), .Q(dpath_mulcore_pc[73]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[44](.D(dpath_mulcore_pcout_dff_n61), .CLK(n9623), .Q(dpath_mulcore_pc[74]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[45](.D(dpath_mulcore_pcout_dff_n59), .CLK(n9623), .Q(dpath_mulcore_pc[75]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[46](.D(dpath_mulcore_pcout_dff_n57), .CLK(n9622), .Q(dpath_mulcore_pc[76]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[47](.D(dpath_mulcore_pcout_dff_n53), .CLK(n9622), .Q(dpath_mulcore_pc[77]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[48](.D(dpath_mulcore_pcout_dff_n51), .CLK(n9622), .Q(dpath_mulcore_pc[78]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[49](.D(dpath_mulcore_pcout_dff_n49), .CLK(n9622), .Q(dpath_mulcore_pc[79]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[50](.D(dpath_mulcore_pcout_dff_n47), .CLK(n9622), .Q(dpath_mulcore_pc[80]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[51](.D(dpath_mulcore_pcout_dff_n45), .CLK(n9622), .Q(dpath_mulcore_pc[81]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[52](.D(dpath_mulcore_pcout_dff_n43), .CLK(n9622), .Q(dpath_mulcore_pc[82]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[53](.D(dpath_mulcore_pcout_dff_n41), .CLK(n9622), .Q(dpath_mulcore_pc[83]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[54](.D(dpath_mulcore_pcout_dff_n39), .CLK(n9622), .Q(dpath_mulcore_pc[84]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[55](.D(dpath_mulcore_pcout_dff_n37), .CLK(n9622), .Q(dpath_mulcore_pc[85]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[56](.D(dpath_mulcore_pcout_dff_n35), .CLK(n9622), .Q(dpath_mulcore_pc[86]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[57](.D(dpath_mulcore_pcout_dff_n31), .CLK(n9622), .Q(dpath_mulcore_pc[87]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[58](.D(dpath_mulcore_pcout_dff_n29), .CLK(n9622), .Q(dpath_mulcore_pc[88]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[59](.D(dpath_mulcore_pcout_dff_n27), .CLK(n9621), .Q(dpath_mulcore_pc[89]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[60](.D(dpath_mulcore_pcout_dff_n25), .CLK(n9621), .Q(dpath_mulcore_pc[90]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[61](.D(dpath_mulcore_pcout_dff_n23), .CLK(n9621), .Q(dpath_mulcore_pc[91]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[62](.D(dpath_mulcore_pcout_dff_n21), .CLK(n9621), .Q(dpath_mulcore_pc[92]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[63](.D(dpath_mulcore_pcout_dff_n19), .CLK(n9621), .Q(dpath_mulcore_pc[93]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[64](.D(dpath_mulcore_pcout_dff_n17), .CLK(n9621), .Q(dpath_mulcore_pc[94]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[65](.D(dpath_mulcore_pcout_dff_n15), .CLK(n9621), .Q(dpath_mulcore_pc[95]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[66](.D(dpath_mulcore_pcout_dff_n13), .CLK(n9621), .Q(dpath_mulcore_pc[96]));
DFFPOSX1 dpath_mulcore_pcout_dff_q_reg[67](.D(dpath_mulcore_pcout_dff_n9), .CLK(n9621), .Q(dpath_mulcore_pc[97]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[0](.D(dpath_mulcore_out_dff_n155), .CLK(n9621), .Q(dpath_mout[32]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[1](.D(dpath_mulcore_out_dff_n133), .CLK(n9621), .Q(dpath_mout[33]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[2](.D(dpath_mulcore_out_dff_n111), .CLK(n9621), .Q(dpath_mout[34]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[3](.D(dpath_mulcore_out_dff_n89), .CLK(n9620), .Q(dpath_mout[35]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[4](.D(dpath_mulcore_out_dff_n67), .CLK(n9620), .Q(dpath_mout[36]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[5](.D(dpath_mulcore_out_dff_n45), .CLK(n9620), .Q(dpath_mout[37]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[6](.D(dpath_mulcore_out_dff_n23), .CLK(n9620), .Q(dpath_mout[38]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[7](.D(dpath_mulcore_out_dff_n209), .CLK(n9620), .Q(dpath_mout[39]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[8](.D(dpath_mulcore_out_dff_n193), .CLK(n9620), .Q(dpath_mout[40]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[9](.D(dpath_mulcore_out_dff_n191), .CLK(n9620), .Q(dpath_mout[41]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[10](.D(dpath_mulcore_out_dff_n189), .CLK(n9620), .Q(dpath_mout[42]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[11](.D(dpath_mulcore_out_dff_n187), .CLK(n9620), .Q(dpath_mout[43]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[12](.D(dpath_mulcore_out_dff_n185), .CLK(n9620), .Q(dpath_mout[44]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[13](.D(dpath_mulcore_out_dff_n183), .CLK(n9620), .Q(dpath_mout[45]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[14](.D(dpath_mulcore_out_dff_n181), .CLK(n9620), .Q(dpath_mout[46]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[15](.D(dpath_mulcore_out_dff_n179), .CLK(n9620), .Q(dpath_mout[47]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[16](.D(dpath_mulcore_out_dff_n177), .CLK(n9619), .Q(dpath_mout[48]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[17](.D(dpath_mulcore_out_dff_n175), .CLK(n9619), .Q(dpath_mout[49]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[18](.D(dpath_mulcore_out_dff_n173), .CLK(n9619), .Q(dpath_mout[50]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[19](.D(dpath_mulcore_out_dff_n171), .CLK(n9619), .Q(dpath_mout[51]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[20](.D(dpath_mulcore_out_dff_n169), .CLK(n9619), .Q(dpath_mout[52]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[21](.D(dpath_mulcore_out_dff_n167), .CLK(n9619), .Q(dpath_mout[53]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[22](.D(dpath_mulcore_out_dff_n165), .CLK(n9619), .Q(dpath_mout[54]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[23](.D(dpath_mulcore_out_dff_n163), .CLK(n9619), .Q(dpath_mout[55]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[24](.D(dpath_mulcore_out_dff_n161), .CLK(n9619), .Q(dpath_mout[56]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[25](.D(dpath_mulcore_out_dff_n159), .CLK(n9619), .Q(dpath_mout[57]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[26](.D(dpath_mulcore_out_dff_n157), .CLK(n9619), .Q(dpath_mout[58]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[27](.D(dpath_mulcore_out_dff_n153), .CLK(n9619), .Q(dpath_mout[59]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[28](.D(dpath_mulcore_out_dff_n151), .CLK(n9619), .Q(dpath_mout[60]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[29](.D(dpath_mulcore_out_dff_n149), .CLK(n9618), .Q(dpath_mout[61]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[30](.D(dpath_mulcore_out_dff_n147), .CLK(n9618), .Q(dpath_mout[62]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[31](.D(dpath_mulcore_out_dff_n145), .CLK(n9618), .Q(dpath_mout[63]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[32](.D(dpath_mulcore_out_dff_n143), .CLK(n9618), .Q(dpath_mout[64]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[33](.D(dpath_mulcore_out_dff_n141), .CLK(n9618), .Q(dpath_mout[65]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[34](.D(dpath_mulcore_out_dff_n139), .CLK(n9618), .Q(dpath_mout[66]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[35](.D(dpath_mulcore_out_dff_n137), .CLK(n9618), .Q(dpath_mout[67]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[36](.D(dpath_mulcore_out_dff_n135), .CLK(n9618), .Q(dpath_mout[68]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[37](.D(dpath_mulcore_out_dff_n131), .CLK(n9618), .Q(dpath_mout[69]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[38](.D(dpath_mulcore_out_dff_n129), .CLK(n9618), .Q(dpath_mout[70]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[39](.D(dpath_mulcore_out_dff_n127), .CLK(n9618), .Q(dpath_mout[71]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[40](.D(dpath_mulcore_out_dff_n125), .CLK(n9618), .Q(dpath_mout[72]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[41](.D(dpath_mulcore_out_dff_n123), .CLK(n9618), .Q(dpath_mout[73]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[42](.D(dpath_mulcore_out_dff_n121), .CLK(n9617), .Q(dpath_mout[74]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[43](.D(dpath_mulcore_out_dff_n119), .CLK(n9617), .Q(dpath_mout[75]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[44](.D(dpath_mulcore_out_dff_n117), .CLK(n9617), .Q(dpath_mout[76]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[45](.D(dpath_mulcore_out_dff_n115), .CLK(n9617), .Q(dpath_mout[77]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[46](.D(dpath_mulcore_out_dff_n113), .CLK(n9617), .Q(dpath_mout[78]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[47](.D(dpath_mulcore_out_dff_n109), .CLK(n9617), .Q(dpath_mout[79]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[48](.D(dpath_mulcore_out_dff_n107), .CLK(n9617), .Q(dpath_mout[80]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[49](.D(dpath_mulcore_out_dff_n105), .CLK(n9617), .Q(dpath_mout[81]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[50](.D(dpath_mulcore_out_dff_n103), .CLK(n9617), .Q(dpath_mout[82]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[51](.D(dpath_mulcore_out_dff_n101), .CLK(n9617), .Q(dpath_mout[83]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[52](.D(dpath_mulcore_out_dff_n99), .CLK(n9617), .Q(dpath_mout[84]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[53](.D(dpath_mulcore_out_dff_n97), .CLK(n9617), .Q(dpath_mout[85]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[54](.D(dpath_mulcore_out_dff_n95), .CLK(n9617), .Q(dpath_mout[86]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[55](.D(dpath_mulcore_out_dff_n93), .CLK(n9616), .Q(dpath_mout[87]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[56](.D(dpath_mulcore_out_dff_n91), .CLK(n9616), .Q(dpath_mout[88]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[57](.D(dpath_mulcore_out_dff_n87), .CLK(n9616), .Q(dpath_mout[89]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[58](.D(dpath_mulcore_out_dff_n85), .CLK(n9616), .Q(dpath_mout[90]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[59](.D(dpath_mulcore_out_dff_n83), .CLK(n9616), .Q(dpath_mout[91]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[60](.D(dpath_mulcore_out_dff_n81), .CLK(n9616), .Q(dpath_mout[92]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[61](.D(dpath_mulcore_out_dff_n79), .CLK(n9616), .Q(dpath_mout[93]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[62](.D(dpath_mulcore_out_dff_n77), .CLK(n9616), .Q(dpath_mout[94]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[63](.D(dpath_mulcore_out_dff_n75), .CLK(n9616), .Q(dpath_mout[95]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[64](.D(dpath_mulcore_out_dff_n73), .CLK(n9616), .Q(dpath_mout[96]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[65](.D(dpath_mulcore_out_dff_n71), .CLK(n9616), .Q(dpath_mout[97]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[66](.D(dpath_mulcore_out_dff_n69), .CLK(n9616), .Q(dpath_mout[98]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[67](.D(dpath_mulcore_out_dff_n65), .CLK(n9616), .Q(dpath_mout[99]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[68](.D(dpath_mulcore_out_dff_n63), .CLK(n9615), .Q(dpath_mout[100]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[69](.D(dpath_mulcore_out_dff_n61), .CLK(n9615), .Q(dpath_mout[101]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[70](.D(dpath_mulcore_out_dff_n59), .CLK(n9615), .Q(dpath_mout[102]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[71](.D(dpath_mulcore_out_dff_n57), .CLK(n9615), .Q(dpath_mout[103]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[72](.D(dpath_mulcore_out_dff_n55), .CLK(n9615), .Q(dpath_mout[104]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[73](.D(dpath_mulcore_out_dff_n53), .CLK(n9615), .Q(dpath_mout[105]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[74](.D(dpath_mulcore_out_dff_n51), .CLK(n9615), .Q(dpath_mout[106]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[75](.D(dpath_mulcore_out_dff_n49), .CLK(n9615), .Q(dpath_mout[107]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[76](.D(dpath_mulcore_out_dff_n47), .CLK(n9615), .Q(dpath_mout[108]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[77](.D(dpath_mulcore_out_dff_n43), .CLK(n9615), .Q(dpath_mout[109]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[78](.D(dpath_mulcore_out_dff_n41), .CLK(n9615), .Q(dpath_mout[110]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[79](.D(dpath_mulcore_out_dff_n39), .CLK(n9615), .Q(dpath_mout[111]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[80](.D(dpath_mulcore_out_dff_n37), .CLK(n9615), .Q(dpath_mout[112]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[81](.D(dpath_mulcore_out_dff_n35), .CLK(n9614), .Q(dpath_mout[113]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[82](.D(dpath_mulcore_out_dff_n33), .CLK(n9614), .Q(dpath_mout[114]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[83](.D(dpath_mulcore_out_dff_n31), .CLK(n9614), .Q(dpath_mout[115]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[84](.D(dpath_mulcore_out_dff_n29), .CLK(n9614), .Q(dpath_mout[116]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[85](.D(dpath_mulcore_out_dff_n27), .CLK(n9614), .Q(dpath_mout[117]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[86](.D(dpath_mulcore_out_dff_n25), .CLK(n9614), .Q(dpath_mout[118]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[87](.D(dpath_mulcore_out_dff_n21), .CLK(n9614), .Q(dpath_mout[119]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[88](.D(dpath_mulcore_out_dff_n19), .CLK(n9614), .Q(dpath_mout[120]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[89](.D(dpath_mulcore_out_dff_n17), .CLK(n9614), .Q(dpath_mout[121]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[90](.D(dpath_mulcore_out_dff_n15), .CLK(n9614), .Q(dpath_mout[122]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[91](.D(dpath_mulcore_out_dff_n13), .CLK(n9614), .Q(dpath_mout[123]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[92](.D(dpath_mulcore_out_dff_n11), .CLK(n9614), .Q(dpath_mout[124]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[93](.D(dpath_mulcore_out_dff_n9), .CLK(n9614), .Q(dpath_mout[125]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[94](.D(dpath_mulcore_out_dff_n7), .CLK(n9613), .Q(dpath_mout[126]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[95](.D(dpath_mulcore_out_dff_n5), .CLK(n9613), .Q(dpath_mout[127]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[96](.D(dpath_mulcore_out_dff_n3), .CLK(n9613), .Q(dpath_mout[128]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[97](.D(dpath_mulcore_out_dff_n207), .CLK(n9613), .Q(dpath_mout[129]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[98](.D(dpath_mulcore_out_dff_n205), .CLK(n9613), .Q(dpath_mout[130]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[99](.D(dpath_mulcore_out_dff_n203), .CLK(n9613), .Q(dpath_mout[131]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[100](.D(dpath_mulcore_out_dff_n201), .CLK(n9613), .Q(dpath_mout[132]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[101](.D(dpath_mulcore_out_dff_n199), .CLK(n9613), .Q(dpath_mout[133]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[102](.D(dpath_mulcore_out_dff_n197), .CLK(n9613), .Q(dpath_mout[134]));
DFFPOSX1 dpath_mulcore_out_dff_q_reg[103](.D(dpath_mulcore_out_dff_n195), .CLK(n9613), .Q(dpath_mout[135]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[0](.D(dpath_mulcore_pip_dff_n25), .CLK(n9613), .Q(dpath_mout[0]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[1](.D(dpath_mulcore_pip_dff_n13), .CLK(n9613), .Q(dpath_mout[1]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[2](.D(dpath_mulcore_pip_dff_n11), .CLK(n9613), .Q(dpath_mout[2]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[3](.D(dpath_mulcore_pip_dff_n9), .CLK(n9612), .Q(dpath_mout[3]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[4](.D(dpath_mulcore_pip_dff_n7), .CLK(n9612), .Q(dpath_mout[4]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[5](.D(dpath_mulcore_pip_dff_n5), .CLK(n9612), .Q(dpath_mout[5]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[6](.D(dpath_mulcore_pip_dff_n3), .CLK(n9612), .Q(dpath_mout[6]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[7](.D(dpath_mulcore_pip_dff_n65), .CLK(n9612), .Q(dpath_mout[7]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[8](.D(dpath_mulcore_pip_dff_n63), .CLK(n9612), .Q(dpath_mout[8]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[9](.D(dpath_mulcore_pip_dff_n61), .CLK(n9612), .Q(dpath_mout[9]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[10](.D(dpath_mulcore_pip_dff_n59), .CLK(n9612), .Q(dpath_mout[10]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[11](.D(dpath_mulcore_pip_dff_n57), .CLK(n9612), .Q(dpath_mout[11]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[12](.D(dpath_mulcore_pip_dff_n55), .CLK(n9612), .Q(dpath_mout[12]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[13](.D(dpath_mulcore_pip_dff_n53), .CLK(n9612), .Q(dpath_mout[13]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[14](.D(dpath_mulcore_pip_dff_n51), .CLK(n9612), .Q(dpath_mout[14]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[15](.D(dpath_mulcore_pip_dff_n49), .CLK(n9612), .Q(dpath_mout[15]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[16](.D(dpath_mulcore_pip_dff_n47), .CLK(n9611), .Q(dpath_mout[16]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[17](.D(dpath_mulcore_pip_dff_n45), .CLK(n9611), .Q(dpath_mout[17]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[18](.D(dpath_mulcore_pip_dff_n43), .CLK(n9611), .Q(dpath_mout[18]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[19](.D(dpath_mulcore_pip_dff_n41), .CLK(n9611), .Q(dpath_mout[19]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[20](.D(dpath_mulcore_pip_dff_n39), .CLK(n9611), .Q(dpath_mout[20]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[21](.D(dpath_mulcore_pip_dff_n37), .CLK(n9611), .Q(dpath_mout[21]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[22](.D(dpath_mulcore_pip_dff_n35), .CLK(n9611), .Q(dpath_mout[22]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[23](.D(dpath_mulcore_pip_dff_n33), .CLK(n9611), .Q(dpath_mout[23]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[24](.D(dpath_mulcore_pip_dff_n31), .CLK(n9611), .Q(dpath_mout[24]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[25](.D(dpath_mulcore_pip_dff_n29), .CLK(n9611), .Q(dpath_mout[25]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[26](.D(dpath_mulcore_pip_dff_n27), .CLK(n9611), .Q(dpath_mout[26]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[27](.D(dpath_mulcore_pip_dff_n23), .CLK(n9611), .Q(dpath_mout[27]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[28](.D(dpath_mulcore_pip_dff_n21), .CLK(n9611), .Q(dpath_mout[28]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[29](.D(dpath_mulcore_pip_dff_n19), .CLK(n9610), .Q(dpath_mout[29]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[30](.D(dpath_mulcore_pip_dff_n17), .CLK(n9610), .Q(dpath_mout[30]));
DFFPOSX1 dpath_mulcore_pip_dff_q_reg[31](.D(dpath_mulcore_pip_dff_n15), .CLK(n9610), .Q(dpath_mout[31]));
DFFPOSX1 dpath_mulcore_booth_out_dff0_q_reg[0](.D(dpath_mulcore_booth_out_dff0_n7), .CLK(n9584), .Q(dpath_mulcore_b0[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff0_q_reg[1](.D(dpath_mulcore_booth_out_dff0_n5), .CLK(n9584), .Q(dpath_mulcore_b0[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff0_q_reg[2](.D(dpath_mulcore_booth_out_dff0_n3), .CLK(n9584), .Q(dpath_mulcore_b0[2]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_71__U12(.A(dpath_mulcore_ary1_a0_sc3_71__n8), .B(dpath_mulcore_ary1_a0_sc3_71__n7), .Y(dpath_mulcore_ary1_a0_sc3_71__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_71__U11(.A(dpath_mulcore_ary1_a0_s_2[71]), .B(dpath_mulcore_ary1_a0_s1[65]), .Y(dpath_mulcore_ary1_a0_sc3_71__n7));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_71__U10(.A(dpath_mulcore_ary1_a0_s1[64]), .B(n9147), .Y(dpath_mulcore_ary1_a0_sc3_71__n8));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_71__U9(.A(n7227), .B(dpath_mulcore_ary1_a0_sc3_71__z), .Y(dpath_mulcore_a0sum[71]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_70__U4(.A(n13754), .B(n13755), .Y(dpath_mulcore_ary1_a0_sc2_2_70__n1));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_70__U1(.A(n8068), .B(dpath_mulcore_ary1_a0_sc2_2_70__n1), .Y(dpath_mulcore_ary1_a0_s_2[70]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_10__U2(.A(n7203), .B(dpath_mulcore_ary1_a0_s0[10]), .Y(dpath_mulcore_ary1_a0_s_1[10]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_U4(.A(n9854), .B(n7416), .Y(dpath_mulcore_ary1_a0_s2[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff16_q_reg[0](.D(n18337), .CLK(n9584), .Q(dpath_mulcore_b16));
DFFPOSX1 dpath_mulcore_booth_hld_dff0_q_reg[0](.D(n18336), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b[31]));
DFFPOSX1 dpath_mulcore_co31_dff_q_reg[0](.D(n18335), .CLK(n9610), .Q(dpath_mulcore_addin_cin));
LATCH dpath_mulcore_booth_ckbuf_1_clken_reg(.D(n9785), .CLK(n3), .Q(dpath_mulcore_booth_ckbuf_1_clken));
LATCH dpath_mulcore_ckbuf_1_clken_reg(.D(n9785), .CLK(n3), .Q(dpath_mulcore_ckbuf_1_clken));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[0](.D(n18314), .CLK(n9590), .Q(dpath_mulcore_booth_b[32]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[1](.D(n18308), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b0_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[2](.D(n18307), .CLK(n9590), .Q(dpath_mulcore_booth_b[34]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[3](.D(n18306), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b1_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[4](.D(n18305), .CLK(n9590), .Q(dpath_mulcore_booth_b[36]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[5](.D(n18304), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b2_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[6](.D(n18303), .CLK(n9590), .Q(dpath_mulcore_booth_b[38]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[7](.D(n18334), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b3_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[8](.D(n18333), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b[40]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[9](.D(n18332), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b4_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[10](.D(n18331), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b[42]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[11](.D(n18330), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b5_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[12](.D(n18329), .CLK(n9590), .Q(dpath_mulcore_booth_b[44]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[13](.D(n18328), .CLK(n9590), .Q(dpath_mulcore_booth_b6_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[14](.D(n18327), .CLK(n9590), .Q(dpath_mulcore_booth_b[46]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[15](.D(n18326), .CLK(n9590), .Q(dpath_mulcore_booth_b7_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[16](.D(n18325), .CLK(n9590), .Q(dpath_mulcore_booth_b[48]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[17](.D(n18324), .CLK(n9590), .Q(dpath_mulcore_booth_b8_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[18](.D(n18323), .CLK(n9590), .Q(dpath_mulcore_booth_b[50]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[19](.D(n18322), .CLK(n9590), .Q(dpath_mulcore_booth_b9_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[20](.D(n18321), .CLK(n9590), .Q(dpath_mulcore_booth_b[52]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[21](.D(n18320), .CLK(n9590), .Q(dpath_mulcore_booth_b10_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[22](.D(n18319), .CLK(n9590), .Q(dpath_mulcore_booth_b[54]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[23](.D(n18318), .CLK(n9590), .Q(dpath_mulcore_booth_b11_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[24](.D(n18317), .CLK(n9590), .Q(dpath_mulcore_booth_b[56]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[25](.D(n18316), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b12_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[26](.D(n18315), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b[58]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[27](.D(n18313), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b13_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[28](.D(n18312), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b[60]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[29](.D(n18311), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b14_in1[2]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[30](.D(n18310), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b[62]));
DFFPOSX1 dpath_mulcore_booth_hld_dff_q_reg[31](.D(n18309), .CLK(dpath_mulcore_booth_clk_enb1), .Q(dpath_mulcore_booth_b15_in1[2]));
DFFPOSX1 dpath_mulcore_x2c3_dff_q_reg[0](.D(n18302), .CLK(n9610), .Q(dpath_mulcore_x2_c3));
DFFPOSX1 dpath_mulcore_x2c2_dff_q_reg[0](.D(n18301), .CLK(n9610), .Q(dpath_mulcore_x2_c2));
DFFPOSX1 dpath_mulcore_x2c1_dff_q_reg[0](.D(n18300), .CLK(n9610), .Q(dpath_mulcore_x2_c1));
DFFPOSX1 dpath_mulcore_cyc3_dff_q_reg[0](.D(n18299), .CLK(n9610), .Q(dpath_mulcore_psum[98]));
DFFPOSX1 dpath_mulcore_cyc2_dff_q_reg[0](.D(n18298), .CLK(n9610), .Q(dpath_mulcore_cyc2));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[0](.D(n18277), .CLK(n9610), .Q(dpath_mulcore_a1c[4]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[1](.D(n18266), .CLK(n9610), .Q(dpath_mulcore_a1c[5]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[2](.D(n18255), .CLK(n9610), .Q(dpath_mulcore_a1c[6]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[3](.D(n18244), .CLK(n9610), .Q(dpath_mulcore_a1c[7]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[4](.D(n18233), .CLK(n9609), .Q(dpath_mulcore_a1c[8]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[5](.D(n18222), .CLK(n9609), .Q(dpath_mulcore_a1c[9]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[6](.D(n18221), .CLK(n9609), .Q(dpath_mulcore_a1c[10]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[7](.D(n18297), .CLK(n9609), .Q(dpath_mulcore_a1c[11]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[8](.D(n18296), .CLK(n9609), .Q(dpath_mulcore_a1c[12]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[9](.D(n18295), .CLK(n9609), .Q(dpath_mulcore_a1c[13]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[10](.D(n18294), .CLK(n9609), .Q(dpath_mulcore_a1c[14]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[11](.D(n18293), .CLK(n9609), .Q(dpath_mulcore_a1c[15]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[12](.D(n18292), .CLK(n9609), .Q(dpath_mulcore_a1c[16]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[13](.D(n18291), .CLK(n9609), .Q(dpath_mulcore_a1c[17]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[14](.D(n18290), .CLK(n9609), .Q(dpath_mulcore_a1c[18]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[15](.D(n18289), .CLK(n9609), .Q(dpath_mulcore_a1c[19]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[16](.D(n18288), .CLK(n9609), .Q(dpath_mulcore_a1c[20]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[17](.D(n18287), .CLK(n9608), .Q(dpath_mulcore_a1c[21]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[18](.D(n18286), .CLK(n9608), .Q(dpath_mulcore_a1c[22]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[19](.D(n18285), .CLK(n9608), .Q(dpath_mulcore_a1c[23]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[20](.D(n18284), .CLK(n9608), .Q(dpath_mulcore_a1c[24]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[21](.D(n18283), .CLK(n9608), .Q(dpath_mulcore_a1c[25]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[22](.D(n18282), .CLK(n9608), .Q(dpath_mulcore_a1c[26]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[23](.D(n18281), .CLK(n9608), .Q(dpath_mulcore_a1c[27]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[24](.D(n18280), .CLK(n9608), .Q(dpath_mulcore_a1c[28]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[25](.D(n18279), .CLK(n9608), .Q(dpath_mulcore_a1c[29]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[26](.D(n18278), .CLK(n9608), .Q(dpath_mulcore_a1c[30]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[27](.D(n18276), .CLK(n9608), .Q(dpath_mulcore_a1c[31]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[28](.D(n18275), .CLK(n9608), .Q(dpath_mulcore_a1c[32]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[29](.D(n18274), .CLK(n9608), .Q(dpath_mulcore_a1c[33]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[30](.D(n18273), .CLK(n9607), .Q(dpath_mulcore_a1c[34]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[31](.D(n18272), .CLK(n9607), .Q(dpath_mulcore_a1c[35]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[32](.D(n18271), .CLK(n9607), .Q(dpath_mulcore_a1c[36]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[33](.D(n18270), .CLK(n9607), .Q(dpath_mulcore_a1c[37]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[34](.D(n18269), .CLK(n9607), .Q(dpath_mulcore_a1c[38]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[35](.D(n18268), .CLK(n9607), .Q(dpath_mulcore_a1c[39]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[36](.D(n18267), .CLK(n9607), .Q(dpath_mulcore_a1c[40]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[37](.D(n18265), .CLK(n9607), .Q(dpath_mulcore_a1c[41]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[38](.D(n18264), .CLK(n9607), .Q(dpath_mulcore_a1c[42]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[39](.D(n18263), .CLK(n9607), .Q(dpath_mulcore_a1c[43]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[40](.D(n18262), .CLK(n9607), .Q(dpath_mulcore_a1c[44]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[41](.D(n18261), .CLK(n9607), .Q(dpath_mulcore_a1c[45]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[42](.D(n18260), .CLK(n9607), .Q(dpath_mulcore_a1c[46]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[43](.D(n18259), .CLK(n9606), .Q(dpath_mulcore_a1c[47]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[44](.D(n18258), .CLK(n9606), .Q(dpath_mulcore_a1c[48]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[45](.D(n18257), .CLK(n9606), .Q(dpath_mulcore_a1c[49]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[46](.D(n18256), .CLK(n9606), .Q(dpath_mulcore_a1c[50]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[47](.D(n18254), .CLK(n9606), .Q(dpath_mulcore_a1c[51]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[48](.D(n18253), .CLK(n9606), .Q(dpath_mulcore_a1c[52]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[49](.D(n18252), .CLK(n9606), .Q(dpath_mulcore_a1c[53]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[50](.D(n18251), .CLK(n9606), .Q(dpath_mulcore_a1c[54]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[51](.D(n18250), .CLK(n9606), .Q(dpath_mulcore_a1c[55]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[52](.D(n18249), .CLK(n9606), .Q(dpath_mulcore_a1c[56]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[53](.D(n18248), .CLK(n9606), .Q(dpath_mulcore_a1c[57]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[54](.D(n18247), .CLK(n9606), .Q(dpath_mulcore_a1c[58]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[55](.D(n18246), .CLK(n9606), .Q(dpath_mulcore_a1c[59]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[56](.D(n18245), .CLK(n9605), .Q(dpath_mulcore_a1c[60]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[57](.D(n18243), .CLK(n9605), .Q(dpath_mulcore_a1c[61]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[58](.D(n18242), .CLK(n9605), .Q(dpath_mulcore_a1c[62]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[59](.D(n18241), .CLK(n9605), .Q(dpath_mulcore_a1c[63]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[60](.D(n18240), .CLK(n9605), .Q(dpath_mulcore_a1c[64]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[61](.D(n18239), .CLK(n9605), .Q(dpath_mulcore_a1c[65]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[62](.D(n18238), .CLK(n9605), .Q(dpath_mulcore_a1c[66]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[63](.D(n18237), .CLK(n9605), .Q(dpath_mulcore_a1c[67]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[64](.D(n18236), .CLK(n9605), .Q(dpath_mulcore_a1c[68]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[65](.D(n18235), .CLK(n9605), .Q(dpath_mulcore_a1c[69]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[66](.D(n18234), .CLK(n9605), .Q(dpath_mulcore_a1c[70]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[67](.D(n18232), .CLK(n9605), .Q(dpath_mulcore_a1c[71]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[68](.D(n18231), .CLK(n9605), .Q(dpath_mulcore_a1c[72]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[69](.D(n18230), .CLK(n9604), .Q(dpath_mulcore_a1c[73]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[70](.D(n18229), .CLK(n9604), .Q(dpath_mulcore_a1c[74]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[71](.D(n18228), .CLK(n9604), .Q(dpath_mulcore_a1c[75]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[72](.D(n18227), .CLK(n9604), .Q(dpath_mulcore_a1c[76]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[73](.D(n18226), .CLK(n9604), .Q(dpath_mulcore_a1c[77]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[74](.D(n18225), .CLK(n9604), .Q(dpath_mulcore_a1c[78]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[75](.D(n18224), .CLK(n9604), .Q(dpath_mulcore_a1c[79]));
DFFPOSX1 dpath_mulcore_a1cot_dff_q_reg[76](.D(n18223), .CLK(n9604), .Q(dpath_mulcore_a1c[80]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[0](.D(n18200), .CLK(n9604), .Q(dpath_mulcore_a1s[0]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[1](.D(n18189), .CLK(n9604), .Q(dpath_mulcore_a1s[1]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[2](.D(n18178), .CLK(n9604), .Q(dpath_mulcore_a1s[2]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[3](.D(n18167), .CLK(n9604), .Q(dpath_mulcore_a1s[3]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[4](.D(n18156), .CLK(n9603), .Q(dpath_mulcore_a1s[4]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[5](.D(n18145), .CLK(n9603), .Q(dpath_mulcore_a1s[5]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[6](.D(n18139), .CLK(n9603), .Q(dpath_mulcore_a1s[6]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[7](.D(n18220), .CLK(n9603), .Q(dpath_mulcore_a1s[7]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[8](.D(n18219), .CLK(n9603), .Q(dpath_mulcore_a1s[8]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[9](.D(n18218), .CLK(n9603), .Q(dpath_mulcore_a1s[9]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[10](.D(n18217), .CLK(n9603), .Q(dpath_mulcore_a1s[10]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[11](.D(n18216), .CLK(n9603), .Q(dpath_mulcore_a1s[11]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[12](.D(n18215), .CLK(n9603), .Q(dpath_mulcore_a1s[12]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[13](.D(n18214), .CLK(n9603), .Q(dpath_mulcore_a1s[13]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[14](.D(n18213), .CLK(n9603), .Q(dpath_mulcore_a1s[14]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[15](.D(n18212), .CLK(n9603), .Q(dpath_mulcore_a1s[15]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[16](.D(n18211), .CLK(n9603), .Q(dpath_mulcore_a1s[16]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[17](.D(n18210), .CLK(n9602), .Q(dpath_mulcore_a1s[17]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[18](.D(n18209), .CLK(n9602), .Q(dpath_mulcore_a1s[18]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[19](.D(n18208), .CLK(n9602), .Q(dpath_mulcore_a1s[19]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[20](.D(n18207), .CLK(n9602), .Q(dpath_mulcore_a1s[20]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[21](.D(n18206), .CLK(n9602), .Q(dpath_mulcore_a1s[21]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[22](.D(n18205), .CLK(n9602), .Q(dpath_mulcore_a1s[22]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[23](.D(n18204), .CLK(n9602), .Q(dpath_mulcore_a1s[23]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[24](.D(n18203), .CLK(n9602), .Q(dpath_mulcore_a1s[24]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[25](.D(n18202), .CLK(n9602), .Q(dpath_mulcore_a1s[25]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[26](.D(n18201), .CLK(n9602), .Q(dpath_mulcore_a1s[26]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[27](.D(n18199), .CLK(n9602), .Q(dpath_mulcore_a1s[27]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[28](.D(n18198), .CLK(n9602), .Q(dpath_mulcore_a1s[28]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[29](.D(n18197), .CLK(n9602), .Q(dpath_mulcore_a1s[29]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[30](.D(n18196), .CLK(n9601), .Q(dpath_mulcore_a1s[30]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[31](.D(n18195), .CLK(n9601), .Q(dpath_mulcore_a1s[31]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[32](.D(n18194), .CLK(n9601), .Q(dpath_mulcore_a1s[32]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[33](.D(n18193), .CLK(n9601), .Q(dpath_mulcore_a1s[33]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[34](.D(n18192), .CLK(n9601), .Q(dpath_mulcore_a1s[34]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[35](.D(n18191), .CLK(n9601), .Q(dpath_mulcore_a1s[35]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[36](.D(n18190), .CLK(n9601), .Q(dpath_mulcore_a1s[36]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[37](.D(n18188), .CLK(n9601), .Q(dpath_mulcore_a1s[37]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[38](.D(n18187), .CLK(n9601), .Q(dpath_mulcore_a1s[38]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[39](.D(n18186), .CLK(n9601), .Q(dpath_mulcore_a1s[39]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[40](.D(n18185), .CLK(n9601), .Q(dpath_mulcore_a1s[40]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[41](.D(n18184), .CLK(n9601), .Q(dpath_mulcore_a1s[41]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[42](.D(n18183), .CLK(n9601), .Q(dpath_mulcore_a1s[42]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[43](.D(n18182), .CLK(n9600), .Q(dpath_mulcore_a1s[43]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[44](.D(n18181), .CLK(n9600), .Q(dpath_mulcore_a1s[44]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[45](.D(n18180), .CLK(n9600), .Q(dpath_mulcore_a1s[45]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[46](.D(n18179), .CLK(n9600), .Q(dpath_mulcore_a1s[46]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[47](.D(n18177), .CLK(n9600), .Q(dpath_mulcore_a1s[47]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[48](.D(n18176), .CLK(n9600), .Q(dpath_mulcore_a1s[48]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[49](.D(n18175), .CLK(n9600), .Q(dpath_mulcore_a1s[49]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[50](.D(n18174), .CLK(n9600), .Q(dpath_mulcore_a1s[50]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[51](.D(n18173), .CLK(n9600), .Q(dpath_mulcore_a1s[51]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[52](.D(n18172), .CLK(n9600), .Q(dpath_mulcore_a1s[52]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[53](.D(n18171), .CLK(n9600), .Q(dpath_mulcore_a1s[53]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[54](.D(n18170), .CLK(n9600), .Q(dpath_mulcore_a1s[54]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[55](.D(n18169), .CLK(n9600), .Q(dpath_mulcore_a1s[55]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[56](.D(n18168), .CLK(n9599), .Q(dpath_mulcore_a1s[56]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[57](.D(n18166), .CLK(n9599), .Q(dpath_mulcore_a1s[57]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[58](.D(n18165), .CLK(n9599), .Q(dpath_mulcore_a1s[58]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[59](.D(n18164), .CLK(n9599), .Q(dpath_mulcore_a1s[59]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[60](.D(n18163), .CLK(n9599), .Q(dpath_mulcore_a1s[60]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[61](.D(n18162), .CLK(n9599), .Q(dpath_mulcore_a1s[61]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[62](.D(n18161), .CLK(n9599), .Q(dpath_mulcore_a1s[62]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[63](.D(n18160), .CLK(n9599), .Q(dpath_mulcore_a1s[63]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[64](.D(n18159), .CLK(n9599), .Q(dpath_mulcore_a1s[64]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[65](.D(n18158), .CLK(n9599), .Q(dpath_mulcore_a1s[65]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[66](.D(n18157), .CLK(n9599), .Q(dpath_mulcore_a1s[66]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[67](.D(n18155), .CLK(n9599), .Q(dpath_mulcore_a1s[67]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[68](.D(n18154), .CLK(n9599), .Q(dpath_mulcore_a1s[68]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[69](.D(n18153), .CLK(n9598), .Q(dpath_mulcore_a1s[69]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[70](.D(n18152), .CLK(n9598), .Q(dpath_mulcore_a1s[70]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[71](.D(n18151), .CLK(n9598), .Q(dpath_mulcore_a1s[71]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[72](.D(n18150), .CLK(n9598), .Q(dpath_mulcore_a1s[72]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[73](.D(n18149), .CLK(n9598), .Q(dpath_mulcore_a1s[73]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[74](.D(n18148), .CLK(n9598), .Q(dpath_mulcore_a1s[74]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[75](.D(n18147), .CLK(n9598), .Q(dpath_mulcore_a1s[75]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[76](.D(n18146), .CLK(n9598), .Q(dpath_mulcore_a1s[76]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[77](.D(n18144), .CLK(n9598), .Q(dpath_mulcore_a1s[77]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[78](.D(n18143), .CLK(n9598), .Q(dpath_mulcore_a1s[78]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[79](.D(n18142), .CLK(n9598), .Q(dpath_mulcore_a1s[79]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[80](.D(n18141), .CLK(n9598), .Q(dpath_mulcore_a1s[80]));
DFFPOSX1 dpath_mulcore_a1sum_dff_q_reg[81](.D(n18140), .CLK(n9598), .Q(dpath_mulcore_a1s[81]));
DFFPOSX1 dpath_mulcore_booth_out_dff15_q_reg[0](.D(n17857), .CLK(n9584), .Q(dpath_mulcore_b15[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff15_q_reg[1](.D(n17856), .CLK(n9584), .Q(dpath_mulcore_b15[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff15_q_reg[2](.D(n17855), .CLK(n9584), .Q(dpath_mulcore_b15[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff14_q_reg[0](.D(n17854), .CLK(n9584), .Q(dpath_mulcore_b14[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff14_q_reg[1](.D(n17853), .CLK(n9584), .Q(dpath_mulcore_b14[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff14_q_reg[2](.D(n17852), .CLK(n9584), .Q(dpath_mulcore_b14[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff13_q_reg[0](.D(n17851), .CLK(n9584), .Q(dpath_mulcore_b13[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff13_q_reg[1](.D(n17850), .CLK(n9584), .Q(dpath_mulcore_b13[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff13_q_reg[2](.D(n17849), .CLK(n9584), .Q(dpath_mulcore_b13[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff12_q_reg[0](.D(n17848), .CLK(n9585), .Q(dpath_mulcore_b12[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff12_q_reg[1](.D(n17847), .CLK(n9585), .Q(dpath_mulcore_b12[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff12_q_reg[2](.D(n17846), .CLK(n9585), .Q(dpath_mulcore_b12[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff11_q_reg[0](.D(n17845), .CLK(n9585), .Q(dpath_mulcore_b11[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff11_q_reg[1](.D(n17844), .CLK(n9585), .Q(dpath_mulcore_b11[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff11_q_reg[2](.D(n17843), .CLK(n9585), .Q(dpath_mulcore_b11[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff10_q_reg[0](.D(n17842), .CLK(n9585), .Q(dpath_mulcore_b10[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff10_q_reg[1](.D(n17841), .CLK(n9585), .Q(dpath_mulcore_b10[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff10_q_reg[2](.D(n17840), .CLK(n9585), .Q(dpath_mulcore_b10[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff9_q_reg[0](.D(n17839), .CLK(n9585), .Q(dpath_mulcore_b9[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff9_q_reg[1](.D(n17838), .CLK(n9585), .Q(dpath_mulcore_b9[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff9_q_reg[2](.D(n17837), .CLK(n9585), .Q(dpath_mulcore_b9[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff8_q_reg[0](.D(n17836), .CLK(n9585), .Q(dpath_mulcore_b8[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff8_q_reg[1](.D(n17835), .CLK(n9586), .Q(dpath_mulcore_b8[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff8_q_reg[2](.D(n17834), .CLK(n9586), .Q(dpath_mulcore_b8[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff7_q_reg[0](.D(n17833), .CLK(n9586), .Q(dpath_mulcore_b7[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff7_q_reg[1](.D(n17832), .CLK(n9586), .Q(dpath_mulcore_b7[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff7_q_reg[2](.D(n17831), .CLK(n9586), .Q(dpath_mulcore_b7[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff6_q_reg[0](.D(n17830), .CLK(n9586), .Q(dpath_mulcore_b6[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff6_q_reg[1](.D(n17829), .CLK(n9586), .Q(dpath_mulcore_b6[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff6_q_reg[2](.D(n17828), .CLK(n9586), .Q(dpath_mulcore_b6[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff5_q_reg[0](.D(n17827), .CLK(n9586), .Q(dpath_mulcore_b5[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff5_q_reg[1](.D(n17826), .CLK(n9586), .Q(dpath_mulcore_b5[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff5_q_reg[2](.D(n17825), .CLK(n9586), .Q(dpath_mulcore_b5[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff4_q_reg[0](.D(n17824), .CLK(n9586), .Q(dpath_mulcore_b4[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff4_q_reg[1](.D(n17823), .CLK(n9586), .Q(dpath_mulcore_b4[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff4_q_reg[2](.D(n17822), .CLK(n9587), .Q(dpath_mulcore_b4[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff3_q_reg[0](.D(n17821), .CLK(n9587), .Q(dpath_mulcore_b3[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff3_q_reg[1](.D(n17820), .CLK(n9587), .Q(dpath_mulcore_b3[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff3_q_reg[2](.D(n17819), .CLK(n9587), .Q(dpath_mulcore_b3[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff2_q_reg[0](.D(n17818), .CLK(n9587), .Q(dpath_mulcore_b2[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff2_q_reg[1](.D(n17817), .CLK(n9587), .Q(dpath_mulcore_b2[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff2_q_reg[2](.D(n17816), .CLK(n9587), .Q(dpath_mulcore_b2[2]));
DFFPOSX1 dpath_mulcore_booth_out_dff1_q_reg[0](.D(n17815), .CLK(n9587), .Q(dpath_mulcore_b1[0]));
DFFPOSX1 dpath_mulcore_booth_out_dff1_q_reg[1](.D(n17814), .CLK(n9587), .Q(dpath_mulcore_b1[1]));
DFFPOSX1 dpath_mulcore_booth_out_dff1_q_reg[2](.D(n17813), .CLK(n9587), .Q(dpath_mulcore_b1[2]));
XOR2X1 mul_dpath_mulcore_array2_sc3_20__U12(.A(n17802), .B(n17801), .Y(dpath_mulcore_array2_sc3_20__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_20__U11(.A(n9428), .B(n9099), .Y(n17801));
XOR2X1 mul_dpath_mulcore_array2_sc3_20__U10(.A(dpath_mulcore_array2_s1[20]), .B(dpath_mulcore_array2_s2[20]), .Y(n17802));
XOR2X1 mul_dpath_mulcore_array2_sc3_21__U12(.A(n17796), .B(n17795), .Y(dpath_mulcore_array2_sc3_21__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_21__U11(.A(n16368), .B(n9146), .Y(n17795));
XOR2X1 mul_dpath_mulcore_array2_sc3_21__U10(.A(dpath_mulcore_array2_s1[21]), .B(dpath_mulcore_array2_s2[21]), .Y(n17796));
XOR2X1 mul_dpath_mulcore_array2_sc3_21__U9(.A(n7394), .B(dpath_mulcore_array2_sc3_21__z), .Y(dpath_mulcore_array2_s3[21]));
XOR2X1 mul_dpath_mulcore_array2_sc3_22__U12(.A(n17789), .B(n17788), .Y(dpath_mulcore_array2_sc3_22__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_22__U11(.A(n9473), .B(n9145), .Y(n17788));
XOR2X1 mul_dpath_mulcore_array2_sc3_22__U10(.A(dpath_mulcore_array2_s1[22]), .B(dpath_mulcore_array2_s2[22]), .Y(n17789));
XOR2X1 mul_dpath_mulcore_array2_sc3_22__U9(.A(n7393), .B(dpath_mulcore_array2_sc3_22__z), .Y(dpath_mulcore_array2_s3[22]));
XOR2X1 mul_dpath_mulcore_array2_sc3_23__U12(.A(n17782), .B(n17781), .Y(dpath_mulcore_array2_sc3_23__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_23__U11(.A(n9472), .B(n9144), .Y(n17781));
XOR2X1 mul_dpath_mulcore_array2_sc3_23__U10(.A(dpath_mulcore_array2_s1[23]), .B(dpath_mulcore_array2_s2[23]), .Y(n17782));
XOR2X1 mul_dpath_mulcore_array2_sc3_23__U9(.A(n7392), .B(dpath_mulcore_array2_sc3_23__z), .Y(dpath_mulcore_array2_s3[23]));
XOR2X1 mul_dpath_mulcore_array2_sc3_24__U12(.A(n17775), .B(n17774), .Y(dpath_mulcore_array2_sc3_24__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_24__U11(.A(n9471), .B(n9143), .Y(n17774));
XOR2X1 mul_dpath_mulcore_array2_sc3_24__U10(.A(dpath_mulcore_array2_s1[24]), .B(dpath_mulcore_array2_s2[24]), .Y(n17775));
XOR2X1 mul_dpath_mulcore_array2_sc3_24__U9(.A(n7391), .B(dpath_mulcore_array2_sc3_24__z), .Y(dpath_mulcore_array2_s3[24]));
XOR2X1 mul_dpath_mulcore_array2_sc3_25__U12(.A(n17768), .B(n17767), .Y(dpath_mulcore_array2_sc3_25__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_25__U11(.A(n9470), .B(n9142), .Y(n17767));
XOR2X1 mul_dpath_mulcore_array2_sc3_25__U10(.A(dpath_mulcore_array2_s1[25]), .B(dpath_mulcore_array2_s2[25]), .Y(n17768));
XOR2X1 mul_dpath_mulcore_array2_sc3_25__U9(.A(n7390), .B(dpath_mulcore_array2_sc3_25__z), .Y(dpath_mulcore_array2_s3[25]));
XOR2X1 mul_dpath_mulcore_array2_sc3_26__U12(.A(n17761), .B(n17760), .Y(dpath_mulcore_array2_sc3_26__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_26__U11(.A(n9469), .B(n9141), .Y(n17760));
XOR2X1 mul_dpath_mulcore_array2_sc3_26__U10(.A(dpath_mulcore_array2_s1[26]), .B(dpath_mulcore_array2_s2[26]), .Y(n17761));
XOR2X1 mul_dpath_mulcore_array2_sc3_26__U9(.A(n7389), .B(dpath_mulcore_array2_sc3_26__z), .Y(dpath_mulcore_array2_s3[26]));
XOR2X1 mul_dpath_mulcore_array2_sc3_27__U12(.A(n17754), .B(n17753), .Y(dpath_mulcore_array2_sc3_27__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_27__U11(.A(n9468), .B(n9140), .Y(n17753));
XOR2X1 mul_dpath_mulcore_array2_sc3_27__U10(.A(dpath_mulcore_array2_s1[27]), .B(dpath_mulcore_array2_s2[27]), .Y(n17754));
XOR2X1 mul_dpath_mulcore_array2_sc3_27__U9(.A(n7388), .B(dpath_mulcore_array2_sc3_27__z), .Y(dpath_mulcore_array2_s3[27]));
XOR2X1 mul_dpath_mulcore_array2_sc3_28__U12(.A(n17747), .B(n17746), .Y(dpath_mulcore_array2_sc3_28__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_28__U11(.A(n9467), .B(n9139), .Y(n17746));
XOR2X1 mul_dpath_mulcore_array2_sc3_28__U10(.A(dpath_mulcore_array2_s1[28]), .B(dpath_mulcore_array2_s2[28]), .Y(n17747));
XOR2X1 mul_dpath_mulcore_array2_sc3_28__U9(.A(n7387), .B(dpath_mulcore_array2_sc3_28__z), .Y(dpath_mulcore_array2_s3[28]));
XOR2X1 mul_dpath_mulcore_array2_sc3_29__U12(.A(n17740), .B(n17739), .Y(dpath_mulcore_array2_sc3_29__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_29__U11(.A(n9466), .B(n9138), .Y(n17739));
XOR2X1 mul_dpath_mulcore_array2_sc3_29__U10(.A(dpath_mulcore_array2_s1[29]), .B(dpath_mulcore_array2_s2[29]), .Y(n17740));
XOR2X1 mul_dpath_mulcore_array2_sc3_29__U9(.A(n7386), .B(dpath_mulcore_array2_sc3_29__z), .Y(dpath_mulcore_array2_s3[29]));
XOR2X1 mul_dpath_mulcore_array2_sc3_30__U12(.A(n17733), .B(n17732), .Y(dpath_mulcore_array2_sc3_30__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_30__U11(.A(n9465), .B(n9137), .Y(n17732));
XOR2X1 mul_dpath_mulcore_array2_sc3_30__U10(.A(dpath_mulcore_array2_s1[30]), .B(dpath_mulcore_array2_s2[30]), .Y(n17733));
XOR2X1 mul_dpath_mulcore_array2_sc3_30__U9(.A(n7385), .B(dpath_mulcore_array2_sc3_30__z), .Y(dpath_mulcore_array2_s3[30]));
XOR2X1 mul_dpath_mulcore_array2_sc3_31__U12(.A(n17726), .B(n17725), .Y(dpath_mulcore_array2_sc3_31__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_31__U11(.A(n9464), .B(n9136), .Y(n17725));
XOR2X1 mul_dpath_mulcore_array2_sc3_31__U10(.A(dpath_mulcore_array2_s1[31]), .B(dpath_mulcore_array2_s2[31]), .Y(n17726));
XOR2X1 mul_dpath_mulcore_array2_sc3_31__U9(.A(n7384), .B(dpath_mulcore_array2_sc3_31__z), .Y(dpath_mulcore_array2_s3[31]));
XOR2X1 mul_dpath_mulcore_array2_sc3_32__U12(.A(n17719), .B(n17718), .Y(dpath_mulcore_array2_sc3_32__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_32__U11(.A(n9463), .B(n9135), .Y(n17718));
XOR2X1 mul_dpath_mulcore_array2_sc3_32__U10(.A(dpath_mulcore_array2_s1[32]), .B(dpath_mulcore_array2_s2[32]), .Y(n17719));
XOR2X1 mul_dpath_mulcore_array2_sc3_32__U9(.A(n7383), .B(dpath_mulcore_array2_sc3_32__z), .Y(dpath_mulcore_array2_s3[32]));
XOR2X1 mul_dpath_mulcore_array2_sc3_33__U12(.A(n17712), .B(n17711), .Y(dpath_mulcore_array2_sc3_33__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_33__U11(.A(n9462), .B(n9134), .Y(n17711));
XOR2X1 mul_dpath_mulcore_array2_sc3_33__U10(.A(dpath_mulcore_array2_s1[33]), .B(dpath_mulcore_array2_s2[33]), .Y(n17712));
XOR2X1 mul_dpath_mulcore_array2_sc3_33__U9(.A(n7382), .B(dpath_mulcore_array2_sc3_33__z), .Y(dpath_mulcore_array2_s3[33]));
XOR2X1 mul_dpath_mulcore_array2_sc3_34__U12(.A(n17705), .B(n17704), .Y(dpath_mulcore_array2_sc3_34__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_34__U11(.A(n9461), .B(n9133), .Y(n17704));
XOR2X1 mul_dpath_mulcore_array2_sc3_34__U10(.A(dpath_mulcore_array2_s1[34]), .B(dpath_mulcore_array2_s2[34]), .Y(n17705));
XOR2X1 mul_dpath_mulcore_array2_sc3_34__U9(.A(n7381), .B(dpath_mulcore_array2_sc3_34__z), .Y(dpath_mulcore_array2_s3[34]));
XOR2X1 mul_dpath_mulcore_array2_sc3_35__U12(.A(n17698), .B(n17697), .Y(dpath_mulcore_array2_sc3_35__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_35__U11(.A(n9460), .B(n9132), .Y(n17697));
XOR2X1 mul_dpath_mulcore_array2_sc3_35__U10(.A(dpath_mulcore_array2_s1[35]), .B(dpath_mulcore_array2_s2[35]), .Y(n17698));
XOR2X1 mul_dpath_mulcore_array2_sc3_35__U9(.A(n7380), .B(dpath_mulcore_array2_sc3_35__z), .Y(dpath_mulcore_array2_s3[35]));
XOR2X1 mul_dpath_mulcore_array2_sc3_36__U12(.A(n17691), .B(n17690), .Y(dpath_mulcore_array2_sc3_36__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_36__U11(.A(n9459), .B(n9131), .Y(n17690));
XOR2X1 mul_dpath_mulcore_array2_sc3_36__U10(.A(dpath_mulcore_array2_s1[36]), .B(dpath_mulcore_array2_s2[36]), .Y(n17691));
XOR2X1 mul_dpath_mulcore_array2_sc3_36__U9(.A(n7379), .B(dpath_mulcore_array2_sc3_36__z), .Y(dpath_mulcore_array2_s3[36]));
XOR2X1 mul_dpath_mulcore_array2_sc3_37__U12(.A(n17684), .B(n17683), .Y(dpath_mulcore_array2_sc3_37__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_37__U11(.A(n9458), .B(n9130), .Y(n17683));
XOR2X1 mul_dpath_mulcore_array2_sc3_37__U10(.A(dpath_mulcore_array2_s1[37]), .B(dpath_mulcore_array2_s2[37]), .Y(n17684));
XOR2X1 mul_dpath_mulcore_array2_sc3_37__U9(.A(n7378), .B(dpath_mulcore_array2_sc3_37__z), .Y(dpath_mulcore_array2_s3[37]));
XOR2X1 mul_dpath_mulcore_array2_sc3_38__U12(.A(n17677), .B(n17676), .Y(dpath_mulcore_array2_sc3_38__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_38__U11(.A(n9457), .B(n9129), .Y(n17676));
XOR2X1 mul_dpath_mulcore_array2_sc3_38__U10(.A(dpath_mulcore_array2_s1[38]), .B(dpath_mulcore_array2_s2[38]), .Y(n17677));
XOR2X1 mul_dpath_mulcore_array2_sc3_38__U9(.A(n7377), .B(dpath_mulcore_array2_sc3_38__z), .Y(dpath_mulcore_array2_s3[38]));
XOR2X1 mul_dpath_mulcore_array2_sc3_39__U12(.A(n17670), .B(n17669), .Y(dpath_mulcore_array2_sc3_39__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_39__U11(.A(n9456), .B(n9128), .Y(n17669));
XOR2X1 mul_dpath_mulcore_array2_sc3_39__U10(.A(dpath_mulcore_array2_s1[39]), .B(dpath_mulcore_array2_s2[39]), .Y(n17670));
XOR2X1 mul_dpath_mulcore_array2_sc3_39__U9(.A(n7376), .B(dpath_mulcore_array2_sc3_39__z), .Y(dpath_mulcore_array2_s3[39]));
XOR2X1 mul_dpath_mulcore_array2_sc3_40__U12(.A(n17663), .B(n17662), .Y(dpath_mulcore_array2_sc3_40__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_40__U11(.A(n9455), .B(n9127), .Y(n17662));
XOR2X1 mul_dpath_mulcore_array2_sc3_40__U10(.A(dpath_mulcore_array2_s1[40]), .B(dpath_mulcore_array2_s2[40]), .Y(n17663));
XOR2X1 mul_dpath_mulcore_array2_sc3_40__U9(.A(n7375), .B(dpath_mulcore_array2_sc3_40__z), .Y(dpath_mulcore_array2_s3[40]));
XOR2X1 mul_dpath_mulcore_array2_sc3_41__U12(.A(n17656), .B(n17655), .Y(dpath_mulcore_array2_sc3_41__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_41__U11(.A(n9454), .B(n9126), .Y(n17655));
XOR2X1 mul_dpath_mulcore_array2_sc3_41__U10(.A(dpath_mulcore_array2_s1[41]), .B(dpath_mulcore_array2_s2[41]), .Y(n17656));
XOR2X1 mul_dpath_mulcore_array2_sc3_41__U9(.A(n7374), .B(dpath_mulcore_array2_sc3_41__z), .Y(dpath_mulcore_array2_s3[41]));
XOR2X1 mul_dpath_mulcore_array2_sc3_42__U12(.A(n17649), .B(n17648), .Y(dpath_mulcore_array2_sc3_42__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_42__U11(.A(n9453), .B(n9125), .Y(n17648));
XOR2X1 mul_dpath_mulcore_array2_sc3_42__U10(.A(dpath_mulcore_array2_s1[42]), .B(dpath_mulcore_array2_s2[42]), .Y(n17649));
XOR2X1 mul_dpath_mulcore_array2_sc3_42__U9(.A(n7373), .B(dpath_mulcore_array2_sc3_42__z), .Y(dpath_mulcore_array2_s3[42]));
XOR2X1 mul_dpath_mulcore_array2_sc3_43__U12(.A(n17642), .B(n17641), .Y(dpath_mulcore_array2_sc3_43__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_43__U11(.A(n9452), .B(n9124), .Y(n17641));
XOR2X1 mul_dpath_mulcore_array2_sc3_43__U10(.A(dpath_mulcore_array2_s1[43]), .B(dpath_mulcore_array2_s2[43]), .Y(n17642));
XOR2X1 mul_dpath_mulcore_array2_sc3_43__U9(.A(n7372), .B(dpath_mulcore_array2_sc3_43__z), .Y(dpath_mulcore_array2_s3[43]));
XOR2X1 mul_dpath_mulcore_array2_sc3_44__U12(.A(n17635), .B(n17634), .Y(dpath_mulcore_array2_sc3_44__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_44__U11(.A(n9451), .B(n9123), .Y(n17634));
XOR2X1 mul_dpath_mulcore_array2_sc3_44__U10(.A(dpath_mulcore_array2_s1[44]), .B(dpath_mulcore_array2_s2[44]), .Y(n17635));
XOR2X1 mul_dpath_mulcore_array2_sc3_44__U9(.A(n7371), .B(dpath_mulcore_array2_sc3_44__z), .Y(dpath_mulcore_array2_s3[44]));
XOR2X1 mul_dpath_mulcore_array2_sc3_45__U12(.A(n17628), .B(n17627), .Y(dpath_mulcore_array2_sc3_45__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_45__U11(.A(n9450), .B(n9122), .Y(n17627));
XOR2X1 mul_dpath_mulcore_array2_sc3_45__U10(.A(dpath_mulcore_array2_s1[45]), .B(dpath_mulcore_array2_s2[45]), .Y(n17628));
XOR2X1 mul_dpath_mulcore_array2_sc3_45__U9(.A(n7370), .B(dpath_mulcore_array2_sc3_45__z), .Y(dpath_mulcore_array2_s3[45]));
XOR2X1 mul_dpath_mulcore_array2_sc3_46__U12(.A(n17621), .B(n17620), .Y(dpath_mulcore_array2_sc3_46__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_46__U11(.A(n9449), .B(n9121), .Y(n17620));
XOR2X1 mul_dpath_mulcore_array2_sc3_46__U10(.A(dpath_mulcore_array2_s1[46]), .B(dpath_mulcore_array2_s2[46]), .Y(n17621));
XOR2X1 mul_dpath_mulcore_array2_sc3_46__U9(.A(n7369), .B(dpath_mulcore_array2_sc3_46__z), .Y(dpath_mulcore_array2_s3[46]));
XOR2X1 mul_dpath_mulcore_array2_sc3_47__U12(.A(n17614), .B(n17613), .Y(dpath_mulcore_array2_sc3_47__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_47__U11(.A(n9448), .B(n9120), .Y(n17613));
XOR2X1 mul_dpath_mulcore_array2_sc3_47__U10(.A(dpath_mulcore_array2_s1[47]), .B(dpath_mulcore_array2_s2[47]), .Y(n17614));
XOR2X1 mul_dpath_mulcore_array2_sc3_47__U9(.A(n7368), .B(dpath_mulcore_array2_sc3_47__z), .Y(dpath_mulcore_array2_s3[47]));
XOR2X1 mul_dpath_mulcore_array2_sc3_48__U12(.A(n17607), .B(n17606), .Y(dpath_mulcore_array2_sc3_48__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_48__U11(.A(n9447), .B(n9119), .Y(n17606));
XOR2X1 mul_dpath_mulcore_array2_sc3_48__U10(.A(dpath_mulcore_array2_s1[48]), .B(dpath_mulcore_array2_s2[48]), .Y(n17607));
XOR2X1 mul_dpath_mulcore_array2_sc3_48__U9(.A(n7367), .B(dpath_mulcore_array2_sc3_48__z), .Y(dpath_mulcore_array2_s3[48]));
XOR2X1 mul_dpath_mulcore_array2_sc3_49__U12(.A(n17600), .B(n17599), .Y(dpath_mulcore_array2_sc3_49__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_49__U11(.A(n9446), .B(n9118), .Y(n17599));
XOR2X1 mul_dpath_mulcore_array2_sc3_49__U10(.A(dpath_mulcore_array2_s1[49]), .B(dpath_mulcore_array2_s2[49]), .Y(n17600));
XOR2X1 mul_dpath_mulcore_array2_sc3_49__U9(.A(n7366), .B(dpath_mulcore_array2_sc3_49__z), .Y(dpath_mulcore_array2_s3[49]));
XOR2X1 mul_dpath_mulcore_array2_sc3_50__U12(.A(n17593), .B(n17592), .Y(dpath_mulcore_array2_sc3_50__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_50__U11(.A(n9445), .B(n9117), .Y(n17592));
XOR2X1 mul_dpath_mulcore_array2_sc3_50__U10(.A(dpath_mulcore_array2_s1[50]), .B(dpath_mulcore_array2_s2[50]), .Y(n17593));
XOR2X1 mul_dpath_mulcore_array2_sc3_50__U9(.A(n7365), .B(dpath_mulcore_array2_sc3_50__z), .Y(dpath_mulcore_array2_s3[50]));
XOR2X1 mul_dpath_mulcore_array2_sc3_51__U12(.A(n17586), .B(n17585), .Y(dpath_mulcore_array2_sc3_51__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_51__U11(.A(n9444), .B(n9116), .Y(n17585));
XOR2X1 mul_dpath_mulcore_array2_sc3_51__U10(.A(dpath_mulcore_array2_s1[51]), .B(dpath_mulcore_array2_s2[51]), .Y(n17586));
XOR2X1 mul_dpath_mulcore_array2_sc3_51__U9(.A(n7364), .B(dpath_mulcore_array2_sc3_51__z), .Y(dpath_mulcore_array2_s3[51]));
XOR2X1 mul_dpath_mulcore_array2_sc3_52__U12(.A(n17579), .B(n17578), .Y(dpath_mulcore_array2_sc3_52__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_52__U11(.A(n9443), .B(n9115), .Y(n17578));
XOR2X1 mul_dpath_mulcore_array2_sc3_52__U10(.A(dpath_mulcore_array2_s1[52]), .B(dpath_mulcore_array2_s2[52]), .Y(n17579));
XOR2X1 mul_dpath_mulcore_array2_sc3_52__U9(.A(n7363), .B(dpath_mulcore_array2_sc3_52__z), .Y(dpath_mulcore_array2_s3[52]));
XOR2X1 mul_dpath_mulcore_array2_sc3_53__U12(.A(n17572), .B(n17571), .Y(dpath_mulcore_array2_sc3_53__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_53__U11(.A(n9442), .B(n9114), .Y(n17571));
XOR2X1 mul_dpath_mulcore_array2_sc3_53__U10(.A(dpath_mulcore_array2_s1[53]), .B(dpath_mulcore_array2_s2[53]), .Y(n17572));
XOR2X1 mul_dpath_mulcore_array2_sc3_53__U9(.A(n7362), .B(dpath_mulcore_array2_sc3_53__z), .Y(dpath_mulcore_array2_s3[53]));
XOR2X1 mul_dpath_mulcore_array2_sc3_54__U12(.A(n17565), .B(n17564), .Y(dpath_mulcore_array2_sc3_54__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_54__U11(.A(n9441), .B(n9113), .Y(n17564));
XOR2X1 mul_dpath_mulcore_array2_sc3_54__U10(.A(dpath_mulcore_array2_s1[54]), .B(dpath_mulcore_array2_s2[54]), .Y(n17565));
XOR2X1 mul_dpath_mulcore_array2_sc3_54__U9(.A(n7361), .B(dpath_mulcore_array2_sc3_54__z), .Y(dpath_mulcore_array2_s3[54]));
XOR2X1 mul_dpath_mulcore_array2_sc3_55__U12(.A(n17558), .B(n17557), .Y(dpath_mulcore_array2_sc3_55__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_55__U11(.A(n9440), .B(n9112), .Y(n17557));
XOR2X1 mul_dpath_mulcore_array2_sc3_55__U10(.A(dpath_mulcore_array2_s1[55]), .B(dpath_mulcore_array2_s2[55]), .Y(n17558));
XOR2X1 mul_dpath_mulcore_array2_sc3_55__U9(.A(n7360), .B(dpath_mulcore_array2_sc3_55__z), .Y(dpath_mulcore_array2_s3[55]));
XOR2X1 mul_dpath_mulcore_array2_sc3_56__U12(.A(n17551), .B(n17550), .Y(dpath_mulcore_array2_sc3_56__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_56__U11(.A(n9439), .B(n9111), .Y(n17550));
XOR2X1 mul_dpath_mulcore_array2_sc3_56__U10(.A(dpath_mulcore_array2_s1[56]), .B(dpath_mulcore_array2_s2[56]), .Y(n17551));
XOR2X1 mul_dpath_mulcore_array2_sc3_56__U9(.A(n7359), .B(dpath_mulcore_array2_sc3_56__z), .Y(dpath_mulcore_array2_s3[56]));
XOR2X1 mul_dpath_mulcore_array2_sc3_57__U12(.A(n17544), .B(n17543), .Y(dpath_mulcore_array2_sc3_57__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_57__U11(.A(n9438), .B(n9110), .Y(n17543));
XOR2X1 mul_dpath_mulcore_array2_sc3_57__U10(.A(dpath_mulcore_array2_s1[57]), .B(dpath_mulcore_array2_s2[57]), .Y(n17544));
XOR2X1 mul_dpath_mulcore_array2_sc3_57__U9(.A(n7358), .B(dpath_mulcore_array2_sc3_57__z), .Y(dpath_mulcore_array2_s3[57]));
XOR2X1 mul_dpath_mulcore_array2_sc3_58__U12(.A(n17537), .B(n17536), .Y(dpath_mulcore_array2_sc3_58__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_58__U11(.A(n9437), .B(n9109), .Y(n17536));
XOR2X1 mul_dpath_mulcore_array2_sc3_58__U10(.A(dpath_mulcore_array2_s1[58]), .B(dpath_mulcore_array2_s2[58]), .Y(n17537));
XOR2X1 mul_dpath_mulcore_array2_sc3_58__U9(.A(n7357), .B(dpath_mulcore_array2_sc3_58__z), .Y(dpath_mulcore_array2_s3[58]));
XOR2X1 mul_dpath_mulcore_array2_sc3_59__U12(.A(n17530), .B(n17529), .Y(dpath_mulcore_array2_sc3_59__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_59__U11(.A(n9436), .B(n9108), .Y(n17529));
XOR2X1 mul_dpath_mulcore_array2_sc3_59__U10(.A(dpath_mulcore_array2_s1[59]), .B(dpath_mulcore_array2_s2[59]), .Y(n17530));
XOR2X1 mul_dpath_mulcore_array2_sc3_59__U9(.A(n7356), .B(dpath_mulcore_array2_sc3_59__z), .Y(dpath_mulcore_array2_s3[59]));
XOR2X1 mul_dpath_mulcore_array2_sc3_60__U12(.A(n17523), .B(n17522), .Y(dpath_mulcore_array2_sc3_60__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_60__U11(.A(n9435), .B(n9107), .Y(n17522));
XOR2X1 mul_dpath_mulcore_array2_sc3_60__U10(.A(dpath_mulcore_array2_s1[60]), .B(dpath_mulcore_array2_s2[60]), .Y(n17523));
XOR2X1 mul_dpath_mulcore_array2_sc3_60__U9(.A(n7355), .B(dpath_mulcore_array2_sc3_60__z), .Y(dpath_mulcore_array2_s3[60]));
XOR2X1 mul_dpath_mulcore_array2_sc3_61__U12(.A(n17516), .B(n17515), .Y(dpath_mulcore_array2_sc3_61__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_61__U11(.A(n9434), .B(n9106), .Y(n17515));
XOR2X1 mul_dpath_mulcore_array2_sc3_61__U10(.A(dpath_mulcore_array2_s1[61]), .B(dpath_mulcore_array2_s2[61]), .Y(n17516));
XOR2X1 mul_dpath_mulcore_array2_sc3_61__U9(.A(n7354), .B(dpath_mulcore_array2_sc3_61__z), .Y(dpath_mulcore_array2_s3[61]));
XOR2X1 mul_dpath_mulcore_array2_sc3_62__U12(.A(n17509), .B(n17508), .Y(dpath_mulcore_array2_sc3_62__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_62__U11(.A(n9433), .B(n9105), .Y(n17508));
XOR2X1 mul_dpath_mulcore_array2_sc3_62__U10(.A(dpath_mulcore_array2_s1[62]), .B(dpath_mulcore_array2_s2[62]), .Y(n17509));
XOR2X1 mul_dpath_mulcore_array2_sc3_62__U9(.A(n7353), .B(dpath_mulcore_array2_sc3_62__z), .Y(dpath_mulcore_array2_s3[62]));
XOR2X1 mul_dpath_mulcore_array2_sc3_63__U12(.A(n17502), .B(n17501), .Y(dpath_mulcore_array2_sc3_63__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_63__U11(.A(n9432), .B(n9104), .Y(n17501));
XOR2X1 mul_dpath_mulcore_array2_sc3_63__U10(.A(dpath_mulcore_array2_s1[63]), .B(dpath_mulcore_array2_s2[63]), .Y(n17502));
XOR2X1 mul_dpath_mulcore_array2_sc3_63__U9(.A(n7352), .B(dpath_mulcore_array2_sc3_63__z), .Y(dpath_mulcore_array2_s3[63]));
XOR2X1 mul_dpath_mulcore_array2_sc3_64__U12(.A(n17495), .B(n17494), .Y(dpath_mulcore_array2_sc3_64__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_64__U11(.A(n9431), .B(n9103), .Y(n17494));
XOR2X1 mul_dpath_mulcore_array2_sc3_64__U10(.A(dpath_mulcore_array2_s1[64]), .B(dpath_mulcore_array2_s2[64]), .Y(n17495));
XOR2X1 mul_dpath_mulcore_array2_sc3_64__U9(.A(n7351), .B(dpath_mulcore_array2_sc3_64__z), .Y(dpath_mulcore_array2_s3[64]));
XOR2X1 mul_dpath_mulcore_array2_sc3_65__U12(.A(n17488), .B(n17487), .Y(dpath_mulcore_array2_sc3_65__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_65__U11(.A(n9430), .B(n9102), .Y(n17487));
XOR2X1 mul_dpath_mulcore_array2_sc3_65__U10(.A(dpath_mulcore_array2_s1[65]), .B(dpath_mulcore_array2_s2[65]), .Y(n17488));
XOR2X1 mul_dpath_mulcore_array2_sc3_65__U9(.A(n7350), .B(dpath_mulcore_array2_sc3_65__z), .Y(dpath_mulcore_array2_s3[65]));
XOR2X1 mul_dpath_mulcore_array2_sc3_66__U12(.A(n17481), .B(n17480), .Y(dpath_mulcore_array2_sc3_66__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_66__U11(.A(n9429), .B(n9101), .Y(n17480));
XOR2X1 mul_dpath_mulcore_array2_sc3_66__U10(.A(dpath_mulcore_array2_s1[66]), .B(dpath_mulcore_array2_s2[66]), .Y(n17481));
XOR2X1 mul_dpath_mulcore_array2_sc3_66__U9(.A(n7349), .B(dpath_mulcore_array2_sc3_66__z), .Y(dpath_mulcore_array2_s3[66]));
XOR2X1 mul_dpath_mulcore_array2_sc3_67__U12(.A(n17474), .B(n9100), .Y(dpath_mulcore_array2_sc3_67__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_67__U10(.A(dpath_mulcore_array2_s1[67]), .B(dpath_mulcore_array2_s2[67]), .Y(n17474));
XOR2X1 mul_dpath_mulcore_array2_sc3_67__U9(.A(n7348), .B(dpath_mulcore_array2_sc3_67__z), .Y(dpath_mulcore_array2_s3[67]));
XOR2X1 mul_dpath_mulcore_array2_sc3_68__U12(.A(dpath_mulcore_array2_s2[68]), .B(n6071), .Y(dpath_mulcore_array2_sc3_68__z));
XOR2X1 mul_dpath_mulcore_array2_sc3_68__U9(.A(n17471), .B(dpath_mulcore_array2_sc3_68__z), .Y(dpath_mulcore_array2_s3[68]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_11__U12(.A(n17468), .B(n17467), .Y(dpath_mulcore_ary1_a1_sc3_11__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_11__U11(.A(dpath_mulcore_ary1_a1_s_2[11]), .B(dpath_mulcore_ary1_a1_s_1[11]), .Y(n17467));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_11__U10(.A(dpath_mulcore_ary1_a1_c_1[10]), .B(n9098), .Y(n17468));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_12__U12(.A(n17462), .B(n17461), .Y(dpath_mulcore_ary1_a1_sc3_12__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_12__U11(.A(dpath_mulcore_ary1_a1_s_2[12]), .B(dpath_mulcore_ary1_a1_s_1[12]), .Y(n17461));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_12__U10(.A(dpath_mulcore_ary1_a1_c_1[11]), .B(n9097), .Y(n17462));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_12__U9(.A(n7347), .B(dpath_mulcore_ary1_a1_sc3_12__z), .Y(dpath_mulcore_a1sum[12]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_13__U12(.A(n17455), .B(n17454), .Y(dpath_mulcore_ary1_a1_sc3_13__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_13__U11(.A(dpath_mulcore_ary1_a1_s_2[13]), .B(dpath_mulcore_ary1_a1_s_1[13]), .Y(n17454));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_13__U10(.A(dpath_mulcore_ary1_a1_c_1[12]), .B(n9096), .Y(n17455));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_13__U9(.A(n7346), .B(dpath_mulcore_ary1_a1_sc3_13__z), .Y(dpath_mulcore_a1sum[13]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_14__U12(.A(n17448), .B(n17447), .Y(dpath_mulcore_ary1_a1_sc3_14__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_14__U11(.A(dpath_mulcore_ary1_a1_s_2[14]), .B(dpath_mulcore_ary1_a1_s_1[14]), .Y(n17447));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_14__U10(.A(dpath_mulcore_ary1_a1_c_1[13]), .B(n9095), .Y(n17448));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_14__U9(.A(n7345), .B(dpath_mulcore_ary1_a1_sc3_14__z), .Y(dpath_mulcore_a1sum[14]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_15__U12(.A(n17441), .B(n17440), .Y(dpath_mulcore_ary1_a1_sc3_15__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_15__U11(.A(dpath_mulcore_ary1_a1_s_2[15]), .B(dpath_mulcore_ary1_a1_s_1[15]), .Y(n17440));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_15__U10(.A(n9424), .B(n9094), .Y(n17441));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_15__U9(.A(n7344), .B(dpath_mulcore_ary1_a1_sc3_15__z), .Y(dpath_mulcore_a1sum[15]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_16__U12(.A(n17434), .B(n17433), .Y(dpath_mulcore_ary1_a1_sc3_16__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_16__U11(.A(dpath_mulcore_ary1_a1_s_2[16]), .B(dpath_mulcore_ary1_a1_s_1[16]), .Y(n17433));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_16__U10(.A(n9423), .B(n9093), .Y(n17434));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_16__U9(.A(n7343), .B(dpath_mulcore_ary1_a1_sc3_16__z), .Y(dpath_mulcore_a1sum[16]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_17__U12(.A(n17427), .B(n17426), .Y(dpath_mulcore_ary1_a1_sc3_17__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_17__U11(.A(dpath_mulcore_ary1_a1_s_2[17]), .B(dpath_mulcore_ary1_a1_s_1[17]), .Y(n17426));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_17__U10(.A(n9422), .B(n9092), .Y(n17427));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_17__U9(.A(n7342), .B(dpath_mulcore_ary1_a1_sc3_17__z), .Y(dpath_mulcore_a1sum[17]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_18__U12(.A(n17420), .B(n17419), .Y(dpath_mulcore_ary1_a1_sc3_18__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_18__U11(.A(dpath_mulcore_ary1_a1_s_2[18]), .B(dpath_mulcore_ary1_a1_s_1[18]), .Y(n17419));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_18__U10(.A(n9421), .B(n9091), .Y(n17420));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_18__U9(.A(n7341), .B(dpath_mulcore_ary1_a1_sc3_18__z), .Y(dpath_mulcore_a1sum[18]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_19__U12(.A(n17413), .B(n17412), .Y(dpath_mulcore_ary1_a1_sc3_19__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_19__U11(.A(dpath_mulcore_ary1_a1_s_2[19]), .B(dpath_mulcore_ary1_a1_s_1[19]), .Y(n17412));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_19__U10(.A(n9420), .B(n9090), .Y(n17413));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_19__U9(.A(n7340), .B(dpath_mulcore_ary1_a1_sc3_19__z), .Y(dpath_mulcore_a1sum[19]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_20__U12(.A(n17406), .B(n17405), .Y(dpath_mulcore_ary1_a1_sc3_20__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_20__U11(.A(dpath_mulcore_ary1_a1_s_2[20]), .B(dpath_mulcore_ary1_a1_s_1[20]), .Y(n17405));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_20__U10(.A(n9419), .B(n9089), .Y(n17406));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_20__U9(.A(n7339), .B(dpath_mulcore_ary1_a1_sc3_20__z), .Y(dpath_mulcore_a1sum[20]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_21__U12(.A(n17399), .B(n17398), .Y(dpath_mulcore_ary1_a1_sc3_21__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_21__U11(.A(dpath_mulcore_ary1_a1_s_2[21]), .B(dpath_mulcore_ary1_a1_s_1[21]), .Y(n17398));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_21__U10(.A(n9418), .B(n9088), .Y(n17399));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_21__U9(.A(n7338), .B(dpath_mulcore_ary1_a1_sc3_21__z), .Y(dpath_mulcore_a1sum[21]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_22__U12(.A(n17392), .B(n17391), .Y(dpath_mulcore_ary1_a1_sc3_22__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_22__U11(.A(dpath_mulcore_ary1_a1_s_2[22]), .B(dpath_mulcore_ary1_a1_s_1[22]), .Y(n17391));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_22__U10(.A(n9417), .B(n9087), .Y(n17392));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_22__U9(.A(n7337), .B(dpath_mulcore_ary1_a1_sc3_22__z), .Y(dpath_mulcore_a1sum[22]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_23__U12(.A(n17385), .B(n17384), .Y(dpath_mulcore_ary1_a1_sc3_23__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_23__U11(.A(dpath_mulcore_ary1_a1_s_2[23]), .B(dpath_mulcore_ary1_a1_s_1[23]), .Y(n17384));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_23__U10(.A(n9416), .B(n9086), .Y(n17385));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_23__U9(.A(n7336), .B(dpath_mulcore_ary1_a1_sc3_23__z), .Y(dpath_mulcore_a1sum[23]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_24__U12(.A(n17378), .B(n17377), .Y(dpath_mulcore_ary1_a1_sc3_24__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_24__U11(.A(dpath_mulcore_ary1_a1_s_2[24]), .B(dpath_mulcore_ary1_a1_s_1[24]), .Y(n17377));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_24__U10(.A(n9415), .B(n9085), .Y(n17378));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_24__U9(.A(n7335), .B(dpath_mulcore_ary1_a1_sc3_24__z), .Y(dpath_mulcore_a1sum[24]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_25__U12(.A(n17371), .B(n17370), .Y(dpath_mulcore_ary1_a1_sc3_25__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_25__U11(.A(dpath_mulcore_ary1_a1_s_2[25]), .B(dpath_mulcore_ary1_a1_s_1[25]), .Y(n17370));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_25__U10(.A(n9414), .B(n9084), .Y(n17371));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_25__U9(.A(n7334), .B(dpath_mulcore_ary1_a1_sc3_25__z), .Y(dpath_mulcore_a1sum[25]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_26__U12(.A(n17364), .B(n17363), .Y(dpath_mulcore_ary1_a1_sc3_26__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_26__U11(.A(dpath_mulcore_ary1_a1_s_2[26]), .B(dpath_mulcore_ary1_a1_s_1[26]), .Y(n17363));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_26__U10(.A(n9413), .B(n9083), .Y(n17364));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_26__U9(.A(n7333), .B(dpath_mulcore_ary1_a1_sc3_26__z), .Y(dpath_mulcore_a1sum[26]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_27__U12(.A(n17357), .B(n17356), .Y(dpath_mulcore_ary1_a1_sc3_27__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_27__U11(.A(dpath_mulcore_ary1_a1_s_2[27]), .B(dpath_mulcore_ary1_a1_s_1[27]), .Y(n17356));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_27__U10(.A(n9412), .B(n9082), .Y(n17357));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_27__U9(.A(n7332), .B(dpath_mulcore_ary1_a1_sc3_27__z), .Y(dpath_mulcore_a1sum[27]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_28__U12(.A(n17350), .B(n17349), .Y(dpath_mulcore_ary1_a1_sc3_28__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_28__U11(.A(dpath_mulcore_ary1_a1_s_2[28]), .B(dpath_mulcore_ary1_a1_s_1[28]), .Y(n17349));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_28__U10(.A(n9411), .B(n9081), .Y(n17350));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_28__U9(.A(n7331), .B(dpath_mulcore_ary1_a1_sc3_28__z), .Y(dpath_mulcore_a1sum[28]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_29__U12(.A(n17343), .B(n17342), .Y(dpath_mulcore_ary1_a1_sc3_29__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_29__U11(.A(dpath_mulcore_ary1_a1_s_2[29]), .B(dpath_mulcore_ary1_a1_s_1[29]), .Y(n17342));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_29__U10(.A(n9410), .B(n9080), .Y(n17343));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_29__U9(.A(n7330), .B(dpath_mulcore_ary1_a1_sc3_29__z), .Y(dpath_mulcore_a1sum[29]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_30__U12(.A(n17336), .B(n17335), .Y(dpath_mulcore_ary1_a1_sc3_30__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_30__U11(.A(dpath_mulcore_ary1_a1_s_2[30]), .B(dpath_mulcore_ary1_a1_s_1[30]), .Y(n17335));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_30__U10(.A(n9409), .B(n9079), .Y(n17336));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_30__U9(.A(n7329), .B(dpath_mulcore_ary1_a1_sc3_30__z), .Y(dpath_mulcore_a1sum[30]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_31__U12(.A(n17329), .B(n17328), .Y(dpath_mulcore_ary1_a1_sc3_31__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_31__U11(.A(dpath_mulcore_ary1_a1_s_2[31]), .B(dpath_mulcore_ary1_a1_s_1[31]), .Y(n17328));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_31__U10(.A(n9408), .B(n9078), .Y(n17329));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_31__U9(.A(n7328), .B(dpath_mulcore_ary1_a1_sc3_31__z), .Y(dpath_mulcore_a1sum[31]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_32__U12(.A(n17322), .B(n17321), .Y(dpath_mulcore_ary1_a1_sc3_32__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_32__U11(.A(dpath_mulcore_ary1_a1_s_2[32]), .B(dpath_mulcore_ary1_a1_s_1[32]), .Y(n17321));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_32__U10(.A(n9407), .B(n9077), .Y(n17322));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_32__U9(.A(n7327), .B(dpath_mulcore_ary1_a1_sc3_32__z), .Y(dpath_mulcore_a1sum[32]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_33__U12(.A(n17315), .B(n17314), .Y(dpath_mulcore_ary1_a1_sc3_33__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_33__U11(.A(dpath_mulcore_ary1_a1_s_2[33]), .B(dpath_mulcore_ary1_a1_s_1[33]), .Y(n17314));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_33__U10(.A(n9406), .B(n9076), .Y(n17315));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_33__U9(.A(n7326), .B(dpath_mulcore_ary1_a1_sc3_33__z), .Y(dpath_mulcore_a1sum[33]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_34__U12(.A(n17308), .B(n17307), .Y(dpath_mulcore_ary1_a1_sc3_34__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_34__U11(.A(dpath_mulcore_ary1_a1_s_2[34]), .B(dpath_mulcore_ary1_a1_s_1[34]), .Y(n17307));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_34__U10(.A(n9405), .B(n9075), .Y(n17308));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_34__U9(.A(n7325), .B(dpath_mulcore_ary1_a1_sc3_34__z), .Y(dpath_mulcore_a1sum[34]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_35__U12(.A(n17301), .B(n17300), .Y(dpath_mulcore_ary1_a1_sc3_35__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_35__U11(.A(dpath_mulcore_ary1_a1_s_2[35]), .B(dpath_mulcore_ary1_a1_s_1[35]), .Y(n17300));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_35__U10(.A(n9404), .B(n9074), .Y(n17301));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_35__U9(.A(n7324), .B(dpath_mulcore_ary1_a1_sc3_35__z), .Y(dpath_mulcore_a1sum[35]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_36__U12(.A(n17294), .B(n17293), .Y(dpath_mulcore_ary1_a1_sc3_36__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_36__U11(.A(dpath_mulcore_ary1_a1_s_2[36]), .B(dpath_mulcore_ary1_a1_s_1[36]), .Y(n17293));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_36__U10(.A(n9403), .B(n9073), .Y(n17294));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_36__U9(.A(n7323), .B(dpath_mulcore_ary1_a1_sc3_36__z), .Y(dpath_mulcore_a1sum[36]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_37__U12(.A(n17287), .B(n17286), .Y(dpath_mulcore_ary1_a1_sc3_37__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_37__U11(.A(dpath_mulcore_ary1_a1_s_2[37]), .B(dpath_mulcore_ary1_a1_s_1[37]), .Y(n17286));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_37__U10(.A(n9402), .B(n9072), .Y(n17287));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_37__U9(.A(n7322), .B(dpath_mulcore_ary1_a1_sc3_37__z), .Y(dpath_mulcore_a1sum[37]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_38__U12(.A(n17280), .B(n17279), .Y(dpath_mulcore_ary1_a1_sc3_38__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_38__U11(.A(dpath_mulcore_ary1_a1_s_2[38]), .B(dpath_mulcore_ary1_a1_s_1[38]), .Y(n17279));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_38__U10(.A(n9401), .B(n9071), .Y(n17280));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_38__U9(.A(n7321), .B(dpath_mulcore_ary1_a1_sc3_38__z), .Y(dpath_mulcore_a1sum[38]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_39__U12(.A(n17273), .B(n17272), .Y(dpath_mulcore_ary1_a1_sc3_39__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_39__U11(.A(dpath_mulcore_ary1_a1_s_2[39]), .B(dpath_mulcore_ary1_a1_s_1[39]), .Y(n17272));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_39__U10(.A(n9400), .B(n9070), .Y(n17273));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_39__U9(.A(n7320), .B(dpath_mulcore_ary1_a1_sc3_39__z), .Y(dpath_mulcore_a1sum[39]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_40__U12(.A(n17266), .B(n17265), .Y(dpath_mulcore_ary1_a1_sc3_40__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_40__U11(.A(dpath_mulcore_ary1_a1_s_2[40]), .B(dpath_mulcore_ary1_a1_s_1[40]), .Y(n17265));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_40__U10(.A(n9399), .B(n9069), .Y(n17266));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_40__U9(.A(n7319), .B(dpath_mulcore_ary1_a1_sc3_40__z), .Y(dpath_mulcore_a1sum[40]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_41__U12(.A(n17259), .B(n17258), .Y(dpath_mulcore_ary1_a1_sc3_41__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_41__U11(.A(dpath_mulcore_ary1_a1_s_2[41]), .B(dpath_mulcore_ary1_a1_s_1[41]), .Y(n17258));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_41__U10(.A(n9398), .B(n9068), .Y(n17259));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_41__U9(.A(n7318), .B(dpath_mulcore_ary1_a1_sc3_41__z), .Y(dpath_mulcore_a1sum[41]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_42__U12(.A(n17252), .B(n17251), .Y(dpath_mulcore_ary1_a1_sc3_42__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_42__U11(.A(dpath_mulcore_ary1_a1_s_2[42]), .B(dpath_mulcore_ary1_a1_s_1[42]), .Y(n17251));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_42__U10(.A(n9397), .B(n9067), .Y(n17252));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_42__U9(.A(n7317), .B(dpath_mulcore_ary1_a1_sc3_42__z), .Y(dpath_mulcore_a1sum[42]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_43__U12(.A(n17245), .B(n17244), .Y(dpath_mulcore_ary1_a1_sc3_43__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_43__U11(.A(dpath_mulcore_ary1_a1_s_2[43]), .B(dpath_mulcore_ary1_a1_s_1[43]), .Y(n17244));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_43__U10(.A(n9396), .B(n9066), .Y(n17245));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_43__U9(.A(n7316), .B(dpath_mulcore_ary1_a1_sc3_43__z), .Y(dpath_mulcore_a1sum[43]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_44__U12(.A(n17238), .B(n17237), .Y(dpath_mulcore_ary1_a1_sc3_44__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_44__U11(.A(dpath_mulcore_ary1_a1_s_2[44]), .B(dpath_mulcore_ary1_a1_s_1[44]), .Y(n17237));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_44__U10(.A(n9395), .B(n9065), .Y(n17238));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_44__U9(.A(n7315), .B(dpath_mulcore_ary1_a1_sc3_44__z), .Y(dpath_mulcore_a1sum[44]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_45__U12(.A(n17231), .B(n17230), .Y(dpath_mulcore_ary1_a1_sc3_45__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_45__U11(.A(dpath_mulcore_ary1_a1_s_2[45]), .B(dpath_mulcore_ary1_a1_s_1[45]), .Y(n17230));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_45__U10(.A(n9394), .B(n9064), .Y(n17231));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_45__U9(.A(n7314), .B(dpath_mulcore_ary1_a1_sc3_45__z), .Y(dpath_mulcore_a1sum[45]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_46__U12(.A(n17224), .B(n17223), .Y(dpath_mulcore_ary1_a1_sc3_46__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_46__U11(.A(dpath_mulcore_ary1_a1_s_2[46]), .B(dpath_mulcore_ary1_a1_s_1[46]), .Y(n17223));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_46__U10(.A(n9393), .B(n9063), .Y(n17224));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_46__U9(.A(n7313), .B(dpath_mulcore_ary1_a1_sc3_46__z), .Y(dpath_mulcore_a1sum[46]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_47__U12(.A(n17217), .B(n17216), .Y(dpath_mulcore_ary1_a1_sc3_47__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_47__U11(.A(dpath_mulcore_ary1_a1_s_2[47]), .B(dpath_mulcore_ary1_a1_s_1[47]), .Y(n17216));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_47__U10(.A(n9392), .B(n9062), .Y(n17217));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_47__U9(.A(n7312), .B(dpath_mulcore_ary1_a1_sc3_47__z), .Y(dpath_mulcore_a1sum[47]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_48__U12(.A(n17210), .B(n17209), .Y(dpath_mulcore_ary1_a1_sc3_48__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_48__U11(.A(dpath_mulcore_ary1_a1_s_2[48]), .B(dpath_mulcore_ary1_a1_s_1[48]), .Y(n17209));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_48__U10(.A(n9391), .B(n9061), .Y(n17210));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_48__U9(.A(n7311), .B(dpath_mulcore_ary1_a1_sc3_48__z), .Y(dpath_mulcore_a1sum[48]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_49__U12(.A(n17203), .B(n17202), .Y(dpath_mulcore_ary1_a1_sc3_49__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_49__U11(.A(dpath_mulcore_ary1_a1_s_2[49]), .B(dpath_mulcore_ary1_a1_s_1[49]), .Y(n17202));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_49__U10(.A(n9390), .B(n9060), .Y(n17203));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_49__U9(.A(n7310), .B(dpath_mulcore_ary1_a1_sc3_49__z), .Y(dpath_mulcore_a1sum[49]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_50__U12(.A(n17196), .B(n17195), .Y(dpath_mulcore_ary1_a1_sc3_50__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_50__U11(.A(dpath_mulcore_ary1_a1_s_2[50]), .B(dpath_mulcore_ary1_a1_s_1[50]), .Y(n17195));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_50__U10(.A(n9389), .B(n9059), .Y(n17196));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_50__U9(.A(n7309), .B(dpath_mulcore_ary1_a1_sc3_50__z), .Y(dpath_mulcore_a1sum[50]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_51__U12(.A(n17189), .B(n17188), .Y(dpath_mulcore_ary1_a1_sc3_51__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_51__U11(.A(dpath_mulcore_ary1_a1_s_2[51]), .B(dpath_mulcore_ary1_a1_s_1[51]), .Y(n17188));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_51__U10(.A(n9388), .B(n9058), .Y(n17189));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_51__U9(.A(n7308), .B(dpath_mulcore_ary1_a1_sc3_51__z), .Y(dpath_mulcore_a1sum[51]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_52__U12(.A(n17182), .B(n17181), .Y(dpath_mulcore_ary1_a1_sc3_52__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_52__U11(.A(dpath_mulcore_ary1_a1_s_2[52]), .B(dpath_mulcore_ary1_a1_s_1[52]), .Y(n17181));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_52__U10(.A(n9387), .B(n9057), .Y(n17182));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_52__U9(.A(n7307), .B(dpath_mulcore_ary1_a1_sc3_52__z), .Y(dpath_mulcore_a1sum[52]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_53__U12(.A(n17175), .B(n17174), .Y(dpath_mulcore_ary1_a1_sc3_53__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_53__U11(.A(dpath_mulcore_ary1_a1_s_2[53]), .B(dpath_mulcore_ary1_a1_s_1[53]), .Y(n17174));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_53__U10(.A(n9386), .B(n9056), .Y(n17175));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_53__U9(.A(n7306), .B(dpath_mulcore_ary1_a1_sc3_53__z), .Y(dpath_mulcore_a1sum[53]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_54__U12(.A(n17168), .B(n17167), .Y(dpath_mulcore_ary1_a1_sc3_54__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_54__U11(.A(dpath_mulcore_ary1_a1_s_2[54]), .B(dpath_mulcore_ary1_a1_s_1[54]), .Y(n17167));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_54__U10(.A(n9385), .B(n9055), .Y(n17168));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_54__U9(.A(n7305), .B(dpath_mulcore_ary1_a1_sc3_54__z), .Y(dpath_mulcore_a1sum[54]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_55__U12(.A(n17161), .B(n17160), .Y(dpath_mulcore_ary1_a1_sc3_55__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_55__U11(.A(dpath_mulcore_ary1_a1_s_2[55]), .B(dpath_mulcore_ary1_a1_s_1[55]), .Y(n17160));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_55__U10(.A(n9384), .B(n9054), .Y(n17161));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_55__U9(.A(n7304), .B(dpath_mulcore_ary1_a1_sc3_55__z), .Y(dpath_mulcore_a1sum[55]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_56__U12(.A(n17154), .B(n17153), .Y(dpath_mulcore_ary1_a1_sc3_56__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_56__U11(.A(dpath_mulcore_ary1_a1_s_2[56]), .B(dpath_mulcore_ary1_a1_s_1[56]), .Y(n17153));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_56__U10(.A(n9383), .B(n9053), .Y(n17154));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_56__U9(.A(n7303), .B(dpath_mulcore_ary1_a1_sc3_56__z), .Y(dpath_mulcore_a1sum[56]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_57__U12(.A(n17147), .B(n17146), .Y(dpath_mulcore_ary1_a1_sc3_57__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_57__U11(.A(dpath_mulcore_ary1_a1_s_2[57]), .B(dpath_mulcore_ary1_a1_s_1[57]), .Y(n17146));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_57__U10(.A(n9382), .B(n9052), .Y(n17147));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_57__U9(.A(n7302), .B(dpath_mulcore_ary1_a1_sc3_57__z), .Y(dpath_mulcore_a1sum[57]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_58__U12(.A(n17140), .B(n17139), .Y(dpath_mulcore_ary1_a1_sc3_58__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_58__U11(.A(dpath_mulcore_ary1_a1_s_2[58]), .B(dpath_mulcore_ary1_a1_s_1[58]), .Y(n17139));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_58__U10(.A(n9381), .B(n9051), .Y(n17140));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_58__U9(.A(n7301), .B(dpath_mulcore_ary1_a1_sc3_58__z), .Y(dpath_mulcore_a1sum[58]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_59__U12(.A(n17133), .B(n17132), .Y(dpath_mulcore_ary1_a1_sc3_59__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_59__U11(.A(dpath_mulcore_ary1_a1_s_2[59]), .B(dpath_mulcore_ary1_a1_s_1[59]), .Y(n17132));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_59__U10(.A(n9380), .B(n9050), .Y(n17133));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_59__U9(.A(n7300), .B(dpath_mulcore_ary1_a1_sc3_59__z), .Y(dpath_mulcore_a1sum[59]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_60__U12(.A(n17126), .B(n17125), .Y(dpath_mulcore_ary1_a1_sc3_60__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_60__U11(.A(dpath_mulcore_ary1_a1_s_2[60]), .B(dpath_mulcore_ary1_a1_s_1[60]), .Y(n17125));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_60__U10(.A(n9379), .B(n9049), .Y(n17126));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_60__U9(.A(n7299), .B(dpath_mulcore_ary1_a1_sc3_60__z), .Y(dpath_mulcore_a1sum[60]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_61__U12(.A(n17119), .B(n17118), .Y(dpath_mulcore_ary1_a1_sc3_61__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_61__U11(.A(dpath_mulcore_ary1_a1_s_2[61]), .B(dpath_mulcore_ary1_a1_s_1[61]), .Y(n17118));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_61__U10(.A(n9378), .B(n9048), .Y(n17119));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_61__U9(.A(n7298), .B(dpath_mulcore_ary1_a1_sc3_61__z), .Y(dpath_mulcore_a1sum[61]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_62__U12(.A(n17112), .B(n17111), .Y(dpath_mulcore_ary1_a1_sc3_62__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_62__U11(.A(dpath_mulcore_ary1_a1_s_2[62]), .B(dpath_mulcore_ary1_a1_s_1[62]), .Y(n17111));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_62__U10(.A(n9377), .B(n9047), .Y(n17112));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_62__U9(.A(n7297), .B(dpath_mulcore_ary1_a1_sc3_62__z), .Y(dpath_mulcore_a1sum[62]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_63__U12(.A(n17105), .B(n17104), .Y(dpath_mulcore_ary1_a1_sc3_63__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_63__U11(.A(dpath_mulcore_ary1_a1_s_2[63]), .B(dpath_mulcore_ary1_a1_s_1[63]), .Y(n17104));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_63__U10(.A(n9376), .B(n9046), .Y(n17105));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_63__U9(.A(n7296), .B(dpath_mulcore_ary1_a1_sc3_63__z), .Y(dpath_mulcore_a1sum[63]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_64__U12(.A(n17098), .B(n17097), .Y(dpath_mulcore_ary1_a1_sc3_64__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_64__U11(.A(dpath_mulcore_ary1_a1_s_2[64]), .B(dpath_mulcore_ary1_a1_s_1[64]), .Y(n17097));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_64__U10(.A(n9375), .B(n9045), .Y(n17098));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_64__U9(.A(n7295), .B(dpath_mulcore_ary1_a1_sc3_64__z), .Y(dpath_mulcore_a1sum[64]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_65__U12(.A(n17091), .B(n17090), .Y(dpath_mulcore_ary1_a1_sc3_65__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_65__U11(.A(dpath_mulcore_ary1_a1_s_2[65]), .B(dpath_mulcore_ary1_a1_s_1[65]), .Y(n17090));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_65__U10(.A(n9374), .B(n9044), .Y(n17091));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_65__U9(.A(n7294), .B(dpath_mulcore_ary1_a1_sc3_65__z), .Y(dpath_mulcore_a1sum[65]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_66__U12(.A(n17084), .B(n17083), .Y(dpath_mulcore_ary1_a1_sc3_66__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_66__U11(.A(dpath_mulcore_ary1_a1_s_2[66]), .B(dpath_mulcore_ary1_a1_s_1[66]), .Y(n17083));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_66__U10(.A(n9373), .B(n9043), .Y(n17084));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_66__U9(.A(n7293), .B(dpath_mulcore_ary1_a1_sc3_66__z), .Y(dpath_mulcore_a1sum[66]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_67__U12(.A(n17077), .B(n17076), .Y(dpath_mulcore_ary1_a1_sc3_67__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_67__U11(.A(dpath_mulcore_ary1_a1_s_2[67]), .B(dpath_mulcore_ary1_a1_s_1[67]), .Y(n17076));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_67__U10(.A(n9372), .B(n9042), .Y(n17077));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_67__U9(.A(n7292), .B(dpath_mulcore_ary1_a1_sc3_67__z), .Y(dpath_mulcore_a1sum[67]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_68__U12(.A(n17070), .B(n17069), .Y(dpath_mulcore_ary1_a1_sc3_68__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_68__U11(.A(dpath_mulcore_ary1_a1_s_2[68]), .B(dpath_mulcore_ary1_a1_s_1[68]), .Y(n17069));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_68__U10(.A(n9371), .B(n9041), .Y(n17070));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_68__U9(.A(n7291), .B(dpath_mulcore_ary1_a1_sc3_68__z), .Y(dpath_mulcore_a1sum[68]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_69__U12(.A(n17063), .B(n17062), .Y(dpath_mulcore_ary1_a1_sc3_69__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_69__U11(.A(dpath_mulcore_ary1_a1_s_2[69]), .B(dpath_mulcore_ary1_a1_s_1[69]), .Y(n17062));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_69__U10(.A(n9370), .B(n9040), .Y(n17063));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_69__U9(.A(n7290), .B(dpath_mulcore_ary1_a1_sc3_69__z), .Y(dpath_mulcore_a1sum[69]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_70__U12(.A(n17056), .B(n17055), .Y(dpath_mulcore_ary1_a1_sc3_70__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_70__U11(.A(dpath_mulcore_ary1_a1_s_2[70]), .B(n10025), .Y(n17055));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_70__U10(.A(n9369), .B(n9039), .Y(n17056));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_70__U9(.A(n7289), .B(dpath_mulcore_ary1_a1_sc3_70__z), .Y(dpath_mulcore_a1sum[70]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_76__U12(.A(n8298), .B(n2), .Y(dpath_mulcore_ary1_a1_sc3_76__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_76__U9(.A(n17032), .B(dpath_mulcore_ary1_a1_sc3_76__z), .Y(dpath_mulcore_a1sum[76]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_72__U12(.A(n8297), .B(n17047), .Y(dpath_mulcore_ary1_a1_sc3_72__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_72__U11(.A(dpath_mulcore_ary1_a1_s_2[72]), .B(dpath_mulcore_ary1_a1_s1[66]), .Y(n17047));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_72__U9(.A(n7287), .B(dpath_mulcore_ary1_a1_sc3_72__z), .Y(dpath_mulcore_a1sum[72]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_73__U12(.A(n8301), .B(n17043), .Y(dpath_mulcore_ary1_a1_sc3_73__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_73__U11(.A(dpath_mulcore_ary1_a1_s_2[73]), .B(dpath_mulcore_ary1_a1_s1[67]), .Y(n17043));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_73__U9(.A(n17044), .B(dpath_mulcore_ary1_a1_sc3_73__z), .Y(dpath_mulcore_a1sum[73]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_74__U12(.A(n8300), .B(n17039), .Y(dpath_mulcore_ary1_a1_sc3_74__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_74__U11(.A(dpath_mulcore_ary1_a1_s_2[74]), .B(dpath_mulcore_ary1_a1_I1_I2_net073), .Y(n17039));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_74__U9(.A(n17040), .B(dpath_mulcore_ary1_a1_sc3_74__z), .Y(dpath_mulcore_a1sum[74]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_75__U12(.A(n8299), .B(n17035), .Y(dpath_mulcore_ary1_a1_sc3_75__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_75__U11(.A(dpath_mulcore_ary1_a1_s_2[75]), .B(n9485), .Y(n17035));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_75__U9(.A(n17036), .B(dpath_mulcore_ary1_a1_sc3_75__z), .Y(dpath_mulcore_a1sum[75]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_71__U12(.A(n17031), .B(n17030), .Y(dpath_mulcore_ary1_a1_sc3_71__z));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_71__U11(.A(dpath_mulcore_ary1_a1_s_2[71]), .B(dpath_mulcore_ary1_a1_s1[65]), .Y(n17030));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_71__U10(.A(dpath_mulcore_ary1_a1_s1[64]), .B(n9038), .Y(n17031));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_71__U9(.A(n7288), .B(dpath_mulcore_ary1_a1_sc3_71__z), .Y(dpath_mulcore_a1sum[71]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_11__U12(.A(n17024), .B(n17023), .Y(dpath_mulcore_ary1_a0_sc3_11__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_11__U11(.A(dpath_mulcore_ary1_a0_s_2[11]), .B(dpath_mulcore_ary1_a0_s_1[11]), .Y(n17023));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_11__U10(.A(dpath_mulcore_ary1_a0_c_1[10]), .B(n9037), .Y(n17024));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_12__U12(.A(n17018), .B(n17017), .Y(dpath_mulcore_ary1_a0_sc3_12__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_12__U11(.A(dpath_mulcore_ary1_a0_s_2[12]), .B(dpath_mulcore_ary1_a0_s_1[12]), .Y(n17017));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_12__U10(.A(dpath_mulcore_ary1_a0_c_1[11]), .B(n9036), .Y(n17018));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_12__U9(.A(n7286), .B(dpath_mulcore_ary1_a0_sc3_12__z), .Y(dpath_mulcore_a0sum[12]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_13__U12(.A(n17011), .B(n17010), .Y(dpath_mulcore_ary1_a0_sc3_13__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_13__U11(.A(dpath_mulcore_ary1_a0_s_2[13]), .B(dpath_mulcore_ary1_a0_s_1[13]), .Y(n17010));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_13__U10(.A(dpath_mulcore_ary1_a0_c_1[12]), .B(n9035), .Y(n17011));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_13__U9(.A(n7285), .B(dpath_mulcore_ary1_a0_sc3_13__z), .Y(dpath_mulcore_a0sum[13]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_14__U12(.A(n17004), .B(n17003), .Y(dpath_mulcore_ary1_a0_sc3_14__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_14__U11(.A(dpath_mulcore_ary1_a0_s_2[14]), .B(dpath_mulcore_ary1_a0_s_1[14]), .Y(n17003));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_14__U10(.A(dpath_mulcore_ary1_a0_c_1[13]), .B(n9034), .Y(n17004));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_14__U9(.A(n7284), .B(dpath_mulcore_ary1_a0_sc3_14__z), .Y(dpath_mulcore_a0sum[14]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_15__U12(.A(n16997), .B(n16996), .Y(dpath_mulcore_ary1_a0_sc3_15__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_15__U11(.A(dpath_mulcore_ary1_a0_s_2[15]), .B(dpath_mulcore_ary1_a0_s_1[15]), .Y(n16996));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_15__U10(.A(n9368), .B(n9033), .Y(n16997));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_15__U9(.A(n7283), .B(dpath_mulcore_ary1_a0_sc3_15__z), .Y(dpath_mulcore_a0sum[15]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_16__U12(.A(n16990), .B(n16989), .Y(dpath_mulcore_ary1_a0_sc3_16__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_16__U11(.A(dpath_mulcore_ary1_a0_s_2[16]), .B(dpath_mulcore_ary1_a0_s_1[16]), .Y(n16989));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_16__U10(.A(n9367), .B(n9032), .Y(n16990));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_16__U9(.A(n7282), .B(dpath_mulcore_ary1_a0_sc3_16__z), .Y(dpath_mulcore_a0sum[16]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_17__U12(.A(n16983), .B(n16982), .Y(dpath_mulcore_ary1_a0_sc3_17__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_17__U11(.A(dpath_mulcore_ary1_a0_s_2[17]), .B(dpath_mulcore_ary1_a0_s_1[17]), .Y(n16982));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_17__U10(.A(n9366), .B(n9031), .Y(n16983));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_17__U9(.A(n7281), .B(dpath_mulcore_ary1_a0_sc3_17__z), .Y(dpath_mulcore_a0sum[17]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_18__U12(.A(n16976), .B(n16975), .Y(dpath_mulcore_ary1_a0_sc3_18__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_18__U11(.A(dpath_mulcore_ary1_a0_s_2[18]), .B(dpath_mulcore_ary1_a0_s_1[18]), .Y(n16975));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_18__U10(.A(n9365), .B(n9030), .Y(n16976));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_18__U9(.A(n7280), .B(dpath_mulcore_ary1_a0_sc3_18__z), .Y(dpath_mulcore_a0sum[18]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_19__U12(.A(n16969), .B(n16968), .Y(dpath_mulcore_ary1_a0_sc3_19__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_19__U11(.A(dpath_mulcore_ary1_a0_s_2[19]), .B(dpath_mulcore_ary1_a0_s_1[19]), .Y(n16968));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_19__U10(.A(n9364), .B(n9029), .Y(n16969));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_19__U9(.A(n7279), .B(dpath_mulcore_ary1_a0_sc3_19__z), .Y(dpath_mulcore_a0sum[19]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_20__U12(.A(n16962), .B(n16961), .Y(dpath_mulcore_ary1_a0_sc3_20__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_20__U11(.A(dpath_mulcore_ary1_a0_s_2[20]), .B(dpath_mulcore_ary1_a0_s_1[20]), .Y(n16961));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_20__U10(.A(n9363), .B(n9028), .Y(n16962));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_20__U9(.A(n7278), .B(dpath_mulcore_ary1_a0_sc3_20__z), .Y(dpath_mulcore_a0sum[20]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_21__U12(.A(n16955), .B(n16954), .Y(dpath_mulcore_ary1_a0_sc3_21__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_21__U11(.A(dpath_mulcore_ary1_a0_s_2[21]), .B(dpath_mulcore_ary1_a0_s_1[21]), .Y(n16954));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_21__U10(.A(n9362), .B(n9027), .Y(n16955));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_21__U9(.A(n7277), .B(dpath_mulcore_ary1_a0_sc3_21__z), .Y(dpath_mulcore_a0sum[21]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_22__U12(.A(n16948), .B(n16947), .Y(dpath_mulcore_ary1_a0_sc3_22__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_22__U11(.A(dpath_mulcore_ary1_a0_s_2[22]), .B(dpath_mulcore_ary1_a0_s_1[22]), .Y(n16947));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_22__U10(.A(n9361), .B(n9026), .Y(n16948));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_22__U9(.A(n7276), .B(dpath_mulcore_ary1_a0_sc3_22__z), .Y(dpath_mulcore_a0sum[22]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_23__U12(.A(n16941), .B(n16940), .Y(dpath_mulcore_ary1_a0_sc3_23__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_23__U11(.A(dpath_mulcore_ary1_a0_s_2[23]), .B(dpath_mulcore_ary1_a0_s_1[23]), .Y(n16940));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_23__U10(.A(n9360), .B(n9025), .Y(n16941));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_23__U9(.A(n7275), .B(dpath_mulcore_ary1_a0_sc3_23__z), .Y(dpath_mulcore_a0sum[23]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_24__U12(.A(n16934), .B(n16933), .Y(dpath_mulcore_ary1_a0_sc3_24__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_24__U11(.A(dpath_mulcore_ary1_a0_s_2[24]), .B(dpath_mulcore_ary1_a0_s_1[24]), .Y(n16933));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_24__U10(.A(n9359), .B(n9024), .Y(n16934));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_24__U9(.A(n7274), .B(dpath_mulcore_ary1_a0_sc3_24__z), .Y(dpath_mulcore_a0sum[24]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_25__U12(.A(n16927), .B(n16926), .Y(dpath_mulcore_ary1_a0_sc3_25__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_25__U11(.A(dpath_mulcore_ary1_a0_s_2[25]), .B(dpath_mulcore_ary1_a0_s_1[25]), .Y(n16926));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_25__U10(.A(n9358), .B(n9023), .Y(n16927));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_25__U9(.A(n7273), .B(dpath_mulcore_ary1_a0_sc3_25__z), .Y(dpath_mulcore_a0sum[25]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_26__U12(.A(n16920), .B(n16919), .Y(dpath_mulcore_ary1_a0_sc3_26__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_26__U11(.A(dpath_mulcore_ary1_a0_s_2[26]), .B(dpath_mulcore_ary1_a0_s_1[26]), .Y(n16919));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_26__U10(.A(n9357), .B(n9022), .Y(n16920));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_26__U9(.A(n7272), .B(dpath_mulcore_ary1_a0_sc3_26__z), .Y(dpath_mulcore_a0sum[26]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_27__U12(.A(n16913), .B(n16912), .Y(dpath_mulcore_ary1_a0_sc3_27__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_27__U11(.A(dpath_mulcore_ary1_a0_s_2[27]), .B(dpath_mulcore_ary1_a0_s_1[27]), .Y(n16912));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_27__U10(.A(n9356), .B(n9021), .Y(n16913));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_27__U9(.A(n7271), .B(dpath_mulcore_ary1_a0_sc3_27__z), .Y(dpath_mulcore_a0sum[27]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_28__U12(.A(n16906), .B(n16905), .Y(dpath_mulcore_ary1_a0_sc3_28__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_28__U11(.A(dpath_mulcore_ary1_a0_s_2[28]), .B(dpath_mulcore_ary1_a0_s_1[28]), .Y(n16905));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_28__U10(.A(n9355), .B(n9020), .Y(n16906));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_28__U9(.A(n7270), .B(dpath_mulcore_ary1_a0_sc3_28__z), .Y(dpath_mulcore_a0sum[28]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_29__U12(.A(n16899), .B(n16898), .Y(dpath_mulcore_ary1_a0_sc3_29__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_29__U11(.A(dpath_mulcore_ary1_a0_s_2[29]), .B(dpath_mulcore_ary1_a0_s_1[29]), .Y(n16898));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_29__U10(.A(n9354), .B(n9019), .Y(n16899));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_29__U9(.A(n7269), .B(dpath_mulcore_ary1_a0_sc3_29__z), .Y(dpath_mulcore_a0sum[29]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_30__U12(.A(n16892), .B(n16891), .Y(dpath_mulcore_ary1_a0_sc3_30__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_30__U11(.A(dpath_mulcore_ary1_a0_s_2[30]), .B(dpath_mulcore_ary1_a0_s_1[30]), .Y(n16891));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_30__U10(.A(n9353), .B(n9018), .Y(n16892));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_30__U9(.A(n7268), .B(dpath_mulcore_ary1_a0_sc3_30__z), .Y(dpath_mulcore_a0sum[30]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_31__U12(.A(n16885), .B(n16884), .Y(dpath_mulcore_ary1_a0_sc3_31__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_31__U11(.A(dpath_mulcore_ary1_a0_s_2[31]), .B(dpath_mulcore_ary1_a0_s_1[31]), .Y(n16884));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_31__U10(.A(n9352), .B(n9017), .Y(n16885));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_31__U9(.A(n7267), .B(dpath_mulcore_ary1_a0_sc3_31__z), .Y(dpath_mulcore_a0sum[31]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_32__U12(.A(n16878), .B(n16877), .Y(dpath_mulcore_ary1_a0_sc3_32__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_32__U11(.A(dpath_mulcore_ary1_a0_s_2[32]), .B(dpath_mulcore_ary1_a0_s_1[32]), .Y(n16877));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_32__U10(.A(n9351), .B(n9016), .Y(n16878));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_32__U9(.A(n7266), .B(dpath_mulcore_ary1_a0_sc3_32__z), .Y(dpath_mulcore_a0sum[32]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_33__U12(.A(n16871), .B(n16870), .Y(dpath_mulcore_ary1_a0_sc3_33__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_33__U11(.A(dpath_mulcore_ary1_a0_s_2[33]), .B(dpath_mulcore_ary1_a0_s_1[33]), .Y(n16870));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_33__U10(.A(n9350), .B(n9015), .Y(n16871));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_33__U9(.A(n7265), .B(dpath_mulcore_ary1_a0_sc3_33__z), .Y(dpath_mulcore_a0sum[33]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_34__U12(.A(n16864), .B(n16863), .Y(dpath_mulcore_ary1_a0_sc3_34__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_34__U11(.A(dpath_mulcore_ary1_a0_s_2[34]), .B(dpath_mulcore_ary1_a0_s_1[34]), .Y(n16863));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_34__U10(.A(n9349), .B(n9014), .Y(n16864));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_34__U9(.A(n7264), .B(dpath_mulcore_ary1_a0_sc3_34__z), .Y(dpath_mulcore_a0sum[34]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_35__U12(.A(n16857), .B(n16856), .Y(dpath_mulcore_ary1_a0_sc3_35__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_35__U11(.A(dpath_mulcore_ary1_a0_s_2[35]), .B(dpath_mulcore_ary1_a0_s_1[35]), .Y(n16856));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_35__U10(.A(n9348), .B(n9013), .Y(n16857));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_35__U9(.A(n7263), .B(dpath_mulcore_ary1_a0_sc3_35__z), .Y(dpath_mulcore_a0sum[35]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_36__U12(.A(n16850), .B(n16849), .Y(dpath_mulcore_ary1_a0_sc3_36__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_36__U11(.A(dpath_mulcore_ary1_a0_s_2[36]), .B(dpath_mulcore_ary1_a0_s_1[36]), .Y(n16849));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_36__U10(.A(n9347), .B(n9012), .Y(n16850));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_36__U9(.A(n7262), .B(dpath_mulcore_ary1_a0_sc3_36__z), .Y(dpath_mulcore_a0sum[36]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_37__U12(.A(n16843), .B(n16842), .Y(dpath_mulcore_ary1_a0_sc3_37__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_37__U11(.A(dpath_mulcore_ary1_a0_s_2[37]), .B(dpath_mulcore_ary1_a0_s_1[37]), .Y(n16842));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_37__U10(.A(n9346), .B(n9011), .Y(n16843));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_37__U9(.A(n7261), .B(dpath_mulcore_ary1_a0_sc3_37__z), .Y(dpath_mulcore_a0sum[37]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_38__U12(.A(n16836), .B(n16835), .Y(dpath_mulcore_ary1_a0_sc3_38__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_38__U11(.A(dpath_mulcore_ary1_a0_s_2[38]), .B(dpath_mulcore_ary1_a0_s_1[38]), .Y(n16835));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_38__U10(.A(n9345), .B(n9010), .Y(n16836));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_38__U9(.A(n7260), .B(dpath_mulcore_ary1_a0_sc3_38__z), .Y(dpath_mulcore_a0sum[38]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_39__U12(.A(n16829), .B(n16828), .Y(dpath_mulcore_ary1_a0_sc3_39__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_39__U11(.A(dpath_mulcore_ary1_a0_s_2[39]), .B(dpath_mulcore_ary1_a0_s_1[39]), .Y(n16828));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_39__U10(.A(n9344), .B(n9009), .Y(n16829));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_39__U9(.A(n7259), .B(dpath_mulcore_ary1_a0_sc3_39__z), .Y(dpath_mulcore_a0sum[39]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_40__U12(.A(n16822), .B(n16821), .Y(dpath_mulcore_ary1_a0_sc3_40__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_40__U11(.A(dpath_mulcore_ary1_a0_s_2[40]), .B(dpath_mulcore_ary1_a0_s_1[40]), .Y(n16821));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_40__U10(.A(n9343), .B(n9008), .Y(n16822));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_40__U9(.A(n7258), .B(dpath_mulcore_ary1_a0_sc3_40__z), .Y(dpath_mulcore_a0sum[40]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_41__U12(.A(n16815), .B(n16814), .Y(dpath_mulcore_ary1_a0_sc3_41__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_41__U11(.A(dpath_mulcore_ary1_a0_s_2[41]), .B(dpath_mulcore_ary1_a0_s_1[41]), .Y(n16814));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_41__U10(.A(n9342), .B(n9007), .Y(n16815));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_41__U9(.A(n7257), .B(dpath_mulcore_ary1_a0_sc3_41__z), .Y(dpath_mulcore_a0sum[41]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_42__U12(.A(n16808), .B(n16807), .Y(dpath_mulcore_ary1_a0_sc3_42__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_42__U11(.A(dpath_mulcore_ary1_a0_s_2[42]), .B(dpath_mulcore_ary1_a0_s_1[42]), .Y(n16807));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_42__U10(.A(n9341), .B(n9006), .Y(n16808));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_42__U9(.A(n7256), .B(dpath_mulcore_ary1_a0_sc3_42__z), .Y(dpath_mulcore_a0sum[42]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_43__U12(.A(n16801), .B(n16800), .Y(dpath_mulcore_ary1_a0_sc3_43__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_43__U11(.A(dpath_mulcore_ary1_a0_s_2[43]), .B(dpath_mulcore_ary1_a0_s_1[43]), .Y(n16800));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_43__U10(.A(n9340), .B(n9005), .Y(n16801));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_43__U9(.A(n7255), .B(dpath_mulcore_ary1_a0_sc3_43__z), .Y(dpath_mulcore_a0sum[43]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_44__U12(.A(n16794), .B(n16793), .Y(dpath_mulcore_ary1_a0_sc3_44__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_44__U11(.A(dpath_mulcore_ary1_a0_s_2[44]), .B(dpath_mulcore_ary1_a0_s_1[44]), .Y(n16793));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_44__U10(.A(n9339), .B(n9004), .Y(n16794));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_44__U9(.A(n7254), .B(dpath_mulcore_ary1_a0_sc3_44__z), .Y(dpath_mulcore_a0sum[44]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_45__U12(.A(n16787), .B(n16786), .Y(dpath_mulcore_ary1_a0_sc3_45__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_45__U11(.A(dpath_mulcore_ary1_a0_s_2[45]), .B(dpath_mulcore_ary1_a0_s_1[45]), .Y(n16786));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_45__U10(.A(n9338), .B(n9003), .Y(n16787));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_45__U9(.A(n7253), .B(dpath_mulcore_ary1_a0_sc3_45__z), .Y(dpath_mulcore_a0sum[45]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_46__U12(.A(n16780), .B(n16779), .Y(dpath_mulcore_ary1_a0_sc3_46__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_46__U11(.A(dpath_mulcore_ary1_a0_s_2[46]), .B(dpath_mulcore_ary1_a0_s_1[46]), .Y(n16779));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_46__U10(.A(n9337), .B(n9002), .Y(n16780));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_46__U9(.A(n7252), .B(dpath_mulcore_ary1_a0_sc3_46__z), .Y(dpath_mulcore_a0sum[46]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_47__U12(.A(n16773), .B(n16772), .Y(dpath_mulcore_ary1_a0_sc3_47__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_47__U11(.A(dpath_mulcore_ary1_a0_s_2[47]), .B(dpath_mulcore_ary1_a0_s_1[47]), .Y(n16772));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_47__U10(.A(n9336), .B(n9001), .Y(n16773));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_47__U9(.A(n7251), .B(dpath_mulcore_ary1_a0_sc3_47__z), .Y(dpath_mulcore_a0sum[47]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_48__U12(.A(n16766), .B(n16765), .Y(dpath_mulcore_ary1_a0_sc3_48__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_48__U11(.A(dpath_mulcore_ary1_a0_s_2[48]), .B(dpath_mulcore_ary1_a0_s_1[48]), .Y(n16765));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_48__U10(.A(n9335), .B(n9000), .Y(n16766));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_48__U9(.A(n7250), .B(dpath_mulcore_ary1_a0_sc3_48__z), .Y(dpath_mulcore_a0sum[48]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_49__U12(.A(n16759), .B(n16758), .Y(dpath_mulcore_ary1_a0_sc3_49__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_49__U11(.A(dpath_mulcore_ary1_a0_s_2[49]), .B(dpath_mulcore_ary1_a0_s_1[49]), .Y(n16758));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_49__U10(.A(n9334), .B(n8999), .Y(n16759));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_49__U9(.A(n7249), .B(dpath_mulcore_ary1_a0_sc3_49__z), .Y(dpath_mulcore_a0sum[49]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_50__U12(.A(n16752), .B(n16751), .Y(dpath_mulcore_ary1_a0_sc3_50__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_50__U11(.A(dpath_mulcore_ary1_a0_s_2[50]), .B(dpath_mulcore_ary1_a0_s_1[50]), .Y(n16751));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_50__U10(.A(n9333), .B(n8998), .Y(n16752));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_50__U9(.A(n7248), .B(dpath_mulcore_ary1_a0_sc3_50__z), .Y(dpath_mulcore_a0sum[50]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_51__U12(.A(n16745), .B(n16744), .Y(dpath_mulcore_ary1_a0_sc3_51__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_51__U11(.A(dpath_mulcore_ary1_a0_s_2[51]), .B(dpath_mulcore_ary1_a0_s_1[51]), .Y(n16744));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_51__U10(.A(n9332), .B(n8997), .Y(n16745));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_51__U9(.A(n7247), .B(dpath_mulcore_ary1_a0_sc3_51__z), .Y(dpath_mulcore_a0sum[51]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_52__U12(.A(n16738), .B(n16737), .Y(dpath_mulcore_ary1_a0_sc3_52__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_52__U11(.A(dpath_mulcore_ary1_a0_s_2[52]), .B(dpath_mulcore_ary1_a0_s_1[52]), .Y(n16737));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_52__U10(.A(n9331), .B(n8996), .Y(n16738));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_52__U9(.A(n7246), .B(dpath_mulcore_ary1_a0_sc3_52__z), .Y(dpath_mulcore_a0sum[52]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_53__U12(.A(n16731), .B(n16730), .Y(dpath_mulcore_ary1_a0_sc3_53__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_53__U11(.A(dpath_mulcore_ary1_a0_s_2[53]), .B(dpath_mulcore_ary1_a0_s_1[53]), .Y(n16730));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_53__U10(.A(n9330), .B(n8995), .Y(n16731));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_53__U9(.A(n7245), .B(dpath_mulcore_ary1_a0_sc3_53__z), .Y(dpath_mulcore_a0sum[53]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_54__U12(.A(n16724), .B(n16723), .Y(dpath_mulcore_ary1_a0_sc3_54__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_54__U11(.A(dpath_mulcore_ary1_a0_s_2[54]), .B(dpath_mulcore_ary1_a0_s_1[54]), .Y(n16723));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_54__U10(.A(n9329), .B(n8994), .Y(n16724));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_54__U9(.A(n7244), .B(dpath_mulcore_ary1_a0_sc3_54__z), .Y(dpath_mulcore_a0sum[54]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_55__U12(.A(n16717), .B(n16716), .Y(dpath_mulcore_ary1_a0_sc3_55__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_55__U11(.A(dpath_mulcore_ary1_a0_s_2[55]), .B(dpath_mulcore_ary1_a0_s_1[55]), .Y(n16716));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_55__U10(.A(n9328), .B(n8993), .Y(n16717));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_55__U9(.A(n7243), .B(dpath_mulcore_ary1_a0_sc3_55__z), .Y(dpath_mulcore_a0sum[55]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_56__U12(.A(n16710), .B(n16709), .Y(dpath_mulcore_ary1_a0_sc3_56__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_56__U11(.A(dpath_mulcore_ary1_a0_s_2[56]), .B(dpath_mulcore_ary1_a0_s_1[56]), .Y(n16709));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_56__U10(.A(n9327), .B(n8992), .Y(n16710));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_56__U9(.A(n7242), .B(dpath_mulcore_ary1_a0_sc3_56__z), .Y(dpath_mulcore_a0sum[56]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_57__U12(.A(n16703), .B(n16702), .Y(dpath_mulcore_ary1_a0_sc3_57__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_57__U11(.A(dpath_mulcore_ary1_a0_s_2[57]), .B(dpath_mulcore_ary1_a0_s_1[57]), .Y(n16702));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_57__U10(.A(n9326), .B(n8991), .Y(n16703));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_57__U9(.A(n7241), .B(dpath_mulcore_ary1_a0_sc3_57__z), .Y(dpath_mulcore_a0sum[57]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_58__U12(.A(n16696), .B(n16695), .Y(dpath_mulcore_ary1_a0_sc3_58__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_58__U11(.A(dpath_mulcore_ary1_a0_s_2[58]), .B(dpath_mulcore_ary1_a0_s_1[58]), .Y(n16695));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_58__U10(.A(n9325), .B(n8990), .Y(n16696));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_58__U9(.A(n7240), .B(dpath_mulcore_ary1_a0_sc3_58__z), .Y(dpath_mulcore_a0sum[58]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_59__U12(.A(n16689), .B(n16688), .Y(dpath_mulcore_ary1_a0_sc3_59__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_59__U11(.A(dpath_mulcore_ary1_a0_s_2[59]), .B(dpath_mulcore_ary1_a0_s_1[59]), .Y(n16688));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_59__U10(.A(n9324), .B(n8989), .Y(n16689));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_59__U9(.A(n7239), .B(dpath_mulcore_ary1_a0_sc3_59__z), .Y(dpath_mulcore_a0sum[59]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_60__U12(.A(n16682), .B(n16681), .Y(dpath_mulcore_ary1_a0_sc3_60__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_60__U11(.A(dpath_mulcore_ary1_a0_s_2[60]), .B(dpath_mulcore_ary1_a0_s_1[60]), .Y(n16681));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_60__U10(.A(n9323), .B(n8988), .Y(n16682));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_60__U9(.A(n7238), .B(dpath_mulcore_ary1_a0_sc3_60__z), .Y(dpath_mulcore_a0sum[60]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_61__U12(.A(n16675), .B(n16674), .Y(dpath_mulcore_ary1_a0_sc3_61__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_61__U11(.A(dpath_mulcore_ary1_a0_s_2[61]), .B(dpath_mulcore_ary1_a0_s_1[61]), .Y(n16674));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_61__U10(.A(n9322), .B(n8987), .Y(n16675));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_61__U9(.A(n7237), .B(dpath_mulcore_ary1_a0_sc3_61__z), .Y(dpath_mulcore_a0sum[61]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_62__U12(.A(n16668), .B(n16667), .Y(dpath_mulcore_ary1_a0_sc3_62__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_62__U11(.A(dpath_mulcore_ary1_a0_s_2[62]), .B(dpath_mulcore_ary1_a0_s_1[62]), .Y(n16667));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_62__U10(.A(n9321), .B(n8986), .Y(n16668));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_62__U9(.A(n7236), .B(dpath_mulcore_ary1_a0_sc3_62__z), .Y(dpath_mulcore_a0sum[62]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_63__U12(.A(n16661), .B(n16660), .Y(dpath_mulcore_ary1_a0_sc3_63__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_63__U11(.A(dpath_mulcore_ary1_a0_s_2[63]), .B(dpath_mulcore_ary1_a0_s_1[63]), .Y(n16660));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_63__U10(.A(n9320), .B(n8985), .Y(n16661));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_63__U9(.A(n7235), .B(dpath_mulcore_ary1_a0_sc3_63__z), .Y(dpath_mulcore_a0sum[63]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_64__U12(.A(n16654), .B(n16653), .Y(dpath_mulcore_ary1_a0_sc3_64__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_64__U11(.A(dpath_mulcore_ary1_a0_s_2[64]), .B(dpath_mulcore_ary1_a0_s_1[64]), .Y(n16653));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_64__U10(.A(n9319), .B(n8984), .Y(n16654));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_64__U9(.A(n7234), .B(dpath_mulcore_ary1_a0_sc3_64__z), .Y(dpath_mulcore_a0sum[64]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_65__U12(.A(n16647), .B(n16646), .Y(dpath_mulcore_ary1_a0_sc3_65__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_65__U11(.A(dpath_mulcore_ary1_a0_s_2[65]), .B(dpath_mulcore_ary1_a0_s_1[65]), .Y(n16646));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_65__U10(.A(n9318), .B(n8983), .Y(n16647));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_65__U9(.A(n7233), .B(dpath_mulcore_ary1_a0_sc3_65__z), .Y(dpath_mulcore_a0sum[65]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_66__U12(.A(n16640), .B(n16639), .Y(dpath_mulcore_ary1_a0_sc3_66__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_66__U11(.A(dpath_mulcore_ary1_a0_s_2[66]), .B(dpath_mulcore_ary1_a0_s_1[66]), .Y(n16639));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_66__U10(.A(n9317), .B(n8982), .Y(n16640));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_66__U9(.A(n7232), .B(dpath_mulcore_ary1_a0_sc3_66__z), .Y(dpath_mulcore_a0sum[66]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_67__U12(.A(n16633), .B(n16632), .Y(dpath_mulcore_ary1_a0_sc3_67__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_67__U11(.A(dpath_mulcore_ary1_a0_s_2[67]), .B(dpath_mulcore_ary1_a0_s_1[67]), .Y(n16632));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_67__U10(.A(n9316), .B(n8981), .Y(n16633));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_67__U9(.A(n7231), .B(dpath_mulcore_ary1_a0_sc3_67__z), .Y(dpath_mulcore_a0sum[67]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_68__U12(.A(n16626), .B(n16625), .Y(dpath_mulcore_ary1_a0_sc3_68__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_68__U11(.A(dpath_mulcore_ary1_a0_s_2[68]), .B(dpath_mulcore_ary1_a0_s_1[68]), .Y(n16625));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_68__U10(.A(n9315), .B(n8980), .Y(n16626));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_68__U9(.A(n7230), .B(dpath_mulcore_ary1_a0_sc3_68__z), .Y(dpath_mulcore_a0sum[68]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_69__U12(.A(n16619), .B(n16618), .Y(dpath_mulcore_ary1_a0_sc3_69__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_69__U11(.A(dpath_mulcore_ary1_a0_s_2[69]), .B(dpath_mulcore_ary1_a0_s_1[69]), .Y(n16618));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_69__U10(.A(n9314), .B(n8979), .Y(n16619));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_69__U9(.A(n7229), .B(dpath_mulcore_ary1_a0_sc3_69__z), .Y(dpath_mulcore_a0sum[69]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_70__U12(.A(n16612), .B(n16611), .Y(dpath_mulcore_ary1_a0_sc3_70__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_70__U11(.A(dpath_mulcore_ary1_a0_s_2[70]), .B(n10026), .Y(n16611));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_70__U10(.A(n9313), .B(n8978), .Y(n16612));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_70__U9(.A(n7228), .B(dpath_mulcore_ary1_a0_sc3_70__z), .Y(dpath_mulcore_a0sum[70]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_76__U12(.A(n8289), .B(n1), .Y(dpath_mulcore_ary1_a0_sc3_76__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_76__U9(.A(n16588), .B(dpath_mulcore_ary1_a0_sc3_76__z), .Y(dpath_mulcore_a0sum[76]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_72__U12(.A(n8288), .B(n16603), .Y(dpath_mulcore_ary1_a0_sc3_72__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_72__U11(.A(dpath_mulcore_ary1_a0_s_2[72]), .B(dpath_mulcore_ary1_a0_s1[66]), .Y(n16603));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_72__U9(.A(n7395), .B(dpath_mulcore_ary1_a0_sc3_72__z), .Y(dpath_mulcore_a0sum[72]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_73__U12(.A(n8292), .B(n16599), .Y(dpath_mulcore_ary1_a0_sc3_73__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_73__U11(.A(dpath_mulcore_ary1_a0_s_2[73]), .B(dpath_mulcore_ary1_a0_s1[67]), .Y(n16599));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_73__U9(.A(n16600), .B(dpath_mulcore_ary1_a0_sc3_73__z), .Y(dpath_mulcore_a0sum[73]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_74__U12(.A(n8291), .B(n16595), .Y(dpath_mulcore_ary1_a0_sc3_74__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_74__U11(.A(dpath_mulcore_ary1_a0_s_2[74]), .B(dpath_mulcore_ary1_a0_I1_I2_net073), .Y(n16595));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_74__U9(.A(n16596), .B(dpath_mulcore_ary1_a0_sc3_74__z), .Y(dpath_mulcore_a0sum[74]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_75__U12(.A(n8290), .B(n16591), .Y(dpath_mulcore_ary1_a0_sc3_75__z));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_75__U11(.A(dpath_mulcore_ary1_a0_s_2[75]), .B(n9484), .Y(n16591));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_75__U9(.A(n16592), .B(dpath_mulcore_ary1_a0_sc3_75__z), .Y(dpath_mulcore_a0sum[75]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_sc1_64__U4(.A(n7485), .B(n8754), .Y(n16585));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_sc1_64__U1(.A(n7486), .B(n16585), .Y(dpath_mulcore_ary1_a0_s1[64]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_sc1_65__U4(.A(n7484), .B(n9475), .Y(n16582));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_sc1_65__U1(.A(n7483), .B(n16582), .Y(dpath_mulcore_ary1_a0_s1[65]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_sc1_66__U1(.A(n7482), .B(dpath_mulcore_ary1_a0_I1_I2_net38), .Y(dpath_mulcore_ary1_a0_s1[66]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_sc1_67__U1(.A(n7481), .B(n9476), .Y(dpath_mulcore_ary1_a0_s1[67]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_sc1_3__U4(.A(n7479), .B(n8448), .Y(n16577));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_sc1_3__U1(.A(n8383), .B(n16577), .Y(dpath_mulcore_ary1_a0_s2[3]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_sc1_2__U4(.A(n7480), .B(n9853), .Y(n16574));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_sc1_2__U1(.A(n8384), .B(n16574), .Y(dpath_mulcore_ary1_a0_s2[2]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_63__sc1_U4(.A(n7419), .B(n8388), .Y(n16572));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I2_sc1_64__U4(.A(n7418), .B(n8977), .Y(n16570));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I2_sc1_65__U4(.A(n7417), .B(n9483), .Y(n16568));
XOR2X1 mul_dpath_mulcore_array2_sc1_67__U1(.A(dpath_mulcore_a1c[50]), .B(dpath_mulcore_a1s[51]), .Y(dpath_mulcore_array2_s1[67]));
XOR2X1 mul_dpath_mulcore_array2_sc1_0__U4(.A(dpath_mulcore_ps[32]), .B(dpath_mulcore_pc[31]), .Y(n16564));
XOR2X1 mul_dpath_mulcore_array2_sc1_0__U1(.A(dpath_mulcore_a0s[0]), .B(n16564), .Y(dpath_mulcore_array2_s1[0]));
XOR2X1 mul_dpath_mulcore_array2_acc_15__U4(.A(n8269), .B(dpath_mulcore_array2_s3[15]), .Y(n16562));
XOR2X1 mul_dpath_mulcore_array2_acc_16__U4(.A(n8268), .B(dpath_mulcore_array2_s3[16]), .Y(n16559));
XOR2X1 mul_dpath_mulcore_array2_acc_16__U1(.A(n8312), .B(n16559), .Y(dpath_mulcore_psum[16]));
XOR2X1 mul_dpath_mulcore_array2_acc_17__U4(.A(n8267), .B(dpath_mulcore_array2_s3[17]), .Y(n16556));
XOR2X1 mul_dpath_mulcore_array2_acc_17__U1(.A(n8311), .B(n16556), .Y(dpath_mulcore_psum[17]));
XOR2X1 mul_dpath_mulcore_array2_acc_18__U4(.A(n8266), .B(dpath_mulcore_array2_s3[18]), .Y(n16553));
XOR2X1 mul_dpath_mulcore_array2_acc_18__U1(.A(n8310), .B(n16553), .Y(dpath_mulcore_psum[18]));
XOR2X1 mul_dpath_mulcore_array2_acc_19__U4(.A(n8265), .B(dpath_mulcore_array2_s3[19]), .Y(n16550));
XOR2X1 mul_dpath_mulcore_array2_acc_19__U1(.A(n8309), .B(n16550), .Y(dpath_mulcore_psum[19]));
XOR2X1 mul_dpath_mulcore_array2_sc2_68__U4(.A(dpath_mulcore_array2_s1[68]), .B(n8974), .Y(n16547));
XOR2X1 mul_dpath_mulcore_array2_sc2_68__U1(.A(dpath_mulcore_a0c[67]), .B(n16547), .Y(dpath_mulcore_array2_s2[68]));
XOR2X1 mul_dpath_mulcore_array2_sc2_69__U4(.A(dpath_mulcore_array2_s1[69]), .B(n8961), .Y(n16544));
XOR2X1 mul_dpath_mulcore_array2_sc2_69__U1(.A(dpath_mulcore_a0c[68]), .B(n16544), .Y(dpath_mulcore_array2_s2[69]));
XOR2X1 mul_dpath_mulcore_array2_sc2_70__U4(.A(dpath_mulcore_array2_s1[70]), .B(n8960), .Y(n16541));
XOR2X1 mul_dpath_mulcore_array2_sc2_70__U1(.A(dpath_mulcore_a0c[69]), .B(n16541), .Y(dpath_mulcore_array2_s2[70]));
XOR2X1 mul_dpath_mulcore_array2_sc2_71__U4(.A(dpath_mulcore_array2_s1[71]), .B(n8959), .Y(n16538));
XOR2X1 mul_dpath_mulcore_array2_sc2_71__U1(.A(dpath_mulcore_a0c[70]), .B(n16538), .Y(dpath_mulcore_array2_s2[71]));
XOR2X1 mul_dpath_mulcore_array2_sc2_72__U4(.A(dpath_mulcore_array2_s1[72]), .B(n8958), .Y(n16535));
XOR2X1 mul_dpath_mulcore_array2_sc2_72__U1(.A(dpath_mulcore_a0c[71]), .B(n16535), .Y(dpath_mulcore_array2_s2[72]));
XOR2X1 mul_dpath_mulcore_array2_sc2_73__U4(.A(dpath_mulcore_array2_s1[73]), .B(n8957), .Y(n16532));
XOR2X1 mul_dpath_mulcore_array2_sc2_73__U1(.A(dpath_mulcore_a0c[72]), .B(n16532), .Y(dpath_mulcore_array2_s2[73]));
XOR2X1 mul_dpath_mulcore_array2_sc2_74__U4(.A(dpath_mulcore_array2_s1[74]), .B(n8956), .Y(n16529));
XOR2X1 mul_dpath_mulcore_array2_sc2_74__U1(.A(dpath_mulcore_a0c[73]), .B(n16529), .Y(dpath_mulcore_array2_s2[74]));
XOR2X1 mul_dpath_mulcore_array2_sc2_75__U4(.A(dpath_mulcore_array2_s1[75]), .B(n8955), .Y(n16526));
XOR2X1 mul_dpath_mulcore_array2_sc2_75__U1(.A(dpath_mulcore_a0c[74]), .B(n16526), .Y(dpath_mulcore_array2_s2[75]));
XOR2X1 mul_dpath_mulcore_array2_sc2_76__U4(.A(dpath_mulcore_array2_s1[76]), .B(n8954), .Y(n16523));
XOR2X1 mul_dpath_mulcore_array2_sc2_76__U1(.A(dpath_mulcore_a0c[75]), .B(n16523), .Y(dpath_mulcore_array2_s2[76]));
XOR2X1 mul_dpath_mulcore_array2_sc2_77__U4(.A(dpath_mulcore_array2_s1[77]), .B(n8953), .Y(n16520));
XOR2X1 mul_dpath_mulcore_array2_sc2_77__U1(.A(dpath_mulcore_a0c[76]), .B(n16520), .Y(dpath_mulcore_array2_s2[77]));
XOR2X1 mul_dpath_mulcore_array2_sc2_78__U4(.A(dpath_mulcore_array2_s1[78]), .B(n8952), .Y(n16517));
XOR2X1 mul_dpath_mulcore_array2_sc2_78__U1(.A(dpath_mulcore_a0c[77]), .B(n16517), .Y(dpath_mulcore_array2_s2[78]));
XOR2X1 mul_dpath_mulcore_array2_sc2_79__U4(.A(dpath_mulcore_array2_s1[79]), .B(n8951), .Y(n16514));
XOR2X1 mul_dpath_mulcore_array2_sc2_79__U1(.A(dpath_mulcore_a0c[78]), .B(n16514), .Y(dpath_mulcore_array2_s2[79]));
XOR2X1 mul_dpath_mulcore_array2_sc2_80__U4(.A(dpath_mulcore_array2_s1[80]), .B(n8950), .Y(n16511));
XOR2X1 mul_dpath_mulcore_array2_sc2_80__U1(.A(dpath_mulcore_a0c[79]), .B(n16511), .Y(dpath_mulcore_array2_s2[80]));
XOR2X1 mul_dpath_mulcore_array2_sc2_81__U4(.A(dpath_mulcore_array2_s1[81]), .B(n8949), .Y(dpath_mulcore_array2_s2[81]));
XOR2X1 mul_dpath_mulcore_array2_sc1_20__U4(.A(dpath_mulcore_ps[52]), .B(dpath_mulcore_pc[51]), .Y(n16507));
XOR2X1 mul_dpath_mulcore_array2_sc1_20__U1(.A(dpath_mulcore_a1s[4]), .B(n16507), .Y(dpath_mulcore_array2_s1[20]));
XOR2X1 mul_dpath_mulcore_array2_sc1_21__U4(.A(dpath_mulcore_ps[53]), .B(dpath_mulcore_pc[52]), .Y(n16504));
XOR2X1 mul_dpath_mulcore_array2_sc1_21__U1(.A(dpath_mulcore_a1s[5]), .B(n16504), .Y(dpath_mulcore_array2_s1[21]));
XOR2X1 mul_dpath_mulcore_array2_sc1_22__U4(.A(dpath_mulcore_ps[54]), .B(dpath_mulcore_pc[53]), .Y(n16501));
XOR2X1 mul_dpath_mulcore_array2_sc1_22__U1(.A(dpath_mulcore_a1s[6]), .B(n16501), .Y(dpath_mulcore_array2_s1[22]));
XOR2X1 mul_dpath_mulcore_array2_sc1_23__U4(.A(dpath_mulcore_ps[55]), .B(dpath_mulcore_pc[54]), .Y(n16498));
XOR2X1 mul_dpath_mulcore_array2_sc1_23__U1(.A(dpath_mulcore_a1s[7]), .B(n16498), .Y(dpath_mulcore_array2_s1[23]));
XOR2X1 mul_dpath_mulcore_array2_sc1_24__U4(.A(dpath_mulcore_ps[56]), .B(dpath_mulcore_pc[55]), .Y(n16495));
XOR2X1 mul_dpath_mulcore_array2_sc1_24__U1(.A(dpath_mulcore_a1s[8]), .B(n16495), .Y(dpath_mulcore_array2_s1[24]));
XOR2X1 mul_dpath_mulcore_array2_sc1_25__U4(.A(dpath_mulcore_ps[57]), .B(dpath_mulcore_pc[56]), .Y(n16492));
XOR2X1 mul_dpath_mulcore_array2_sc1_25__U1(.A(dpath_mulcore_a1s[9]), .B(n16492), .Y(dpath_mulcore_array2_s1[25]));
XOR2X1 mul_dpath_mulcore_array2_sc1_26__U4(.A(dpath_mulcore_ps[58]), .B(dpath_mulcore_pc[57]), .Y(n16489));
XOR2X1 mul_dpath_mulcore_array2_sc1_26__U1(.A(dpath_mulcore_a1s[10]), .B(n16489), .Y(dpath_mulcore_array2_s1[26]));
XOR2X1 mul_dpath_mulcore_array2_sc1_27__U4(.A(dpath_mulcore_ps[59]), .B(dpath_mulcore_pc[58]), .Y(n16486));
XOR2X1 mul_dpath_mulcore_array2_sc1_27__U1(.A(dpath_mulcore_a1s[11]), .B(n16486), .Y(dpath_mulcore_array2_s1[27]));
XOR2X1 mul_dpath_mulcore_array2_sc1_28__U4(.A(dpath_mulcore_ps[60]), .B(dpath_mulcore_pc[59]), .Y(n16483));
XOR2X1 mul_dpath_mulcore_array2_sc1_28__U1(.A(dpath_mulcore_a1s[12]), .B(n16483), .Y(dpath_mulcore_array2_s1[28]));
XOR2X1 mul_dpath_mulcore_array2_sc1_29__U4(.A(dpath_mulcore_ps[61]), .B(dpath_mulcore_pc[60]), .Y(n16480));
XOR2X1 mul_dpath_mulcore_array2_sc1_29__U1(.A(dpath_mulcore_a1s[13]), .B(n16480), .Y(dpath_mulcore_array2_s1[29]));
XOR2X1 mul_dpath_mulcore_array2_sc1_30__U4(.A(dpath_mulcore_ps[62]), .B(dpath_mulcore_pc[61]), .Y(n16477));
XOR2X1 mul_dpath_mulcore_array2_sc1_30__U1(.A(dpath_mulcore_a1s[14]), .B(n16477), .Y(dpath_mulcore_array2_s1[30]));
XOR2X1 mul_dpath_mulcore_array2_sc1_31__U4(.A(dpath_mulcore_ps[63]), .B(dpath_mulcore_pc[62]), .Y(n16474));
XOR2X1 mul_dpath_mulcore_array2_sc1_31__U1(.A(dpath_mulcore_a1s[15]), .B(n16474), .Y(dpath_mulcore_array2_s1[31]));
XOR2X1 mul_dpath_mulcore_array2_sc1_32__U4(.A(dpath_mulcore_ps[64]), .B(dpath_mulcore_pc[63]), .Y(n16471));
XOR2X1 mul_dpath_mulcore_array2_sc1_32__U1(.A(dpath_mulcore_a1s[16]), .B(n16471), .Y(dpath_mulcore_array2_s1[32]));
XOR2X1 mul_dpath_mulcore_array2_sc1_33__U4(.A(dpath_mulcore_ps[65]), .B(dpath_mulcore_pc[64]), .Y(n16468));
XOR2X1 mul_dpath_mulcore_array2_sc1_33__U1(.A(dpath_mulcore_a1s[17]), .B(n16468), .Y(dpath_mulcore_array2_s1[33]));
XOR2X1 mul_dpath_mulcore_array2_sc1_34__U4(.A(dpath_mulcore_ps[66]), .B(dpath_mulcore_pc[65]), .Y(n16465));
XOR2X1 mul_dpath_mulcore_array2_sc1_34__U1(.A(dpath_mulcore_a1s[18]), .B(n16465), .Y(dpath_mulcore_array2_s1[34]));
XOR2X1 mul_dpath_mulcore_array2_sc1_35__U4(.A(dpath_mulcore_ps[67]), .B(dpath_mulcore_pc[66]), .Y(n16462));
XOR2X1 mul_dpath_mulcore_array2_sc1_35__U1(.A(dpath_mulcore_a1s[19]), .B(n16462), .Y(dpath_mulcore_array2_s1[35]));
XOR2X1 mul_dpath_mulcore_array2_sc1_36__U4(.A(dpath_mulcore_ps[68]), .B(dpath_mulcore_pc[67]), .Y(n16459));
XOR2X1 mul_dpath_mulcore_array2_sc1_36__U1(.A(dpath_mulcore_a1s[20]), .B(n16459), .Y(dpath_mulcore_array2_s1[36]));
XOR2X1 mul_dpath_mulcore_array2_sc1_37__U4(.A(dpath_mulcore_ps[69]), .B(dpath_mulcore_pc[68]), .Y(n16456));
XOR2X1 mul_dpath_mulcore_array2_sc1_37__U1(.A(dpath_mulcore_a1s[21]), .B(n16456), .Y(dpath_mulcore_array2_s1[37]));
XOR2X1 mul_dpath_mulcore_array2_sc1_38__U4(.A(dpath_mulcore_ps[70]), .B(dpath_mulcore_pc[69]), .Y(n16453));
XOR2X1 mul_dpath_mulcore_array2_sc1_38__U1(.A(dpath_mulcore_a1s[22]), .B(n16453), .Y(dpath_mulcore_array2_s1[38]));
XOR2X1 mul_dpath_mulcore_array2_sc1_39__U4(.A(dpath_mulcore_ps[71]), .B(dpath_mulcore_pc[70]), .Y(n16450));
XOR2X1 mul_dpath_mulcore_array2_sc1_39__U1(.A(dpath_mulcore_a1s[23]), .B(n16450), .Y(dpath_mulcore_array2_s1[39]));
XOR2X1 mul_dpath_mulcore_array2_sc1_40__U4(.A(dpath_mulcore_ps[72]), .B(dpath_mulcore_pc[71]), .Y(n16447));
XOR2X1 mul_dpath_mulcore_array2_sc1_40__U1(.A(dpath_mulcore_a1s[24]), .B(n16447), .Y(dpath_mulcore_array2_s1[40]));
XOR2X1 mul_dpath_mulcore_array2_sc1_41__U4(.A(dpath_mulcore_ps[73]), .B(dpath_mulcore_pc[72]), .Y(n16444));
XOR2X1 mul_dpath_mulcore_array2_sc1_41__U1(.A(dpath_mulcore_a1s[25]), .B(n16444), .Y(dpath_mulcore_array2_s1[41]));
XOR2X1 mul_dpath_mulcore_array2_sc1_42__U4(.A(dpath_mulcore_ps[74]), .B(dpath_mulcore_pc[73]), .Y(n16441));
XOR2X1 mul_dpath_mulcore_array2_sc1_42__U1(.A(dpath_mulcore_a1s[26]), .B(n16441), .Y(dpath_mulcore_array2_s1[42]));
XOR2X1 mul_dpath_mulcore_array2_sc1_43__U4(.A(dpath_mulcore_ps[75]), .B(dpath_mulcore_pc[74]), .Y(n16438));
XOR2X1 mul_dpath_mulcore_array2_sc1_43__U1(.A(dpath_mulcore_a1s[27]), .B(n16438), .Y(dpath_mulcore_array2_s1[43]));
XOR2X1 mul_dpath_mulcore_array2_sc1_44__U4(.A(dpath_mulcore_ps[76]), .B(dpath_mulcore_pc[75]), .Y(n16435));
XOR2X1 mul_dpath_mulcore_array2_sc1_44__U1(.A(dpath_mulcore_a1s[28]), .B(n16435), .Y(dpath_mulcore_array2_s1[44]));
XOR2X1 mul_dpath_mulcore_array2_sc1_45__U4(.A(dpath_mulcore_ps[77]), .B(dpath_mulcore_pc[76]), .Y(n16432));
XOR2X1 mul_dpath_mulcore_array2_sc1_45__U1(.A(dpath_mulcore_a1s[29]), .B(n16432), .Y(dpath_mulcore_array2_s1[45]));
XOR2X1 mul_dpath_mulcore_array2_sc1_46__U4(.A(dpath_mulcore_ps[78]), .B(dpath_mulcore_pc[77]), .Y(n16429));
XOR2X1 mul_dpath_mulcore_array2_sc1_46__U1(.A(dpath_mulcore_a1s[30]), .B(n16429), .Y(dpath_mulcore_array2_s1[46]));
XOR2X1 mul_dpath_mulcore_array2_sc1_47__U4(.A(dpath_mulcore_ps[79]), .B(dpath_mulcore_pc[78]), .Y(n16426));
XOR2X1 mul_dpath_mulcore_array2_sc1_47__U1(.A(dpath_mulcore_a1s[31]), .B(n16426), .Y(dpath_mulcore_array2_s1[47]));
XOR2X1 mul_dpath_mulcore_array2_sc1_48__U4(.A(dpath_mulcore_ps[80]), .B(dpath_mulcore_pc[79]), .Y(n16423));
XOR2X1 mul_dpath_mulcore_array2_sc1_48__U1(.A(dpath_mulcore_a1s[32]), .B(n16423), .Y(dpath_mulcore_array2_s1[48]));
XOR2X1 mul_dpath_mulcore_array2_sc1_49__U4(.A(dpath_mulcore_ps[81]), .B(dpath_mulcore_pc[80]), .Y(n16420));
XOR2X1 mul_dpath_mulcore_array2_sc1_49__U1(.A(dpath_mulcore_a1s[33]), .B(n16420), .Y(dpath_mulcore_array2_s1[49]));
XOR2X1 mul_dpath_mulcore_array2_sc1_50__U4(.A(dpath_mulcore_ps[82]), .B(dpath_mulcore_pc[81]), .Y(n16417));
XOR2X1 mul_dpath_mulcore_array2_sc1_50__U1(.A(dpath_mulcore_a1s[34]), .B(n16417), .Y(dpath_mulcore_array2_s1[50]));
XOR2X1 mul_dpath_mulcore_array2_sc1_51__U4(.A(dpath_mulcore_ps[83]), .B(dpath_mulcore_pc[82]), .Y(n16414));
XOR2X1 mul_dpath_mulcore_array2_sc1_51__U1(.A(dpath_mulcore_a1s[35]), .B(n16414), .Y(dpath_mulcore_array2_s1[51]));
XOR2X1 mul_dpath_mulcore_array2_sc1_52__U4(.A(dpath_mulcore_ps[84]), .B(dpath_mulcore_pc[83]), .Y(n16411));
XOR2X1 mul_dpath_mulcore_array2_sc1_52__U1(.A(dpath_mulcore_a1s[36]), .B(n16411), .Y(dpath_mulcore_array2_s1[52]));
XOR2X1 mul_dpath_mulcore_array2_sc1_53__U4(.A(dpath_mulcore_ps[85]), .B(dpath_mulcore_pc[84]), .Y(n16408));
XOR2X1 mul_dpath_mulcore_array2_sc1_53__U1(.A(dpath_mulcore_a1s[37]), .B(n16408), .Y(dpath_mulcore_array2_s1[53]));
XOR2X1 mul_dpath_mulcore_array2_sc1_54__U4(.A(dpath_mulcore_ps[86]), .B(dpath_mulcore_pc[85]), .Y(n16405));
XOR2X1 mul_dpath_mulcore_array2_sc1_54__U1(.A(dpath_mulcore_a1s[38]), .B(n16405), .Y(dpath_mulcore_array2_s1[54]));
XOR2X1 mul_dpath_mulcore_array2_sc1_55__U4(.A(dpath_mulcore_ps[87]), .B(dpath_mulcore_pc[86]), .Y(n16402));
XOR2X1 mul_dpath_mulcore_array2_sc1_55__U1(.A(dpath_mulcore_a1s[39]), .B(n16402), .Y(dpath_mulcore_array2_s1[55]));
XOR2X1 mul_dpath_mulcore_array2_sc1_56__U4(.A(dpath_mulcore_ps[88]), .B(dpath_mulcore_pc[87]), .Y(n16399));
XOR2X1 mul_dpath_mulcore_array2_sc1_56__U1(.A(dpath_mulcore_a1s[40]), .B(n16399), .Y(dpath_mulcore_array2_s1[56]));
XOR2X1 mul_dpath_mulcore_array2_sc1_57__U4(.A(dpath_mulcore_ps[89]), .B(dpath_mulcore_pc[88]), .Y(n16396));
XOR2X1 mul_dpath_mulcore_array2_sc1_57__U1(.A(dpath_mulcore_a1s[41]), .B(n16396), .Y(dpath_mulcore_array2_s1[57]));
XOR2X1 mul_dpath_mulcore_array2_sc1_58__U4(.A(dpath_mulcore_ps[90]), .B(dpath_mulcore_pc[89]), .Y(n16393));
XOR2X1 mul_dpath_mulcore_array2_sc1_58__U1(.A(dpath_mulcore_a1s[42]), .B(n16393), .Y(dpath_mulcore_array2_s1[58]));
XOR2X1 mul_dpath_mulcore_array2_sc1_59__U4(.A(dpath_mulcore_ps[91]), .B(dpath_mulcore_pc[90]), .Y(n16390));
XOR2X1 mul_dpath_mulcore_array2_sc1_59__U1(.A(dpath_mulcore_a1s[43]), .B(n16390), .Y(dpath_mulcore_array2_s1[59]));
XOR2X1 mul_dpath_mulcore_array2_sc1_60__U4(.A(dpath_mulcore_ps[92]), .B(dpath_mulcore_pc[91]), .Y(n16387));
XOR2X1 mul_dpath_mulcore_array2_sc1_60__U1(.A(dpath_mulcore_a1s[44]), .B(n16387), .Y(dpath_mulcore_array2_s1[60]));
XOR2X1 mul_dpath_mulcore_array2_sc1_61__U4(.A(dpath_mulcore_ps[93]), .B(dpath_mulcore_pc[92]), .Y(n16384));
XOR2X1 mul_dpath_mulcore_array2_sc1_61__U1(.A(dpath_mulcore_a1s[45]), .B(n16384), .Y(dpath_mulcore_array2_s1[61]));
XOR2X1 mul_dpath_mulcore_array2_sc1_62__U4(.A(dpath_mulcore_ps[94]), .B(dpath_mulcore_pc[93]), .Y(n16381));
XOR2X1 mul_dpath_mulcore_array2_sc1_62__U1(.A(dpath_mulcore_a1s[46]), .B(n16381), .Y(dpath_mulcore_array2_s1[62]));
XOR2X1 mul_dpath_mulcore_array2_sc1_63__U4(.A(dpath_mulcore_ps[95]), .B(dpath_mulcore_pc[94]), .Y(n16378));
XOR2X1 mul_dpath_mulcore_array2_sc1_63__U1(.A(dpath_mulcore_a1s[47]), .B(n16378), .Y(dpath_mulcore_array2_s1[63]));
XOR2X1 mul_dpath_mulcore_array2_sc1_64__U4(.A(dpath_mulcore_ps[96]), .B(dpath_mulcore_pc[95]), .Y(n16375));
XOR2X1 mul_dpath_mulcore_array2_sc1_64__U1(.A(dpath_mulcore_a1s[48]), .B(n16375), .Y(dpath_mulcore_array2_s1[64]));
XOR2X1 mul_dpath_mulcore_array2_sc1_65__U4(.A(dpath_mulcore_ps[97]), .B(dpath_mulcore_pc[96]), .Y(n16372));
XOR2X1 mul_dpath_mulcore_array2_sc1_65__U1(.A(dpath_mulcore_a1s[49]), .B(n16372), .Y(dpath_mulcore_array2_s1[65]));
XOR2X1 mul_dpath_mulcore_array2_sc1_66__U4(.A(dpath_mulcore_ps[98]), .B(dpath_mulcore_pc[97]), .Y(n16369));
XOR2X1 mul_dpath_mulcore_array2_sc1_66__U1(.A(dpath_mulcore_a1s[50]), .B(n16369), .Y(dpath_mulcore_array2_s1[66]));
XOR2X1 mul_dpath_mulcore_array2_sc2_20__U1(.A(dpath_mulcore_a0c[19]), .B(dpath_mulcore_a0s[20]), .Y(dpath_mulcore_array2_s2[20]));
XOR2X1 mul_dpath_mulcore_array2_sc2_21__U4(.A(dpath_mulcore_a1c[4]), .B(dpath_mulcore_a0s[21]), .Y(n16365));
XOR2X1 mul_dpath_mulcore_array2_sc2_21__U1(.A(dpath_mulcore_a0c[20]), .B(n16365), .Y(dpath_mulcore_array2_s2[21]));
XOR2X1 mul_dpath_mulcore_array2_sc2_22__U4(.A(dpath_mulcore_a1c[5]), .B(dpath_mulcore_a0s[22]), .Y(n16362));
XOR2X1 mul_dpath_mulcore_array2_sc2_22__U1(.A(dpath_mulcore_a0c[21]), .B(n16362), .Y(dpath_mulcore_array2_s2[22]));
XOR2X1 mul_dpath_mulcore_array2_sc2_23__U4(.A(dpath_mulcore_a1c[6]), .B(dpath_mulcore_a0s[23]), .Y(n16359));
XOR2X1 mul_dpath_mulcore_array2_sc2_23__U1(.A(dpath_mulcore_a0c[22]), .B(n16359), .Y(dpath_mulcore_array2_s2[23]));
XOR2X1 mul_dpath_mulcore_array2_sc2_24__U4(.A(dpath_mulcore_a1c[7]), .B(dpath_mulcore_a0s[24]), .Y(n16356));
XOR2X1 mul_dpath_mulcore_array2_sc2_24__U1(.A(dpath_mulcore_a0c[23]), .B(n16356), .Y(dpath_mulcore_array2_s2[24]));
XOR2X1 mul_dpath_mulcore_array2_sc2_25__U4(.A(dpath_mulcore_a1c[8]), .B(dpath_mulcore_a0s[25]), .Y(n16353));
XOR2X1 mul_dpath_mulcore_array2_sc2_25__U1(.A(dpath_mulcore_a0c[24]), .B(n16353), .Y(dpath_mulcore_array2_s2[25]));
XOR2X1 mul_dpath_mulcore_array2_sc2_26__U4(.A(dpath_mulcore_a1c[9]), .B(dpath_mulcore_a0s[26]), .Y(n16350));
XOR2X1 mul_dpath_mulcore_array2_sc2_26__U1(.A(dpath_mulcore_a0c[25]), .B(n16350), .Y(dpath_mulcore_array2_s2[26]));
XOR2X1 mul_dpath_mulcore_array2_sc2_27__U4(.A(dpath_mulcore_a1c[10]), .B(dpath_mulcore_a0s[27]), .Y(n16347));
XOR2X1 mul_dpath_mulcore_array2_sc2_27__U1(.A(dpath_mulcore_a0c[26]), .B(n16347), .Y(dpath_mulcore_array2_s2[27]));
XOR2X1 mul_dpath_mulcore_array2_sc2_28__U4(.A(dpath_mulcore_a1c[11]), .B(dpath_mulcore_a0s[28]), .Y(n16344));
XOR2X1 mul_dpath_mulcore_array2_sc2_28__U1(.A(dpath_mulcore_a0c[27]), .B(n16344), .Y(dpath_mulcore_array2_s2[28]));
XOR2X1 mul_dpath_mulcore_array2_sc2_29__U4(.A(dpath_mulcore_a1c[12]), .B(dpath_mulcore_a0s[29]), .Y(n16341));
XOR2X1 mul_dpath_mulcore_array2_sc2_29__U1(.A(dpath_mulcore_a0c[28]), .B(n16341), .Y(dpath_mulcore_array2_s2[29]));
XOR2X1 mul_dpath_mulcore_array2_sc2_30__U4(.A(dpath_mulcore_a1c[13]), .B(dpath_mulcore_a0s[30]), .Y(n16338));
XOR2X1 mul_dpath_mulcore_array2_sc2_30__U1(.A(dpath_mulcore_a0c[29]), .B(n16338), .Y(dpath_mulcore_array2_s2[30]));
XOR2X1 mul_dpath_mulcore_array2_sc2_31__U4(.A(dpath_mulcore_a1c[14]), .B(dpath_mulcore_a0s[31]), .Y(n16335));
XOR2X1 mul_dpath_mulcore_array2_sc2_31__U1(.A(dpath_mulcore_a0c[30]), .B(n16335), .Y(dpath_mulcore_array2_s2[31]));
XOR2X1 mul_dpath_mulcore_array2_sc2_32__U4(.A(dpath_mulcore_a1c[15]), .B(dpath_mulcore_a0s[32]), .Y(n16332));
XOR2X1 mul_dpath_mulcore_array2_sc2_32__U1(.A(dpath_mulcore_a0c[31]), .B(n16332), .Y(dpath_mulcore_array2_s2[32]));
XOR2X1 mul_dpath_mulcore_array2_sc2_33__U4(.A(dpath_mulcore_a1c[16]), .B(dpath_mulcore_a0s[33]), .Y(n16329));
XOR2X1 mul_dpath_mulcore_array2_sc2_33__U1(.A(dpath_mulcore_a0c[32]), .B(n16329), .Y(dpath_mulcore_array2_s2[33]));
XOR2X1 mul_dpath_mulcore_array2_sc2_34__U4(.A(dpath_mulcore_a1c[17]), .B(dpath_mulcore_a0s[34]), .Y(n16326));
XOR2X1 mul_dpath_mulcore_array2_sc2_34__U1(.A(dpath_mulcore_a0c[33]), .B(n16326), .Y(dpath_mulcore_array2_s2[34]));
XOR2X1 mul_dpath_mulcore_array2_sc2_35__U4(.A(dpath_mulcore_a1c[18]), .B(dpath_mulcore_a0s[35]), .Y(n16323));
XOR2X1 mul_dpath_mulcore_array2_sc2_35__U1(.A(dpath_mulcore_a0c[34]), .B(n16323), .Y(dpath_mulcore_array2_s2[35]));
XOR2X1 mul_dpath_mulcore_array2_sc2_36__U4(.A(dpath_mulcore_a1c[19]), .B(dpath_mulcore_a0s[36]), .Y(n16320));
XOR2X1 mul_dpath_mulcore_array2_sc2_36__U1(.A(dpath_mulcore_a0c[35]), .B(n16320), .Y(dpath_mulcore_array2_s2[36]));
XOR2X1 mul_dpath_mulcore_array2_sc2_37__U4(.A(dpath_mulcore_a1c[20]), .B(dpath_mulcore_a0s[37]), .Y(n16317));
XOR2X1 mul_dpath_mulcore_array2_sc2_37__U1(.A(dpath_mulcore_a0c[36]), .B(n16317), .Y(dpath_mulcore_array2_s2[37]));
XOR2X1 mul_dpath_mulcore_array2_sc2_38__U4(.A(dpath_mulcore_a1c[21]), .B(dpath_mulcore_a0s[38]), .Y(n16314));
XOR2X1 mul_dpath_mulcore_array2_sc2_38__U1(.A(dpath_mulcore_a0c[37]), .B(n16314), .Y(dpath_mulcore_array2_s2[38]));
XOR2X1 mul_dpath_mulcore_array2_sc2_39__U4(.A(dpath_mulcore_a1c[22]), .B(dpath_mulcore_a0s[39]), .Y(n16311));
XOR2X1 mul_dpath_mulcore_array2_sc2_39__U1(.A(dpath_mulcore_a0c[38]), .B(n16311), .Y(dpath_mulcore_array2_s2[39]));
XOR2X1 mul_dpath_mulcore_array2_sc2_40__U4(.A(dpath_mulcore_a1c[23]), .B(dpath_mulcore_a0s[40]), .Y(n16308));
XOR2X1 mul_dpath_mulcore_array2_sc2_40__U1(.A(dpath_mulcore_a0c[39]), .B(n16308), .Y(dpath_mulcore_array2_s2[40]));
XOR2X1 mul_dpath_mulcore_array2_sc2_41__U4(.A(dpath_mulcore_a1c[24]), .B(dpath_mulcore_a0s[41]), .Y(n16305));
XOR2X1 mul_dpath_mulcore_array2_sc2_41__U1(.A(dpath_mulcore_a0c[40]), .B(n16305), .Y(dpath_mulcore_array2_s2[41]));
XOR2X1 mul_dpath_mulcore_array2_sc2_42__U4(.A(dpath_mulcore_a1c[25]), .B(dpath_mulcore_a0s[42]), .Y(n16302));
XOR2X1 mul_dpath_mulcore_array2_sc2_42__U1(.A(dpath_mulcore_a0c[41]), .B(n16302), .Y(dpath_mulcore_array2_s2[42]));
XOR2X1 mul_dpath_mulcore_array2_sc2_43__U4(.A(dpath_mulcore_a1c[26]), .B(dpath_mulcore_a0s[43]), .Y(n16299));
XOR2X1 mul_dpath_mulcore_array2_sc2_43__U1(.A(dpath_mulcore_a0c[42]), .B(n16299), .Y(dpath_mulcore_array2_s2[43]));
XOR2X1 mul_dpath_mulcore_array2_sc2_44__U4(.A(dpath_mulcore_a1c[27]), .B(dpath_mulcore_a0s[44]), .Y(n16296));
XOR2X1 mul_dpath_mulcore_array2_sc2_44__U1(.A(dpath_mulcore_a0c[43]), .B(n16296), .Y(dpath_mulcore_array2_s2[44]));
XOR2X1 mul_dpath_mulcore_array2_sc2_45__U4(.A(dpath_mulcore_a1c[28]), .B(dpath_mulcore_a0s[45]), .Y(n16293));
XOR2X1 mul_dpath_mulcore_array2_sc2_45__U1(.A(dpath_mulcore_a0c[44]), .B(n16293), .Y(dpath_mulcore_array2_s2[45]));
XOR2X1 mul_dpath_mulcore_array2_sc2_46__U4(.A(dpath_mulcore_a1c[29]), .B(dpath_mulcore_a0s[46]), .Y(n16290));
XOR2X1 mul_dpath_mulcore_array2_sc2_46__U1(.A(dpath_mulcore_a0c[45]), .B(n16290), .Y(dpath_mulcore_array2_s2[46]));
XOR2X1 mul_dpath_mulcore_array2_sc2_47__U4(.A(dpath_mulcore_a1c[30]), .B(dpath_mulcore_a0s[47]), .Y(n16287));
XOR2X1 mul_dpath_mulcore_array2_sc2_47__U1(.A(dpath_mulcore_a0c[46]), .B(n16287), .Y(dpath_mulcore_array2_s2[47]));
XOR2X1 mul_dpath_mulcore_array2_sc2_48__U4(.A(dpath_mulcore_a1c[31]), .B(dpath_mulcore_a0s[48]), .Y(n16284));
XOR2X1 mul_dpath_mulcore_array2_sc2_48__U1(.A(dpath_mulcore_a0c[47]), .B(n16284), .Y(dpath_mulcore_array2_s2[48]));
XOR2X1 mul_dpath_mulcore_array2_sc2_49__U4(.A(dpath_mulcore_a1c[32]), .B(dpath_mulcore_a0s[49]), .Y(n16281));
XOR2X1 mul_dpath_mulcore_array2_sc2_49__U1(.A(dpath_mulcore_a0c[48]), .B(n16281), .Y(dpath_mulcore_array2_s2[49]));
XOR2X1 mul_dpath_mulcore_array2_sc2_50__U4(.A(dpath_mulcore_a1c[33]), .B(dpath_mulcore_a0s[50]), .Y(n16278));
XOR2X1 mul_dpath_mulcore_array2_sc2_50__U1(.A(dpath_mulcore_a0c[49]), .B(n16278), .Y(dpath_mulcore_array2_s2[50]));
XOR2X1 mul_dpath_mulcore_array2_sc2_51__U4(.A(dpath_mulcore_a1c[34]), .B(dpath_mulcore_a0s[51]), .Y(n16275));
XOR2X1 mul_dpath_mulcore_array2_sc2_51__U1(.A(dpath_mulcore_a0c[50]), .B(n16275), .Y(dpath_mulcore_array2_s2[51]));
XOR2X1 mul_dpath_mulcore_array2_sc2_52__U4(.A(dpath_mulcore_a1c[35]), .B(dpath_mulcore_a0s[52]), .Y(n16272));
XOR2X1 mul_dpath_mulcore_array2_sc2_52__U1(.A(dpath_mulcore_a0c[51]), .B(n16272), .Y(dpath_mulcore_array2_s2[52]));
XOR2X1 mul_dpath_mulcore_array2_sc2_53__U4(.A(dpath_mulcore_a1c[36]), .B(dpath_mulcore_a0s[53]), .Y(n16269));
XOR2X1 mul_dpath_mulcore_array2_sc2_53__U1(.A(dpath_mulcore_a0c[52]), .B(n16269), .Y(dpath_mulcore_array2_s2[53]));
XOR2X1 mul_dpath_mulcore_array2_sc2_54__U4(.A(dpath_mulcore_a1c[37]), .B(dpath_mulcore_a0s[54]), .Y(n16266));
XOR2X1 mul_dpath_mulcore_array2_sc2_54__U1(.A(dpath_mulcore_a0c[53]), .B(n16266), .Y(dpath_mulcore_array2_s2[54]));
XOR2X1 mul_dpath_mulcore_array2_sc2_55__U4(.A(dpath_mulcore_a1c[38]), .B(dpath_mulcore_a0s[55]), .Y(n16263));
XOR2X1 mul_dpath_mulcore_array2_sc2_55__U1(.A(dpath_mulcore_a0c[54]), .B(n16263), .Y(dpath_mulcore_array2_s2[55]));
XOR2X1 mul_dpath_mulcore_array2_sc2_56__U4(.A(dpath_mulcore_a1c[39]), .B(dpath_mulcore_a0s[56]), .Y(n16260));
XOR2X1 mul_dpath_mulcore_array2_sc2_56__U1(.A(dpath_mulcore_a0c[55]), .B(n16260), .Y(dpath_mulcore_array2_s2[56]));
XOR2X1 mul_dpath_mulcore_array2_sc2_57__U4(.A(dpath_mulcore_a1c[40]), .B(dpath_mulcore_a0s[57]), .Y(n16257));
XOR2X1 mul_dpath_mulcore_array2_sc2_57__U1(.A(dpath_mulcore_a0c[56]), .B(n16257), .Y(dpath_mulcore_array2_s2[57]));
XOR2X1 mul_dpath_mulcore_array2_sc2_58__U4(.A(dpath_mulcore_a1c[41]), .B(dpath_mulcore_a0s[58]), .Y(n16254));
XOR2X1 mul_dpath_mulcore_array2_sc2_58__U1(.A(dpath_mulcore_a0c[57]), .B(n16254), .Y(dpath_mulcore_array2_s2[58]));
XOR2X1 mul_dpath_mulcore_array2_sc2_59__U4(.A(dpath_mulcore_a1c[42]), .B(dpath_mulcore_a0s[59]), .Y(n16251));
XOR2X1 mul_dpath_mulcore_array2_sc2_59__U1(.A(dpath_mulcore_a0c[58]), .B(n16251), .Y(dpath_mulcore_array2_s2[59]));
XOR2X1 mul_dpath_mulcore_array2_sc2_60__U4(.A(dpath_mulcore_a1c[43]), .B(dpath_mulcore_a0s[60]), .Y(n16248));
XOR2X1 mul_dpath_mulcore_array2_sc2_60__U1(.A(dpath_mulcore_a0c[59]), .B(n16248), .Y(dpath_mulcore_array2_s2[60]));
XOR2X1 mul_dpath_mulcore_array2_sc2_61__U4(.A(dpath_mulcore_a1c[44]), .B(dpath_mulcore_a0s[61]), .Y(n16245));
XOR2X1 mul_dpath_mulcore_array2_sc2_61__U1(.A(dpath_mulcore_a0c[60]), .B(n16245), .Y(dpath_mulcore_array2_s2[61]));
XOR2X1 mul_dpath_mulcore_array2_sc2_62__U4(.A(dpath_mulcore_a1c[45]), .B(dpath_mulcore_a0s[62]), .Y(n16242));
XOR2X1 mul_dpath_mulcore_array2_sc2_62__U1(.A(dpath_mulcore_a0c[61]), .B(n16242), .Y(dpath_mulcore_array2_s2[62]));
XOR2X1 mul_dpath_mulcore_array2_sc2_63__U4(.A(dpath_mulcore_a1c[46]), .B(dpath_mulcore_a0s[63]), .Y(n16239));
XOR2X1 mul_dpath_mulcore_array2_sc2_63__U1(.A(dpath_mulcore_a0c[62]), .B(n16239), .Y(dpath_mulcore_array2_s2[63]));
XOR2X1 mul_dpath_mulcore_array2_sc2_64__U4(.A(dpath_mulcore_a1c[47]), .B(dpath_mulcore_a0s[64]), .Y(n16236));
XOR2X1 mul_dpath_mulcore_array2_sc2_64__U1(.A(dpath_mulcore_a0c[63]), .B(n16236), .Y(dpath_mulcore_array2_s2[64]));
XOR2X1 mul_dpath_mulcore_array2_sc2_65__U4(.A(dpath_mulcore_a1c[48]), .B(dpath_mulcore_a0s[65]), .Y(n16233));
XOR2X1 mul_dpath_mulcore_array2_sc2_65__U1(.A(dpath_mulcore_a0c[64]), .B(n16233), .Y(dpath_mulcore_array2_s2[65]));
XOR2X1 mul_dpath_mulcore_array2_sc2_66__U4(.A(dpath_mulcore_a1c[49]), .B(dpath_mulcore_a0s[66]), .Y(n16230));
XOR2X1 mul_dpath_mulcore_array2_sc2_66__U1(.A(dpath_mulcore_a0c[65]), .B(n16230), .Y(dpath_mulcore_array2_s2[66]));
XOR2X1 mul_dpath_mulcore_array2_sc1_1__U4(.A(dpath_mulcore_ps[33]), .B(dpath_mulcore_pc[32]), .Y(n16227));
XOR2X1 mul_dpath_mulcore_array2_sc1_1__U1(.A(dpath_mulcore_a0s[1]), .B(n16227), .Y(dpath_mulcore_array2_s1[1]));
XOR2X1 mul_dpath_mulcore_array2_sc1_2__U4(.A(dpath_mulcore_ps[34]), .B(dpath_mulcore_pc[33]), .Y(n16224));
XOR2X1 mul_dpath_mulcore_array2_sc1_2__U1(.A(dpath_mulcore_a0s[2]), .B(n16224), .Y(dpath_mulcore_array2_s1[2]));
XOR2X1 mul_dpath_mulcore_array2_sc1_3__U4(.A(dpath_mulcore_ps[35]), .B(dpath_mulcore_pc[34]), .Y(n16221));
XOR2X1 mul_dpath_mulcore_array2_sc1_3__U1(.A(dpath_mulcore_a0s[3]), .B(n16221), .Y(dpath_mulcore_array2_s1[3]));
XOR2X1 mul_dpath_mulcore_array2_sc1_4__U4(.A(dpath_mulcore_ps[36]), .B(dpath_mulcore_pc[35]), .Y(n16218));
XOR2X1 mul_dpath_mulcore_array2_sc1_4__U1(.A(dpath_mulcore_a0s[4]), .B(n16218), .Y(dpath_mulcore_array2_s1[4]));
XOR2X1 mul_dpath_mulcore_array2_sc2_82__U4(.A(dpath_mulcore_array2_s1[82]), .B(n8948), .Y(n16215));
XOR2X1 mul_dpath_mulcore_array2_sc2_82__U1(.A(n8325), .B(n16215), .Y(dpath_mulcore_array2_s2[82]));
XOR2X1 mul_dpath_mulcore_array2_sc2_5__U4(.A(dpath_mulcore_array2_s1[5]), .B(n8972), .Y(n16212));
XOR2X1 mul_dpath_mulcore_array2_sc2_5__U1(.A(dpath_mulcore_a0c[4]), .B(n16212), .Y(dpath_mulcore_array2_s2[5]));
XOR2X1 mul_dpath_mulcore_array2_sc2_6__U4(.A(dpath_mulcore_array2_s1[6]), .B(n8971), .Y(n16209));
XOR2X1 mul_dpath_mulcore_array2_sc2_6__U1(.A(dpath_mulcore_a0c[5]), .B(n16209), .Y(dpath_mulcore_array2_s2[6]));
XOR2X1 mul_dpath_mulcore_array2_sc2_7__U4(.A(dpath_mulcore_array2_s1[7]), .B(n8970), .Y(n16206));
XOR2X1 mul_dpath_mulcore_array2_sc2_7__U1(.A(dpath_mulcore_a0c[6]), .B(n16206), .Y(dpath_mulcore_array2_s2[7]));
XOR2X1 mul_dpath_mulcore_array2_sc2_8__U4(.A(dpath_mulcore_array2_s1[8]), .B(n8969), .Y(n16203));
XOR2X1 mul_dpath_mulcore_array2_sc2_8__U1(.A(dpath_mulcore_a0c[7]), .B(n16203), .Y(dpath_mulcore_array2_s2[8]));
XOR2X1 mul_dpath_mulcore_array2_sc2_9__U4(.A(dpath_mulcore_array2_s1[9]), .B(n8968), .Y(n16200));
XOR2X1 mul_dpath_mulcore_array2_sc2_9__U1(.A(dpath_mulcore_a0c[8]), .B(n16200), .Y(dpath_mulcore_array2_s2[9]));
XOR2X1 mul_dpath_mulcore_array2_sc2_10__U4(.A(dpath_mulcore_array2_s1[10]), .B(n8967), .Y(n16197));
XOR2X1 mul_dpath_mulcore_array2_sc2_10__U1(.A(dpath_mulcore_a0c[9]), .B(n16197), .Y(dpath_mulcore_array2_s2[10]));
XOR2X1 mul_dpath_mulcore_array2_sc2_11__U4(.A(dpath_mulcore_array2_s1[11]), .B(n8966), .Y(n16194));
XOR2X1 mul_dpath_mulcore_array2_sc2_11__U1(.A(dpath_mulcore_a0c[10]), .B(n16194), .Y(dpath_mulcore_array2_s2[11]));
XOR2X1 mul_dpath_mulcore_array2_sc2_12__U4(.A(dpath_mulcore_array2_s1[12]), .B(n8965), .Y(n16191));
XOR2X1 mul_dpath_mulcore_array2_sc2_12__U1(.A(dpath_mulcore_a0c[11]), .B(n16191), .Y(dpath_mulcore_array2_s2[12]));
XOR2X1 mul_dpath_mulcore_array2_sc2_13__U4(.A(dpath_mulcore_array2_s1[13]), .B(n8964), .Y(n16188));
XOR2X1 mul_dpath_mulcore_array2_sc2_13__U1(.A(dpath_mulcore_a0c[12]), .B(n16188), .Y(dpath_mulcore_array2_s2[13]));
XOR2X1 mul_dpath_mulcore_array2_sc2_14__U4(.A(dpath_mulcore_array2_s1[14]), .B(n8963), .Y(n16185));
XOR2X1 mul_dpath_mulcore_array2_sc2_14__U1(.A(dpath_mulcore_a0c[13]), .B(n16185), .Y(dpath_mulcore_array2_s2[14]));
XOR2X1 mul_dpath_mulcore_array2_sc1_5__U4(.A(dpath_mulcore_ps[37]), .B(dpath_mulcore_pc[36]), .Y(n16182));
XOR2X1 mul_dpath_mulcore_array2_sc1_5__U1(.A(dpath_mulcore_a0s[5]), .B(n16182), .Y(dpath_mulcore_array2_s1[5]));
XOR2X1 mul_dpath_mulcore_array2_sc1_6__U4(.A(dpath_mulcore_ps[38]), .B(dpath_mulcore_pc[37]), .Y(n16179));
XOR2X1 mul_dpath_mulcore_array2_sc1_6__U1(.A(dpath_mulcore_a0s[6]), .B(n16179), .Y(dpath_mulcore_array2_s1[6]));
XOR2X1 mul_dpath_mulcore_array2_sc1_7__U4(.A(dpath_mulcore_ps[39]), .B(dpath_mulcore_pc[38]), .Y(n16176));
XOR2X1 mul_dpath_mulcore_array2_sc1_7__U1(.A(dpath_mulcore_a0s[7]), .B(n16176), .Y(dpath_mulcore_array2_s1[7]));
XOR2X1 mul_dpath_mulcore_array2_sc1_8__U4(.A(dpath_mulcore_ps[40]), .B(dpath_mulcore_pc[39]), .Y(n16173));
XOR2X1 mul_dpath_mulcore_array2_sc1_8__U1(.A(dpath_mulcore_a0s[8]), .B(n16173), .Y(dpath_mulcore_array2_s1[8]));
XOR2X1 mul_dpath_mulcore_array2_sc1_9__U4(.A(dpath_mulcore_ps[41]), .B(dpath_mulcore_pc[40]), .Y(n16170));
XOR2X1 mul_dpath_mulcore_array2_sc1_9__U1(.A(dpath_mulcore_a0s[9]), .B(n16170), .Y(dpath_mulcore_array2_s1[9]));
XOR2X1 mul_dpath_mulcore_array2_sc1_10__U4(.A(dpath_mulcore_ps[42]), .B(dpath_mulcore_pc[41]), .Y(n16167));
XOR2X1 mul_dpath_mulcore_array2_sc1_10__U1(.A(dpath_mulcore_a0s[10]), .B(n16167), .Y(dpath_mulcore_array2_s1[10]));
XOR2X1 mul_dpath_mulcore_array2_sc1_11__U4(.A(dpath_mulcore_ps[43]), .B(dpath_mulcore_pc[42]), .Y(n16164));
XOR2X1 mul_dpath_mulcore_array2_sc1_11__U1(.A(dpath_mulcore_a0s[11]), .B(n16164), .Y(dpath_mulcore_array2_s1[11]));
XOR2X1 mul_dpath_mulcore_array2_sc1_12__U4(.A(dpath_mulcore_ps[44]), .B(dpath_mulcore_pc[43]), .Y(n16161));
XOR2X1 mul_dpath_mulcore_array2_sc1_12__U1(.A(dpath_mulcore_a0s[12]), .B(n16161), .Y(dpath_mulcore_array2_s1[12]));
XOR2X1 mul_dpath_mulcore_array2_sc1_13__U4(.A(dpath_mulcore_ps[45]), .B(dpath_mulcore_pc[44]), .Y(n16158));
XOR2X1 mul_dpath_mulcore_array2_sc1_13__U1(.A(dpath_mulcore_a0s[13]), .B(n16158), .Y(dpath_mulcore_array2_s1[13]));
XOR2X1 mul_dpath_mulcore_array2_sc1_14__U4(.A(dpath_mulcore_ps[46]), .B(dpath_mulcore_pc[45]), .Y(n16155));
XOR2X1 mul_dpath_mulcore_array2_sc1_14__U1(.A(dpath_mulcore_a0s[14]), .B(n16155), .Y(dpath_mulcore_array2_s1[14]));
XOR2X1 mul_dpath_mulcore_array2_sc2_67__U4(.A(dpath_mulcore_a0s[67]), .B(n8973), .Y(n16152));
XOR2X1 mul_dpath_mulcore_array2_sc2_67__U1(.A(dpath_mulcore_a0c[66]), .B(n16152), .Y(dpath_mulcore_array2_s2[67]));
XOR2X1 mul_dpath_mulcore_array2_acc_5__U4(.A(n8284), .B(dpath_mulcore_array2_s2[5]), .Y(n16149));
XOR2X1 mul_dpath_mulcore_array2_acc_5__U1(.A(dpath_mulcore_array2_c2[4]), .B(n16149), .Y(dpath_mulcore_psum[5]));
XOR2X1 mul_dpath_mulcore_array2_acc_6__U4(.A(n8283), .B(dpath_mulcore_array2_s2[6]), .Y(n16146));
XOR2X1 mul_dpath_mulcore_array2_acc_6__U1(.A(n8323), .B(n16146), .Y(dpath_mulcore_psum[6]));
XOR2X1 mul_dpath_mulcore_array2_acc_7__U4(.A(n8282), .B(dpath_mulcore_array2_s2[7]), .Y(n16143));
XOR2X1 mul_dpath_mulcore_array2_acc_7__U1(.A(n8322), .B(n16143), .Y(dpath_mulcore_psum[7]));
XOR2X1 mul_dpath_mulcore_array2_acc_8__U4(.A(n8281), .B(dpath_mulcore_array2_s2[8]), .Y(n16140));
XOR2X1 mul_dpath_mulcore_array2_acc_8__U1(.A(n8321), .B(n16140), .Y(dpath_mulcore_psum[8]));
XOR2X1 mul_dpath_mulcore_array2_acc_9__U4(.A(n8280), .B(dpath_mulcore_array2_s2[9]), .Y(n16137));
XOR2X1 mul_dpath_mulcore_array2_acc_9__U1(.A(n8320), .B(n16137), .Y(dpath_mulcore_psum[9]));
XOR2X1 mul_dpath_mulcore_array2_acc_10__U4(.A(n8279), .B(dpath_mulcore_array2_s2[10]), .Y(n16134));
XOR2X1 mul_dpath_mulcore_array2_acc_10__U1(.A(n8319), .B(n16134), .Y(dpath_mulcore_psum[10]));
XOR2X1 mul_dpath_mulcore_array2_acc_11__U4(.A(n8278), .B(dpath_mulcore_array2_s2[11]), .Y(n16131));
XOR2X1 mul_dpath_mulcore_array2_acc_11__U1(.A(n8318), .B(n16131), .Y(dpath_mulcore_psum[11]));
XOR2X1 mul_dpath_mulcore_array2_acc_12__U4(.A(n8277), .B(dpath_mulcore_array2_s2[12]), .Y(n16128));
XOR2X1 mul_dpath_mulcore_array2_acc_12__U1(.A(n8317), .B(n16128), .Y(dpath_mulcore_psum[12]));
XOR2X1 mul_dpath_mulcore_array2_acc_13__U4(.A(n8276), .B(dpath_mulcore_array2_s2[13]), .Y(n16125));
XOR2X1 mul_dpath_mulcore_array2_acc_13__U1(.A(n8316), .B(n16125), .Y(dpath_mulcore_psum[13]));
XOR2X1 mul_dpath_mulcore_array2_acc_14__U4(.A(n8275), .B(dpath_mulcore_array2_s2[14]), .Y(n16122));
XOR2X1 mul_dpath_mulcore_array2_acc_14__U1(.A(n8315), .B(n16122), .Y(dpath_mulcore_psum[14]));
XOR2X1 mul_dpath_mulcore_array2_sc1_82__U4(.A(dpath_mulcore_a1s[66]), .B(dpath_mulcore_a1c[65]), .Y(dpath_mulcore_array2_s1[82]));
XOR2X1 mul_dpath_mulcore_array2_sc3_15__U4(.A(dpath_mulcore_array2_s2[15]), .B(n8962), .Y(n16118));
XOR2X1 mul_dpath_mulcore_array2_sc3_15__U1(.A(n8314), .B(n16118), .Y(dpath_mulcore_array2_s3[15]));
XOR2X1 mul_dpath_mulcore_array2_sc3_16__U4(.A(dpath_mulcore_array2_s2[16]), .B(n16044), .Y(n16115));
XOR2X1 mul_dpath_mulcore_array2_sc3_16__U1(.A(n8307), .B(n16115), .Y(dpath_mulcore_array2_s3[16]));
XOR2X1 mul_dpath_mulcore_array2_sc3_17__U4(.A(dpath_mulcore_array2_s2[17]), .B(n8947), .Y(n16112));
XOR2X1 mul_dpath_mulcore_array2_sc3_17__U1(.A(n8306), .B(n16112), .Y(dpath_mulcore_array2_s3[17]));
XOR2X1 mul_dpath_mulcore_array2_sc3_18__U4(.A(dpath_mulcore_array2_s2[18]), .B(n8946), .Y(n16109));
XOR2X1 mul_dpath_mulcore_array2_sc3_18__U1(.A(n8305), .B(n16109), .Y(dpath_mulcore_array2_s3[18]));
XOR2X1 mul_dpath_mulcore_array2_sc3_19__U4(.A(dpath_mulcore_array2_s2[19]), .B(n8945), .Y(n16106));
XOR2X1 mul_dpath_mulcore_array2_sc3_19__U1(.A(n8304), .B(n16106), .Y(dpath_mulcore_array2_s3[19]));
XOR2X1 mul_dpath_mulcore_array2_sc1_68__U4(.A(dpath_mulcore_a1s[52]), .B(dpath_mulcore_a1c[51]), .Y(n16103));
XOR2X1 mul_dpath_mulcore_array2_sc1_68__U1(.A(dpath_mulcore_a0s[68]), .B(n16103), .Y(dpath_mulcore_array2_s1[68]));
XOR2X1 mul_dpath_mulcore_array2_sc1_69__U4(.A(dpath_mulcore_a1s[53]), .B(dpath_mulcore_a1c[52]), .Y(n16100));
XOR2X1 mul_dpath_mulcore_array2_sc1_69__U1(.A(dpath_mulcore_a0s[69]), .B(n16100), .Y(dpath_mulcore_array2_s1[69]));
XOR2X1 mul_dpath_mulcore_array2_sc1_70__U4(.A(dpath_mulcore_a1s[54]), .B(dpath_mulcore_a1c[53]), .Y(n16097));
XOR2X1 mul_dpath_mulcore_array2_sc1_70__U1(.A(dpath_mulcore_a0s[70]), .B(n16097), .Y(dpath_mulcore_array2_s1[70]));
XOR2X1 mul_dpath_mulcore_array2_sc1_71__U4(.A(dpath_mulcore_a1s[55]), .B(dpath_mulcore_a1c[54]), .Y(n16094));
XOR2X1 mul_dpath_mulcore_array2_sc1_71__U1(.A(dpath_mulcore_a0s[71]), .B(n16094), .Y(dpath_mulcore_array2_s1[71]));
XOR2X1 mul_dpath_mulcore_array2_sc1_72__U4(.A(dpath_mulcore_a1s[56]), .B(dpath_mulcore_a1c[55]), .Y(n16091));
XOR2X1 mul_dpath_mulcore_array2_sc1_72__U1(.A(dpath_mulcore_a0s[72]), .B(n16091), .Y(dpath_mulcore_array2_s1[72]));
XOR2X1 mul_dpath_mulcore_array2_sc1_73__U4(.A(dpath_mulcore_a1s[57]), .B(dpath_mulcore_a1c[56]), .Y(n16088));
XOR2X1 mul_dpath_mulcore_array2_sc1_73__U1(.A(dpath_mulcore_a0s[73]), .B(n16088), .Y(dpath_mulcore_array2_s1[73]));
XOR2X1 mul_dpath_mulcore_array2_sc1_74__U4(.A(dpath_mulcore_a1s[58]), .B(dpath_mulcore_a1c[57]), .Y(n16085));
XOR2X1 mul_dpath_mulcore_array2_sc1_74__U1(.A(dpath_mulcore_a0s[74]), .B(n16085), .Y(dpath_mulcore_array2_s1[74]));
XOR2X1 mul_dpath_mulcore_array2_sc1_75__U4(.A(dpath_mulcore_a1s[59]), .B(dpath_mulcore_a1c[58]), .Y(n16082));
XOR2X1 mul_dpath_mulcore_array2_sc1_75__U1(.A(dpath_mulcore_a0s[75]), .B(n16082), .Y(dpath_mulcore_array2_s1[75]));
XOR2X1 mul_dpath_mulcore_array2_sc1_76__U4(.A(dpath_mulcore_a1s[60]), .B(dpath_mulcore_a1c[59]), .Y(n16079));
XOR2X1 mul_dpath_mulcore_array2_sc1_76__U1(.A(dpath_mulcore_a0s[76]), .B(n16079), .Y(dpath_mulcore_array2_s1[76]));
XOR2X1 mul_dpath_mulcore_array2_sc1_77__U4(.A(dpath_mulcore_a1s[61]), .B(dpath_mulcore_a1c[60]), .Y(n16076));
XOR2X1 mul_dpath_mulcore_array2_sc1_77__U1(.A(dpath_mulcore_a0s[77]), .B(n16076), .Y(dpath_mulcore_array2_s1[77]));
XOR2X1 mul_dpath_mulcore_array2_sc1_78__U4(.A(dpath_mulcore_a1s[62]), .B(dpath_mulcore_a1c[61]), .Y(n16073));
XOR2X1 mul_dpath_mulcore_array2_sc1_78__U1(.A(dpath_mulcore_a0s[78]), .B(n16073), .Y(dpath_mulcore_array2_s1[78]));
XOR2X1 mul_dpath_mulcore_array2_sc1_79__U4(.A(dpath_mulcore_a1s[63]), .B(dpath_mulcore_a1c[62]), .Y(n16070));
XOR2X1 mul_dpath_mulcore_array2_sc1_79__U1(.A(dpath_mulcore_a0s[79]), .B(n16070), .Y(dpath_mulcore_array2_s1[79]));
XOR2X1 mul_dpath_mulcore_array2_sc1_80__U4(.A(dpath_mulcore_a1s[64]), .B(dpath_mulcore_a1c[63]), .Y(n16067));
XOR2X1 mul_dpath_mulcore_array2_sc1_80__U1(.A(dpath_mulcore_a0s[80]), .B(n16067), .Y(dpath_mulcore_array2_s1[80]));
XOR2X1 mul_dpath_mulcore_array2_sc1_81__U4(.A(dpath_mulcore_a1s[65]), .B(dpath_mulcore_a1c[64]), .Y(dpath_mulcore_array2_s1[81]));
XOR2X1 mul_dpath_mulcore_array2_sc2_15__U4(.A(n16043), .B(dpath_mulcore_a0s[15]), .Y(n16063));
XOR2X1 mul_dpath_mulcore_array2_sc2_15__U1(.A(dpath_mulcore_a0c[14]), .B(n16063), .Y(dpath_mulcore_array2_s2[15]));
XOR2X1 mul_dpath_mulcore_array2_sc2_16__U4(.A(dpath_mulcore_array2_s1[16]), .B(dpath_mulcore_a0s[16]), .Y(n16060));
XOR2X1 mul_dpath_mulcore_array2_sc2_16__U1(.A(dpath_mulcore_a0c[15]), .B(n16060), .Y(dpath_mulcore_array2_s2[16]));
XOR2X1 mul_dpath_mulcore_array2_sc2_17__U4(.A(dpath_mulcore_array2_s1[17]), .B(dpath_mulcore_a0s[17]), .Y(n16057));
XOR2X1 mul_dpath_mulcore_array2_sc2_17__U1(.A(dpath_mulcore_a0c[16]), .B(n16057), .Y(dpath_mulcore_array2_s2[17]));
XOR2X1 mul_dpath_mulcore_array2_sc2_18__U4(.A(dpath_mulcore_array2_s1[18]), .B(dpath_mulcore_a0s[18]), .Y(n16054));
XOR2X1 mul_dpath_mulcore_array2_sc2_18__U1(.A(dpath_mulcore_a0c[17]), .B(n16054), .Y(dpath_mulcore_array2_s2[18]));
XOR2X1 mul_dpath_mulcore_array2_sc2_19__U4(.A(dpath_mulcore_array2_s1[19]), .B(dpath_mulcore_a0s[19]), .Y(n16051));
XOR2X1 mul_dpath_mulcore_array2_sc2_19__U1(.A(dpath_mulcore_a0c[18]), .B(n16051), .Y(dpath_mulcore_array2_s2[19]));
XOR2X1 mul_dpath_mulcore_array2_sc2_83__U4(.A(dpath_mulcore_a1s[67]), .B(dpath_mulcore_a1c[66]), .Y(n16048));
XOR2X1 mul_dpath_mulcore_array2_sc2_83__U1(.A(n8313), .B(n16048), .Y(dpath_mulcore_array2_s2[83]));
XOR2X1 mul_dpath_mulcore_array2_sc4_83__U4(.A(n8274), .B(dpath_mulcore_array2_s2[83]), .Y(n16045));
XOR2X1 mul_dpath_mulcore_array2_sc4_83__U1(.A(n8324), .B(n16045), .Y(dpath_mulcore_psum[83]));
XOR2X1 mul_dpath_mulcore_array2_sc1_15__U4(.A(dpath_mulcore_ps[47]), .B(dpath_mulcore_pc[46]), .Y(n16043));
XOR2X1 mul_dpath_mulcore_array2_sc1_16__U4(.A(dpath_mulcore_ps[48]), .B(dpath_mulcore_pc[47]), .Y(n16040));
XOR2X1 mul_dpath_mulcore_array2_sc1_16__U1(.A(dpath_mulcore_a1s[0]), .B(n16040), .Y(dpath_mulcore_array2_s1[16]));
XOR2X1 mul_dpath_mulcore_array2_sc1_17__U4(.A(dpath_mulcore_ps[49]), .B(dpath_mulcore_pc[48]), .Y(n16037));
XOR2X1 mul_dpath_mulcore_array2_sc1_17__U1(.A(dpath_mulcore_a1s[1]), .B(n16037), .Y(dpath_mulcore_array2_s1[17]));
XOR2X1 mul_dpath_mulcore_array2_sc1_18__U4(.A(dpath_mulcore_ps[50]), .B(dpath_mulcore_pc[49]), .Y(n16034));
XOR2X1 mul_dpath_mulcore_array2_sc1_18__U1(.A(dpath_mulcore_a1s[2]), .B(n16034), .Y(dpath_mulcore_array2_s1[18]));
XOR2X1 mul_dpath_mulcore_array2_sc1_19__U4(.A(dpath_mulcore_ps[51]), .B(dpath_mulcore_pc[50]), .Y(n16031));
XOR2X1 mul_dpath_mulcore_array2_sc1_19__U1(.A(dpath_mulcore_a1s[3]), .B(n16031), .Y(dpath_mulcore_array2_s1[19]));
XOR2X1 mul_dpath_mulcore_array2_sc3_97__U4(.A(dpath_mulcore_a1s[81]), .B(dpath_mulcore_a1c[80]), .Y(n16028));
XOR2X1 mul_dpath_mulcore_array2_sc3_97__U1(.A(dpath_mulcore_array2_c2[96]), .B(n16028), .Y(dpath_mulcore_psum[97]));
XOR2X1 mul_dpath_mulcore_array2_acc_1__U4(.A(n8273), .B(dpath_mulcore_array2_s2[1]), .Y(n16025));
XOR2X1 mul_dpath_mulcore_array2_acc_1__U1(.A(dpath_mulcore_array2_c2[0]), .B(n16025), .Y(dpath_mulcore_psum[1]));
XOR2X1 mul_dpath_mulcore_array2_acc_2__U4(.A(n8272), .B(dpath_mulcore_array2_s2[2]), .Y(n16022));
XOR2X1 mul_dpath_mulcore_array2_acc_2__U1(.A(dpath_mulcore_array2_c2[1]), .B(n16022), .Y(dpath_mulcore_psum[2]));
XOR2X1 mul_dpath_mulcore_array2_acc_3__U4(.A(n8271), .B(dpath_mulcore_array2_s2[3]), .Y(n16019));
XOR2X1 mul_dpath_mulcore_array2_acc_3__U1(.A(dpath_mulcore_array2_c2[2]), .B(n16019), .Y(dpath_mulcore_psum[3]));
XOR2X1 mul_dpath_mulcore_array2_acc_4__U4(.A(n8270), .B(dpath_mulcore_array2_s2[4]), .Y(n16016));
XOR2X1 mul_dpath_mulcore_array2_acc_4__U1(.A(dpath_mulcore_array2_c2[3]), .B(n16016), .Y(dpath_mulcore_psum[4]));
XOR2X1 mul_dpath_mulcore_array2_sc4_69__U4(.A(n8264), .B(dpath_mulcore_array2_s3[69]), .Y(n16013));
XOR2X1 mul_dpath_mulcore_array2_sc4_69__U1(.A(n8329), .B(n16013), .Y(dpath_mulcore_psum[69]));
XOR2X1 mul_dpath_mulcore_array2_sc4_70__U4(.A(n8263), .B(dpath_mulcore_array2_s3[70]), .Y(n16010));
XOR2X1 mul_dpath_mulcore_array2_sc4_70__U1(.A(dpath_mulcore_array2_c3[69]), .B(n16010), .Y(dpath_mulcore_psum[70]));
XOR2X1 mul_dpath_mulcore_array2_sc4_71__U4(.A(n8262), .B(dpath_mulcore_array2_s3[71]), .Y(n16007));
XOR2X1 mul_dpath_mulcore_array2_sc4_71__U1(.A(dpath_mulcore_array2_c3[70]), .B(n16007), .Y(dpath_mulcore_psum[71]));
XOR2X1 mul_dpath_mulcore_array2_sc4_72__U4(.A(n8261), .B(dpath_mulcore_array2_s3[72]), .Y(n16004));
XOR2X1 mul_dpath_mulcore_array2_sc4_72__U1(.A(dpath_mulcore_array2_c3[71]), .B(n16004), .Y(dpath_mulcore_psum[72]));
XOR2X1 mul_dpath_mulcore_array2_sc4_73__U4(.A(n8260), .B(dpath_mulcore_array2_s3[73]), .Y(n16001));
XOR2X1 mul_dpath_mulcore_array2_sc4_73__U1(.A(dpath_mulcore_array2_c3[72]), .B(n16001), .Y(dpath_mulcore_psum[73]));
XOR2X1 mul_dpath_mulcore_array2_sc4_74__U4(.A(n8259), .B(dpath_mulcore_array2_s3[74]), .Y(n15998));
XOR2X1 mul_dpath_mulcore_array2_sc4_74__U1(.A(dpath_mulcore_array2_c3[73]), .B(n15998), .Y(dpath_mulcore_psum[74]));
XOR2X1 mul_dpath_mulcore_array2_sc4_75__U4(.A(n8258), .B(dpath_mulcore_array2_s3[75]), .Y(n15995));
XOR2X1 mul_dpath_mulcore_array2_sc4_75__U1(.A(dpath_mulcore_array2_c3[74]), .B(n15995), .Y(dpath_mulcore_psum[75]));
XOR2X1 mul_dpath_mulcore_array2_sc4_76__U4(.A(n8257), .B(dpath_mulcore_array2_s3[76]), .Y(n15992));
XOR2X1 mul_dpath_mulcore_array2_sc4_76__U1(.A(dpath_mulcore_array2_c3[75]), .B(n15992), .Y(dpath_mulcore_psum[76]));
XOR2X1 mul_dpath_mulcore_array2_sc4_77__U4(.A(n8256), .B(dpath_mulcore_array2_s3[77]), .Y(n15989));
XOR2X1 mul_dpath_mulcore_array2_sc4_77__U1(.A(dpath_mulcore_array2_c3[76]), .B(n15989), .Y(dpath_mulcore_psum[77]));
XOR2X1 mul_dpath_mulcore_array2_sc4_78__U4(.A(n8255), .B(dpath_mulcore_array2_s3[78]), .Y(n15986));
XOR2X1 mul_dpath_mulcore_array2_sc4_78__U1(.A(dpath_mulcore_array2_c3[77]), .B(n15986), .Y(dpath_mulcore_psum[78]));
XOR2X1 mul_dpath_mulcore_array2_sc4_79__U4(.A(n8254), .B(dpath_mulcore_array2_s3[79]), .Y(n15983));
XOR2X1 mul_dpath_mulcore_array2_sc4_79__U1(.A(dpath_mulcore_array2_c3[78]), .B(n15983), .Y(dpath_mulcore_psum[79]));
XOR2X1 mul_dpath_mulcore_array2_sc4_80__U4(.A(n8253), .B(dpath_mulcore_array2_s3[80]), .Y(n15980));
XOR2X1 mul_dpath_mulcore_array2_sc4_80__U1(.A(dpath_mulcore_array2_c3[79]), .B(n15980), .Y(dpath_mulcore_psum[80]));
XOR2X1 mul_dpath_mulcore_array2_sc4_81__U4(.A(n8252), .B(dpath_mulcore_array2_s3[81]), .Y(n15977));
XOR2X1 mul_dpath_mulcore_array2_sc4_81__U1(.A(dpath_mulcore_array2_c3[80]), .B(n15977), .Y(dpath_mulcore_psum[81]));
XOR2X1 mul_dpath_mulcore_array2_sc4_84__U4(.A(n8251), .B(dpath_mulcore_array2_s2[84]), .Y(n15974));
XOR2X1 mul_dpath_mulcore_array2_sc4_84__U1(.A(n8303), .B(n15974), .Y(dpath_mulcore_psum[84]));
XOR2X1 mul_dpath_mulcore_array2_sc4_85__U4(.A(n8250), .B(dpath_mulcore_array2_s2[85]), .Y(n15971));
XOR2X1 mul_dpath_mulcore_array2_sc4_85__U1(.A(dpath_mulcore_array2_c2[84]), .B(n15971), .Y(dpath_mulcore_psum[85]));
XOR2X1 mul_dpath_mulcore_array2_sc4_86__U4(.A(n8249), .B(dpath_mulcore_array2_s2[86]), .Y(n15968));
XOR2X1 mul_dpath_mulcore_array2_sc4_86__U1(.A(dpath_mulcore_array2_c2[85]), .B(n15968), .Y(dpath_mulcore_psum[86]));
XOR2X1 mul_dpath_mulcore_array2_sc4_87__U4(.A(n8248), .B(dpath_mulcore_array2_s2[87]), .Y(n15965));
XOR2X1 mul_dpath_mulcore_array2_sc4_87__U1(.A(dpath_mulcore_array2_c2[86]), .B(n15965), .Y(dpath_mulcore_psum[87]));
XOR2X1 mul_dpath_mulcore_array2_sc4_88__U4(.A(n8247), .B(dpath_mulcore_array2_s2[88]), .Y(n15962));
XOR2X1 mul_dpath_mulcore_array2_sc4_88__U1(.A(dpath_mulcore_array2_c2[87]), .B(n15962), .Y(dpath_mulcore_psum[88]));
XOR2X1 mul_dpath_mulcore_array2_sc4_89__U4(.A(n8246), .B(dpath_mulcore_array2_s2[89]), .Y(n15959));
XOR2X1 mul_dpath_mulcore_array2_sc4_89__U1(.A(dpath_mulcore_array2_c2[88]), .B(n15959), .Y(dpath_mulcore_psum[89]));
XOR2X1 mul_dpath_mulcore_array2_sc4_90__U4(.A(n8245), .B(dpath_mulcore_array2_s2[90]), .Y(n15956));
XOR2X1 mul_dpath_mulcore_array2_sc4_90__U1(.A(dpath_mulcore_array2_c2[89]), .B(n15956), .Y(dpath_mulcore_psum[90]));
XOR2X1 mul_dpath_mulcore_array2_sc4_91__U4(.A(n8244), .B(dpath_mulcore_array2_s2[91]), .Y(n15953));
XOR2X1 mul_dpath_mulcore_array2_sc4_91__U1(.A(dpath_mulcore_array2_c2[90]), .B(n15953), .Y(dpath_mulcore_psum[91]));
XOR2X1 mul_dpath_mulcore_array2_sc4_92__U4(.A(n8243), .B(dpath_mulcore_array2_s2[92]), .Y(n15950));
XOR2X1 mul_dpath_mulcore_array2_sc4_92__U1(.A(dpath_mulcore_array2_c2[91]), .B(n15950), .Y(dpath_mulcore_psum[92]));
XOR2X1 mul_dpath_mulcore_array2_sc4_93__U4(.A(n8242), .B(dpath_mulcore_array2_s2[93]), .Y(n15947));
XOR2X1 mul_dpath_mulcore_array2_sc4_93__U1(.A(dpath_mulcore_array2_c2[92]), .B(n15947), .Y(dpath_mulcore_psum[93]));
XOR2X1 mul_dpath_mulcore_array2_sc4_94__U4(.A(n8241), .B(dpath_mulcore_array2_s2[94]), .Y(n15944));
XOR2X1 mul_dpath_mulcore_array2_sc4_94__U1(.A(dpath_mulcore_array2_c2[93]), .B(n15944), .Y(dpath_mulcore_psum[94]));
XOR2X1 mul_dpath_mulcore_array2_sc4_95__U4(.A(n8240), .B(dpath_mulcore_array2_s2[95]), .Y(n15941));
XOR2X1 mul_dpath_mulcore_array2_sc4_95__U1(.A(dpath_mulcore_array2_c2[94]), .B(n15941), .Y(dpath_mulcore_psum[95]));
XOR2X1 mul_dpath_mulcore_array2_sc4_96__U4(.A(n14897), .B(dpath_mulcore_array2_s2[96]), .Y(n15938));
XOR2X1 mul_dpath_mulcore_array2_sc4_96__U1(.A(dpath_mulcore_array2_c2[95]), .B(n15938), .Y(dpath_mulcore_psum[96]));
XOR2X1 mul_dpath_mulcore_array2_sc4_20__U4(.A(n8239), .B(dpath_mulcore_array2_sc3_20__z), .Y(n15935));
XOR2X1 mul_dpath_mulcore_array2_sc4_20__U1(.A(n8308), .B(n15935), .Y(dpath_mulcore_psum[20]));
XOR2X1 mul_dpath_mulcore_array2_sc4_21__U4(.A(n8238), .B(dpath_mulcore_array2_s3[21]), .Y(n15932));
XOR2X1 mul_dpath_mulcore_array2_sc4_21__U1(.A(n17800), .B(n15932), .Y(dpath_mulcore_psum[21]));
XOR2X1 mul_dpath_mulcore_array2_sc4_22__U4(.A(n8237), .B(dpath_mulcore_array2_s3[22]), .Y(n15929));
XOR2X1 mul_dpath_mulcore_array2_sc4_22__U1(.A(n8376), .B(n15929), .Y(dpath_mulcore_psum[22]));
XOR2X1 mul_dpath_mulcore_array2_sc4_23__U4(.A(n8236), .B(dpath_mulcore_array2_s3[23]), .Y(n15926));
XOR2X1 mul_dpath_mulcore_array2_sc4_23__U1(.A(n8375), .B(n15926), .Y(dpath_mulcore_psum[23]));
XOR2X1 mul_dpath_mulcore_array2_sc4_24__U4(.A(n8235), .B(dpath_mulcore_array2_s3[24]), .Y(n15923));
XOR2X1 mul_dpath_mulcore_array2_sc4_24__U1(.A(n8374), .B(n15923), .Y(dpath_mulcore_psum[24]));
XOR2X1 mul_dpath_mulcore_array2_sc4_25__U4(.A(n8234), .B(dpath_mulcore_array2_s3[25]), .Y(n15920));
XOR2X1 mul_dpath_mulcore_array2_sc4_25__U1(.A(n8373), .B(n15920), .Y(dpath_mulcore_psum[25]));
XOR2X1 mul_dpath_mulcore_array2_sc4_26__U4(.A(n8233), .B(dpath_mulcore_array2_s3[26]), .Y(n15917));
XOR2X1 mul_dpath_mulcore_array2_sc4_26__U1(.A(n8372), .B(n15917), .Y(dpath_mulcore_psum[26]));
XOR2X1 mul_dpath_mulcore_array2_sc4_27__U4(.A(n8232), .B(dpath_mulcore_array2_s3[27]), .Y(n15914));
XOR2X1 mul_dpath_mulcore_array2_sc4_27__U1(.A(n8371), .B(n15914), .Y(dpath_mulcore_psum[27]));
XOR2X1 mul_dpath_mulcore_array2_sc4_28__U4(.A(n8231), .B(dpath_mulcore_array2_s3[28]), .Y(n15911));
XOR2X1 mul_dpath_mulcore_array2_sc4_28__U1(.A(n8370), .B(n15911), .Y(dpath_mulcore_psum[28]));
XOR2X1 mul_dpath_mulcore_array2_sc4_29__U4(.A(n8230), .B(dpath_mulcore_array2_s3[29]), .Y(n15908));
XOR2X1 mul_dpath_mulcore_array2_sc4_29__U1(.A(n8369), .B(n15908), .Y(dpath_mulcore_psum[29]));
XOR2X1 mul_dpath_mulcore_array2_sc4_30__U4(.A(n8229), .B(dpath_mulcore_array2_s3[30]), .Y(n15905));
XOR2X1 mul_dpath_mulcore_array2_sc4_30__U1(.A(n8368), .B(n15905), .Y(dpath_mulcore_psum[30]));
XOR2X1 mul_dpath_mulcore_array2_sc4_31__U4(.A(n8228), .B(dpath_mulcore_array2_s3[31]), .Y(n15902));
XOR2X1 mul_dpath_mulcore_array2_sc4_31__U1(.A(n8367), .B(n15902), .Y(dpath_mulcore_psum[31]));
XOR2X1 mul_dpath_mulcore_array2_sc4_32__U4(.A(n8227), .B(dpath_mulcore_array2_s3[32]), .Y(n15899));
XOR2X1 mul_dpath_mulcore_array2_sc4_32__U1(.A(n8366), .B(n15899), .Y(dpath_mulcore_psum[32]));
XOR2X1 mul_dpath_mulcore_array2_sc4_33__U4(.A(n8226), .B(dpath_mulcore_array2_s3[33]), .Y(n15896));
XOR2X1 mul_dpath_mulcore_array2_sc4_33__U1(.A(n8365), .B(n15896), .Y(dpath_mulcore_psum[33]));
XOR2X1 mul_dpath_mulcore_array2_sc4_34__U4(.A(n8225), .B(dpath_mulcore_array2_s3[34]), .Y(n15893));
XOR2X1 mul_dpath_mulcore_array2_sc4_34__U1(.A(n8364), .B(n15893), .Y(dpath_mulcore_psum[34]));
XOR2X1 mul_dpath_mulcore_array2_sc4_35__U4(.A(n8224), .B(dpath_mulcore_array2_s3[35]), .Y(n15890));
XOR2X1 mul_dpath_mulcore_array2_sc4_35__U1(.A(n8363), .B(n15890), .Y(dpath_mulcore_psum[35]));
XOR2X1 mul_dpath_mulcore_array2_sc4_36__U4(.A(n8223), .B(dpath_mulcore_array2_s3[36]), .Y(n15887));
XOR2X1 mul_dpath_mulcore_array2_sc4_36__U1(.A(n8362), .B(n15887), .Y(dpath_mulcore_psum[36]));
XOR2X1 mul_dpath_mulcore_array2_sc4_37__U4(.A(n8222), .B(dpath_mulcore_array2_s3[37]), .Y(n15884));
XOR2X1 mul_dpath_mulcore_array2_sc4_37__U1(.A(n8361), .B(n15884), .Y(dpath_mulcore_psum[37]));
XOR2X1 mul_dpath_mulcore_array2_sc4_38__U4(.A(n8221), .B(dpath_mulcore_array2_s3[38]), .Y(n15881));
XOR2X1 mul_dpath_mulcore_array2_sc4_38__U1(.A(n8360), .B(n15881), .Y(dpath_mulcore_psum[38]));
XOR2X1 mul_dpath_mulcore_array2_sc4_39__U4(.A(n8220), .B(dpath_mulcore_array2_s3[39]), .Y(n15878));
XOR2X1 mul_dpath_mulcore_array2_sc4_39__U1(.A(n8359), .B(n15878), .Y(dpath_mulcore_psum[39]));
XOR2X1 mul_dpath_mulcore_array2_sc4_40__U4(.A(n8219), .B(dpath_mulcore_array2_s3[40]), .Y(n15875));
XOR2X1 mul_dpath_mulcore_array2_sc4_40__U1(.A(n8358), .B(n15875), .Y(dpath_mulcore_psum[40]));
XOR2X1 mul_dpath_mulcore_array2_sc4_41__U4(.A(n8218), .B(dpath_mulcore_array2_s3[41]), .Y(n15872));
XOR2X1 mul_dpath_mulcore_array2_sc4_41__U1(.A(n8357), .B(n15872), .Y(dpath_mulcore_psum[41]));
XOR2X1 mul_dpath_mulcore_array2_sc4_42__U4(.A(n8217), .B(dpath_mulcore_array2_s3[42]), .Y(n15869));
XOR2X1 mul_dpath_mulcore_array2_sc4_42__U1(.A(n8356), .B(n15869), .Y(dpath_mulcore_psum[42]));
XOR2X1 mul_dpath_mulcore_array2_sc4_43__U4(.A(n8216), .B(dpath_mulcore_array2_s3[43]), .Y(n15866));
XOR2X1 mul_dpath_mulcore_array2_sc4_43__U1(.A(n8355), .B(n15866), .Y(dpath_mulcore_psum[43]));
XOR2X1 mul_dpath_mulcore_array2_sc4_44__U4(.A(n8215), .B(dpath_mulcore_array2_s3[44]), .Y(n15863));
XOR2X1 mul_dpath_mulcore_array2_sc4_44__U1(.A(n8354), .B(n15863), .Y(dpath_mulcore_psum[44]));
XOR2X1 mul_dpath_mulcore_array2_sc4_45__U4(.A(n8214), .B(dpath_mulcore_array2_s3[45]), .Y(n15860));
XOR2X1 mul_dpath_mulcore_array2_sc4_45__U1(.A(n8353), .B(n15860), .Y(dpath_mulcore_psum[45]));
XOR2X1 mul_dpath_mulcore_array2_sc4_46__U4(.A(n8213), .B(dpath_mulcore_array2_s3[46]), .Y(n15857));
XOR2X1 mul_dpath_mulcore_array2_sc4_46__U1(.A(n8352), .B(n15857), .Y(dpath_mulcore_psum[46]));
XOR2X1 mul_dpath_mulcore_array2_sc4_47__U4(.A(n8212), .B(dpath_mulcore_array2_s3[47]), .Y(n15854));
XOR2X1 mul_dpath_mulcore_array2_sc4_47__U1(.A(n8351), .B(n15854), .Y(dpath_mulcore_psum[47]));
XOR2X1 mul_dpath_mulcore_array2_sc4_48__U4(.A(n8211), .B(dpath_mulcore_array2_s3[48]), .Y(n15851));
XOR2X1 mul_dpath_mulcore_array2_sc4_48__U1(.A(n8350), .B(n15851), .Y(dpath_mulcore_psum[48]));
XOR2X1 mul_dpath_mulcore_array2_sc4_49__U4(.A(n8210), .B(dpath_mulcore_array2_s3[49]), .Y(n15848));
XOR2X1 mul_dpath_mulcore_array2_sc4_49__U1(.A(n8349), .B(n15848), .Y(dpath_mulcore_psum[49]));
XOR2X1 mul_dpath_mulcore_array2_sc4_50__U4(.A(n8209), .B(dpath_mulcore_array2_s3[50]), .Y(n15845));
XOR2X1 mul_dpath_mulcore_array2_sc4_50__U1(.A(n8348), .B(n15845), .Y(dpath_mulcore_psum[50]));
XOR2X1 mul_dpath_mulcore_array2_sc4_51__U4(.A(n8208), .B(dpath_mulcore_array2_s3[51]), .Y(n15842));
XOR2X1 mul_dpath_mulcore_array2_sc4_51__U1(.A(n8347), .B(n15842), .Y(dpath_mulcore_psum[51]));
XOR2X1 mul_dpath_mulcore_array2_sc4_52__U4(.A(n8207), .B(dpath_mulcore_array2_s3[52]), .Y(n15839));
XOR2X1 mul_dpath_mulcore_array2_sc4_52__U1(.A(n8346), .B(n15839), .Y(dpath_mulcore_psum[52]));
XOR2X1 mul_dpath_mulcore_array2_sc4_53__U4(.A(n8206), .B(dpath_mulcore_array2_s3[53]), .Y(n15836));
XOR2X1 mul_dpath_mulcore_array2_sc4_53__U1(.A(n8345), .B(n15836), .Y(dpath_mulcore_psum[53]));
XOR2X1 mul_dpath_mulcore_array2_sc4_54__U4(.A(n8205), .B(dpath_mulcore_array2_s3[54]), .Y(n15833));
XOR2X1 mul_dpath_mulcore_array2_sc4_54__U1(.A(n8344), .B(n15833), .Y(dpath_mulcore_psum[54]));
XOR2X1 mul_dpath_mulcore_array2_sc4_55__U4(.A(n8204), .B(dpath_mulcore_array2_s3[55]), .Y(n15830));
XOR2X1 mul_dpath_mulcore_array2_sc4_55__U1(.A(n8343), .B(n15830), .Y(dpath_mulcore_psum[55]));
XOR2X1 mul_dpath_mulcore_array2_sc4_56__U4(.A(n8203), .B(dpath_mulcore_array2_s3[56]), .Y(n15827));
XOR2X1 mul_dpath_mulcore_array2_sc4_56__U1(.A(n8342), .B(n15827), .Y(dpath_mulcore_psum[56]));
XOR2X1 mul_dpath_mulcore_array2_sc4_57__U4(.A(n8202), .B(dpath_mulcore_array2_s3[57]), .Y(n15824));
XOR2X1 mul_dpath_mulcore_array2_sc4_57__U1(.A(n8341), .B(n15824), .Y(dpath_mulcore_psum[57]));
XOR2X1 mul_dpath_mulcore_array2_sc4_58__U4(.A(n8201), .B(dpath_mulcore_array2_s3[58]), .Y(n15821));
XOR2X1 mul_dpath_mulcore_array2_sc4_58__U1(.A(n8340), .B(n15821), .Y(dpath_mulcore_psum[58]));
XOR2X1 mul_dpath_mulcore_array2_sc4_59__U4(.A(n8200), .B(dpath_mulcore_array2_s3[59]), .Y(n15818));
XOR2X1 mul_dpath_mulcore_array2_sc4_59__U1(.A(n8339), .B(n15818), .Y(dpath_mulcore_psum[59]));
XOR2X1 mul_dpath_mulcore_array2_sc4_60__U4(.A(n8199), .B(dpath_mulcore_array2_s3[60]), .Y(n15815));
XOR2X1 mul_dpath_mulcore_array2_sc4_60__U1(.A(n8338), .B(n15815), .Y(dpath_mulcore_psum[60]));
XOR2X1 mul_dpath_mulcore_array2_sc4_61__U4(.A(n8198), .B(dpath_mulcore_array2_s3[61]), .Y(n15812));
XOR2X1 mul_dpath_mulcore_array2_sc4_61__U1(.A(n8337), .B(n15812), .Y(dpath_mulcore_psum[61]));
XOR2X1 mul_dpath_mulcore_array2_sc4_62__U4(.A(n8197), .B(dpath_mulcore_array2_s3[62]), .Y(n15809));
XOR2X1 mul_dpath_mulcore_array2_sc4_62__U1(.A(n8336), .B(n15809), .Y(dpath_mulcore_psum[62]));
XOR2X1 mul_dpath_mulcore_array2_sc4_63__U4(.A(n8196), .B(dpath_mulcore_array2_s3[63]), .Y(n15806));
XOR2X1 mul_dpath_mulcore_array2_sc4_63__U1(.A(n8335), .B(n15806), .Y(dpath_mulcore_psum[63]));
XOR2X1 mul_dpath_mulcore_array2_sc4_64__U4(.A(n8195), .B(dpath_mulcore_array2_s3[64]), .Y(n15803));
XOR2X1 mul_dpath_mulcore_array2_sc4_64__U1(.A(n8334), .B(n15803), .Y(dpath_mulcore_psum[64]));
XOR2X1 mul_dpath_mulcore_array2_sc4_65__U4(.A(n8194), .B(dpath_mulcore_array2_s3[65]), .Y(n15800));
XOR2X1 mul_dpath_mulcore_array2_sc4_65__U1(.A(n8333), .B(n15800), .Y(dpath_mulcore_psum[65]));
XOR2X1 mul_dpath_mulcore_array2_sc4_66__U4(.A(n8193), .B(dpath_mulcore_array2_s3[66]), .Y(n15797));
XOR2X1 mul_dpath_mulcore_array2_sc4_66__U1(.A(n8332), .B(n15797), .Y(dpath_mulcore_psum[66]));
XOR2X1 mul_dpath_mulcore_array2_sc4_67__U4(.A(n8192), .B(dpath_mulcore_array2_s3[67]), .Y(n15794));
XOR2X1 mul_dpath_mulcore_array2_sc4_67__U1(.A(n8331), .B(n15794), .Y(dpath_mulcore_psum[67]));
XOR2X1 mul_dpath_mulcore_array2_sc4_68__U4(.A(n8191), .B(dpath_mulcore_array2_s3[68]), .Y(n15791));
XOR2X1 mul_dpath_mulcore_array2_sc4_68__U1(.A(n8330), .B(n15791), .Y(dpath_mulcore_psum[68]));
XOR2X1 mul_dpath_mulcore_array2_sc4_82__U4(.A(n8385), .B(dpath_mulcore_array2_s2[82]), .Y(n15788));
XOR2X1 mul_dpath_mulcore_array2_sc4_82__U1(.A(dpath_mulcore_array2_c3[81]), .B(n15788), .Y(dpath_mulcore_psum[82]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_4__U4(.A(dpath_mulcore_ary1_a1_s0[4]), .B(n8763), .Y(n15785));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_4__U1(.A(n8382), .B(n15785), .Y(dpath_mulcore_ary1_a1_s_1[4]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_5__U4(.A(dpath_mulcore_ary1_a1_s0[5]), .B(n8936), .Y(n15782));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_5__U1(.A(n8381), .B(n15782), .Y(dpath_mulcore_ary1_a1_s_1[5]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_6__U4(.A(dpath_mulcore_ary1_a1_s0[6]), .B(n8935), .Y(n15779));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_6__U1(.A(dpath_mulcore_ary1_a1_s1[0]), .B(n15779), .Y(dpath_mulcore_ary1_a1_s_1[6]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_7__U4(.A(dpath_mulcore_ary1_a1_s0[7]), .B(n8934), .Y(n15776));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_7__U1(.A(dpath_mulcore_ary1_a1_s1[1]), .B(n15776), .Y(dpath_mulcore_ary1_a1_s_1[7]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_14__U4(.A(dpath_mulcore_ary1_a1_s0[14]), .B(n8931), .Y(n15773));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_14__U1(.A(dpath_mulcore_ary1_a1_s1[8]), .B(n15773), .Y(dpath_mulcore_ary1_a1_s_1[14]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_15__U4(.A(dpath_mulcore_ary1_a1_s0[15]), .B(n8930), .Y(n15770));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_15__U1(.A(dpath_mulcore_ary1_a1_s1[9]), .B(n15770), .Y(dpath_mulcore_ary1_a1_s_1[15]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_16__U4(.A(dpath_mulcore_ary1_a1_s0[16]), .B(n8929), .Y(n15767));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_16__U1(.A(dpath_mulcore_ary1_a1_s1[10]), .B(n15767), .Y(dpath_mulcore_ary1_a1_s_1[16]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_17__U4(.A(dpath_mulcore_ary1_a1_s0[17]), .B(n8928), .Y(n15764));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_17__U1(.A(dpath_mulcore_ary1_a1_s1[11]), .B(n15764), .Y(dpath_mulcore_ary1_a1_s_1[17]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_18__U4(.A(dpath_mulcore_ary1_a1_s0[18]), .B(n8927), .Y(n15761));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_18__U1(.A(dpath_mulcore_ary1_a1_s1[12]), .B(n15761), .Y(dpath_mulcore_ary1_a1_s_1[18]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_19__U4(.A(dpath_mulcore_ary1_a1_s0[19]), .B(n8926), .Y(n15758));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_19__U1(.A(dpath_mulcore_ary1_a1_s1[13]), .B(n15758), .Y(dpath_mulcore_ary1_a1_s_1[19]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_20__U4(.A(dpath_mulcore_ary1_a1_s0[20]), .B(n8925), .Y(n15755));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_20__U1(.A(dpath_mulcore_ary1_a1_s1[14]), .B(n15755), .Y(dpath_mulcore_ary1_a1_s_1[20]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_21__U4(.A(dpath_mulcore_ary1_a1_s0[21]), .B(n8924), .Y(n15752));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_21__U1(.A(dpath_mulcore_ary1_a1_s1[15]), .B(n15752), .Y(dpath_mulcore_ary1_a1_s_1[21]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_22__U4(.A(dpath_mulcore_ary1_a1_s0[22]), .B(n8923), .Y(n15749));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_22__U1(.A(dpath_mulcore_ary1_a1_s1[16]), .B(n15749), .Y(dpath_mulcore_ary1_a1_s_1[22]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_23__U4(.A(dpath_mulcore_ary1_a1_s0[23]), .B(n8922), .Y(n15746));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_23__U1(.A(dpath_mulcore_ary1_a1_s1[17]), .B(n15746), .Y(dpath_mulcore_ary1_a1_s_1[23]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_24__U4(.A(dpath_mulcore_ary1_a1_s0[24]), .B(n8921), .Y(n15743));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_24__U1(.A(dpath_mulcore_ary1_a1_s1[18]), .B(n15743), .Y(dpath_mulcore_ary1_a1_s_1[24]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_25__U4(.A(dpath_mulcore_ary1_a1_s0[25]), .B(n8920), .Y(n15740));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_25__U1(.A(dpath_mulcore_ary1_a1_s1[19]), .B(n15740), .Y(dpath_mulcore_ary1_a1_s_1[25]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_26__U4(.A(dpath_mulcore_ary1_a1_s0[26]), .B(n8919), .Y(n15737));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_26__U1(.A(dpath_mulcore_ary1_a1_s1[20]), .B(n15737), .Y(dpath_mulcore_ary1_a1_s_1[26]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_27__U4(.A(dpath_mulcore_ary1_a1_s0[27]), .B(n8918), .Y(n15734));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_27__U1(.A(dpath_mulcore_ary1_a1_s1[21]), .B(n15734), .Y(dpath_mulcore_ary1_a1_s_1[27]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_28__U4(.A(dpath_mulcore_ary1_a1_s0[28]), .B(n8917), .Y(n15731));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_28__U1(.A(dpath_mulcore_ary1_a1_s1[22]), .B(n15731), .Y(dpath_mulcore_ary1_a1_s_1[28]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_29__U4(.A(dpath_mulcore_ary1_a1_s0[29]), .B(n8916), .Y(n15728));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_29__U1(.A(dpath_mulcore_ary1_a1_s1[23]), .B(n15728), .Y(dpath_mulcore_ary1_a1_s_1[29]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_30__U4(.A(dpath_mulcore_ary1_a1_s0[30]), .B(n8915), .Y(n15725));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_30__U1(.A(dpath_mulcore_ary1_a1_s1[24]), .B(n15725), .Y(dpath_mulcore_ary1_a1_s_1[30]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_31__U4(.A(dpath_mulcore_ary1_a1_s0[31]), .B(n8914), .Y(n15722));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_31__U1(.A(dpath_mulcore_ary1_a1_s1[25]), .B(n15722), .Y(dpath_mulcore_ary1_a1_s_1[31]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_32__U4(.A(dpath_mulcore_ary1_a1_s0[32]), .B(n8913), .Y(n15719));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_32__U1(.A(dpath_mulcore_ary1_a1_s1[26]), .B(n15719), .Y(dpath_mulcore_ary1_a1_s_1[32]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_33__U4(.A(dpath_mulcore_ary1_a1_s0[33]), .B(n8912), .Y(n15716));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_33__U1(.A(dpath_mulcore_ary1_a1_s1[27]), .B(n15716), .Y(dpath_mulcore_ary1_a1_s_1[33]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_34__U4(.A(dpath_mulcore_ary1_a1_s0[34]), .B(n8911), .Y(n15713));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_34__U1(.A(dpath_mulcore_ary1_a1_s1[28]), .B(n15713), .Y(dpath_mulcore_ary1_a1_s_1[34]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_35__U4(.A(dpath_mulcore_ary1_a1_s0[35]), .B(n8910), .Y(n15710));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_35__U1(.A(dpath_mulcore_ary1_a1_s1[29]), .B(n15710), .Y(dpath_mulcore_ary1_a1_s_1[35]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_36__U4(.A(dpath_mulcore_ary1_a1_s0[36]), .B(n8909), .Y(n15707));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_36__U1(.A(dpath_mulcore_ary1_a1_s1[30]), .B(n15707), .Y(dpath_mulcore_ary1_a1_s_1[36]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_37__U4(.A(dpath_mulcore_ary1_a1_s0[37]), .B(n8908), .Y(n15704));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_37__U1(.A(dpath_mulcore_ary1_a1_s1[31]), .B(n15704), .Y(dpath_mulcore_ary1_a1_s_1[37]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_38__U4(.A(dpath_mulcore_ary1_a1_s0[38]), .B(n8907), .Y(n15701));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_38__U1(.A(dpath_mulcore_ary1_a1_s1[32]), .B(n15701), .Y(dpath_mulcore_ary1_a1_s_1[38]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_39__U4(.A(dpath_mulcore_ary1_a1_s0[39]), .B(n8906), .Y(n15698));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_39__U1(.A(dpath_mulcore_ary1_a1_s1[33]), .B(n15698), .Y(dpath_mulcore_ary1_a1_s_1[39]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_40__U4(.A(dpath_mulcore_ary1_a1_s0[40]), .B(n8905), .Y(n15695));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_40__U1(.A(dpath_mulcore_ary1_a1_s1[34]), .B(n15695), .Y(dpath_mulcore_ary1_a1_s_1[40]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_41__U4(.A(dpath_mulcore_ary1_a1_s0[41]), .B(n8904), .Y(n15692));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_41__U1(.A(dpath_mulcore_ary1_a1_s1[35]), .B(n15692), .Y(dpath_mulcore_ary1_a1_s_1[41]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_42__U4(.A(dpath_mulcore_ary1_a1_s0[42]), .B(n8903), .Y(n15689));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_42__U1(.A(dpath_mulcore_ary1_a1_s1[36]), .B(n15689), .Y(dpath_mulcore_ary1_a1_s_1[42]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_43__U4(.A(dpath_mulcore_ary1_a1_s0[43]), .B(n8902), .Y(n15686));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_43__U1(.A(dpath_mulcore_ary1_a1_s1[37]), .B(n15686), .Y(dpath_mulcore_ary1_a1_s_1[43]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_44__U4(.A(dpath_mulcore_ary1_a1_s0[44]), .B(n8901), .Y(n15683));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_44__U1(.A(dpath_mulcore_ary1_a1_s1[38]), .B(n15683), .Y(dpath_mulcore_ary1_a1_s_1[44]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_45__U4(.A(dpath_mulcore_ary1_a1_s0[45]), .B(n8900), .Y(n15680));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_45__U1(.A(dpath_mulcore_ary1_a1_s1[39]), .B(n15680), .Y(dpath_mulcore_ary1_a1_s_1[45]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_46__U4(.A(dpath_mulcore_ary1_a1_s0[46]), .B(n8899), .Y(n15677));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_46__U1(.A(dpath_mulcore_ary1_a1_s1[40]), .B(n15677), .Y(dpath_mulcore_ary1_a1_s_1[46]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_47__U4(.A(dpath_mulcore_ary1_a1_s0[47]), .B(n8898), .Y(n15674));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_47__U1(.A(dpath_mulcore_ary1_a1_s1[41]), .B(n15674), .Y(dpath_mulcore_ary1_a1_s_1[47]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_48__U4(.A(dpath_mulcore_ary1_a1_s0[48]), .B(n8897), .Y(n15671));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_48__U1(.A(dpath_mulcore_ary1_a1_s1[42]), .B(n15671), .Y(dpath_mulcore_ary1_a1_s_1[48]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_49__U4(.A(dpath_mulcore_ary1_a1_s0[49]), .B(n8896), .Y(n15668));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_49__U1(.A(dpath_mulcore_ary1_a1_s1[43]), .B(n15668), .Y(dpath_mulcore_ary1_a1_s_1[49]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_50__U4(.A(dpath_mulcore_ary1_a1_s0[50]), .B(n8895), .Y(n15665));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_50__U1(.A(dpath_mulcore_ary1_a1_s1[44]), .B(n15665), .Y(dpath_mulcore_ary1_a1_s_1[50]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_51__U4(.A(dpath_mulcore_ary1_a1_s0[51]), .B(n8894), .Y(n15662));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_51__U1(.A(dpath_mulcore_ary1_a1_s1[45]), .B(n15662), .Y(dpath_mulcore_ary1_a1_s_1[51]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_52__U4(.A(dpath_mulcore_ary1_a1_s0[52]), .B(n8893), .Y(n15659));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_52__U1(.A(dpath_mulcore_ary1_a1_s1[46]), .B(n15659), .Y(dpath_mulcore_ary1_a1_s_1[52]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_53__U4(.A(dpath_mulcore_ary1_a1_s0[53]), .B(n8892), .Y(n15656));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_53__U1(.A(dpath_mulcore_ary1_a1_s1[47]), .B(n15656), .Y(dpath_mulcore_ary1_a1_s_1[53]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_54__U4(.A(dpath_mulcore_ary1_a1_s0[54]), .B(n8891), .Y(n15653));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_54__U1(.A(dpath_mulcore_ary1_a1_s1[48]), .B(n15653), .Y(dpath_mulcore_ary1_a1_s_1[54]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_55__U4(.A(dpath_mulcore_ary1_a1_s0[55]), .B(n8890), .Y(n15650));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_55__U1(.A(dpath_mulcore_ary1_a1_s1[49]), .B(n15650), .Y(dpath_mulcore_ary1_a1_s_1[55]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_56__U4(.A(dpath_mulcore_ary1_a1_s0[56]), .B(n8889), .Y(n15647));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_56__U1(.A(dpath_mulcore_ary1_a1_s1[50]), .B(n15647), .Y(dpath_mulcore_ary1_a1_s_1[56]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_57__U4(.A(dpath_mulcore_ary1_a1_s0[57]), .B(n8888), .Y(n15644));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_57__U1(.A(dpath_mulcore_ary1_a1_s1[51]), .B(n15644), .Y(dpath_mulcore_ary1_a1_s_1[57]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_58__U4(.A(dpath_mulcore_ary1_a1_s0[58]), .B(n8887), .Y(n15641));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_58__U1(.A(dpath_mulcore_ary1_a1_s1[52]), .B(n15641), .Y(dpath_mulcore_ary1_a1_s_1[58]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_59__U4(.A(dpath_mulcore_ary1_a1_s0[59]), .B(n8886), .Y(n15638));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_59__U1(.A(dpath_mulcore_ary1_a1_s1[53]), .B(n15638), .Y(dpath_mulcore_ary1_a1_s_1[59]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_60__U4(.A(dpath_mulcore_ary1_a1_s0[60]), .B(n8885), .Y(n15635));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_60__U1(.A(dpath_mulcore_ary1_a1_s1[54]), .B(n15635), .Y(dpath_mulcore_ary1_a1_s_1[60]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_61__U4(.A(dpath_mulcore_ary1_a1_s0[61]), .B(n8884), .Y(n15632));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_61__U1(.A(dpath_mulcore_ary1_a1_s1[55]), .B(n15632), .Y(dpath_mulcore_ary1_a1_s_1[61]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_62__U4(.A(dpath_mulcore_ary1_a1_s0[62]), .B(n8883), .Y(n15629));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_62__U1(.A(dpath_mulcore_ary1_a1_s1[56]), .B(n15629), .Y(dpath_mulcore_ary1_a1_s_1[62]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_63__U4(.A(dpath_mulcore_ary1_a1_s0[63]), .B(n8882), .Y(n15626));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_63__U1(.A(dpath_mulcore_ary1_a1_s1[57]), .B(n15626), .Y(dpath_mulcore_ary1_a1_s_1[63]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_64__U4(.A(dpath_mulcore_ary1_a1_s0[64]), .B(n8881), .Y(n15623));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_64__U1(.A(dpath_mulcore_ary1_a1_s1[58]), .B(n15623), .Y(dpath_mulcore_ary1_a1_s_1[64]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_65__U4(.A(dpath_mulcore_ary1_a1_s0[65]), .B(n8942), .Y(n15620));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_65__U1(.A(dpath_mulcore_ary1_a1_s1[59]), .B(n15620), .Y(dpath_mulcore_ary1_a1_s_1[65]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_66__U4(.A(dpath_mulcore_ary1_a1_s0[66]), .B(n8943), .Y(n15617));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_66__U1(.A(dpath_mulcore_ary1_a1_s1[60]), .B(n15617), .Y(dpath_mulcore_ary1_a1_s_1[66]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_67__U4(.A(dpath_mulcore_ary1_a1_s0[67]), .B(n8944), .Y(n15614));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_67__U1(.A(dpath_mulcore_ary1_a1_s1[61]), .B(n15614), .Y(dpath_mulcore_ary1_a1_s_1[67]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_68__U4(.A(dpath_mulcore_ary1_a1_I0_I2_net073), .B(n14798), .Y(n15611));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_68__U1(.A(dpath_mulcore_ary1_a1_s1[62]), .B(n15611), .Y(dpath_mulcore_ary1_a1_s_1[68]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_69__U4(.A(n9427), .B(n9489), .Y(n15608));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_69__U1(.A(dpath_mulcore_ary1_a1_s1[63]), .B(n15608), .Y(dpath_mulcore_ary1_a1_s_1[69]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_72__U4(.A(dpath_mulcore_ary1_a1_s2[60]), .B(n8825), .Y(n15605));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_72__U1(.A(n8189), .B(n15605), .Y(dpath_mulcore_ary1_a1_s_2[72]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_73__U4(.A(dpath_mulcore_ary1_a1_s2[61]), .B(n8824), .Y(n15602));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_73__U1(.A(n8190), .B(n15602), .Y(dpath_mulcore_ary1_a1_s_2[73]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_74__U4(.A(dpath_mulcore_ary1_a1_s2[62]), .B(n8823), .Y(n15599));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_74__U1(.A(n14790), .B(n15599), .Y(dpath_mulcore_ary1_a1_s_2[74]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_75__U4(.A(dpath_mulcore_ary1_a1_s2[63]), .B(n8822), .Y(n15596));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_75__U1(.A(n9487), .B(n15596), .Y(dpath_mulcore_ary1_a1_s_2[75]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_71__U4(.A(dpath_mulcore_ary1_a1_s2[59]), .B(n8826), .Y(n15593));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_71__U1(.A(n8188), .B(n15593), .Y(dpath_mulcore_ary1_a1_s_2[71]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_8__U4(.A(n8302), .B(dpath_mulcore_ary1_a1_s_1[8]), .Y(n15590));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_8__U1(.A(dpath_mulcore_ary1_a1_c1[1]), .B(n15590), .Y(dpath_mulcore_a1sum[8]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_9__U4(.A(n8296), .B(dpath_mulcore_ary1_a1_s_1[9]), .Y(n15587));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_9__U1(.A(n8065), .B(n15587), .Y(dpath_mulcore_a1sum[9]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_10__U4(.A(n8295), .B(dpath_mulcore_ary1_a1_s_1[10]), .Y(n15584));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_10__U1(.A(dpath_mulcore_ary1_a1_s_2[10]), .B(n15584), .Y(dpath_mulcore_a1sum[10]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_3__U4(.A(dpath_mulcore_ary1_a1_s0[3]), .B(n8764), .Y(n15581));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_3__U1(.A(dpath_mulcore_ary1_a1_c_1[2]), .B(n15581), .Y(dpath_mulcore_a1sum[3]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_8__U4(.A(dpath_mulcore_ary1_a1_s0[8]), .B(n8933), .Y(n15578));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_8__U1(.A(dpath_mulcore_ary1_a1_s1[2]), .B(n15578), .Y(dpath_mulcore_ary1_a1_s_1[8]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_9__U4(.A(dpath_mulcore_ary1_a1_s0[9]), .B(n8932), .Y(n15575));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_9__U1(.A(dpath_mulcore_ary1_a1_s1[3]), .B(n15575), .Y(dpath_mulcore_ary1_a1_s_1[9]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_77__U4(.A(dpath_mulcore_ary1_a1_s2[65]), .B(n8941), .Y(n15572));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_77__U1(.A(n8294), .B(n15572), .Y(dpath_mulcore_a1sum[77]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_10__U4(.A(n8380), .B(dpath_mulcore_ary1_a1_s1[4]), .Y(n15568));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_10__U1(.A(n8064), .B(n15568), .Y(dpath_mulcore_ary1_a1_s_2[10]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_11__U4(.A(n8379), .B(dpath_mulcore_ary1_a1_s1[5]), .Y(n15565));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_11__U1(.A(n8187), .B(n15565), .Y(dpath_mulcore_ary1_a1_s_2[11]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_12__U4(.A(dpath_mulcore_ary1_a1_s2[0]), .B(dpath_mulcore_ary1_a1_s1[6]), .Y(n15562));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_12__U1(.A(n8186), .B(n15562), .Y(dpath_mulcore_ary1_a1_s_2[12]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_13__U4(.A(dpath_mulcore_ary1_a1_s2[1]), .B(dpath_mulcore_ary1_a1_s1[7]), .Y(n15559));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_13__U1(.A(n8185), .B(n15559), .Y(dpath_mulcore_ary1_a1_s_2[13]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_14__U4(.A(dpath_mulcore_ary1_a1_s2[2]), .B(dpath_mulcore_ary1_a1_c2[1]), .Y(n15556));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_14__U1(.A(n8184), .B(n15556), .Y(dpath_mulcore_ary1_a1_s_2[14]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_15__U4(.A(dpath_mulcore_ary1_a1_s2[3]), .B(n8762), .Y(n15553));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_15__U1(.A(n8183), .B(n15553), .Y(dpath_mulcore_ary1_a1_s_2[15]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_16__U4(.A(dpath_mulcore_ary1_a1_s2[4]), .B(n8761), .Y(n15550));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_16__U1(.A(n8182), .B(n15550), .Y(dpath_mulcore_ary1_a1_s_2[16]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_17__U4(.A(dpath_mulcore_ary1_a1_s2[5]), .B(n8880), .Y(n15547));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_17__U1(.A(n8181), .B(n15547), .Y(dpath_mulcore_ary1_a1_s_2[17]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_18__U4(.A(dpath_mulcore_ary1_a1_s2[6]), .B(n8879), .Y(n15544));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_18__U1(.A(n8180), .B(n15544), .Y(dpath_mulcore_ary1_a1_s_2[18]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_19__U4(.A(dpath_mulcore_ary1_a1_s2[7]), .B(n8878), .Y(n15541));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_19__U1(.A(n8179), .B(n15541), .Y(dpath_mulcore_ary1_a1_s_2[19]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_20__U4(.A(dpath_mulcore_ary1_a1_s2[8]), .B(n8877), .Y(n15538));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_20__U1(.A(n8178), .B(n15538), .Y(dpath_mulcore_ary1_a1_s_2[20]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_21__U4(.A(dpath_mulcore_ary1_a1_s2[9]), .B(n8876), .Y(n15535));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_21__U1(.A(n8177), .B(n15535), .Y(dpath_mulcore_ary1_a1_s_2[21]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_22__U4(.A(dpath_mulcore_ary1_a1_s2[10]), .B(n8875), .Y(n15532));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_22__U1(.A(n8176), .B(n15532), .Y(dpath_mulcore_ary1_a1_s_2[22]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_23__U4(.A(dpath_mulcore_ary1_a1_s2[11]), .B(n8874), .Y(n15529));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_23__U1(.A(n8175), .B(n15529), .Y(dpath_mulcore_ary1_a1_s_2[23]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_24__U4(.A(dpath_mulcore_ary1_a1_s2[12]), .B(n8873), .Y(n15526));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_24__U1(.A(n8174), .B(n15526), .Y(dpath_mulcore_ary1_a1_s_2[24]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_25__U4(.A(dpath_mulcore_ary1_a1_s2[13]), .B(n8872), .Y(n15523));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_25__U1(.A(n8173), .B(n15523), .Y(dpath_mulcore_ary1_a1_s_2[25]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_26__U4(.A(dpath_mulcore_ary1_a1_s2[14]), .B(n8871), .Y(n15520));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_26__U1(.A(n8172), .B(n15520), .Y(dpath_mulcore_ary1_a1_s_2[26]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_27__U4(.A(dpath_mulcore_ary1_a1_s2[15]), .B(n8870), .Y(n15517));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_27__U1(.A(n8171), .B(n15517), .Y(dpath_mulcore_ary1_a1_s_2[27]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_28__U4(.A(dpath_mulcore_ary1_a1_s2[16]), .B(n8869), .Y(n15514));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_28__U1(.A(n8170), .B(n15514), .Y(dpath_mulcore_ary1_a1_s_2[28]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_29__U4(.A(dpath_mulcore_ary1_a1_s2[17]), .B(n8868), .Y(n15511));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_29__U1(.A(n8169), .B(n15511), .Y(dpath_mulcore_ary1_a1_s_2[29]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_30__U4(.A(dpath_mulcore_ary1_a1_s2[18]), .B(n8867), .Y(n15508));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_30__U1(.A(n8168), .B(n15508), .Y(dpath_mulcore_ary1_a1_s_2[30]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_31__U4(.A(dpath_mulcore_ary1_a1_s2[19]), .B(n8866), .Y(n15505));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_31__U1(.A(n8167), .B(n15505), .Y(dpath_mulcore_ary1_a1_s_2[31]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_32__U4(.A(dpath_mulcore_ary1_a1_s2[20]), .B(n8865), .Y(n15502));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_32__U1(.A(n8166), .B(n15502), .Y(dpath_mulcore_ary1_a1_s_2[32]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_33__U4(.A(dpath_mulcore_ary1_a1_s2[21]), .B(n8864), .Y(n15499));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_33__U1(.A(n8165), .B(n15499), .Y(dpath_mulcore_ary1_a1_s_2[33]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_34__U4(.A(dpath_mulcore_ary1_a1_s2[22]), .B(n8863), .Y(n15496));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_34__U1(.A(n8164), .B(n15496), .Y(dpath_mulcore_ary1_a1_s_2[34]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_35__U4(.A(dpath_mulcore_ary1_a1_s2[23]), .B(n8862), .Y(n15493));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_35__U1(.A(n8163), .B(n15493), .Y(dpath_mulcore_ary1_a1_s_2[35]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_36__U4(.A(dpath_mulcore_ary1_a1_s2[24]), .B(n8861), .Y(n15490));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_36__U1(.A(n8162), .B(n15490), .Y(dpath_mulcore_ary1_a1_s_2[36]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_37__U4(.A(dpath_mulcore_ary1_a1_s2[25]), .B(n8860), .Y(n15487));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_37__U1(.A(n8161), .B(n15487), .Y(dpath_mulcore_ary1_a1_s_2[37]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_38__U4(.A(dpath_mulcore_ary1_a1_s2[26]), .B(n8859), .Y(n15484));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_38__U1(.A(n8160), .B(n15484), .Y(dpath_mulcore_ary1_a1_s_2[38]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_39__U4(.A(dpath_mulcore_ary1_a1_s2[27]), .B(n8858), .Y(n15481));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_39__U1(.A(n8159), .B(n15481), .Y(dpath_mulcore_ary1_a1_s_2[39]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_40__U4(.A(dpath_mulcore_ary1_a1_s2[28]), .B(n8857), .Y(n15478));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_40__U1(.A(n8158), .B(n15478), .Y(dpath_mulcore_ary1_a1_s_2[40]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_41__U4(.A(dpath_mulcore_ary1_a1_s2[29]), .B(n8856), .Y(n15475));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_41__U1(.A(n8157), .B(n15475), .Y(dpath_mulcore_ary1_a1_s_2[41]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_42__U4(.A(dpath_mulcore_ary1_a1_s2[30]), .B(n8855), .Y(n15472));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_42__U1(.A(n8156), .B(n15472), .Y(dpath_mulcore_ary1_a1_s_2[42]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_43__U4(.A(dpath_mulcore_ary1_a1_s2[31]), .B(n8854), .Y(n15469));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_43__U1(.A(n8155), .B(n15469), .Y(dpath_mulcore_ary1_a1_s_2[43]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_44__U4(.A(dpath_mulcore_ary1_a1_s2[32]), .B(n8853), .Y(n15466));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_44__U1(.A(n8154), .B(n15466), .Y(dpath_mulcore_ary1_a1_s_2[44]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_45__U4(.A(dpath_mulcore_ary1_a1_s2[33]), .B(n8852), .Y(n15463));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_45__U1(.A(n8153), .B(n15463), .Y(dpath_mulcore_ary1_a1_s_2[45]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_46__U4(.A(dpath_mulcore_ary1_a1_s2[34]), .B(n8851), .Y(n15460));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_46__U1(.A(n8152), .B(n15460), .Y(dpath_mulcore_ary1_a1_s_2[46]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_47__U4(.A(dpath_mulcore_ary1_a1_s2[35]), .B(n8850), .Y(n15457));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_47__U1(.A(n8151), .B(n15457), .Y(dpath_mulcore_ary1_a1_s_2[47]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_48__U4(.A(dpath_mulcore_ary1_a1_s2[36]), .B(n8849), .Y(n15454));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_48__U1(.A(n8150), .B(n15454), .Y(dpath_mulcore_ary1_a1_s_2[48]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_49__U4(.A(dpath_mulcore_ary1_a1_s2[37]), .B(n8848), .Y(n15451));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_49__U1(.A(n8149), .B(n15451), .Y(dpath_mulcore_ary1_a1_s_2[49]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_50__U4(.A(dpath_mulcore_ary1_a1_s2[38]), .B(n8847), .Y(n15448));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_50__U1(.A(n8148), .B(n15448), .Y(dpath_mulcore_ary1_a1_s_2[50]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_51__U4(.A(dpath_mulcore_ary1_a1_s2[39]), .B(n8846), .Y(n15445));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_51__U1(.A(n8147), .B(n15445), .Y(dpath_mulcore_ary1_a1_s_2[51]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_52__U4(.A(dpath_mulcore_ary1_a1_s2[40]), .B(n8845), .Y(n15442));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_52__U1(.A(n8146), .B(n15442), .Y(dpath_mulcore_ary1_a1_s_2[52]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_53__U4(.A(dpath_mulcore_ary1_a1_s2[41]), .B(n8844), .Y(n15439));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_53__U1(.A(n8145), .B(n15439), .Y(dpath_mulcore_ary1_a1_s_2[53]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_54__U4(.A(dpath_mulcore_ary1_a1_s2[42]), .B(n8843), .Y(n15436));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_54__U1(.A(n8144), .B(n15436), .Y(dpath_mulcore_ary1_a1_s_2[54]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_55__U4(.A(dpath_mulcore_ary1_a1_s2[43]), .B(n8842), .Y(n15433));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_55__U1(.A(n8143), .B(n15433), .Y(dpath_mulcore_ary1_a1_s_2[55]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_56__U4(.A(dpath_mulcore_ary1_a1_s2[44]), .B(n8841), .Y(n15430));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_56__U1(.A(n8142), .B(n15430), .Y(dpath_mulcore_ary1_a1_s_2[56]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_57__U4(.A(dpath_mulcore_ary1_a1_s2[45]), .B(n8840), .Y(n15427));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_57__U1(.A(n8141), .B(n15427), .Y(dpath_mulcore_ary1_a1_s_2[57]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_58__U4(.A(dpath_mulcore_ary1_a1_s2[46]), .B(n8839), .Y(n15424));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_58__U1(.A(n8140), .B(n15424), .Y(dpath_mulcore_ary1_a1_s_2[58]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_59__U4(.A(dpath_mulcore_ary1_a1_s2[47]), .B(n8838), .Y(n15421));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_59__U1(.A(n8139), .B(n15421), .Y(dpath_mulcore_ary1_a1_s_2[59]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_60__U4(.A(dpath_mulcore_ary1_a1_s2[48]), .B(n8837), .Y(n15418));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_60__U1(.A(n8138), .B(n15418), .Y(dpath_mulcore_ary1_a1_s_2[60]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_61__U4(.A(dpath_mulcore_ary1_a1_s2[49]), .B(n8836), .Y(n15415));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_61__U1(.A(n8137), .B(n15415), .Y(dpath_mulcore_ary1_a1_s_2[61]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_62__U4(.A(dpath_mulcore_ary1_a1_s2[50]), .B(n8835), .Y(n15412));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_62__U1(.A(n8136), .B(n15412), .Y(dpath_mulcore_ary1_a1_s_2[62]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_63__U4(.A(dpath_mulcore_ary1_a1_s2[51]), .B(n8834), .Y(n15409));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_63__U1(.A(n8135), .B(n15409), .Y(dpath_mulcore_ary1_a1_s_2[63]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_64__U4(.A(dpath_mulcore_ary1_a1_s2[52]), .B(n8833), .Y(n15406));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_64__U1(.A(n8134), .B(n15406), .Y(dpath_mulcore_ary1_a1_s_2[64]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_65__U4(.A(dpath_mulcore_ary1_a1_s2[53]), .B(n8832), .Y(n15403));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_65__U1(.A(n8133), .B(n15403), .Y(dpath_mulcore_ary1_a1_s_2[65]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_66__U4(.A(dpath_mulcore_ary1_a1_s2[54]), .B(n8831), .Y(n15400));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_66__U1(.A(n8132), .B(n15400), .Y(dpath_mulcore_ary1_a1_s_2[66]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_67__U4(.A(dpath_mulcore_ary1_a1_s2[55]), .B(n8830), .Y(n15397));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_67__U1(.A(n8131), .B(n15397), .Y(dpath_mulcore_ary1_a1_s_2[67]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_68__U4(.A(dpath_mulcore_ary1_a1_s2[56]), .B(n8829), .Y(n15394));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_68__U1(.A(n8130), .B(n15394), .Y(dpath_mulcore_ary1_a1_s_2[68]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_69__U4(.A(dpath_mulcore_ary1_a1_s2[57]), .B(n8828), .Y(n15391));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_69__U1(.A(n8129), .B(n15391), .Y(dpath_mulcore_ary1_a1_s_2[69]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_70__U4(.A(dpath_mulcore_ary1_a1_s2[58]), .B(n8827), .Y(n15388));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_70__U1(.A(n8128), .B(n15388), .Y(dpath_mulcore_ary1_a1_s_2[70]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_4__U4(.A(dpath_mulcore_ary1_a0_s0[4]), .B(n8759), .Y(n15385));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_4__U1(.A(n8378), .B(n15385), .Y(dpath_mulcore_ary1_a0_s_1[4]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_5__U4(.A(dpath_mulcore_ary1_a0_s0[5]), .B(n8820), .Y(n15382));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_5__U1(.A(n8377), .B(n15382), .Y(dpath_mulcore_ary1_a0_s_1[5]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_6__U4(.A(dpath_mulcore_ary1_a0_s0[6]), .B(n8819), .Y(n15379));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_6__U1(.A(dpath_mulcore_ary1_a0_s1[0]), .B(n15379), .Y(dpath_mulcore_ary1_a0_s_1[6]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_7__U4(.A(dpath_mulcore_ary1_a0_s0[7]), .B(n8818), .Y(n15376));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_7__U1(.A(dpath_mulcore_ary1_a0_s1[1]), .B(n15376), .Y(dpath_mulcore_ary1_a0_s_1[7]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_14__U4(.A(dpath_mulcore_ary1_a0_s0[14]), .B(n8815), .Y(n15373));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_14__U1(.A(dpath_mulcore_ary1_a0_s1[8]), .B(n15373), .Y(dpath_mulcore_ary1_a0_s_1[14]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_15__U4(.A(dpath_mulcore_ary1_a0_s0[15]), .B(n8814), .Y(n15370));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_15__U1(.A(dpath_mulcore_ary1_a0_s1[9]), .B(n15370), .Y(dpath_mulcore_ary1_a0_s_1[15]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_16__U4(.A(dpath_mulcore_ary1_a0_s0[16]), .B(n8813), .Y(n15367));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_16__U1(.A(dpath_mulcore_ary1_a0_s1[10]), .B(n15367), .Y(dpath_mulcore_ary1_a0_s_1[16]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_17__U4(.A(dpath_mulcore_ary1_a0_s0[17]), .B(n8812), .Y(n15364));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_17__U1(.A(dpath_mulcore_ary1_a0_s1[11]), .B(n15364), .Y(dpath_mulcore_ary1_a0_s_1[17]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_18__U4(.A(dpath_mulcore_ary1_a0_s0[18]), .B(n8811), .Y(n15361));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_18__U1(.A(dpath_mulcore_ary1_a0_s1[12]), .B(n15361), .Y(dpath_mulcore_ary1_a0_s_1[18]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_19__U4(.A(dpath_mulcore_ary1_a0_s0[19]), .B(n8810), .Y(n15358));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_19__U1(.A(dpath_mulcore_ary1_a0_s1[13]), .B(n15358), .Y(dpath_mulcore_ary1_a0_s_1[19]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_20__U4(.A(dpath_mulcore_ary1_a0_s0[20]), .B(n8809), .Y(n15355));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_20__U1(.A(dpath_mulcore_ary1_a0_s1[14]), .B(n15355), .Y(dpath_mulcore_ary1_a0_s_1[20]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_21__U4(.A(dpath_mulcore_ary1_a0_s0[21]), .B(n8808), .Y(n15352));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_21__U1(.A(dpath_mulcore_ary1_a0_s1[15]), .B(n15352), .Y(dpath_mulcore_ary1_a0_s_1[21]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_22__U4(.A(dpath_mulcore_ary1_a0_s0[22]), .B(n8807), .Y(n15349));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_22__U1(.A(dpath_mulcore_ary1_a0_s1[16]), .B(n15349), .Y(dpath_mulcore_ary1_a0_s_1[22]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_23__U4(.A(dpath_mulcore_ary1_a0_s0[23]), .B(n8806), .Y(n15346));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_23__U1(.A(dpath_mulcore_ary1_a0_s1[17]), .B(n15346), .Y(dpath_mulcore_ary1_a0_s_1[23]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_24__U4(.A(dpath_mulcore_ary1_a0_s0[24]), .B(n8805), .Y(n15343));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_24__U1(.A(dpath_mulcore_ary1_a0_s1[18]), .B(n15343), .Y(dpath_mulcore_ary1_a0_s_1[24]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_25__U4(.A(dpath_mulcore_ary1_a0_s0[25]), .B(n8804), .Y(n15340));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_25__U1(.A(dpath_mulcore_ary1_a0_s1[19]), .B(n15340), .Y(dpath_mulcore_ary1_a0_s_1[25]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_26__U4(.A(dpath_mulcore_ary1_a0_s0[26]), .B(n8803), .Y(n15337));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_26__U1(.A(dpath_mulcore_ary1_a0_s1[20]), .B(n15337), .Y(dpath_mulcore_ary1_a0_s_1[26]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_27__U4(.A(dpath_mulcore_ary1_a0_s0[27]), .B(n8802), .Y(n15334));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_27__U1(.A(dpath_mulcore_ary1_a0_s1[21]), .B(n15334), .Y(dpath_mulcore_ary1_a0_s_1[27]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_28__U4(.A(dpath_mulcore_ary1_a0_s0[28]), .B(n8801), .Y(n15331));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_28__U1(.A(dpath_mulcore_ary1_a0_s1[22]), .B(n15331), .Y(dpath_mulcore_ary1_a0_s_1[28]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_29__U4(.A(dpath_mulcore_ary1_a0_s0[29]), .B(n8800), .Y(n15328));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_29__U1(.A(dpath_mulcore_ary1_a0_s1[23]), .B(n15328), .Y(dpath_mulcore_ary1_a0_s_1[29]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_30__U4(.A(dpath_mulcore_ary1_a0_s0[30]), .B(n8799), .Y(n15325));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_30__U1(.A(dpath_mulcore_ary1_a0_s1[24]), .B(n15325), .Y(dpath_mulcore_ary1_a0_s_1[30]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_31__U4(.A(dpath_mulcore_ary1_a0_s0[31]), .B(n8798), .Y(n15322));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_31__U1(.A(dpath_mulcore_ary1_a0_s1[25]), .B(n15322), .Y(dpath_mulcore_ary1_a0_s_1[31]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_32__U4(.A(dpath_mulcore_ary1_a0_s0[32]), .B(n8797), .Y(n15319));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_32__U1(.A(dpath_mulcore_ary1_a0_s1[26]), .B(n15319), .Y(dpath_mulcore_ary1_a0_s_1[32]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_33__U4(.A(dpath_mulcore_ary1_a0_s0[33]), .B(n8796), .Y(n15316));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_33__U1(.A(dpath_mulcore_ary1_a0_s1[27]), .B(n15316), .Y(dpath_mulcore_ary1_a0_s_1[33]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_34__U4(.A(dpath_mulcore_ary1_a0_s0[34]), .B(n8795), .Y(n15313));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_34__U1(.A(dpath_mulcore_ary1_a0_s1[28]), .B(n15313), .Y(dpath_mulcore_ary1_a0_s_1[34]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_35__U4(.A(dpath_mulcore_ary1_a0_s0[35]), .B(n8794), .Y(n15310));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_35__U1(.A(dpath_mulcore_ary1_a0_s1[29]), .B(n15310), .Y(dpath_mulcore_ary1_a0_s_1[35]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_36__U4(.A(dpath_mulcore_ary1_a0_s0[36]), .B(n8793), .Y(n15307));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_36__U1(.A(dpath_mulcore_ary1_a0_s1[30]), .B(n15307), .Y(dpath_mulcore_ary1_a0_s_1[36]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_37__U4(.A(dpath_mulcore_ary1_a0_s0[37]), .B(n8792), .Y(n15304));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_37__U1(.A(dpath_mulcore_ary1_a0_s1[31]), .B(n15304), .Y(dpath_mulcore_ary1_a0_s_1[37]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_38__U4(.A(dpath_mulcore_ary1_a0_s0[38]), .B(n8791), .Y(n15301));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_38__U1(.A(dpath_mulcore_ary1_a0_s1[32]), .B(n15301), .Y(dpath_mulcore_ary1_a0_s_1[38]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_39__U4(.A(dpath_mulcore_ary1_a0_s0[39]), .B(n8790), .Y(n15298));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_39__U1(.A(dpath_mulcore_ary1_a0_s1[33]), .B(n15298), .Y(dpath_mulcore_ary1_a0_s_1[39]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_40__U4(.A(dpath_mulcore_ary1_a0_s0[40]), .B(n8789), .Y(n15295));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_40__U1(.A(dpath_mulcore_ary1_a0_s1[34]), .B(n15295), .Y(dpath_mulcore_ary1_a0_s_1[40]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_41__U4(.A(dpath_mulcore_ary1_a0_s0[41]), .B(n8788), .Y(n15292));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_41__U1(.A(dpath_mulcore_ary1_a0_s1[35]), .B(n15292), .Y(dpath_mulcore_ary1_a0_s_1[41]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_42__U4(.A(dpath_mulcore_ary1_a0_s0[42]), .B(n8787), .Y(n15289));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_42__U1(.A(dpath_mulcore_ary1_a0_s1[36]), .B(n15289), .Y(dpath_mulcore_ary1_a0_s_1[42]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_43__U4(.A(dpath_mulcore_ary1_a0_s0[43]), .B(n8786), .Y(n15286));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_43__U1(.A(dpath_mulcore_ary1_a0_s1[37]), .B(n15286), .Y(dpath_mulcore_ary1_a0_s_1[43]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_44__U4(.A(dpath_mulcore_ary1_a0_s0[44]), .B(n8785), .Y(n15283));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_44__U1(.A(dpath_mulcore_ary1_a0_s1[38]), .B(n15283), .Y(dpath_mulcore_ary1_a0_s_1[44]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_45__U4(.A(dpath_mulcore_ary1_a0_s0[45]), .B(n8784), .Y(n15280));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_45__U1(.A(dpath_mulcore_ary1_a0_s1[39]), .B(n15280), .Y(dpath_mulcore_ary1_a0_s_1[45]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_46__U4(.A(dpath_mulcore_ary1_a0_s0[46]), .B(n8783), .Y(n15277));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_46__U1(.A(dpath_mulcore_ary1_a0_s1[40]), .B(n15277), .Y(dpath_mulcore_ary1_a0_s_1[46]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_47__U4(.A(dpath_mulcore_ary1_a0_s0[47]), .B(n8782), .Y(n15274));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_47__U1(.A(dpath_mulcore_ary1_a0_s1[41]), .B(n15274), .Y(dpath_mulcore_ary1_a0_s_1[47]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_48__U4(.A(dpath_mulcore_ary1_a0_s0[48]), .B(n8781), .Y(n15271));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_48__U1(.A(dpath_mulcore_ary1_a0_s1[42]), .B(n15271), .Y(dpath_mulcore_ary1_a0_s_1[48]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_49__U4(.A(dpath_mulcore_ary1_a0_s0[49]), .B(n8780), .Y(n15268));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_49__U1(.A(dpath_mulcore_ary1_a0_s1[43]), .B(n15268), .Y(dpath_mulcore_ary1_a0_s_1[49]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_50__U4(.A(dpath_mulcore_ary1_a0_s0[50]), .B(n8779), .Y(n15265));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_50__U1(.A(dpath_mulcore_ary1_a0_s1[44]), .B(n15265), .Y(dpath_mulcore_ary1_a0_s_1[50]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_51__U4(.A(dpath_mulcore_ary1_a0_s0[51]), .B(n8778), .Y(n15262));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_51__U1(.A(dpath_mulcore_ary1_a0_s1[45]), .B(n15262), .Y(dpath_mulcore_ary1_a0_s_1[51]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_52__U4(.A(dpath_mulcore_ary1_a0_s0[52]), .B(n8777), .Y(n15259));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_52__U1(.A(dpath_mulcore_ary1_a0_s1[46]), .B(n15259), .Y(dpath_mulcore_ary1_a0_s_1[52]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_53__U4(.A(dpath_mulcore_ary1_a0_s0[53]), .B(n8776), .Y(n15256));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_53__U1(.A(dpath_mulcore_ary1_a0_s1[47]), .B(n15256), .Y(dpath_mulcore_ary1_a0_s_1[53]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_54__U4(.A(dpath_mulcore_ary1_a0_s0[54]), .B(n8775), .Y(n15253));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_54__U1(.A(dpath_mulcore_ary1_a0_s1[48]), .B(n15253), .Y(dpath_mulcore_ary1_a0_s_1[54]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_55__U4(.A(dpath_mulcore_ary1_a0_s0[55]), .B(n8774), .Y(n15250));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_55__U1(.A(dpath_mulcore_ary1_a0_s1[49]), .B(n15250), .Y(dpath_mulcore_ary1_a0_s_1[55]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_56__U4(.A(dpath_mulcore_ary1_a0_s0[56]), .B(n8773), .Y(n15247));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_56__U1(.A(dpath_mulcore_ary1_a0_s1[50]), .B(n15247), .Y(dpath_mulcore_ary1_a0_s_1[56]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_57__U4(.A(dpath_mulcore_ary1_a0_s0[57]), .B(n8772), .Y(n15244));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_57__U1(.A(dpath_mulcore_ary1_a0_s1[51]), .B(n15244), .Y(dpath_mulcore_ary1_a0_s_1[57]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_58__U4(.A(dpath_mulcore_ary1_a0_s0[58]), .B(n8771), .Y(n15241));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_58__U1(.A(dpath_mulcore_ary1_a0_s1[52]), .B(n15241), .Y(dpath_mulcore_ary1_a0_s_1[58]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_59__U4(.A(dpath_mulcore_ary1_a0_s0[59]), .B(n8770), .Y(n15238));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_59__U1(.A(dpath_mulcore_ary1_a0_s1[53]), .B(n15238), .Y(dpath_mulcore_ary1_a0_s_1[59]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_60__U4(.A(dpath_mulcore_ary1_a0_s0[60]), .B(n8769), .Y(n15235));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_60__U1(.A(dpath_mulcore_ary1_a0_s1[54]), .B(n15235), .Y(dpath_mulcore_ary1_a0_s_1[60]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_61__U4(.A(dpath_mulcore_ary1_a0_s0[61]), .B(n8768), .Y(n15232));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_61__U1(.A(dpath_mulcore_ary1_a0_s1[55]), .B(n15232), .Y(dpath_mulcore_ary1_a0_s_1[61]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_62__U4(.A(dpath_mulcore_ary1_a0_s0[62]), .B(n8767), .Y(n15229));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_62__U1(.A(dpath_mulcore_ary1_a0_s1[56]), .B(n15229), .Y(dpath_mulcore_ary1_a0_s_1[62]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_63__U4(.A(dpath_mulcore_ary1_a0_s0[63]), .B(n8766), .Y(n15226));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_63__U1(.A(dpath_mulcore_ary1_a0_s1[57]), .B(n15226), .Y(dpath_mulcore_ary1_a0_s_1[63]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_64__U4(.A(dpath_mulcore_ary1_a0_s0[64]), .B(n8765), .Y(n15223));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_64__U1(.A(dpath_mulcore_ary1_a0_s1[58]), .B(n15223), .Y(dpath_mulcore_ary1_a0_s_1[64]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_65__U4(.A(dpath_mulcore_ary1_a0_s0[65]), .B(n8937), .Y(n15220));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_65__U1(.A(dpath_mulcore_ary1_a0_s1[59]), .B(n15220), .Y(dpath_mulcore_ary1_a0_s_1[65]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_66__U4(.A(dpath_mulcore_ary1_a0_s0[66]), .B(n8938), .Y(n15217));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_66__U1(.A(dpath_mulcore_ary1_a0_s1[60]), .B(n15217), .Y(dpath_mulcore_ary1_a0_s_1[66]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_67__U4(.A(dpath_mulcore_ary1_a0_s0[67]), .B(n8939), .Y(n15214));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_67__U1(.A(dpath_mulcore_ary1_a0_s1[61]), .B(n15214), .Y(dpath_mulcore_ary1_a0_s_1[67]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_68__U4(.A(dpath_mulcore_ary1_a0_I0_I2_net073), .B(n8940), .Y(n15211));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_68__U1(.A(dpath_mulcore_ary1_a0_s1[62]), .B(n15211), .Y(dpath_mulcore_ary1_a0_s_1[68]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_69__U4(.A(n9425), .B(n9488), .Y(n15208));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_69__U1(.A(dpath_mulcore_ary1_a0_s1[63]), .B(n15208), .Y(dpath_mulcore_ary1_a0_s_1[69]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_72__U4(.A(n13750), .B(n13751), .Y(n15205));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_72__U1(.A(n8327), .B(n15205), .Y(dpath_mulcore_ary1_a0_s_2[72]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_73__U4(.A(n13748), .B(n13749), .Y(n15202));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_73__U1(.A(n8326), .B(n15202), .Y(dpath_mulcore_ary1_a0_s_2[73]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_74__U4(.A(n13746), .B(n13747), .Y(n15199));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_74__U1(.A(n16580), .B(n15199), .Y(dpath_mulcore_ary1_a0_s_2[74]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_75__U4(.A(n16572), .B(n13745), .Y(n15196));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_75__U1(.A(n9486), .B(n15196), .Y(dpath_mulcore_ary1_a0_s_2[75]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_71__U4(.A(n13752), .B(n13753), .Y(n15193));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_71__U1(.A(n8328), .B(n15193), .Y(dpath_mulcore_ary1_a0_s_2[71]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_8__U4(.A(n8293), .B(dpath_mulcore_ary1_a0_s_1[8]), .Y(n15190));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_8__U1(.A(dpath_mulcore_ary1_a0_c1[1]), .B(n15190), .Y(dpath_mulcore_a0sum[8]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_9__U4(.A(n8287), .B(dpath_mulcore_ary1_a0_s_1[9]), .Y(n15187));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_9__U1(.A(n8057), .B(n15187), .Y(dpath_mulcore_a0sum[9]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_10__U4(.A(n8286), .B(dpath_mulcore_ary1_a0_s_1[10]), .Y(n15184));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_10__U1(.A(dpath_mulcore_ary1_a0_s_2[10]), .B(n15184), .Y(dpath_mulcore_a0sum[10]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_3__U4(.A(dpath_mulcore_ary1_a0_s0[3]), .B(n8760), .Y(n15181));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_3__U1(.A(dpath_mulcore_ary1_a0_c_1[2]), .B(n15181), .Y(dpath_mulcore_a0sum[3]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_8__U4(.A(dpath_mulcore_ary1_a0_s0[8]), .B(n8817), .Y(n15178));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_8__U1(.A(dpath_mulcore_ary1_a0_s1[2]), .B(n15178), .Y(dpath_mulcore_ary1_a0_s_1[8]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_9__U4(.A(dpath_mulcore_ary1_a0_s0[9]), .B(n8816), .Y(n15175));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_9__U1(.A(dpath_mulcore_ary1_a0_s1[3]), .B(n15175), .Y(dpath_mulcore_ary1_a0_s_1[9]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_77__U4(.A(n16568), .B(n16571), .Y(n15172));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_77__U1(.A(n8285), .B(n15172), .Y(dpath_mulcore_a0sum[77]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_10__U4(.A(n8387), .B(dpath_mulcore_ary1_a0_s1[4]), .Y(n15168));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_10__U1(.A(n8056), .B(n15168), .Y(dpath_mulcore_ary1_a0_s_2[10]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_11__U4(.A(n8386), .B(dpath_mulcore_ary1_a0_s1[5]), .Y(n15165));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_11__U1(.A(n8127), .B(n15165), .Y(dpath_mulcore_ary1_a0_s_2[11]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_12__U4(.A(dpath_mulcore_ary1_a0_s2[0]), .B(dpath_mulcore_ary1_a0_s1[6]), .Y(n15162));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_12__U1(.A(n8126), .B(n15162), .Y(dpath_mulcore_ary1_a0_s_2[12]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_13__U4(.A(dpath_mulcore_ary1_a0_s2[1]), .B(dpath_mulcore_ary1_a0_s1[7]), .Y(n15159));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_13__U1(.A(n8125), .B(n15159), .Y(dpath_mulcore_ary1_a0_s_2[13]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_14__U4(.A(dpath_mulcore_ary1_a0_s2[2]), .B(dpath_mulcore_ary1_a0_c2[1]), .Y(n15156));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_14__U1(.A(n8124), .B(n15156), .Y(dpath_mulcore_ary1_a0_s_2[14]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_15__U4(.A(dpath_mulcore_ary1_a0_s2[3]), .B(n8975), .Y(n15153));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_15__U1(.A(n8123), .B(n15153), .Y(dpath_mulcore_ary1_a0_s_2[15]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_16__U4(.A(n13862), .B(n8976), .Y(n15150));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_16__U1(.A(n8122), .B(n15150), .Y(dpath_mulcore_ary1_a0_s_2[16]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_17__U4(.A(n13860), .B(n13861), .Y(n15147));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_17__U1(.A(n8121), .B(n15147), .Y(dpath_mulcore_ary1_a0_s_2[17]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_18__U4(.A(n13858), .B(n13859), .Y(n15144));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_18__U1(.A(n8120), .B(n15144), .Y(dpath_mulcore_ary1_a0_s_2[18]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_19__U4(.A(n13856), .B(n13857), .Y(n15141));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_19__U1(.A(n8119), .B(n15141), .Y(dpath_mulcore_ary1_a0_s_2[19]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_20__U4(.A(n13854), .B(n13855), .Y(n15138));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_20__U1(.A(n8118), .B(n15138), .Y(dpath_mulcore_ary1_a0_s_2[20]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_21__U4(.A(n13852), .B(n13853), .Y(n15135));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_21__U1(.A(n8117), .B(n15135), .Y(dpath_mulcore_ary1_a0_s_2[21]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_22__U4(.A(n13850), .B(n13851), .Y(n15132));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_22__U1(.A(n8116), .B(n15132), .Y(dpath_mulcore_ary1_a0_s_2[22]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_23__U4(.A(n13848), .B(n13849), .Y(n15129));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_23__U1(.A(n8115), .B(n15129), .Y(dpath_mulcore_ary1_a0_s_2[23]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_24__U4(.A(n13846), .B(n13847), .Y(n15126));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_24__U1(.A(n8114), .B(n15126), .Y(dpath_mulcore_ary1_a0_s_2[24]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_25__U4(.A(n13844), .B(n13845), .Y(n15123));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_25__U1(.A(n8113), .B(n15123), .Y(dpath_mulcore_ary1_a0_s_2[25]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_26__U4(.A(n13842), .B(n13843), .Y(n15120));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_26__U1(.A(n8112), .B(n15120), .Y(dpath_mulcore_ary1_a0_s_2[26]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_27__U4(.A(n13840), .B(n13841), .Y(n15117));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_27__U1(.A(n8111), .B(n15117), .Y(dpath_mulcore_ary1_a0_s_2[27]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_28__U4(.A(n13838), .B(n13839), .Y(n15114));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_28__U1(.A(n8110), .B(n15114), .Y(dpath_mulcore_ary1_a0_s_2[28]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_29__U4(.A(n13836), .B(n13837), .Y(n15111));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_29__U1(.A(n8109), .B(n15111), .Y(dpath_mulcore_ary1_a0_s_2[29]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_30__U4(.A(n13834), .B(n13835), .Y(n15108));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_30__U1(.A(n8108), .B(n15108), .Y(dpath_mulcore_ary1_a0_s_2[30]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_31__U4(.A(n13832), .B(n13833), .Y(n15105));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_31__U1(.A(n8107), .B(n15105), .Y(dpath_mulcore_ary1_a0_s_2[31]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_32__U4(.A(n13830), .B(n13831), .Y(n15102));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_32__U1(.A(n8106), .B(n15102), .Y(dpath_mulcore_ary1_a0_s_2[32]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_33__U4(.A(n13828), .B(n13829), .Y(n15099));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_33__U1(.A(n8105), .B(n15099), .Y(dpath_mulcore_ary1_a0_s_2[33]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_34__U4(.A(n13826), .B(n13827), .Y(n15096));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_34__U1(.A(n8104), .B(n15096), .Y(dpath_mulcore_ary1_a0_s_2[34]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_35__U4(.A(n13824), .B(n13825), .Y(n15093));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_35__U1(.A(n8103), .B(n15093), .Y(dpath_mulcore_ary1_a0_s_2[35]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_36__U4(.A(n13822), .B(n13823), .Y(n15090));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_36__U1(.A(n8102), .B(n15090), .Y(dpath_mulcore_ary1_a0_s_2[36]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_37__U4(.A(n13820), .B(n13821), .Y(n15087));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_37__U1(.A(n8101), .B(n15087), .Y(dpath_mulcore_ary1_a0_s_2[37]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_38__U4(.A(n13818), .B(n13819), .Y(n15084));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_38__U1(.A(n8100), .B(n15084), .Y(dpath_mulcore_ary1_a0_s_2[38]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_39__U4(.A(n13816), .B(n13817), .Y(n15081));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_39__U1(.A(n8099), .B(n15081), .Y(dpath_mulcore_ary1_a0_s_2[39]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_40__U4(.A(n13814), .B(n13815), .Y(n15078));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_40__U1(.A(n8098), .B(n15078), .Y(dpath_mulcore_ary1_a0_s_2[40]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_41__U4(.A(n13812), .B(n13813), .Y(n15075));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_41__U1(.A(n8097), .B(n15075), .Y(dpath_mulcore_ary1_a0_s_2[41]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_42__U4(.A(n13810), .B(n13811), .Y(n15072));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_42__U1(.A(n8096), .B(n15072), .Y(dpath_mulcore_ary1_a0_s_2[42]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_43__U4(.A(n13808), .B(n13809), .Y(n15069));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_43__U1(.A(n8095), .B(n15069), .Y(dpath_mulcore_ary1_a0_s_2[43]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_44__U4(.A(n13806), .B(n13807), .Y(n15066));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_44__U1(.A(n8094), .B(n15066), .Y(dpath_mulcore_ary1_a0_s_2[44]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_45__U4(.A(n13804), .B(n13805), .Y(n15063));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_45__U1(.A(n8093), .B(n15063), .Y(dpath_mulcore_ary1_a0_s_2[45]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_46__U4(.A(n13802), .B(n13803), .Y(n15060));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_46__U1(.A(n8092), .B(n15060), .Y(dpath_mulcore_ary1_a0_s_2[46]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_47__U4(.A(n13800), .B(n13801), .Y(n15057));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_47__U1(.A(n8091), .B(n15057), .Y(dpath_mulcore_ary1_a0_s_2[47]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_48__U4(.A(n13798), .B(n13799), .Y(n15054));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_48__U1(.A(n8090), .B(n15054), .Y(dpath_mulcore_ary1_a0_s_2[48]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_49__U4(.A(n13796), .B(n13797), .Y(n15051));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_49__U1(.A(n8089), .B(n15051), .Y(dpath_mulcore_ary1_a0_s_2[49]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_50__U4(.A(n13794), .B(n13795), .Y(n15048));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_50__U1(.A(n8088), .B(n15048), .Y(dpath_mulcore_ary1_a0_s_2[50]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_51__U4(.A(n13792), .B(n13793), .Y(n15045));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_51__U1(.A(n8087), .B(n15045), .Y(dpath_mulcore_ary1_a0_s_2[51]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_52__U4(.A(n13790), .B(n13791), .Y(n15042));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_52__U1(.A(n8086), .B(n15042), .Y(dpath_mulcore_ary1_a0_s_2[52]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_53__U4(.A(n13788), .B(n13789), .Y(n15039));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_53__U1(.A(n8085), .B(n15039), .Y(dpath_mulcore_ary1_a0_s_2[53]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_54__U4(.A(n13786), .B(n13787), .Y(n15036));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_54__U1(.A(n8084), .B(n15036), .Y(dpath_mulcore_ary1_a0_s_2[54]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_55__U4(.A(n13784), .B(n13785), .Y(n15033));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_55__U1(.A(n8083), .B(n15033), .Y(dpath_mulcore_ary1_a0_s_2[55]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_56__U4(.A(n13782), .B(n13783), .Y(n15030));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_56__U1(.A(n8082), .B(n15030), .Y(dpath_mulcore_ary1_a0_s_2[56]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_57__U4(.A(n13780), .B(n13781), .Y(n15027));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_57__U1(.A(n8081), .B(n15027), .Y(dpath_mulcore_ary1_a0_s_2[57]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_58__U4(.A(n13778), .B(n13779), .Y(n15024));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_58__U1(.A(n8080), .B(n15024), .Y(dpath_mulcore_ary1_a0_s_2[58]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_59__U4(.A(n13776), .B(n13777), .Y(n15021));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_59__U1(.A(n8079), .B(n15021), .Y(dpath_mulcore_ary1_a0_s_2[59]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_60__U4(.A(n13774), .B(n13775), .Y(n15018));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_60__U1(.A(n8078), .B(n15018), .Y(dpath_mulcore_ary1_a0_s_2[60]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_61__U4(.A(n13772), .B(n13773), .Y(n15015));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_61__U1(.A(n8077), .B(n15015), .Y(dpath_mulcore_ary1_a0_s_2[61]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_62__U4(.A(n13770), .B(n13771), .Y(n15012));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_62__U1(.A(n8076), .B(n15012), .Y(dpath_mulcore_ary1_a0_s_2[62]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_63__U4(.A(n13768), .B(n13769), .Y(n15009));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_63__U1(.A(n8075), .B(n15009), .Y(dpath_mulcore_ary1_a0_s_2[63]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_64__U4(.A(n13766), .B(n13767), .Y(n15006));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_64__U1(.A(n8074), .B(n15006), .Y(dpath_mulcore_ary1_a0_s_2[64]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_65__U4(.A(n13764), .B(n13765), .Y(n15003));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_65__U1(.A(n8073), .B(n15003), .Y(dpath_mulcore_ary1_a0_s_2[65]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_66__U4(.A(n13762), .B(n13763), .Y(n15000));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_66__U1(.A(n8072), .B(n15000), .Y(dpath_mulcore_ary1_a0_s_2[66]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_67__U4(.A(n13760), .B(n13761), .Y(n14997));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_67__U1(.A(n8071), .B(n14997), .Y(dpath_mulcore_ary1_a0_s_2[67]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_68__U4(.A(n13758), .B(n13759), .Y(n14994));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_68__U1(.A(n8070), .B(n14994), .Y(dpath_mulcore_ary1_a0_s_2[68]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_69__U4(.A(n13756), .B(n13757), .Y(n14991));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_69__U1(.A(n8069), .B(n14991), .Y(dpath_mulcore_ary1_a0_s_2[69]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_sc1_1__U2(.A(dpath_mulcore_ary1_a0_I2_I0_b0n), .B(n7396), .Y(dpath_mulcore_ary1_a0_s2[1]));
XOR2X1 mul_dpath_mulcore_array2_sc1x2_U2(.A(dpath_mulcore_pc[30]), .B(dpath_mulcore_ps[31]), .Y(dpath_mulcore_array2_s1x2));
XOR2X1 mul_dpath_mulcore_array2_sc2_0__U2(.A(dpath_mulcore_array2_c1x2), .B(dpath_mulcore_array2_s1[0]), .Y(dpath_mulcore_array2_s2[0]));
XOR2X1 mul_dpath_mulcore_array2_sc2_1__U2(.A(n7226), .B(dpath_mulcore_array2_s1[1]), .Y(dpath_mulcore_array2_s2[1]));
XOR2X1 mul_dpath_mulcore_array2_sc2_2__U2(.A(n7212), .B(dpath_mulcore_array2_s1[2]), .Y(dpath_mulcore_array2_s2[2]));
XOR2X1 mul_dpath_mulcore_array2_sc2_3__U2(.A(n7211), .B(dpath_mulcore_array2_s1[3]), .Y(dpath_mulcore_array2_s2[3]));
XOR2X1 mul_dpath_mulcore_array2_sc2_4__U2(.A(n7210), .B(dpath_mulcore_array2_s1[4]), .Y(dpath_mulcore_array2_s2[4]));
XOR2X1 mul_dpath_mulcore_array2_accx2_U2(.A(dpath_mulcore_array2_s1x2), .B(n14968), .Y(dpath_mulcore_psumx2));
XOR2X1 mul_dpath_mulcore_array2_sc3_69__U2(.A(n7225), .B(dpath_mulcore_array2_s2[69]), .Y(dpath_mulcore_array2_s3[69]));
XOR2X1 mul_dpath_mulcore_array2_sc3_70__U2(.A(n7224), .B(dpath_mulcore_array2_s2[70]), .Y(dpath_mulcore_array2_s3[70]));
XOR2X1 mul_dpath_mulcore_array2_sc3_71__U2(.A(n7223), .B(dpath_mulcore_array2_s2[71]), .Y(dpath_mulcore_array2_s3[71]));
XOR2X1 mul_dpath_mulcore_array2_sc3_72__U2(.A(n7222), .B(dpath_mulcore_array2_s2[72]), .Y(dpath_mulcore_array2_s3[72]));
XOR2X1 mul_dpath_mulcore_array2_sc3_73__U2(.A(n7221), .B(dpath_mulcore_array2_s2[73]), .Y(dpath_mulcore_array2_s3[73]));
XOR2X1 mul_dpath_mulcore_array2_sc3_74__U2(.A(n7220), .B(dpath_mulcore_array2_s2[74]), .Y(dpath_mulcore_array2_s3[74]));
XOR2X1 mul_dpath_mulcore_array2_sc3_75__U2(.A(n7219), .B(dpath_mulcore_array2_s2[75]), .Y(dpath_mulcore_array2_s3[75]));
XOR2X1 mul_dpath_mulcore_array2_sc3_76__U2(.A(n7218), .B(dpath_mulcore_array2_s2[76]), .Y(dpath_mulcore_array2_s3[76]));
XOR2X1 mul_dpath_mulcore_array2_sc3_77__U2(.A(n7217), .B(dpath_mulcore_array2_s2[77]), .Y(dpath_mulcore_array2_s3[77]));
XOR2X1 mul_dpath_mulcore_array2_sc3_78__U2(.A(n7216), .B(dpath_mulcore_array2_s2[78]), .Y(dpath_mulcore_array2_s3[78]));
XOR2X1 mul_dpath_mulcore_array2_sc3_79__U2(.A(n7215), .B(dpath_mulcore_array2_s2[79]), .Y(dpath_mulcore_array2_s3[79]));
XOR2X1 mul_dpath_mulcore_array2_sc3_80__U2(.A(n7214), .B(dpath_mulcore_array2_s2[80]), .Y(dpath_mulcore_array2_s3[80]));
XOR2X1 mul_dpath_mulcore_array2_sc3_81__U2(.A(n7213), .B(dpath_mulcore_array2_s2[81]), .Y(dpath_mulcore_array2_s3[81]));
XOR2X1 mul_dpath_mulcore_array2_sc2_84__U2(.A(dpath_mulcore_a1c[67]), .B(dpath_mulcore_a1s[68]), .Y(dpath_mulcore_array2_s2[84]));
XOR2X1 mul_dpath_mulcore_array2_sc2_85__U2(.A(dpath_mulcore_a1c[68]), .B(dpath_mulcore_a1s[69]), .Y(dpath_mulcore_array2_s2[85]));
XOR2X1 mul_dpath_mulcore_array2_sc2_86__U2(.A(dpath_mulcore_a1c[69]), .B(dpath_mulcore_a1s[70]), .Y(dpath_mulcore_array2_s2[86]));
XOR2X1 mul_dpath_mulcore_array2_sc2_87__U2(.A(dpath_mulcore_a1c[70]), .B(dpath_mulcore_a1s[71]), .Y(dpath_mulcore_array2_s2[87]));
XOR2X1 mul_dpath_mulcore_array2_sc2_88__U2(.A(dpath_mulcore_a1c[71]), .B(dpath_mulcore_a1s[72]), .Y(dpath_mulcore_array2_s2[88]));
XOR2X1 mul_dpath_mulcore_array2_sc2_89__U2(.A(dpath_mulcore_a1c[72]), .B(dpath_mulcore_a1s[73]), .Y(dpath_mulcore_array2_s2[89]));
XOR2X1 mul_dpath_mulcore_array2_sc2_90__U2(.A(dpath_mulcore_a1c[73]), .B(dpath_mulcore_a1s[74]), .Y(dpath_mulcore_array2_s2[90]));
XOR2X1 mul_dpath_mulcore_array2_sc2_91__U2(.A(dpath_mulcore_a1c[74]), .B(dpath_mulcore_a1s[75]), .Y(dpath_mulcore_array2_s2[91]));
XOR2X1 mul_dpath_mulcore_array2_sc2_92__U2(.A(dpath_mulcore_a1c[75]), .B(dpath_mulcore_a1s[76]), .Y(dpath_mulcore_array2_s2[92]));
XOR2X1 mul_dpath_mulcore_array2_sc2_93__U2(.A(dpath_mulcore_a1c[76]), .B(dpath_mulcore_a1s[77]), .Y(dpath_mulcore_array2_s2[93]));
XOR2X1 mul_dpath_mulcore_array2_sc2_94__U2(.A(dpath_mulcore_a1c[77]), .B(dpath_mulcore_a1s[78]), .Y(dpath_mulcore_array2_s2[94]));
XOR2X1 mul_dpath_mulcore_array2_sc2_95__U2(.A(dpath_mulcore_a1c[78]), .B(dpath_mulcore_a1s[79]), .Y(dpath_mulcore_array2_s2[95]));
XOR2X1 mul_dpath_mulcore_array2_sc2_96__U2(.A(dpath_mulcore_a1c[79]), .B(dpath_mulcore_a1s[80]), .Y(dpath_mulcore_array2_s2[96]));
XOR2X1 mul_dpath_mulcore_array2_acc_0__U2(.A(dpath_mulcore_array2_s2[0]), .B(n7407), .Y(dpath_mulcore_psum[0]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_11__U2(.A(n7206), .B(dpath_mulcore_ary1_a1_s0[11]), .Y(dpath_mulcore_ary1_a1_s_1[11]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_12__U2(.A(n7205), .B(dpath_mulcore_ary1_a1_s0[12]), .Y(dpath_mulcore_ary1_a1_s_1[12]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_13__U2(.A(n7204), .B(dpath_mulcore_ary1_a1_s0[13]), .Y(dpath_mulcore_ary1_a1_s_1[13]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_2__U2(.A(dpath_mulcore_ary1_a1_c0[1]), .B(dpath_mulcore_ary1_a1_s0[2]), .Y(dpath_mulcore_a1sum[2]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_78__U2(.A(n7208), .B(dpath_mulcore_ary1_a1_s2[66]), .Y(dpath_mulcore_a1sum[78]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_2_79__U2(.A(n7209), .B(dpath_mulcore_ary1_a1_s2[67]), .Y(dpath_mulcore_a1sum[79]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_4__U2(.A(dpath_mulcore_ary1_a1_s_1[4]), .B(n7412), .Y(dpath_mulcore_a1sum[4]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_5__U2(.A(dpath_mulcore_ary1_a1_s_1[5]), .B(n7415), .Y(dpath_mulcore_a1sum[5]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_6__U2(.A(dpath_mulcore_ary1_a1_s_1[6]), .B(n7414), .Y(dpath_mulcore_a1sum[6]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc3_7__U2(.A(dpath_mulcore_ary1_a1_s_1[7]), .B(n7413), .Y(dpath_mulcore_a1sum[7]));
XOR2X1 mul_dpath_mulcore_ary1_a1_sc2_1_10__U2(.A(n7207), .B(dpath_mulcore_ary1_a1_s0[10]), .Y(dpath_mulcore_ary1_a1_s_1[10]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_11__U2(.A(n7202), .B(dpath_mulcore_ary1_a0_s0[11]), .Y(dpath_mulcore_ary1_a0_s_1[11]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_12__U2(.A(n7201), .B(dpath_mulcore_ary1_a0_s0[12]), .Y(dpath_mulcore_ary1_a0_s_1[12]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_13__U2(.A(n7200), .B(dpath_mulcore_ary1_a0_s0[13]), .Y(dpath_mulcore_ary1_a0_s_1[13]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_1_2__U2(.A(dpath_mulcore_ary1_a0_c0[1]), .B(dpath_mulcore_ary1_a0_s0[2]), .Y(dpath_mulcore_a0sum[2]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_78__U2(.A(n16569), .B(dpath_mulcore_ary1_a0_I2_I2_net38), .Y(dpath_mulcore_a0sum[78]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc2_2_79__U2(.A(n9474), .B(n9312), .Y(dpath_mulcore_a0sum[79]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_4__U2(.A(dpath_mulcore_ary1_a0_s_1[4]), .B(n7408), .Y(dpath_mulcore_a0sum[4]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_5__U2(.A(dpath_mulcore_ary1_a0_s_1[5]), .B(n7411), .Y(dpath_mulcore_a0sum[5]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_6__U2(.A(dpath_mulcore_ary1_a0_s_1[6]), .B(n7410), .Y(dpath_mulcore_a0sum[6]));
XOR2X1 mul_dpath_mulcore_ary1_a0_sc3_7__U2(.A(dpath_mulcore_ary1_a0_s_1[7]), .B(n7409), .Y(dpath_mulcore_a0sum[7]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_sc1_67__U1(.A(n7926), .B(n9482), .Y(dpath_mulcore_ary1_a1_s0[67]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_sc1_66__U1(.A(n7927), .B(dpath_mulcore_ary1_a1_I0_I2_net38), .Y(dpath_mulcore_ary1_a1_s0[66]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_sc1_65__U1(.A(n7928), .B(n14796), .Y(dpath_mulcore_ary1_a1_s0[65]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_sc1_65__U4(.A(n7929), .B(n9481), .Y(n14796));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_sc1_64__U1(.A(n7931), .B(n14793), .Y(dpath_mulcore_ary1_a1_s0[64]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_sc1_64__U4(.A(n7930), .B(n8758), .Y(n14793));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_sc1_67__U1(.A(n7799), .B(n9480), .Y(dpath_mulcore_ary1_a1_s1[67]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_sc1_66__U1(.A(n7800), .B(dpath_mulcore_ary1_a1_I1_I2_net38), .Y(dpath_mulcore_ary1_a1_s1[66]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_sc1_65__U1(.A(n7801), .B(n14788), .Y(dpath_mulcore_ary1_a1_s1[65]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_sc1_65__U4(.A(n7802), .B(n9479), .Y(n14788));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_sc1_64__U1(.A(n7804), .B(n14785), .Y(dpath_mulcore_ary1_a1_s1[64]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_sc1_64__U4(.A(n7803), .B(n8757), .Y(n14785));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I2_sc1_67__U1(.A(dpath_mulcore_ary1_a1_I2_I2_p2_l_67), .B(n9478), .Y(dpath_mulcore_ary1_a1_s2[67]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I2_sc1_66__U1(.A(dpath_mulcore_ary1_a1_I2_I2_p2_l_66), .B(dpath_mulcore_ary1_a1_I2_I2_net38), .Y(dpath_mulcore_ary1_a1_s2[66]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I2_sc1_65__U1(.A(dpath_mulcore_ary1_a1_I2_I2_p2_l_65), .B(n14780), .Y(dpath_mulcore_ary1_a1_s2[65]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I2_sc1_65__U4(.A(n7735), .B(n9477), .Y(n14780));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I2_sc1_64__U1(.A(dpath_mulcore_ary1_a1_I2_I2_p2_l_64), .B(n14777), .Y(dpath_mulcore_ary1_a1_s2[64]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I2_sc1_64__U4(.A(n7736), .B(n8756), .Y(n14777));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_sc1_67__U1(.A(n7608), .B(n14774), .Y(dpath_mulcore_ary1_a0_s0[67]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_sc1_67__U4(.A(n9426), .B(dpath_mulcore_ary1_a0_I0_I2_sc1_66__b), .Y(n14774));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_sc1_66__U1(.A(n7609), .B(n14771), .Y(dpath_mulcore_ary1_a0_s0[66]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_sc1_66__U4(.A(n8053), .B(n9490), .Y(n14771));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_sc1_65__U1(.A(n7610), .B(n14768), .Y(dpath_mulcore_ary1_a0_s0[65]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_sc1_65__U4(.A(n7611), .B(dpath_mulcore_ary1_a0_I0_I2_net42), .Y(n14768));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_sc1_64__U1(.A(n7613), .B(n14765), .Y(dpath_mulcore_ary1_a0_s0[64]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_sc1_64__U4(.A(n7612), .B(n8755), .Y(n14765));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_U4(.A(n9217), .B(dpath_mulcore_cyc1), .Y(dpath_mulcore_ary1_a0_I0_I2_net42));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_4__sc1_U1(.A(n9829), .B(n14762), .Y(dpath_mulcore_ary1_a1_s0[4]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_4__sc1_U4(.A(n8050), .B(n8752), .Y(n14762));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_5__sc1_U1(.A(n8048), .B(n14759), .Y(dpath_mulcore_ary1_a1_s0[5]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_5__sc1_U4(.A(n8049), .B(n8751), .Y(n14759));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_6__sc1_U1(.A(n8046), .B(n14756), .Y(dpath_mulcore_ary1_a1_s0[6]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_6__sc1_U4(.A(n8047), .B(n8750), .Y(n14756));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_7__sc1_U1(.A(n8044), .B(n14753), .Y(dpath_mulcore_ary1_a1_s0[7]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_7__sc1_U4(.A(n8045), .B(n8749), .Y(n14753));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_8__sc1_U1(.A(n8042), .B(n14750), .Y(dpath_mulcore_ary1_a1_s0[8]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_8__sc1_U4(.A(n8043), .B(n8748), .Y(n14750));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_9__sc1_U1(.A(n8040), .B(n14747), .Y(dpath_mulcore_ary1_a1_s0[9]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_9__sc1_U4(.A(n8041), .B(n8747), .Y(n14747));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_10__sc1_U1(.A(n8038), .B(n14744), .Y(dpath_mulcore_ary1_a1_s0[10]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_10__sc1_U4(.A(n8039), .B(n8746), .Y(n14744));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_11__sc1_U1(.A(n8036), .B(n14741), .Y(dpath_mulcore_ary1_a1_s0[11]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_11__sc1_U4(.A(n8037), .B(n8745), .Y(n14741));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_12__sc1_U1(.A(n8034), .B(n14738), .Y(dpath_mulcore_ary1_a1_s0[12]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_12__sc1_U4(.A(n8035), .B(n8744), .Y(n14738));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_13__sc1_U1(.A(n8032), .B(n14735), .Y(dpath_mulcore_ary1_a1_s0[13]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_13__sc1_U4(.A(n8033), .B(n8743), .Y(n14735));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_14__sc1_U1(.A(n8030), .B(n14732), .Y(dpath_mulcore_ary1_a1_s0[14]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_14__sc1_U4(.A(n8031), .B(n8742), .Y(n14732));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_15__sc1_U1(.A(n8028), .B(n14729), .Y(dpath_mulcore_ary1_a1_s0[15]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_15__sc1_U4(.A(n8029), .B(n8741), .Y(n14729));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_16__sc1_U1(.A(n8026), .B(n14726), .Y(dpath_mulcore_ary1_a1_s0[16]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_16__sc1_U4(.A(n8027), .B(n8740), .Y(n14726));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_17__sc1_U1(.A(n8024), .B(n14723), .Y(dpath_mulcore_ary1_a1_s0[17]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_17__sc1_U4(.A(n8025), .B(n8739), .Y(n14723));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_18__sc1_U1(.A(n8022), .B(n14720), .Y(dpath_mulcore_ary1_a1_s0[18]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_18__sc1_U4(.A(n8023), .B(n8738), .Y(n14720));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_19__sc1_U1(.A(n8020), .B(n14717), .Y(dpath_mulcore_ary1_a1_s0[19]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_19__sc1_U4(.A(n8021), .B(n8737), .Y(n14717));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_20__sc1_U1(.A(n8018), .B(n14714), .Y(dpath_mulcore_ary1_a1_s0[20]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_20__sc1_U4(.A(n8019), .B(n8736), .Y(n14714));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_21__sc1_U1(.A(n8016), .B(n14711), .Y(dpath_mulcore_ary1_a1_s0[21]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_21__sc1_U4(.A(n8017), .B(n8735), .Y(n14711));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_22__sc1_U1(.A(n8014), .B(n14708), .Y(dpath_mulcore_ary1_a1_s0[22]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_22__sc1_U4(.A(n8015), .B(n8734), .Y(n14708));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_23__sc1_U1(.A(n8012), .B(n14705), .Y(dpath_mulcore_ary1_a1_s0[23]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_23__sc1_U4(.A(n8013), .B(n8733), .Y(n14705));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_24__sc1_U1(.A(n8010), .B(n14702), .Y(dpath_mulcore_ary1_a1_s0[24]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_24__sc1_U4(.A(n8011), .B(n8732), .Y(n14702));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_25__sc1_U1(.A(n8008), .B(n14699), .Y(dpath_mulcore_ary1_a1_s0[25]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_25__sc1_U4(.A(n8009), .B(n8731), .Y(n14699));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_26__sc1_U1(.A(n8006), .B(n14696), .Y(dpath_mulcore_ary1_a1_s0[26]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_26__sc1_U4(.A(n8007), .B(n8730), .Y(n14696));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_27__sc1_U1(.A(n8004), .B(n14693), .Y(dpath_mulcore_ary1_a1_s0[27]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_27__sc1_U4(.A(n8005), .B(n8729), .Y(n14693));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_28__sc1_U1(.A(n8002), .B(n14690), .Y(dpath_mulcore_ary1_a1_s0[28]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_28__sc1_U4(.A(n8003), .B(n8728), .Y(n14690));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_29__sc1_U1(.A(n8000), .B(n14687), .Y(dpath_mulcore_ary1_a1_s0[29]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_29__sc1_U4(.A(n8001), .B(n8727), .Y(n14687));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_30__sc1_U1(.A(n7998), .B(n14684), .Y(dpath_mulcore_ary1_a1_s0[30]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_30__sc1_U4(.A(n7999), .B(n8726), .Y(n14684));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_31__sc1_U1(.A(n7996), .B(n14681), .Y(dpath_mulcore_ary1_a1_s0[31]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_31__sc1_U4(.A(n7997), .B(n8725), .Y(n14681));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_32__sc1_U1(.A(n7994), .B(n14678), .Y(dpath_mulcore_ary1_a1_s0[32]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_32__sc1_U4(.A(n7995), .B(n8724), .Y(n14678));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_33__sc1_U1(.A(n7992), .B(n14675), .Y(dpath_mulcore_ary1_a1_s0[33]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_33__sc1_U4(.A(n7993), .B(n8723), .Y(n14675));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_34__sc1_U1(.A(n7990), .B(n14672), .Y(dpath_mulcore_ary1_a1_s0[34]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_34__sc1_U4(.A(n7991), .B(n8722), .Y(n14672));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_35__sc1_U1(.A(n7988), .B(n14669), .Y(dpath_mulcore_ary1_a1_s0[35]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_35__sc1_U4(.A(n7989), .B(n8721), .Y(n14669));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_36__sc1_U1(.A(n7986), .B(n14666), .Y(dpath_mulcore_ary1_a1_s0[36]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_36__sc1_U4(.A(n7987), .B(n8720), .Y(n14666));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_37__sc1_U1(.A(n7984), .B(n14663), .Y(dpath_mulcore_ary1_a1_s0[37]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_37__sc1_U4(.A(n7985), .B(n8719), .Y(n14663));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_38__sc1_U1(.A(n7982), .B(n14660), .Y(dpath_mulcore_ary1_a1_s0[38]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_38__sc1_U4(.A(n7983), .B(n8718), .Y(n14660));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_39__sc1_U1(.A(n7980), .B(n14657), .Y(dpath_mulcore_ary1_a1_s0[39]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_39__sc1_U4(.A(n7981), .B(n8717), .Y(n14657));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_40__sc1_U1(.A(n7978), .B(n14654), .Y(dpath_mulcore_ary1_a1_s0[40]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_40__sc1_U4(.A(n7979), .B(n8716), .Y(n14654));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_41__sc1_U1(.A(n7976), .B(n14651), .Y(dpath_mulcore_ary1_a1_s0[41]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_41__sc1_U4(.A(n7977), .B(n8715), .Y(n14651));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_42__sc1_U1(.A(n7974), .B(n14648), .Y(dpath_mulcore_ary1_a1_s0[42]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_42__sc1_U4(.A(n7975), .B(n8714), .Y(n14648));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_43__sc1_U1(.A(n7972), .B(n14645), .Y(dpath_mulcore_ary1_a1_s0[43]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_43__sc1_U4(.A(n7973), .B(n8713), .Y(n14645));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_44__sc1_U1(.A(n7970), .B(n14642), .Y(dpath_mulcore_ary1_a1_s0[44]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_44__sc1_U4(.A(n7971), .B(n8712), .Y(n14642));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_45__sc1_U1(.A(n7968), .B(n14639), .Y(dpath_mulcore_ary1_a1_s0[45]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_45__sc1_U4(.A(n7969), .B(n8711), .Y(n14639));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_46__sc1_U1(.A(n7966), .B(n14636), .Y(dpath_mulcore_ary1_a1_s0[46]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_46__sc1_U4(.A(n7967), .B(n8710), .Y(n14636));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_47__sc1_U1(.A(n7964), .B(n14633), .Y(dpath_mulcore_ary1_a1_s0[47]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_47__sc1_U4(.A(n7965), .B(n8709), .Y(n14633));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_48__sc1_U1(.A(n7962), .B(n14630), .Y(dpath_mulcore_ary1_a1_s0[48]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_48__sc1_U4(.A(n7963), .B(n8708), .Y(n14630));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_49__sc1_U1(.A(n7960), .B(n14627), .Y(dpath_mulcore_ary1_a1_s0[49]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_49__sc1_U4(.A(n7961), .B(n8707), .Y(n14627));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_50__sc1_U1(.A(n7958), .B(n14624), .Y(dpath_mulcore_ary1_a1_s0[50]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_50__sc1_U4(.A(n7959), .B(n8706), .Y(n14624));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_51__sc1_U1(.A(n7956), .B(n14621), .Y(dpath_mulcore_ary1_a1_s0[51]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_51__sc1_U4(.A(n7957), .B(n8705), .Y(n14621));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_52__sc1_U1(.A(n7954), .B(n14618), .Y(dpath_mulcore_ary1_a1_s0[52]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_52__sc1_U4(.A(n7955), .B(n8704), .Y(n14618));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_53__sc1_U1(.A(n7952), .B(n14615), .Y(dpath_mulcore_ary1_a1_s0[53]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_53__sc1_U4(.A(n7953), .B(n8703), .Y(n14615));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_54__sc1_U1(.A(n7950), .B(n14612), .Y(dpath_mulcore_ary1_a1_s0[54]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_54__sc1_U4(.A(n7951), .B(n8702), .Y(n14612));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_55__sc1_U1(.A(n7948), .B(n14609), .Y(dpath_mulcore_ary1_a1_s0[55]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_55__sc1_U4(.A(n7949), .B(n8701), .Y(n14609));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_56__sc1_U1(.A(n7946), .B(n14606), .Y(dpath_mulcore_ary1_a1_s0[56]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_56__sc1_U4(.A(n7947), .B(n8700), .Y(n14606));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_57__sc1_U1(.A(n7944), .B(n14603), .Y(dpath_mulcore_ary1_a1_s0[57]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_57__sc1_U4(.A(n7945), .B(n8699), .Y(n14603));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_58__sc1_U1(.A(n7942), .B(n14600), .Y(dpath_mulcore_ary1_a1_s0[58]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_58__sc1_U4(.A(n7943), .B(n8698), .Y(n14600));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_59__sc1_U1(.A(n7940), .B(n14597), .Y(dpath_mulcore_ary1_a1_s0[59]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_59__sc1_U4(.A(n7941), .B(n8697), .Y(n14597));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_60__sc1_U1(.A(n7938), .B(n14594), .Y(dpath_mulcore_ary1_a1_s0[60]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_60__sc1_U4(.A(n7939), .B(n8696), .Y(n14594));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_61__sc1_U1(.A(n7936), .B(n14591), .Y(dpath_mulcore_ary1_a1_s0[61]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_61__sc1_U4(.A(n7937), .B(n8695), .Y(n14591));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_62__sc1_U1(.A(n7934), .B(n14588), .Y(dpath_mulcore_ary1_a1_s0[62]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_62__sc1_U4(.A(n7935), .B(n8694), .Y(n14588));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_63__sc1_U1(.A(n7932), .B(n14585), .Y(dpath_mulcore_ary1_a1_s0[63]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_63__sc1_U4(.A(n7933), .B(n8693), .Y(n14585));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_4__sc1_U1(.A(n9835), .B(n14582), .Y(dpath_mulcore_ary1_a1_s1[4]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_4__sc1_U4(.A(n7923), .B(n8691), .Y(n14582));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_5__sc1_U1(.A(n7921), .B(n14579), .Y(dpath_mulcore_ary1_a1_s1[5]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_5__sc1_U4(.A(n7922), .B(n8690), .Y(n14579));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_6__sc1_U1(.A(n7919), .B(n14576), .Y(dpath_mulcore_ary1_a1_s1[6]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_6__sc1_U4(.A(n7920), .B(n8689), .Y(n14576));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_7__sc1_U1(.A(n7917), .B(n14573), .Y(dpath_mulcore_ary1_a1_s1[7]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_7__sc1_U4(.A(n7918), .B(n8688), .Y(n14573));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_8__sc1_U1(.A(n7915), .B(n14570), .Y(dpath_mulcore_ary1_a1_s1[8]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_8__sc1_U4(.A(n7916), .B(n8687), .Y(n14570));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_9__sc1_U1(.A(n7913), .B(n14567), .Y(dpath_mulcore_ary1_a1_s1[9]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_9__sc1_U4(.A(n7914), .B(n8686), .Y(n14567));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_10__sc1_U1(.A(n7911), .B(n14564), .Y(dpath_mulcore_ary1_a1_s1[10]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_10__sc1_U4(.A(n7912), .B(n8685), .Y(n14564));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_11__sc1_U1(.A(n7909), .B(n14561), .Y(dpath_mulcore_ary1_a1_s1[11]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_11__sc1_U4(.A(n7910), .B(n8684), .Y(n14561));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_12__sc1_U1(.A(n7907), .B(n14558), .Y(dpath_mulcore_ary1_a1_s1[12]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_12__sc1_U4(.A(n7908), .B(n8683), .Y(n14558));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_13__sc1_U1(.A(n7905), .B(n14555), .Y(dpath_mulcore_ary1_a1_s1[13]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_13__sc1_U4(.A(n7906), .B(n8682), .Y(n14555));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_14__sc1_U1(.A(n7903), .B(n14552), .Y(dpath_mulcore_ary1_a1_s1[14]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_14__sc1_U4(.A(n7904), .B(n8681), .Y(n14552));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_15__sc1_U1(.A(n7901), .B(n14549), .Y(dpath_mulcore_ary1_a1_s1[15]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_15__sc1_U4(.A(n7902), .B(n8680), .Y(n14549));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_16__sc1_U1(.A(n7899), .B(n14546), .Y(dpath_mulcore_ary1_a1_s1[16]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_16__sc1_U4(.A(n7900), .B(n8679), .Y(n14546));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_17__sc1_U1(.A(n7897), .B(n14543), .Y(dpath_mulcore_ary1_a1_s1[17]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_17__sc1_U4(.A(n7898), .B(n8678), .Y(n14543));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_18__sc1_U1(.A(n7895), .B(n14540), .Y(dpath_mulcore_ary1_a1_s1[18]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_18__sc1_U4(.A(n7896), .B(n8677), .Y(n14540));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_19__sc1_U1(.A(n7893), .B(n14537), .Y(dpath_mulcore_ary1_a1_s1[19]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_19__sc1_U4(.A(n7894), .B(n8676), .Y(n14537));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_20__sc1_U1(.A(n7891), .B(n14534), .Y(dpath_mulcore_ary1_a1_s1[20]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_20__sc1_U4(.A(n7892), .B(n8675), .Y(n14534));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_21__sc1_U1(.A(n7889), .B(n14531), .Y(dpath_mulcore_ary1_a1_s1[21]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_21__sc1_U4(.A(n7890), .B(n8674), .Y(n14531));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_22__sc1_U1(.A(n7887), .B(n14528), .Y(dpath_mulcore_ary1_a1_s1[22]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_22__sc1_U4(.A(n7888), .B(n8673), .Y(n14528));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_23__sc1_U1(.A(n7885), .B(n14525), .Y(dpath_mulcore_ary1_a1_s1[23]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_23__sc1_U4(.A(n7886), .B(n8672), .Y(n14525));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_24__sc1_U1(.A(n7883), .B(n14522), .Y(dpath_mulcore_ary1_a1_s1[24]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_24__sc1_U4(.A(n7884), .B(n8671), .Y(n14522));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_25__sc1_U1(.A(n7881), .B(n14519), .Y(dpath_mulcore_ary1_a1_s1[25]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_25__sc1_U4(.A(n7882), .B(n8670), .Y(n14519));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_26__sc1_U1(.A(n7879), .B(n14516), .Y(dpath_mulcore_ary1_a1_s1[26]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_26__sc1_U4(.A(n7880), .B(n8669), .Y(n14516));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_27__sc1_U1(.A(n7877), .B(n14513), .Y(dpath_mulcore_ary1_a1_s1[27]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_27__sc1_U4(.A(n7878), .B(n8668), .Y(n14513));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_28__sc1_U1(.A(n7875), .B(n14510), .Y(dpath_mulcore_ary1_a1_s1[28]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_28__sc1_U4(.A(n7876), .B(n8667), .Y(n14510));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_29__sc1_U1(.A(n7873), .B(n14507), .Y(dpath_mulcore_ary1_a1_s1[29]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_29__sc1_U4(.A(n7874), .B(n8666), .Y(n14507));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_30__sc1_U1(.A(n7871), .B(n14504), .Y(dpath_mulcore_ary1_a1_s1[30]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_30__sc1_U4(.A(n7872), .B(n8665), .Y(n14504));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_31__sc1_U1(.A(n7869), .B(n14501), .Y(dpath_mulcore_ary1_a1_s1[31]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_31__sc1_U4(.A(n7870), .B(n8664), .Y(n14501));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_32__sc1_U1(.A(n7867), .B(n14498), .Y(dpath_mulcore_ary1_a1_s1[32]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_32__sc1_U4(.A(n7868), .B(n8663), .Y(n14498));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_33__sc1_U1(.A(n7865), .B(n14495), .Y(dpath_mulcore_ary1_a1_s1[33]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_33__sc1_U4(.A(n7866), .B(n8662), .Y(n14495));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_34__sc1_U1(.A(n7863), .B(n14492), .Y(dpath_mulcore_ary1_a1_s1[34]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_34__sc1_U4(.A(n7864), .B(n8661), .Y(n14492));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_35__sc1_U1(.A(n7861), .B(n14489), .Y(dpath_mulcore_ary1_a1_s1[35]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_35__sc1_U4(.A(n7862), .B(n8660), .Y(n14489));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_36__sc1_U1(.A(n7859), .B(n14486), .Y(dpath_mulcore_ary1_a1_s1[36]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_36__sc1_U4(.A(n7860), .B(n8659), .Y(n14486));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_37__sc1_U1(.A(n7857), .B(n14483), .Y(dpath_mulcore_ary1_a1_s1[37]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_37__sc1_U4(.A(n7858), .B(n8658), .Y(n14483));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_38__sc1_U1(.A(n7855), .B(n14480), .Y(dpath_mulcore_ary1_a1_s1[38]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_38__sc1_U4(.A(n7856), .B(n8657), .Y(n14480));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_39__sc1_U1(.A(n7853), .B(n14477), .Y(dpath_mulcore_ary1_a1_s1[39]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_39__sc1_U4(.A(n7854), .B(n8656), .Y(n14477));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_40__sc1_U1(.A(n7851), .B(n14474), .Y(dpath_mulcore_ary1_a1_s1[40]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_40__sc1_U4(.A(n7852), .B(n8655), .Y(n14474));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_41__sc1_U1(.A(n7849), .B(n14471), .Y(dpath_mulcore_ary1_a1_s1[41]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_41__sc1_U4(.A(n7850), .B(n8654), .Y(n14471));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_42__sc1_U1(.A(n7847), .B(n14468), .Y(dpath_mulcore_ary1_a1_s1[42]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_42__sc1_U4(.A(n7848), .B(n8653), .Y(n14468));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_43__sc1_U1(.A(n7845), .B(n14465), .Y(dpath_mulcore_ary1_a1_s1[43]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_43__sc1_U4(.A(n7846), .B(n8652), .Y(n14465));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_44__sc1_U1(.A(n7843), .B(n14462), .Y(dpath_mulcore_ary1_a1_s1[44]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_44__sc1_U4(.A(n7844), .B(n8651), .Y(n14462));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_45__sc1_U1(.A(n7841), .B(n14459), .Y(dpath_mulcore_ary1_a1_s1[45]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_45__sc1_U4(.A(n7842), .B(n8650), .Y(n14459));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_46__sc1_U1(.A(n7839), .B(n14456), .Y(dpath_mulcore_ary1_a1_s1[46]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_46__sc1_U4(.A(n7840), .B(n8649), .Y(n14456));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_47__sc1_U1(.A(n7837), .B(n14453), .Y(dpath_mulcore_ary1_a1_s1[47]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_47__sc1_U4(.A(n7838), .B(n8648), .Y(n14453));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_48__sc1_U1(.A(n7835), .B(n14450), .Y(dpath_mulcore_ary1_a1_s1[48]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_48__sc1_U4(.A(n7836), .B(n8647), .Y(n14450));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_49__sc1_U1(.A(n7833), .B(n14447), .Y(dpath_mulcore_ary1_a1_s1[49]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_49__sc1_U4(.A(n7834), .B(n8646), .Y(n14447));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_50__sc1_U1(.A(n7831), .B(n14444), .Y(dpath_mulcore_ary1_a1_s1[50]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_50__sc1_U4(.A(n7832), .B(n8645), .Y(n14444));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_51__sc1_U1(.A(n7829), .B(n14441), .Y(dpath_mulcore_ary1_a1_s1[51]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_51__sc1_U4(.A(n7830), .B(n8644), .Y(n14441));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_52__sc1_U1(.A(n7827), .B(n14438), .Y(dpath_mulcore_ary1_a1_s1[52]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_52__sc1_U4(.A(n7828), .B(n8643), .Y(n14438));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_53__sc1_U1(.A(n7825), .B(n14435), .Y(dpath_mulcore_ary1_a1_s1[53]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_53__sc1_U4(.A(n7826), .B(n8642), .Y(n14435));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_54__sc1_U1(.A(n7823), .B(n14432), .Y(dpath_mulcore_ary1_a1_s1[54]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_54__sc1_U4(.A(n7824), .B(n8641), .Y(n14432));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_55__sc1_U1(.A(n7821), .B(n14429), .Y(dpath_mulcore_ary1_a1_s1[55]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_55__sc1_U4(.A(n7822), .B(n8640), .Y(n14429));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_56__sc1_U1(.A(n7819), .B(n14426), .Y(dpath_mulcore_ary1_a1_s1[56]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_56__sc1_U4(.A(n7820), .B(n8639), .Y(n14426));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_57__sc1_U1(.A(n7817), .B(n14423), .Y(dpath_mulcore_ary1_a1_s1[57]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_57__sc1_U4(.A(n7818), .B(n8638), .Y(n14423));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_58__sc1_U1(.A(n7815), .B(n14420), .Y(dpath_mulcore_ary1_a1_s1[58]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_58__sc1_U4(.A(n7816), .B(n8637), .Y(n14420));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_59__sc1_U1(.A(n7813), .B(n14417), .Y(dpath_mulcore_ary1_a1_s1[59]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_59__sc1_U4(.A(n7814), .B(n8636), .Y(n14417));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_60__sc1_U1(.A(n7811), .B(n14414), .Y(dpath_mulcore_ary1_a1_s1[60]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_60__sc1_U4(.A(n7812), .B(n8635), .Y(n14414));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_61__sc1_U1(.A(n7809), .B(n14411), .Y(dpath_mulcore_ary1_a1_s1[61]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_61__sc1_U4(.A(n7810), .B(n8634), .Y(n14411));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_62__sc1_U1(.A(n7807), .B(n14408), .Y(dpath_mulcore_ary1_a1_s1[62]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_62__sc1_U4(.A(n7808), .B(n8633), .Y(n14408));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_63__sc1_U1(.A(n7805), .B(n14405), .Y(dpath_mulcore_ary1_a1_s1[63]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_63__sc1_U4(.A(n7806), .B(n8632), .Y(n14405));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_4__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[4]), .B(n14402), .Y(dpath_mulcore_ary1_a1_s2[4]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_4__sc1_U4(.A(n7796), .B(n8630), .Y(n14402));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_5__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[5]), .B(n14399), .Y(dpath_mulcore_ary1_a1_s2[5]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_5__sc1_U4(.A(n7795), .B(n8629), .Y(n14399));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_6__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[6]), .B(n14396), .Y(dpath_mulcore_ary1_a1_s2[6]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_6__sc1_U4(.A(n7794), .B(n8628), .Y(n14396));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_7__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[7]), .B(n14393), .Y(dpath_mulcore_ary1_a1_s2[7]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_7__sc1_U4(.A(n7793), .B(n8627), .Y(n14393));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_8__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[8]), .B(n14390), .Y(dpath_mulcore_ary1_a1_s2[8]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_8__sc1_U4(.A(n7792), .B(n8626), .Y(n14390));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_9__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[9]), .B(n14387), .Y(dpath_mulcore_ary1_a1_s2[9]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_9__sc1_U4(.A(n7791), .B(n8625), .Y(n14387));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_10__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[10]), .B(n14384), .Y(dpath_mulcore_ary1_a1_s2[10]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_10__sc1_U4(.A(n7790), .B(n8624), .Y(n14384));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_11__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[11]), .B(n14381), .Y(dpath_mulcore_ary1_a1_s2[11]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_11__sc1_U4(.A(n7789), .B(n8623), .Y(n14381));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_12__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[12]), .B(n14378), .Y(dpath_mulcore_ary1_a1_s2[12]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_12__sc1_U4(.A(n7788), .B(n8622), .Y(n14378));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_13__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[13]), .B(n14375), .Y(dpath_mulcore_ary1_a1_s2[13]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_13__sc1_U4(.A(n7787), .B(n8621), .Y(n14375));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_14__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[14]), .B(n14372), .Y(dpath_mulcore_ary1_a1_s2[14]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_14__sc1_U4(.A(n7786), .B(n8620), .Y(n14372));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_15__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[15]), .B(n14369), .Y(dpath_mulcore_ary1_a1_s2[15]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_15__sc1_U4(.A(n7785), .B(n8619), .Y(n14369));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_16__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[16]), .B(n14366), .Y(dpath_mulcore_ary1_a1_s2[16]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_16__sc1_U4(.A(n7784), .B(n8618), .Y(n14366));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_17__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[17]), .B(n14363), .Y(dpath_mulcore_ary1_a1_s2[17]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_17__sc1_U4(.A(n7783), .B(n8617), .Y(n14363));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_18__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[18]), .B(n14360), .Y(dpath_mulcore_ary1_a1_s2[18]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_18__sc1_U4(.A(n7782), .B(n8616), .Y(n14360));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_19__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[19]), .B(n14357), .Y(dpath_mulcore_ary1_a1_s2[19]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_19__sc1_U4(.A(n7781), .B(n8615), .Y(n14357));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_20__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[20]), .B(n14354), .Y(dpath_mulcore_ary1_a1_s2[20]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_20__sc1_U4(.A(n7780), .B(n8614), .Y(n14354));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_21__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[21]), .B(n14351), .Y(dpath_mulcore_ary1_a1_s2[21]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_21__sc1_U4(.A(n7779), .B(n8613), .Y(n14351));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_22__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[22]), .B(n14348), .Y(dpath_mulcore_ary1_a1_s2[22]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_22__sc1_U4(.A(n7778), .B(n8612), .Y(n14348));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_23__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[23]), .B(n14345), .Y(dpath_mulcore_ary1_a1_s2[23]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_23__sc1_U4(.A(n7777), .B(n8611), .Y(n14345));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_24__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[24]), .B(n14342), .Y(dpath_mulcore_ary1_a1_s2[24]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_24__sc1_U4(.A(n7776), .B(n8610), .Y(n14342));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_25__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[25]), .B(n14339), .Y(dpath_mulcore_ary1_a1_s2[25]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_25__sc1_U4(.A(n7775), .B(n8609), .Y(n14339));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_26__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[26]), .B(n14336), .Y(dpath_mulcore_ary1_a1_s2[26]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_26__sc1_U4(.A(n7774), .B(n8608), .Y(n14336));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_27__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[27]), .B(n14333), .Y(dpath_mulcore_ary1_a1_s2[27]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_27__sc1_U4(.A(n7773), .B(n8607), .Y(n14333));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_28__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[28]), .B(n14330), .Y(dpath_mulcore_ary1_a1_s2[28]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_28__sc1_U4(.A(n7772), .B(n8606), .Y(n14330));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_29__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[29]), .B(n14327), .Y(dpath_mulcore_ary1_a1_s2[29]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_29__sc1_U4(.A(n7771), .B(n8605), .Y(n14327));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_30__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[30]), .B(n14324), .Y(dpath_mulcore_ary1_a1_s2[30]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_30__sc1_U4(.A(n7770), .B(n8604), .Y(n14324));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_31__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[31]), .B(n14321), .Y(dpath_mulcore_ary1_a1_s2[31]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_31__sc1_U4(.A(n7769), .B(n8603), .Y(n14321));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_32__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[32]), .B(n14318), .Y(dpath_mulcore_ary1_a1_s2[32]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_32__sc1_U4(.A(n7768), .B(n8602), .Y(n14318));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_33__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[33]), .B(n14315), .Y(dpath_mulcore_ary1_a1_s2[33]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_33__sc1_U4(.A(n7767), .B(n8601), .Y(n14315));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_34__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[34]), .B(n14312), .Y(dpath_mulcore_ary1_a1_s2[34]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_34__sc1_U4(.A(n7766), .B(n8600), .Y(n14312));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_35__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[35]), .B(n14309), .Y(dpath_mulcore_ary1_a1_s2[35]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_35__sc1_U4(.A(n7765), .B(n8599), .Y(n14309));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_36__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[36]), .B(n14306), .Y(dpath_mulcore_ary1_a1_s2[36]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_36__sc1_U4(.A(n7764), .B(n8598), .Y(n14306));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_37__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[37]), .B(n14303), .Y(dpath_mulcore_ary1_a1_s2[37]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_37__sc1_U4(.A(n7763), .B(n8597), .Y(n14303));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_38__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[38]), .B(n14300), .Y(dpath_mulcore_ary1_a1_s2[38]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_38__sc1_U4(.A(n7762), .B(n8596), .Y(n14300));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_39__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[39]), .B(n14297), .Y(dpath_mulcore_ary1_a1_s2[39]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_39__sc1_U4(.A(n7761), .B(n8595), .Y(n14297));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_40__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[40]), .B(n14294), .Y(dpath_mulcore_ary1_a1_s2[40]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_40__sc1_U4(.A(n7760), .B(n8594), .Y(n14294));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_41__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[41]), .B(n14291), .Y(dpath_mulcore_ary1_a1_s2[41]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_41__sc1_U4(.A(n7759), .B(n8593), .Y(n14291));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_42__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[42]), .B(n14288), .Y(dpath_mulcore_ary1_a1_s2[42]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_42__sc1_U4(.A(n7758), .B(n8592), .Y(n14288));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_43__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[43]), .B(n14285), .Y(dpath_mulcore_ary1_a1_s2[43]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_43__sc1_U4(.A(n7757), .B(n8591), .Y(n14285));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_44__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[44]), .B(n14282), .Y(dpath_mulcore_ary1_a1_s2[44]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_44__sc1_U4(.A(n7756), .B(n8590), .Y(n14282));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_45__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[45]), .B(n14279), .Y(dpath_mulcore_ary1_a1_s2[45]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_45__sc1_U4(.A(n7755), .B(n8589), .Y(n14279));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_46__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[46]), .B(n14276), .Y(dpath_mulcore_ary1_a1_s2[46]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_46__sc1_U4(.A(n7754), .B(n8588), .Y(n14276));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_47__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[47]), .B(n14273), .Y(dpath_mulcore_ary1_a1_s2[47]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_47__sc1_U4(.A(n7753), .B(n8587), .Y(n14273));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_48__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[48]), .B(n14270), .Y(dpath_mulcore_ary1_a1_s2[48]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_48__sc1_U4(.A(n7752), .B(n8586), .Y(n14270));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_49__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[49]), .B(n14267), .Y(dpath_mulcore_ary1_a1_s2[49]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_49__sc1_U4(.A(n7751), .B(n8585), .Y(n14267));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_50__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[50]), .B(n14264), .Y(dpath_mulcore_ary1_a1_s2[50]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_50__sc1_U4(.A(n7750), .B(n8584), .Y(n14264));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_51__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[51]), .B(n14261), .Y(dpath_mulcore_ary1_a1_s2[51]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_51__sc1_U4(.A(n7749), .B(n8583), .Y(n14261));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_52__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[52]), .B(n14258), .Y(dpath_mulcore_ary1_a1_s2[52]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_52__sc1_U4(.A(n7748), .B(n8582), .Y(n14258));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_53__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[53]), .B(n14255), .Y(dpath_mulcore_ary1_a1_s2[53]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_53__sc1_U4(.A(n7747), .B(n8581), .Y(n14255));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_54__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[54]), .B(n14252), .Y(dpath_mulcore_ary1_a1_s2[54]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_54__sc1_U4(.A(n7746), .B(n8580), .Y(n14252));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_55__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[55]), .B(n14249), .Y(dpath_mulcore_ary1_a1_s2[55]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_55__sc1_U4(.A(n7745), .B(n8579), .Y(n14249));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_56__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[56]), .B(n14246), .Y(dpath_mulcore_ary1_a1_s2[56]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_56__sc1_U4(.A(n7744), .B(n8578), .Y(n14246));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_57__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[57]), .B(n14243), .Y(dpath_mulcore_ary1_a1_s2[57]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_57__sc1_U4(.A(n7743), .B(n8577), .Y(n14243));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_58__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[58]), .B(n14240), .Y(dpath_mulcore_ary1_a1_s2[58]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_58__sc1_U4(.A(n7742), .B(n8576), .Y(n14240));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_59__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[59]), .B(n14237), .Y(dpath_mulcore_ary1_a1_s2[59]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_59__sc1_U4(.A(n7741), .B(n8575), .Y(n14237));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_60__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[60]), .B(n14234), .Y(dpath_mulcore_ary1_a1_s2[60]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_60__sc1_U4(.A(n7740), .B(n8574), .Y(n14234));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_61__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[61]), .B(n14231), .Y(dpath_mulcore_ary1_a1_s2[61]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_61__sc1_U4(.A(n7739), .B(n8573), .Y(n14231));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_62__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[62]), .B(n14228), .Y(dpath_mulcore_ary1_a1_s2[62]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_62__sc1_U4(.A(n7738), .B(n8572), .Y(n14228));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_63__sc1_U1(.A(dpath_mulcore_ary1_a1_I2_p2_l[63]), .B(n14225), .Y(dpath_mulcore_ary1_a1_s2[63]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_63__sc1_U4(.A(n7737), .B(n8571), .Y(n14225));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_4__sc1_U1(.A(n9842), .B(n14222), .Y(dpath_mulcore_ary1_a0_s0[4]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_4__sc1_U4(.A(n7732), .B(n8569), .Y(n14222));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_5__sc1_U1(.A(n7730), .B(n14219), .Y(dpath_mulcore_ary1_a0_s0[5]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_5__sc1_U4(.A(n7731), .B(n8568), .Y(n14219));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_6__sc1_U1(.A(n7728), .B(n14216), .Y(dpath_mulcore_ary1_a0_s0[6]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_6__sc1_U4(.A(n7729), .B(n8567), .Y(n14216));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_7__sc1_U1(.A(n7726), .B(n14213), .Y(dpath_mulcore_ary1_a0_s0[7]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_7__sc1_U4(.A(n7727), .B(n8566), .Y(n14213));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_8__sc1_U1(.A(n7724), .B(n14210), .Y(dpath_mulcore_ary1_a0_s0[8]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_8__sc1_U4(.A(n7725), .B(n8565), .Y(n14210));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_9__sc1_U1(.A(n7722), .B(n14207), .Y(dpath_mulcore_ary1_a0_s0[9]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_9__sc1_U4(.A(n7723), .B(n8564), .Y(n14207));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_10__sc1_U1(.A(n7720), .B(n14204), .Y(dpath_mulcore_ary1_a0_s0[10]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_10__sc1_U4(.A(n7721), .B(n8563), .Y(n14204));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_11__sc1_U1(.A(n7718), .B(n14201), .Y(dpath_mulcore_ary1_a0_s0[11]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_11__sc1_U4(.A(n7719), .B(n8562), .Y(n14201));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_12__sc1_U1(.A(n7716), .B(n14198), .Y(dpath_mulcore_ary1_a0_s0[12]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_12__sc1_U4(.A(n7717), .B(n8561), .Y(n14198));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_13__sc1_U1(.A(n7714), .B(n14195), .Y(dpath_mulcore_ary1_a0_s0[13]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_13__sc1_U4(.A(n7715), .B(n8560), .Y(n14195));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_14__sc1_U1(.A(n7712), .B(n14192), .Y(dpath_mulcore_ary1_a0_s0[14]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_14__sc1_U4(.A(n7713), .B(n8559), .Y(n14192));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_15__sc1_U1(.A(n7710), .B(n14189), .Y(dpath_mulcore_ary1_a0_s0[15]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_15__sc1_U4(.A(n7711), .B(n8558), .Y(n14189));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_16__sc1_U1(.A(n7708), .B(n14186), .Y(dpath_mulcore_ary1_a0_s0[16]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_16__sc1_U4(.A(n7709), .B(n8557), .Y(n14186));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_17__sc1_U1(.A(n7706), .B(n14183), .Y(dpath_mulcore_ary1_a0_s0[17]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_17__sc1_U4(.A(n7707), .B(n8556), .Y(n14183));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_18__sc1_U1(.A(n7704), .B(n14180), .Y(dpath_mulcore_ary1_a0_s0[18]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_18__sc1_U4(.A(n7705), .B(n8555), .Y(n14180));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_19__sc1_U1(.A(n7702), .B(n14177), .Y(dpath_mulcore_ary1_a0_s0[19]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_19__sc1_U4(.A(n7703), .B(n8554), .Y(n14177));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_20__sc1_U1(.A(n7700), .B(n14174), .Y(dpath_mulcore_ary1_a0_s0[20]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_20__sc1_U4(.A(n7701), .B(n8553), .Y(n14174));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_21__sc1_U1(.A(n7698), .B(n14171), .Y(dpath_mulcore_ary1_a0_s0[21]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_21__sc1_U4(.A(n7699), .B(n8552), .Y(n14171));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_22__sc1_U1(.A(n7696), .B(n14168), .Y(dpath_mulcore_ary1_a0_s0[22]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_22__sc1_U4(.A(n7697), .B(n8551), .Y(n14168));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_23__sc1_U1(.A(n7694), .B(n14165), .Y(dpath_mulcore_ary1_a0_s0[23]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_23__sc1_U4(.A(n7695), .B(n8550), .Y(n14165));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_24__sc1_U1(.A(n7692), .B(n14162), .Y(dpath_mulcore_ary1_a0_s0[24]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_24__sc1_U4(.A(n7693), .B(n8549), .Y(n14162));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_25__sc1_U1(.A(n7690), .B(n14159), .Y(dpath_mulcore_ary1_a0_s0[25]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_25__sc1_U4(.A(n7691), .B(n8548), .Y(n14159));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_26__sc1_U1(.A(n7688), .B(n14156), .Y(dpath_mulcore_ary1_a0_s0[26]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_26__sc1_U4(.A(n7689), .B(n8547), .Y(n14156));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_27__sc1_U1(.A(n7686), .B(n14153), .Y(dpath_mulcore_ary1_a0_s0[27]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_27__sc1_U4(.A(n7687), .B(n8546), .Y(n14153));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_28__sc1_U1(.A(n7684), .B(n14150), .Y(dpath_mulcore_ary1_a0_s0[28]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_28__sc1_U4(.A(n7685), .B(n8545), .Y(n14150));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_29__sc1_U1(.A(n7682), .B(n14147), .Y(dpath_mulcore_ary1_a0_s0[29]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_29__sc1_U4(.A(n7683), .B(n8544), .Y(n14147));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_30__sc1_U1(.A(n7680), .B(n14144), .Y(dpath_mulcore_ary1_a0_s0[30]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_30__sc1_U4(.A(n7681), .B(n8543), .Y(n14144));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_31__sc1_U1(.A(n7678), .B(n14141), .Y(dpath_mulcore_ary1_a0_s0[31]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_31__sc1_U4(.A(n7679), .B(n8542), .Y(n14141));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_32__sc1_U1(.A(n7676), .B(n14138), .Y(dpath_mulcore_ary1_a0_s0[32]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_32__sc1_U4(.A(n7677), .B(n8541), .Y(n14138));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_33__sc1_U1(.A(n7674), .B(n14135), .Y(dpath_mulcore_ary1_a0_s0[33]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_33__sc1_U4(.A(n7675), .B(n8540), .Y(n14135));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_34__sc1_U1(.A(n7672), .B(n14132), .Y(dpath_mulcore_ary1_a0_s0[34]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_34__sc1_U4(.A(n7673), .B(n8539), .Y(n14132));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_35__sc1_U1(.A(n7670), .B(n14129), .Y(dpath_mulcore_ary1_a0_s0[35]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_35__sc1_U4(.A(n7671), .B(n8538), .Y(n14129));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_36__sc1_U1(.A(n7668), .B(n14126), .Y(dpath_mulcore_ary1_a0_s0[36]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_36__sc1_U4(.A(n7669), .B(n8537), .Y(n14126));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_37__sc1_U1(.A(n7666), .B(n14123), .Y(dpath_mulcore_ary1_a0_s0[37]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_37__sc1_U4(.A(n7667), .B(n8536), .Y(n14123));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_38__sc1_U1(.A(n7664), .B(n14120), .Y(dpath_mulcore_ary1_a0_s0[38]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_38__sc1_U4(.A(n7665), .B(n8535), .Y(n14120));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_39__sc1_U1(.A(n7662), .B(n14117), .Y(dpath_mulcore_ary1_a0_s0[39]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_39__sc1_U4(.A(n7663), .B(n8534), .Y(n14117));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_40__sc1_U1(.A(n7660), .B(n14114), .Y(dpath_mulcore_ary1_a0_s0[40]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_40__sc1_U4(.A(n7661), .B(n8533), .Y(n14114));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_41__sc1_U1(.A(n7658), .B(n14111), .Y(dpath_mulcore_ary1_a0_s0[41]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_41__sc1_U4(.A(n7659), .B(n8532), .Y(n14111));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_42__sc1_U1(.A(n7656), .B(n14108), .Y(dpath_mulcore_ary1_a0_s0[42]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_42__sc1_U4(.A(n7657), .B(n8531), .Y(n14108));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_43__sc1_U1(.A(n7654), .B(n14105), .Y(dpath_mulcore_ary1_a0_s0[43]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_43__sc1_U4(.A(n7655), .B(n8530), .Y(n14105));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_44__sc1_U1(.A(n7652), .B(n14102), .Y(dpath_mulcore_ary1_a0_s0[44]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_44__sc1_U4(.A(n7653), .B(n8529), .Y(n14102));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_45__sc1_U1(.A(n7650), .B(n14099), .Y(dpath_mulcore_ary1_a0_s0[45]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_45__sc1_U4(.A(n7651), .B(n8528), .Y(n14099));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_46__sc1_U1(.A(n7648), .B(n14096), .Y(dpath_mulcore_ary1_a0_s0[46]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_46__sc1_U4(.A(n7649), .B(n8527), .Y(n14096));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_47__sc1_U1(.A(n7646), .B(n14093), .Y(dpath_mulcore_ary1_a0_s0[47]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_47__sc1_U4(.A(n7647), .B(n8526), .Y(n14093));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_48__sc1_U1(.A(n7644), .B(n14090), .Y(dpath_mulcore_ary1_a0_s0[48]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_48__sc1_U4(.A(n7645), .B(n8525), .Y(n14090));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_49__sc1_U1(.A(n7642), .B(n14087), .Y(dpath_mulcore_ary1_a0_s0[49]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_49__sc1_U4(.A(n7643), .B(n8524), .Y(n14087));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_50__sc1_U1(.A(n7640), .B(n14084), .Y(dpath_mulcore_ary1_a0_s0[50]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_50__sc1_U4(.A(n7641), .B(n8523), .Y(n14084));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_51__sc1_U1(.A(n7638), .B(n14081), .Y(dpath_mulcore_ary1_a0_s0[51]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_51__sc1_U4(.A(n7639), .B(n8522), .Y(n14081));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_52__sc1_U1(.A(n7636), .B(n14078), .Y(dpath_mulcore_ary1_a0_s0[52]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_52__sc1_U4(.A(n7637), .B(n8521), .Y(n14078));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_53__sc1_U1(.A(n7634), .B(n14075), .Y(dpath_mulcore_ary1_a0_s0[53]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_53__sc1_U4(.A(n7635), .B(n8520), .Y(n14075));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_54__sc1_U1(.A(n7632), .B(n14072), .Y(dpath_mulcore_ary1_a0_s0[54]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_54__sc1_U4(.A(n7633), .B(n8519), .Y(n14072));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_55__sc1_U1(.A(n7630), .B(n14069), .Y(dpath_mulcore_ary1_a0_s0[55]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_55__sc1_U4(.A(n7631), .B(n8518), .Y(n14069));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_56__sc1_U1(.A(n7628), .B(n14066), .Y(dpath_mulcore_ary1_a0_s0[56]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_56__sc1_U4(.A(n7629), .B(n8517), .Y(n14066));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_57__sc1_U1(.A(n7626), .B(n14063), .Y(dpath_mulcore_ary1_a0_s0[57]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_57__sc1_U4(.A(n7627), .B(n8516), .Y(n14063));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_58__sc1_U1(.A(n7624), .B(n14060), .Y(dpath_mulcore_ary1_a0_s0[58]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_58__sc1_U4(.A(n7625), .B(n8515), .Y(n14060));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_59__sc1_U1(.A(n7622), .B(n14057), .Y(dpath_mulcore_ary1_a0_s0[59]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_59__sc1_U4(.A(n7623), .B(n8514), .Y(n14057));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_60__sc1_U1(.A(n7620), .B(n14054), .Y(dpath_mulcore_ary1_a0_s0[60]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_60__sc1_U4(.A(n7621), .B(n8513), .Y(n14054));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_61__sc1_U1(.A(n7618), .B(n14051), .Y(dpath_mulcore_ary1_a0_s0[61]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_61__sc1_U4(.A(n7619), .B(n8512), .Y(n14051));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_62__sc1_U1(.A(n7616), .B(n14048), .Y(dpath_mulcore_ary1_a0_s0[62]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_62__sc1_U4(.A(n7617), .B(n8511), .Y(n14048));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_63__sc1_U1(.A(n7614), .B(n14045), .Y(dpath_mulcore_ary1_a0_s0[63]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_63__sc1_U4(.A(n7615), .B(n8510), .Y(n14045));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_4__sc1_U1(.A(n9848), .B(n14042), .Y(dpath_mulcore_ary1_a0_s1[4]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_4__sc1_U4(.A(n7605), .B(n8508), .Y(n14042));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_5__sc1_U1(.A(n7603), .B(n14039), .Y(dpath_mulcore_ary1_a0_s1[5]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_5__sc1_U4(.A(n7604), .B(n8507), .Y(n14039));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_6__sc1_U1(.A(n7601), .B(n14036), .Y(dpath_mulcore_ary1_a0_s1[6]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_6__sc1_U4(.A(n7602), .B(n8506), .Y(n14036));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_7__sc1_U1(.A(n7599), .B(n14033), .Y(dpath_mulcore_ary1_a0_s1[7]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_7__sc1_U4(.A(n7600), .B(n8505), .Y(n14033));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_8__sc1_U1(.A(n7597), .B(n14030), .Y(dpath_mulcore_ary1_a0_s1[8]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_8__sc1_U4(.A(n7598), .B(n8504), .Y(n14030));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_9__sc1_U1(.A(n7595), .B(n14027), .Y(dpath_mulcore_ary1_a0_s1[9]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_9__sc1_U4(.A(n7596), .B(n8503), .Y(n14027));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_10__sc1_U1(.A(n7593), .B(n14024), .Y(dpath_mulcore_ary1_a0_s1[10]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_10__sc1_U4(.A(n7594), .B(n8502), .Y(n14024));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_11__sc1_U1(.A(n7591), .B(n14021), .Y(dpath_mulcore_ary1_a0_s1[11]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_11__sc1_U4(.A(n7592), .B(n8501), .Y(n14021));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_12__sc1_U1(.A(n7589), .B(n14018), .Y(dpath_mulcore_ary1_a0_s1[12]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_12__sc1_U4(.A(n7590), .B(n8500), .Y(n14018));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_13__sc1_U1(.A(n7587), .B(n14015), .Y(dpath_mulcore_ary1_a0_s1[13]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_13__sc1_U4(.A(n7588), .B(n8499), .Y(n14015));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_14__sc1_U1(.A(n7585), .B(n14012), .Y(dpath_mulcore_ary1_a0_s1[14]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_14__sc1_U4(.A(n7586), .B(n8498), .Y(n14012));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_15__sc1_U1(.A(n7583), .B(n14009), .Y(dpath_mulcore_ary1_a0_s1[15]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_15__sc1_U4(.A(n7584), .B(n8497), .Y(n14009));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_16__sc1_U1(.A(n7581), .B(n14006), .Y(dpath_mulcore_ary1_a0_s1[16]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_16__sc1_U4(.A(n7582), .B(n8496), .Y(n14006));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_17__sc1_U1(.A(n7579), .B(n14003), .Y(dpath_mulcore_ary1_a0_s1[17]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_17__sc1_U4(.A(n7580), .B(n8495), .Y(n14003));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_18__sc1_U1(.A(n7577), .B(n14000), .Y(dpath_mulcore_ary1_a0_s1[18]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_18__sc1_U4(.A(n7578), .B(n8494), .Y(n14000));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_19__sc1_U1(.A(n7575), .B(n13997), .Y(dpath_mulcore_ary1_a0_s1[19]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_19__sc1_U4(.A(n7576), .B(n8493), .Y(n13997));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_20__sc1_U1(.A(n7573), .B(n13994), .Y(dpath_mulcore_ary1_a0_s1[20]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_20__sc1_U4(.A(n7574), .B(n8492), .Y(n13994));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_21__sc1_U1(.A(n7571), .B(n13991), .Y(dpath_mulcore_ary1_a0_s1[21]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_21__sc1_U4(.A(n7572), .B(n8491), .Y(n13991));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_22__sc1_U1(.A(n7569), .B(n13988), .Y(dpath_mulcore_ary1_a0_s1[22]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_22__sc1_U4(.A(n7570), .B(n8490), .Y(n13988));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_23__sc1_U1(.A(n7567), .B(n13985), .Y(dpath_mulcore_ary1_a0_s1[23]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_23__sc1_U4(.A(n7568), .B(n8489), .Y(n13985));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_24__sc1_U1(.A(n7565), .B(n13982), .Y(dpath_mulcore_ary1_a0_s1[24]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_24__sc1_U4(.A(n7566), .B(n8488), .Y(n13982));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_25__sc1_U1(.A(n7563), .B(n13979), .Y(dpath_mulcore_ary1_a0_s1[25]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_25__sc1_U4(.A(n7564), .B(n8487), .Y(n13979));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_26__sc1_U1(.A(n7561), .B(n13976), .Y(dpath_mulcore_ary1_a0_s1[26]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_26__sc1_U4(.A(n7562), .B(n8486), .Y(n13976));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_27__sc1_U1(.A(n7559), .B(n13973), .Y(dpath_mulcore_ary1_a0_s1[27]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_27__sc1_U4(.A(n7560), .B(n8485), .Y(n13973));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_28__sc1_U1(.A(n7557), .B(n13970), .Y(dpath_mulcore_ary1_a0_s1[28]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_28__sc1_U4(.A(n7558), .B(n8484), .Y(n13970));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_29__sc1_U1(.A(n7555), .B(n13967), .Y(dpath_mulcore_ary1_a0_s1[29]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_29__sc1_U4(.A(n7556), .B(n8483), .Y(n13967));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_30__sc1_U1(.A(n7553), .B(n13964), .Y(dpath_mulcore_ary1_a0_s1[30]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_30__sc1_U4(.A(n7554), .B(n8482), .Y(n13964));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_31__sc1_U1(.A(n7551), .B(n13961), .Y(dpath_mulcore_ary1_a0_s1[31]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_31__sc1_U4(.A(n7552), .B(n8481), .Y(n13961));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_32__sc1_U1(.A(n7549), .B(n13958), .Y(dpath_mulcore_ary1_a0_s1[32]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_32__sc1_U4(.A(n7550), .B(n8480), .Y(n13958));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_33__sc1_U1(.A(n7547), .B(n13955), .Y(dpath_mulcore_ary1_a0_s1[33]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_33__sc1_U4(.A(n7548), .B(n8479), .Y(n13955));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_34__sc1_U1(.A(n7545), .B(n13952), .Y(dpath_mulcore_ary1_a0_s1[34]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_34__sc1_U4(.A(n7546), .B(n8478), .Y(n13952));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_35__sc1_U1(.A(n7543), .B(n13949), .Y(dpath_mulcore_ary1_a0_s1[35]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_35__sc1_U4(.A(n7544), .B(n8477), .Y(n13949));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_36__sc1_U1(.A(n7541), .B(n13946), .Y(dpath_mulcore_ary1_a0_s1[36]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_36__sc1_U4(.A(n7542), .B(n8476), .Y(n13946));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_37__sc1_U1(.A(n7539), .B(n13943), .Y(dpath_mulcore_ary1_a0_s1[37]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_37__sc1_U4(.A(n7540), .B(n8475), .Y(n13943));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_38__sc1_U1(.A(n7537), .B(n13940), .Y(dpath_mulcore_ary1_a0_s1[38]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_38__sc1_U4(.A(n7538), .B(n8474), .Y(n13940));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_39__sc1_U1(.A(n7535), .B(n13937), .Y(dpath_mulcore_ary1_a0_s1[39]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_39__sc1_U4(.A(n7536), .B(n8473), .Y(n13937));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_40__sc1_U1(.A(n7533), .B(n13934), .Y(dpath_mulcore_ary1_a0_s1[40]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_40__sc1_U4(.A(n7534), .B(n8472), .Y(n13934));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_41__sc1_U1(.A(n7531), .B(n13931), .Y(dpath_mulcore_ary1_a0_s1[41]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_41__sc1_U4(.A(n7532), .B(n8471), .Y(n13931));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_42__sc1_U1(.A(n7529), .B(n13928), .Y(dpath_mulcore_ary1_a0_s1[42]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_42__sc1_U4(.A(n7530), .B(n8470), .Y(n13928));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_43__sc1_U1(.A(n7527), .B(n13925), .Y(dpath_mulcore_ary1_a0_s1[43]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_43__sc1_U4(.A(n7528), .B(n8469), .Y(n13925));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_44__sc1_U1(.A(n7525), .B(n13922), .Y(dpath_mulcore_ary1_a0_s1[44]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_44__sc1_U4(.A(n7526), .B(n8468), .Y(n13922));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_45__sc1_U1(.A(n7523), .B(n13919), .Y(dpath_mulcore_ary1_a0_s1[45]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_45__sc1_U4(.A(n7524), .B(n8467), .Y(n13919));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_46__sc1_U1(.A(n7521), .B(n13916), .Y(dpath_mulcore_ary1_a0_s1[46]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_46__sc1_U4(.A(n7522), .B(n8466), .Y(n13916));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_47__sc1_U1(.A(n7519), .B(n13913), .Y(dpath_mulcore_ary1_a0_s1[47]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_47__sc1_U4(.A(n7520), .B(n8465), .Y(n13913));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_48__sc1_U1(.A(n7517), .B(n13910), .Y(dpath_mulcore_ary1_a0_s1[48]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_48__sc1_U4(.A(n7518), .B(n8464), .Y(n13910));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_49__sc1_U1(.A(n7515), .B(n13907), .Y(dpath_mulcore_ary1_a0_s1[49]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_49__sc1_U4(.A(n7516), .B(n8463), .Y(n13907));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_50__sc1_U1(.A(n7513), .B(n13904), .Y(dpath_mulcore_ary1_a0_s1[50]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_50__sc1_U4(.A(n7514), .B(n8462), .Y(n13904));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_51__sc1_U1(.A(n7511), .B(n13901), .Y(dpath_mulcore_ary1_a0_s1[51]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_51__sc1_U4(.A(n7512), .B(n8461), .Y(n13901));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_52__sc1_U1(.A(n7509), .B(n13898), .Y(dpath_mulcore_ary1_a0_s1[52]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_52__sc1_U4(.A(n7510), .B(n8460), .Y(n13898));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_53__sc1_U1(.A(n7507), .B(n13895), .Y(dpath_mulcore_ary1_a0_s1[53]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_53__sc1_U4(.A(n7508), .B(n8459), .Y(n13895));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_54__sc1_U1(.A(n7505), .B(n13892), .Y(dpath_mulcore_ary1_a0_s1[54]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_54__sc1_U4(.A(n7506), .B(n8458), .Y(n13892));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_55__sc1_U1(.A(n7503), .B(n13889), .Y(dpath_mulcore_ary1_a0_s1[55]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_55__sc1_U4(.A(n7504), .B(n8457), .Y(n13889));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_56__sc1_U1(.A(n7501), .B(n13886), .Y(dpath_mulcore_ary1_a0_s1[56]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_56__sc1_U4(.A(n7502), .B(n8456), .Y(n13886));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_57__sc1_U1(.A(n7499), .B(n13883), .Y(dpath_mulcore_ary1_a0_s1[57]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_57__sc1_U4(.A(n7500), .B(n8455), .Y(n13883));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_58__sc1_U1(.A(n7497), .B(n13880), .Y(dpath_mulcore_ary1_a0_s1[58]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_58__sc1_U4(.A(n7498), .B(n8454), .Y(n13880));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_59__sc1_U1(.A(n7495), .B(n13877), .Y(dpath_mulcore_ary1_a0_s1[59]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_59__sc1_U4(.A(n7496), .B(n8453), .Y(n13877));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_60__sc1_U1(.A(n7493), .B(n13874), .Y(dpath_mulcore_ary1_a0_s1[60]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_60__sc1_U4(.A(n7494), .B(n8452), .Y(n13874));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_61__sc1_U1(.A(n7491), .B(n13871), .Y(dpath_mulcore_ary1_a0_s1[61]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_61__sc1_U4(.A(n7492), .B(n8451), .Y(n13871));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_62__sc1_U1(.A(n7489), .B(n13868), .Y(dpath_mulcore_ary1_a0_s1[62]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_62__sc1_U4(.A(n7490), .B(n8450), .Y(n13868));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_63__sc1_U1(.A(n7487), .B(n13865), .Y(dpath_mulcore_ary1_a0_s1[63]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_63__sc1_U4(.A(n7488), .B(n8449), .Y(n13865));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_4__sc1_U4(.A(n7478), .B(n8447), .Y(n13862));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_5__sc1_U4(.A(n7477), .B(n8446), .Y(n13860));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_6__sc1_U4(.A(n7476), .B(n8445), .Y(n13858));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_7__sc1_U4(.A(n7475), .B(n8444), .Y(n13856));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_8__sc1_U4(.A(n7474), .B(n8443), .Y(n13854));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_9__sc1_U4(.A(n7473), .B(n8442), .Y(n13852));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_10__sc1_U4(.A(n7472), .B(n8441), .Y(n13850));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_11__sc1_U4(.A(n7471), .B(n8440), .Y(n13848));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_12__sc1_U4(.A(n7470), .B(n8439), .Y(n13846));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_13__sc1_U4(.A(n7469), .B(n8438), .Y(n13844));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_14__sc1_U4(.A(n7468), .B(n8437), .Y(n13842));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_15__sc1_U4(.A(n7467), .B(n8436), .Y(n13840));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_16__sc1_U4(.A(n7466), .B(n8435), .Y(n13838));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_17__sc1_U4(.A(n7465), .B(n8434), .Y(n13836));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_18__sc1_U4(.A(n7464), .B(n8433), .Y(n13834));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_19__sc1_U4(.A(n7463), .B(n8432), .Y(n13832));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_20__sc1_U4(.A(n7462), .B(n8431), .Y(n13830));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_21__sc1_U4(.A(n7461), .B(n8430), .Y(n13828));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_22__sc1_U4(.A(n7460), .B(n8429), .Y(n13826));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_23__sc1_U4(.A(n7459), .B(n8428), .Y(n13824));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_24__sc1_U4(.A(n7458), .B(n8427), .Y(n13822));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_25__sc1_U4(.A(n7457), .B(n8426), .Y(n13820));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_26__sc1_U4(.A(n7456), .B(n8425), .Y(n13818));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_27__sc1_U4(.A(n7455), .B(n8424), .Y(n13816));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_28__sc1_U4(.A(n7454), .B(n8423), .Y(n13814));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_29__sc1_U4(.A(n7453), .B(n8422), .Y(n13812));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_30__sc1_U4(.A(n7452), .B(n8421), .Y(n13810));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_31__sc1_U4(.A(n7451), .B(n8420), .Y(n13808));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_32__sc1_U4(.A(n7450), .B(n8419), .Y(n13806));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_33__sc1_U4(.A(n7449), .B(n8418), .Y(n13804));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_34__sc1_U4(.A(n7448), .B(n8417), .Y(n13802));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_35__sc1_U4(.A(n7447), .B(n8416), .Y(n13800));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_36__sc1_U4(.A(n7446), .B(n8415), .Y(n13798));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_37__sc1_U4(.A(n7445), .B(n8414), .Y(n13796));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_38__sc1_U4(.A(n7444), .B(n8413), .Y(n13794));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_39__sc1_U4(.A(n7443), .B(n8412), .Y(n13792));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_40__sc1_U4(.A(n7442), .B(n8411), .Y(n13790));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_41__sc1_U4(.A(n7441), .B(n8410), .Y(n13788));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_42__sc1_U4(.A(n7440), .B(n8409), .Y(n13786));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_43__sc1_U4(.A(n7439), .B(n8408), .Y(n13784));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_44__sc1_U4(.A(n7438), .B(n8407), .Y(n13782));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_45__sc1_U4(.A(n7437), .B(n8406), .Y(n13780));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_46__sc1_U4(.A(n7436), .B(n8405), .Y(n13778));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_47__sc1_U4(.A(n7435), .B(n8404), .Y(n13776));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_48__sc1_U4(.A(n7434), .B(n8403), .Y(n13774));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_49__sc1_U4(.A(n7433), .B(n8402), .Y(n13772));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_50__sc1_U4(.A(n7432), .B(n8401), .Y(n13770));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_51__sc1_U4(.A(n7431), .B(n8400), .Y(n13768));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_52__sc1_U4(.A(n7430), .B(n8399), .Y(n13766));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_53__sc1_U4(.A(n7429), .B(n8398), .Y(n13764));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_54__sc1_U4(.A(n7428), .B(n8397), .Y(n13762));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_55__sc1_U4(.A(n7427), .B(n8396), .Y(n13760));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_56__sc1_U4(.A(n7426), .B(n8395), .Y(n13758));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_57__sc1_U4(.A(n7425), .B(n8394), .Y(n13756));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_58__sc1_U4(.A(n7424), .B(n8393), .Y(n13754));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_59__sc1_U4(.A(n7423), .B(n8392), .Y(n13752));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_60__sc1_U4(.A(n7422), .B(n8391), .Y(n13750));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_61__sc1_U4(.A(n7421), .B(n8390), .Y(n13748));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_62__sc1_U4(.A(n7420), .B(n8389), .Y(n13746));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_sc1_1__U2(.A(dpath_mulcore_ary1_a1_I0_I0_b0n), .B(n7401), .Y(dpath_mulcore_a1sum[1]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_sc1_2__U1(.A(n8066), .B(n13744), .Y(dpath_mulcore_ary1_a1_s0[2]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_sc1_2__U4(.A(n8052), .B(n9827), .Y(n13744));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_sc1_3__U1(.A(n8067), .B(n13741), .Y(dpath_mulcore_ary1_a1_s0[3]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_sc1_3__U4(.A(n8051), .B(n8753), .Y(n13741));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_U4(.A(n9828), .B(n7406), .Y(dpath_mulcore_a1sum[0]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_sc1_1__U2(.A(dpath_mulcore_ary1_a1_I1_I0_b0n), .B(n7400), .Y(dpath_mulcore_ary1_a1_s1[1]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_sc1_2__U1(.A(n8062), .B(n13733), .Y(dpath_mulcore_ary1_a1_s1[2]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_sc1_2__U4(.A(n7925), .B(n9831), .Y(n13733));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_sc1_3__U1(.A(n8063), .B(n13730), .Y(dpath_mulcore_ary1_a1_s1[3]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_sc1_3__U4(.A(n7924), .B(n8692), .Y(n13730));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_U4(.A(n9832), .B(n7405), .Y(dpath_mulcore_ary1_a1_s1[0]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_sc1_1__U2(.A(dpath_mulcore_ary1_a1_I2_I0_b0n), .B(n7399), .Y(dpath_mulcore_ary1_a1_s2[1]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_sc1_2__U1(.A(n8060), .B(n13722), .Y(dpath_mulcore_ary1_a1_s2[2]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_sc1_2__U4(.A(n7798), .B(n9838), .Y(n13722));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_sc1_3__U1(.A(n8061), .B(n13719), .Y(dpath_mulcore_ary1_a1_s2[3]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_sc1_3__U4(.A(n7797), .B(n8631), .Y(n13719));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_U4(.A(n9839), .B(n7404), .Y(dpath_mulcore_ary1_a1_s2[0]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_sc1_1__U2(.A(dpath_mulcore_ary1_a0_I0_I0_b0n), .B(n7398), .Y(dpath_mulcore_a0sum[1]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_sc1_2__U1(.A(n8058), .B(n13711), .Y(dpath_mulcore_ary1_a0_s0[2]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_sc1_2__U4(.A(n7734), .B(n9840), .Y(n13711));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_sc1_3__U1(.A(n8059), .B(n13708), .Y(dpath_mulcore_ary1_a0_s0[3]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_sc1_3__U4(.A(n7733), .B(n8570), .Y(n13708));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_U4(.A(n9841), .B(n7403), .Y(dpath_mulcore_a0sum[0]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_sc1_1__U2(.A(dpath_mulcore_ary1_a0_I1_I0_b0n), .B(n7397), .Y(dpath_mulcore_ary1_a0_s1[1]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_sc1_2__U1(.A(n8054), .B(n13700), .Y(dpath_mulcore_ary1_a0_s1[2]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_sc1_2__U4(.A(n7607), .B(n9844), .Y(n13700));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_sc1_3__U1(.A(n8055), .B(n13697), .Y(dpath_mulcore_ary1_a0_s1[3]));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_sc1_3__U4(.A(n7606), .B(n8509), .Y(n13697));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_U4(.A(n9845), .B(n7402), .Y(dpath_mulcore_ary1_a0_s1[0]));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_p1_2__U6(.A(dpath_mulcore_b9[2]), .B(n9855), .Y(n13659));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_p0_0__U6(.A(dpath_mulcore_b8[2]), .B(n9855), .Y(n13657));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_p0_1__U6(.A(dpath_mulcore_b8[2]), .B(n9858), .Y(n13655));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_p0_2__U6(.A(dpath_mulcore_b8[2]), .B(n9861), .Y(n13652));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_p1_3__U6(.A(dpath_mulcore_b9[2]), .B(n9858), .Y(n13649));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I0_p0_3__U6(.A(dpath_mulcore_b8[2]), .B(n9864), .Y(n13646));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_4__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9867), .Y(n13643));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_4__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9861), .Y(n13640));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_4__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9855), .Y(n13637));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_5__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9870), .Y(n13635));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_5__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9864), .Y(n13632));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_5__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9858), .Y(n13629));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_6__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9873), .Y(n13626));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_6__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9867), .Y(n13623));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_6__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9861), .Y(n13620));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_7__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9876), .Y(n13617));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_7__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9870), .Y(n13614));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_7__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9864), .Y(n13611));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_8__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9879), .Y(n13608));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_8__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9873), .Y(n13605));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_8__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9867), .Y(n13602));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_9__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9882), .Y(n13599));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_9__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9876), .Y(n13596));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_9__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9870), .Y(n13593));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_10__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9885), .Y(n13590));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_10__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9879), .Y(n13587));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_10__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9873), .Y(n13584));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_11__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9888), .Y(n13581));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_11__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9882), .Y(n13578));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_11__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9876), .Y(n13575));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_12__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9891), .Y(n13572));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_12__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9885), .Y(n13569));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_12__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9879), .Y(n13566));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_13__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9894), .Y(n13563));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_13__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9888), .Y(n13560));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_13__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9882), .Y(n13557));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_14__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9897), .Y(n13554));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_14__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9891), .Y(n13551));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_14__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9885), .Y(n13548));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_15__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9900), .Y(n13545));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_15__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9894), .Y(n13542));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_15__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9888), .Y(n13539));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_16__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9903), .Y(n13536));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_16__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9897), .Y(n13533));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_16__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9891), .Y(n13530));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_17__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9906), .Y(n13527));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_17__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9900), .Y(n13524));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_17__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9894), .Y(n13521));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_18__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9909), .Y(n13518));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_18__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9903), .Y(n13515));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_18__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9897), .Y(n13512));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_19__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9912), .Y(n13509));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_19__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9906), .Y(n13506));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_19__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9900), .Y(n13503));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_20__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9915), .Y(n13500));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_20__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9909), .Y(n13497));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_20__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9903), .Y(n13494));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_21__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9918), .Y(n13491));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_21__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9912), .Y(n13488));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_21__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9906), .Y(n13485));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_22__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9921), .Y(n13482));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_22__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9915), .Y(n13479));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_22__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9909), .Y(n13476));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_23__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9924), .Y(n13473));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_23__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9918), .Y(n13470));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_23__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9912), .Y(n13467));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_24__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9927), .Y(n13464));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_24__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9921), .Y(n13461));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_24__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9915), .Y(n13458));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_25__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9930), .Y(n13455));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_25__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9924), .Y(n13452));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_25__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9918), .Y(n13449));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_26__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9933), .Y(n13446));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_26__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9927), .Y(n13443));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_26__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9921), .Y(n13440));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_27__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9936), .Y(n13437));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_27__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9930), .Y(n13434));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_27__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9924), .Y(n13431));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_28__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9939), .Y(n13428));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_28__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9933), .Y(n13425));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_28__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9927), .Y(n13422));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_29__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9942), .Y(n13419));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_29__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9936), .Y(n13416));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_29__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9930), .Y(n13413));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_30__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9945), .Y(n13410));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_30__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9939), .Y(n13407));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_30__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9933), .Y(n13404));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_31__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9948), .Y(n13401));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_31__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9942), .Y(n13398));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_31__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9936), .Y(n13395));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_32__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9951), .Y(n13392));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_32__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9945), .Y(n13389));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_32__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9939), .Y(n13386));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_33__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9954), .Y(n13383));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_33__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9948), .Y(n13380));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_33__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9942), .Y(n13377));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_34__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9957), .Y(n13374));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_34__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9951), .Y(n13371));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_34__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9945), .Y(n13368));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_35__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9960), .Y(n13365));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_35__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9954), .Y(n13362));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_35__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9948), .Y(n13359));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_36__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9963), .Y(n13356));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_36__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9957), .Y(n13353));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_36__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9951), .Y(n13350));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_37__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9966), .Y(n13347));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_37__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9960), .Y(n13344));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_37__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9954), .Y(n13341));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_38__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9969), .Y(n13338));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_38__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9963), .Y(n13335));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_38__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9957), .Y(n13332));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_39__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9972), .Y(n13329));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_39__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9966), .Y(n13326));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_39__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9960), .Y(n13323));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_40__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9975), .Y(n13320));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_40__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9969), .Y(n13317));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_40__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9963), .Y(n13314));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_41__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9978), .Y(n13311));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_41__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9972), .Y(n13308));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_41__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9966), .Y(n13305));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_42__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9981), .Y(n13302));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_42__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9975), .Y(n13299));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_42__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9969), .Y(n13296));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_43__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9984), .Y(n13293));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_43__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9978), .Y(n13290));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_43__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9972), .Y(n13287));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_44__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9987), .Y(n13284));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_44__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9981), .Y(n13281));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_44__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9975), .Y(n13278));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_45__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9990), .Y(n13275));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_45__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9984), .Y(n13272));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_45__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9978), .Y(n13269));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_46__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9993), .Y(n13266));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_46__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9987), .Y(n13263));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_46__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9981), .Y(n13260));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_47__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9996), .Y(n13257));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_47__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9990), .Y(n13254));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_47__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9984), .Y(n13251));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_48__p0_U6(.A(dpath_mulcore_b8[2]), .B(n9998), .Y(n13248));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_48__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9993), .Y(n13245));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_48__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9987), .Y(n13242));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_49__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10000), .Y(n13239));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_49__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9996), .Y(n13236));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_49__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9990), .Y(n13233));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_50__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10002), .Y(n13230));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_50__p1_U6(.A(dpath_mulcore_b9[2]), .B(n9998), .Y(n13227));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_50__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9993), .Y(n13224));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_51__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10004), .Y(n13221));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_51__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10000), .Y(n13218));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_51__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9996), .Y(n13215));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_52__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10006), .Y(n13212));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_52__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10002), .Y(n13209));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_52__p2_U6(.A(dpath_mulcore_b10[2]), .B(n9998), .Y(n13206));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_53__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10009), .Y(n13203));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_53__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10004), .Y(n13200));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_53__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10000), .Y(n13197));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_54__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10012), .Y(n13194));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_54__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10006), .Y(n13191));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_54__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10002), .Y(n13188));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_55__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10015), .Y(n13185));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_55__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10009), .Y(n13182));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_55__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10004), .Y(n13179));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_56__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10018), .Y(n13176));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_56__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10012), .Y(n13173));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_56__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10006), .Y(n13170));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_57__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10021), .Y(n13167));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_57__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10015), .Y(n13164));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_57__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10009), .Y(n13161));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_58__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10024), .Y(n13158));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_58__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10018), .Y(n13155));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_58__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10012), .Y(n13152));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_59__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10028), .Y(n13149));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_59__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10021), .Y(n13146));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_59__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10015), .Y(n13143));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_60__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10029), .Y(n13140));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_60__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10024), .Y(n13137));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_60__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10018), .Y(n13134));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_61__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10030), .Y(n13131));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_61__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10028), .Y(n13128));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_61__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10021), .Y(n13125));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_62__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10031), .Y(n13122));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_62__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10029), .Y(n13119));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_62__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10024), .Y(n13116));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_63__p0_U6(.A(dpath_mulcore_b8[2]), .B(n10032), .Y(n13113));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_63__p1_U6(.A(dpath_mulcore_b9[2]), .B(n10030), .Y(n13110));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I1_63__p2_U6(.A(dpath_mulcore_b10[2]), .B(n10028), .Y(n13107));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_p2_64__U6(.A(dpath_mulcore_b10[2]), .B(n10029), .Y(n13104));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_p1_64__U6(.A(dpath_mulcore_b9[2]), .B(n10031), .Y(n13101));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_p1_65__U6(.A(dpath_mulcore_b9[2]), .B(n10032), .Y(n13098));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_p2_65__U6(.A(dpath_mulcore_b10[2]), .B(n10030), .Y(n13095));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_p2_66__U6(.A(dpath_mulcore_b10[2]), .B(n10031), .Y(n13092));
XOR2X1 mul_dpath_mulcore_ary1_a1_I0_I2_p2_67__U6(.A(dpath_mulcore_b10[2]), .B(n10032), .Y(n13089));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_p1_2__U6(.A(dpath_mulcore_b12[2]), .B(n9855), .Y(n13086));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_p0_0__U6(.A(dpath_mulcore_b11[2]), .B(n9855), .Y(n13084));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_p0_1__U6(.A(dpath_mulcore_b11[2]), .B(n9858), .Y(n13082));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_p0_2__U6(.A(dpath_mulcore_b11[2]), .B(n9861), .Y(n13079));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_p1_3__U6(.A(dpath_mulcore_b12[2]), .B(n9858), .Y(n13076));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I0_p0_3__U6(.A(dpath_mulcore_b11[2]), .B(n9864), .Y(n13073));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_4__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9867), .Y(n13070));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_4__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9861), .Y(n13067));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_4__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9855), .Y(n13064));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_5__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9870), .Y(n13062));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_5__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9864), .Y(n13059));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_5__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9858), .Y(n13056));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_6__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9873), .Y(n13053));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_6__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9867), .Y(n13050));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_6__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9861), .Y(n13047));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_7__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9876), .Y(n13044));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_7__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9870), .Y(n13041));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_7__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9864), .Y(n13038));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_8__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9879), .Y(n13035));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_8__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9873), .Y(n13032));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_8__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9867), .Y(n13029));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_9__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9882), .Y(n13026));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_9__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9876), .Y(n13023));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_9__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9870), .Y(n13020));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_10__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9885), .Y(n13017));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_10__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9879), .Y(n13014));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_10__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9873), .Y(n13011));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_11__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9888), .Y(n13008));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_11__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9882), .Y(n13005));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_11__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9876), .Y(n13002));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_12__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9891), .Y(n12999));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_12__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9885), .Y(n12996));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_12__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9879), .Y(n12993));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_13__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9894), .Y(n12990));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_13__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9888), .Y(n12987));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_13__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9882), .Y(n12984));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_14__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9897), .Y(n12981));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_14__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9891), .Y(n12978));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_14__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9885), .Y(n12975));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_15__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9900), .Y(n12972));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_15__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9894), .Y(n12969));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_15__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9888), .Y(n12966));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_16__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9903), .Y(n12963));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_16__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9897), .Y(n12960));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_16__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9891), .Y(n12957));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_17__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9906), .Y(n12954));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_17__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9900), .Y(n12951));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_17__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9894), .Y(n12948));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_18__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9909), .Y(n12945));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_18__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9903), .Y(n12942));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_18__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9897), .Y(n12939));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_19__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9912), .Y(n12936));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_19__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9906), .Y(n12933));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_19__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9900), .Y(n12930));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_20__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9915), .Y(n12927));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_20__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9909), .Y(n12924));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_20__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9903), .Y(n12921));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_21__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9918), .Y(n12918));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_21__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9912), .Y(n12915));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_21__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9906), .Y(n12912));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_22__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9921), .Y(n12909));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_22__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9915), .Y(n12906));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_22__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9909), .Y(n12903));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_23__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9924), .Y(n12900));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_23__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9918), .Y(n12897));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_23__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9912), .Y(n12894));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_24__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9927), .Y(n12891));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_24__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9921), .Y(n12888));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_24__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9915), .Y(n12885));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_25__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9930), .Y(n12882));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_25__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9924), .Y(n12879));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_25__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9918), .Y(n12876));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_26__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9933), .Y(n12873));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_26__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9927), .Y(n12870));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_26__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9921), .Y(n12867));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_27__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9936), .Y(n12864));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_27__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9930), .Y(n12861));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_27__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9924), .Y(n12858));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_28__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9939), .Y(n12855));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_28__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9933), .Y(n12852));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_28__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9927), .Y(n12849));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_29__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9942), .Y(n12846));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_29__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9936), .Y(n12843));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_29__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9930), .Y(n12840));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_30__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9945), .Y(n12837));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_30__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9939), .Y(n12834));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_30__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9933), .Y(n12831));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_31__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9948), .Y(n12828));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_31__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9942), .Y(n12825));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_31__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9936), .Y(n12822));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_32__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9951), .Y(n12819));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_32__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9945), .Y(n12816));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_32__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9939), .Y(n12813));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_33__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9954), .Y(n12810));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_33__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9948), .Y(n12807));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_33__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9942), .Y(n12804));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_34__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9957), .Y(n12801));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_34__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9951), .Y(n12798));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_34__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9945), .Y(n12795));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_35__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9960), .Y(n12792));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_35__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9954), .Y(n12789));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_35__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9948), .Y(n12786));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_36__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9963), .Y(n12783));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_36__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9957), .Y(n12780));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_36__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9951), .Y(n12777));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_37__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9966), .Y(n12774));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_37__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9960), .Y(n12771));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_37__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9954), .Y(n12768));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_38__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9969), .Y(n12765));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_38__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9963), .Y(n12762));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_38__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9957), .Y(n12759));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_39__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9972), .Y(n12756));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_39__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9966), .Y(n12753));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_39__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9960), .Y(n12750));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_40__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9975), .Y(n12747));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_40__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9969), .Y(n12744));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_40__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9963), .Y(n12741));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_41__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9978), .Y(n12738));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_41__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9972), .Y(n12735));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_41__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9966), .Y(n12732));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_42__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9981), .Y(n12729));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_42__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9975), .Y(n12726));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_42__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9969), .Y(n12723));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_43__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9984), .Y(n12720));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_43__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9978), .Y(n12717));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_43__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9972), .Y(n12714));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_44__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9987), .Y(n12711));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_44__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9981), .Y(n12708));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_44__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9975), .Y(n12705));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_45__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9990), .Y(n12702));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_45__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9984), .Y(n12699));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_45__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9978), .Y(n12696));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_46__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9993), .Y(n12693));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_46__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9987), .Y(n12690));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_46__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9981), .Y(n12687));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_47__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9996), .Y(n12684));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_47__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9990), .Y(n12681));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_47__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9984), .Y(n12678));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_48__p0_U6(.A(dpath_mulcore_b11[2]), .B(n9998), .Y(n12675));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_48__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9993), .Y(n12672));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_48__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9987), .Y(n12669));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_49__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10000), .Y(n12666));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_49__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9996), .Y(n12663));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_49__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9990), .Y(n12660));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_50__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10002), .Y(n12657));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_50__p1_U6(.A(dpath_mulcore_b12[2]), .B(n9998), .Y(n12654));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_50__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9993), .Y(n12651));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_51__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10004), .Y(n12648));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_51__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10000), .Y(n12645));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_51__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9996), .Y(n12642));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_52__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10006), .Y(n12639));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_52__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10002), .Y(n12636));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_52__p2_U6(.A(dpath_mulcore_b13[2]), .B(n9998), .Y(n12633));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_53__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10009), .Y(n12630));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_53__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10004), .Y(n12627));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_53__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10000), .Y(n12624));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_54__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10012), .Y(n12621));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_54__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10006), .Y(n12618));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_54__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10002), .Y(n12615));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_55__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10015), .Y(n12612));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_55__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10009), .Y(n12609));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_55__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10004), .Y(n12606));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_56__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10018), .Y(n12603));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_56__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10012), .Y(n12600));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_56__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10006), .Y(n12597));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_57__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10021), .Y(n12594));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_57__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10015), .Y(n12591));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_57__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10009), .Y(n12588));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_58__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10024), .Y(n12585));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_58__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10018), .Y(n12582));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_58__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10012), .Y(n12579));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_59__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10028), .Y(n12576));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_59__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10021), .Y(n12573));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_59__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10015), .Y(n12570));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_60__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10029), .Y(n12567));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_60__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10024), .Y(n12564));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_60__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10018), .Y(n12561));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_61__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10030), .Y(n12558));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_61__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10028), .Y(n12555));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_61__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10021), .Y(n12552));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_62__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10031), .Y(n12549));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_62__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10029), .Y(n12546));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_62__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10024), .Y(n12543));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_63__p0_U6(.A(dpath_mulcore_b11[2]), .B(n10032), .Y(n12540));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_63__p1_U6(.A(dpath_mulcore_b12[2]), .B(n10030), .Y(n12537));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I1_63__p2_U6(.A(dpath_mulcore_b13[2]), .B(n10028), .Y(n12534));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_p2_64__U6(.A(dpath_mulcore_b13[2]), .B(n10029), .Y(n12531));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_p1_64__U6(.A(dpath_mulcore_b12[2]), .B(n10031), .Y(n12528));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_p1_65__U6(.A(dpath_mulcore_b12[2]), .B(n10032), .Y(n12525));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_p2_65__U6(.A(dpath_mulcore_b13[2]), .B(n10030), .Y(n12522));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_p2_66__U6(.A(dpath_mulcore_b13[2]), .B(n10031), .Y(n12519));
XOR2X1 mul_dpath_mulcore_ary1_a1_I1_I2_p2_67__U6(.A(dpath_mulcore_b13[2]), .B(n10032), .Y(n12516));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_p1_2__U6(.A(dpath_mulcore_b15[2]), .B(n9855), .Y(n12513));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_p0_0__U6(.A(dpath_mulcore_b14[2]), .B(n9855), .Y(n12511));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_p0_1__U6(.A(dpath_mulcore_b14[2]), .B(n9858), .Y(n12509));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_p0_2__U6(.A(dpath_mulcore_b14[2]), .B(n9861), .Y(n12506));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_p1_3__U6(.A(dpath_mulcore_b15[2]), .B(n9858), .Y(n12503));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I0_p0_3__U6(.A(dpath_mulcore_b14[2]), .B(n9864), .Y(n12500));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_4__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9867), .Y(n12497));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_4__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9861), .Y(n12494));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_5__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9870), .Y(n12491));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_5__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9864), .Y(n12488));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_6__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9873), .Y(n12485));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_6__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9867), .Y(n12482));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_7__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9876), .Y(n12479));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_7__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9870), .Y(n12476));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_8__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9879), .Y(n12473));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_8__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9873), .Y(n12470));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_9__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9882), .Y(n12467));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_9__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9876), .Y(n12464));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_10__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9885), .Y(n12461));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_10__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9879), .Y(n12458));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_11__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9888), .Y(n12455));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_11__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9882), .Y(n12452));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_12__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9891), .Y(n12449));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_12__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9885), .Y(n12446));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_13__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9894), .Y(n12443));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_13__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9888), .Y(n12440));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_14__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9897), .Y(n12437));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_14__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9891), .Y(n12434));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_15__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9900), .Y(n12431));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_15__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9894), .Y(n12428));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_16__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9903), .Y(n12425));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_16__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9897), .Y(n12422));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_17__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9906), .Y(n12419));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_17__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9900), .Y(n12416));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_18__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9909), .Y(n12413));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_18__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9903), .Y(n12410));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_19__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9912), .Y(n12407));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_19__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9906), .Y(n12404));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_20__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9915), .Y(n12401));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_20__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9909), .Y(n12398));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_21__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9918), .Y(n12395));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_21__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9912), .Y(n12392));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_22__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9921), .Y(n12389));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_22__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9915), .Y(n12386));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_23__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9924), .Y(n12383));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_23__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9918), .Y(n12380));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_24__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9927), .Y(n12377));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_24__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9921), .Y(n12374));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_25__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9930), .Y(n12371));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_25__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9924), .Y(n12368));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_26__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9933), .Y(n12365));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_26__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9927), .Y(n12362));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_27__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9936), .Y(n12359));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_27__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9930), .Y(n12356));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_28__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9939), .Y(n12353));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_28__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9933), .Y(n12350));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_29__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9942), .Y(n12347));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_29__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9936), .Y(n12344));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_30__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9945), .Y(n12341));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_30__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9939), .Y(n12338));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_31__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9948), .Y(n12335));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_31__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9942), .Y(n12332));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_32__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9951), .Y(n12329));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_32__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9945), .Y(n12326));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_33__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9954), .Y(n12323));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_33__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9948), .Y(n12320));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_34__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9957), .Y(n12317));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_34__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9951), .Y(n12314));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_35__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9960), .Y(n12311));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_35__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9954), .Y(n12308));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_36__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9963), .Y(n12305));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_36__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9957), .Y(n12302));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_37__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9966), .Y(n12299));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_37__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9960), .Y(n12296));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_38__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9969), .Y(n12293));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_38__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9963), .Y(n12290));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_39__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9972), .Y(n12287));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_39__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9966), .Y(n12284));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_40__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9975), .Y(n12281));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_40__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9969), .Y(n12278));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_41__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9978), .Y(n12275));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_41__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9972), .Y(n12272));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_42__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9981), .Y(n12269));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_42__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9975), .Y(n12266));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_43__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9984), .Y(n12263));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_43__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9978), .Y(n12260));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_44__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9987), .Y(n12257));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_44__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9981), .Y(n12254));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_45__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9990), .Y(n12251));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_45__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9984), .Y(n12248));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_46__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9993), .Y(n12245));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_46__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9987), .Y(n12242));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_47__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9996), .Y(n12239));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_47__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9990), .Y(n12236));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_48__p0_U6(.A(dpath_mulcore_b14[2]), .B(n9998), .Y(n12233));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_48__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9993), .Y(n12230));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_49__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10000), .Y(n12227));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_49__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9996), .Y(n12224));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_50__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10002), .Y(n12221));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_50__p1_U6(.A(dpath_mulcore_b15[2]), .B(n9998), .Y(n12218));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_51__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10004), .Y(n12215));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_51__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10000), .Y(n12212));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_52__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10006), .Y(n12209));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_52__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10002), .Y(n12206));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_53__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10009), .Y(n12203));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_53__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10004), .Y(n12200));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_54__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10012), .Y(n12197));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_54__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10006), .Y(n12194));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_55__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10015), .Y(n12191));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_55__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10009), .Y(n12188));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_56__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10018), .Y(n12185));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_56__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10012), .Y(n12182));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_57__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10021), .Y(n12179));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_57__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10015), .Y(n12176));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_58__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10024), .Y(n12173));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_58__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10018), .Y(n12170));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_59__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10028), .Y(n12167));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_59__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10021), .Y(n12164));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_60__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10029), .Y(n12161));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_60__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10024), .Y(n12158));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_61__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10030), .Y(n12155));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_61__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10028), .Y(n12152));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_62__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10031), .Y(n12149));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_62__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10029), .Y(n12146));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_63__p0_U6(.A(dpath_mulcore_b14[2]), .B(n10032), .Y(n12143));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I1_63__p1_U6(.A(dpath_mulcore_b15[2]), .B(n10030), .Y(n12140));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I2_p1_64__U6(.A(dpath_mulcore_b15[2]), .B(n10031), .Y(n12137));
XOR2X1 mul_dpath_mulcore_ary1_a1_I2_I2_p1_65__U6(.A(dpath_mulcore_b15[2]), .B(n10032), .Y(n12134));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_p1_2__U6(.A(dpath_mulcore_b1[2]), .B(n9855), .Y(n12131));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_p0_0__U6(.A(dpath_mulcore_b0[2]), .B(n9855), .Y(n12129));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_p0_1__U6(.A(dpath_mulcore_b0[2]), .B(n9858), .Y(n12127));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_p0_2__U6(.A(dpath_mulcore_b0[2]), .B(n9861), .Y(n12124));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_p1_3__U6(.A(dpath_mulcore_b1[2]), .B(n9858), .Y(n12121));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I0_p0_3__U6(.A(dpath_mulcore_b0[2]), .B(n9864), .Y(n12118));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_4__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9867), .Y(n12115));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_4__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9861), .Y(n12112));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_4__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9855), .Y(n12109));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_5__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9870), .Y(n12107));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_5__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9864), .Y(n12104));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_5__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9858), .Y(n12101));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_6__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9873), .Y(n12098));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_6__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9867), .Y(n12095));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_6__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9861), .Y(n12092));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_7__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9876), .Y(n12089));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_7__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9870), .Y(n12086));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_7__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9864), .Y(n12083));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_8__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9879), .Y(n12080));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_8__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9873), .Y(n12077));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_8__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9867), .Y(n12074));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_9__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9882), .Y(n12071));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_9__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9876), .Y(n12068));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_9__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9870), .Y(n12065));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_10__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9885), .Y(n12062));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_10__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9879), .Y(n12059));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_10__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9873), .Y(n12056));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_11__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9888), .Y(n12053));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_11__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9882), .Y(n12050));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_11__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9876), .Y(n12047));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_12__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9891), .Y(n12044));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_12__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9885), .Y(n12041));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_12__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9879), .Y(n12038));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_13__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9894), .Y(n12035));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_13__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9888), .Y(n12032));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_13__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9882), .Y(n12029));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_14__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9897), .Y(n12026));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_14__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9891), .Y(n12023));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_14__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9885), .Y(n12020));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_15__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9900), .Y(n12017));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_15__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9894), .Y(n12014));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_15__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9888), .Y(n12011));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_16__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9903), .Y(n12008));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_16__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9897), .Y(n12005));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_16__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9891), .Y(n12002));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_17__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9906), .Y(n11999));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_17__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9900), .Y(n11996));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_17__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9894), .Y(n11993));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_18__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9909), .Y(n11990));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_18__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9903), .Y(n11987));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_18__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9897), .Y(n11984));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_19__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9912), .Y(n11981));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_19__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9906), .Y(n11978));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_19__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9900), .Y(n11975));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_20__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9915), .Y(n11972));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_20__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9909), .Y(n11969));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_20__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9903), .Y(n11966));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_21__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9918), .Y(n11963));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_21__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9912), .Y(n11960));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_21__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9906), .Y(n11957));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_22__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9921), .Y(n11954));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_22__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9915), .Y(n11951));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_22__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9909), .Y(n11948));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_23__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9924), .Y(n11945));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_23__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9918), .Y(n11942));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_23__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9912), .Y(n11939));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_24__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9927), .Y(n11936));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_24__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9921), .Y(n11933));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_24__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9915), .Y(n11930));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_25__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9930), .Y(n11927));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_25__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9924), .Y(n11924));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_25__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9918), .Y(n11921));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_26__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9933), .Y(n11918));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_26__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9927), .Y(n11915));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_26__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9921), .Y(n11912));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_27__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9936), .Y(n11909));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_27__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9930), .Y(n11906));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_27__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9924), .Y(n11903));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_28__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9939), .Y(n11900));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_28__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9933), .Y(n11897));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_28__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9927), .Y(n11894));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_29__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9942), .Y(n11891));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_29__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9936), .Y(n11888));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_29__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9930), .Y(n11885));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_30__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9945), .Y(n11882));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_30__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9939), .Y(n11879));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_30__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9933), .Y(n11876));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_31__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9948), .Y(n11873));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_31__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9942), .Y(n11870));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_31__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9936), .Y(n11867));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_32__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9951), .Y(n11864));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_32__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9945), .Y(n11861));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_32__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9939), .Y(n11858));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_33__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9954), .Y(n11855));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_33__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9948), .Y(n11852));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_33__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9942), .Y(n11849));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_34__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9957), .Y(n11846));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_34__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9951), .Y(n11843));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_34__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9945), .Y(n11840));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_35__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9960), .Y(n11837));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_35__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9954), .Y(n11834));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_35__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9948), .Y(n11831));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_36__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9963), .Y(n11828));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_36__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9957), .Y(n11825));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_36__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9951), .Y(n11822));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_37__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9966), .Y(n11819));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_37__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9960), .Y(n11816));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_37__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9954), .Y(n11813));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_38__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9969), .Y(n11810));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_38__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9963), .Y(n11807));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_38__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9957), .Y(n11804));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_39__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9972), .Y(n11801));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_39__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9966), .Y(n11798));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_39__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9960), .Y(n11795));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_40__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9975), .Y(n11792));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_40__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9969), .Y(n11789));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_40__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9963), .Y(n11786));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_41__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9978), .Y(n11783));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_41__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9972), .Y(n11780));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_41__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9966), .Y(n11777));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_42__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9981), .Y(n11774));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_42__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9975), .Y(n11771));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_42__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9969), .Y(n11768));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_43__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9984), .Y(n11765));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_43__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9978), .Y(n11762));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_43__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9972), .Y(n11759));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_44__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9987), .Y(n11756));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_44__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9981), .Y(n11753));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_44__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9975), .Y(n11750));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_45__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9990), .Y(n11747));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_45__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9984), .Y(n11744));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_45__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9978), .Y(n11741));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_46__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9993), .Y(n11738));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_46__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9987), .Y(n11735));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_46__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9981), .Y(n11732));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_47__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9996), .Y(n11729));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_47__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9990), .Y(n11726));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_47__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9984), .Y(n11723));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_48__p0_U6(.A(dpath_mulcore_b0[2]), .B(n9998), .Y(n11720));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_48__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9993), .Y(n11717));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_48__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9987), .Y(n11714));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_49__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10000), .Y(n11711));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_49__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9996), .Y(n11708));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_49__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9990), .Y(n11705));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_50__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10002), .Y(n11702));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_50__p1_U6(.A(dpath_mulcore_b1[2]), .B(n9998), .Y(n11699));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_50__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9993), .Y(n11696));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_51__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10004), .Y(n11693));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_51__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10000), .Y(n11690));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_51__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9996), .Y(n11687));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_52__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10006), .Y(n11684));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_52__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10002), .Y(n11681));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_52__p2_U6(.A(dpath_mulcore_b2[2]), .B(n9998), .Y(n11678));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_53__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10009), .Y(n11675));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_53__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10004), .Y(n11672));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_53__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10000), .Y(n11669));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_54__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10012), .Y(n11666));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_54__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10006), .Y(n11663));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_54__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10002), .Y(n11660));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_55__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10015), .Y(n11657));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_55__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10009), .Y(n11654));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_55__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10004), .Y(n11651));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_56__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10018), .Y(n11648));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_56__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10012), .Y(n11645));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_56__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10006), .Y(n11642));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_57__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10021), .Y(n11639));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_57__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10015), .Y(n11636));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_57__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10009), .Y(n11633));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_58__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10024), .Y(n11630));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_58__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10018), .Y(n11627));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_58__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10012), .Y(n11624));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_59__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10028), .Y(n11621));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_59__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10021), .Y(n11618));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_59__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10015), .Y(n11615));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_60__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10029), .Y(n11612));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_60__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10024), .Y(n11609));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_60__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10018), .Y(n11606));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_61__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10030), .Y(n11603));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_61__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10028), .Y(n11600));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_61__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10021), .Y(n11597));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_62__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10031), .Y(n11594));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_62__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10029), .Y(n11591));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_62__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10024), .Y(n11588));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_63__p0_U6(.A(dpath_mulcore_b0[2]), .B(n10032), .Y(n11585));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_63__p1_U6(.A(dpath_mulcore_b1[2]), .B(n10030), .Y(n11582));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I1_63__p2_U6(.A(dpath_mulcore_b2[2]), .B(n10028), .Y(n11579));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_p2_64__U6(.A(dpath_mulcore_b2[2]), .B(n10029), .Y(n11576));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_p1_64__U6(.A(dpath_mulcore_b1[2]), .B(n10031), .Y(n11573));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_p1_65__U6(.A(dpath_mulcore_b1[2]), .B(n10032), .Y(n11570));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_p2_65__U6(.A(dpath_mulcore_b2[2]), .B(n10030), .Y(n11567));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_p2_66__U6(.A(dpath_mulcore_b2[2]), .B(n10031), .Y(n11564));
XOR2X1 mul_dpath_mulcore_ary1_a0_I0_I2_p2_67__U6(.A(dpath_mulcore_b2[2]), .B(n10032), .Y(n11561));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_p1_2__U6(.A(dpath_mulcore_b4[2]), .B(n9855), .Y(n11558));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_p0_0__U6(.A(dpath_mulcore_b3[2]), .B(n9855), .Y(n11556));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_p0_1__U6(.A(dpath_mulcore_b3[2]), .B(n9858), .Y(n11554));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_p0_2__U6(.A(dpath_mulcore_b3[2]), .B(n9861), .Y(n11551));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_p1_3__U6(.A(dpath_mulcore_b4[2]), .B(n9858), .Y(n11548));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I0_p0_3__U6(.A(dpath_mulcore_b3[2]), .B(n9864), .Y(n11545));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_4__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9867), .Y(n11542));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_4__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9861), .Y(n11539));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_4__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9855), .Y(n11536));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_5__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9870), .Y(n11534));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_5__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9864), .Y(n11531));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_5__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9858), .Y(n11528));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_6__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9873), .Y(n11525));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_6__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9867), .Y(n11522));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_6__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9861), .Y(n11519));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_7__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9876), .Y(n11516));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_7__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9870), .Y(n11513));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_7__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9864), .Y(n11510));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_8__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9879), .Y(n11507));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_8__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9873), .Y(n11504));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_8__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9867), .Y(n11501));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_9__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9882), .Y(n11498));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_9__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9876), .Y(n11495));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_9__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9870), .Y(n11492));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_10__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9885), .Y(n11489));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_10__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9879), .Y(n11486));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_10__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9873), .Y(n11483));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_11__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9888), .Y(n11480));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_11__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9882), .Y(n11477));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_11__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9876), .Y(n11474));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_12__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9891), .Y(n11471));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_12__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9885), .Y(n11468));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_12__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9879), .Y(n11465));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_13__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9894), .Y(n11462));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_13__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9888), .Y(n11459));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_13__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9882), .Y(n11456));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_14__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9897), .Y(n11453));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_14__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9891), .Y(n11450));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_14__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9885), .Y(n11447));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_15__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9900), .Y(n11444));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_15__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9894), .Y(n11441));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_15__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9888), .Y(n11438));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_16__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9903), .Y(n11435));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_16__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9897), .Y(n11432));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_16__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9891), .Y(n11429));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_17__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9906), .Y(n11426));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_17__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9900), .Y(n11423));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_17__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9894), .Y(n11420));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_18__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9909), .Y(n11417));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_18__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9903), .Y(n11414));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_18__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9897), .Y(n11411));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_19__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9912), .Y(n11408));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_19__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9906), .Y(n11405));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_19__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9900), .Y(n11402));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_20__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9915), .Y(n11399));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_20__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9909), .Y(n11396));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_20__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9903), .Y(n11393));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_21__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9918), .Y(n11390));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_21__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9912), .Y(n11387));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_21__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9906), .Y(n11384));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_22__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9921), .Y(n11381));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_22__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9915), .Y(n11378));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_22__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9909), .Y(n11375));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_23__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9924), .Y(n11372));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_23__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9918), .Y(n11369));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_23__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9912), .Y(n11366));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_24__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9927), .Y(n11363));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_24__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9921), .Y(n11360));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_24__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9915), .Y(n11357));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_25__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9930), .Y(n11354));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_25__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9924), .Y(n11351));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_25__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9918), .Y(n11348));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_26__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9933), .Y(n11345));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_26__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9927), .Y(n11342));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_26__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9921), .Y(n11339));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_27__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9936), .Y(n11336));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_27__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9930), .Y(n11333));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_27__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9924), .Y(n11330));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_28__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9939), .Y(n11327));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_28__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9933), .Y(n11324));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_28__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9927), .Y(n11321));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_29__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9942), .Y(n11318));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_29__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9936), .Y(n11315));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_29__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9930), .Y(n11312));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_30__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9945), .Y(n11309));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_30__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9939), .Y(n11306));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_30__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9933), .Y(n11303));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_31__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9948), .Y(n11300));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_31__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9942), .Y(n11297));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_31__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9936), .Y(n11294));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_32__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9951), .Y(n11291));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_32__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9945), .Y(n11288));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_32__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9939), .Y(n11285));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_33__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9954), .Y(n11282));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_33__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9948), .Y(n11279));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_33__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9942), .Y(n11276));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_34__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9957), .Y(n11273));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_34__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9951), .Y(n11270));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_34__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9945), .Y(n11267));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_35__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9960), .Y(n11264));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_35__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9954), .Y(n11261));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_35__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9948), .Y(n11258));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_36__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9963), .Y(n11255));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_36__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9957), .Y(n11252));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_36__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9951), .Y(n11249));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_37__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9966), .Y(n11246));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_37__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9960), .Y(n11243));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_37__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9954), .Y(n11240));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_38__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9969), .Y(n11237));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_38__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9963), .Y(n11234));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_38__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9957), .Y(n11231));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_39__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9972), .Y(n11228));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_39__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9966), .Y(n11225));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_39__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9960), .Y(n11222));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_40__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9975), .Y(n11219));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_40__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9969), .Y(n11216));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_40__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9963), .Y(n11213));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_41__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9978), .Y(n11210));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_41__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9972), .Y(n11207));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_41__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9966), .Y(n11204));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_42__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9981), .Y(n11201));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_42__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9975), .Y(n11198));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_42__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9969), .Y(n11195));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_43__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9984), .Y(n11192));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_43__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9978), .Y(n11189));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_43__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9972), .Y(n11186));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_44__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9987), .Y(n11183));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_44__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9981), .Y(n11180));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_44__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9975), .Y(n11177));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_45__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9990), .Y(n11174));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_45__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9984), .Y(n11171));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_45__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9978), .Y(n11168));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_46__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9993), .Y(n11165));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_46__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9987), .Y(n11162));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_46__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9981), .Y(n11159));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_47__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9996), .Y(n11156));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_47__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9990), .Y(n11153));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_47__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9984), .Y(n11150));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_48__p0_U6(.A(dpath_mulcore_b3[2]), .B(n9998), .Y(n11147));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_48__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9993), .Y(n11144));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_48__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9987), .Y(n11141));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_49__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10000), .Y(n11138));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_49__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9996), .Y(n11135));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_49__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9990), .Y(n11132));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_50__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10002), .Y(n11129));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_50__p1_U6(.A(dpath_mulcore_b4[2]), .B(n9998), .Y(n11126));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_50__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9993), .Y(n11123));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_51__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10004), .Y(n11120));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_51__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10000), .Y(n11117));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_51__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9996), .Y(n11114));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_52__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10006), .Y(n11111));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_52__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10002), .Y(n11108));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_52__p2_U6(.A(dpath_mulcore_b5[2]), .B(n9998), .Y(n11105));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_53__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10009), .Y(n11102));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_53__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10004), .Y(n11099));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_53__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10000), .Y(n11096));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_54__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10012), .Y(n11093));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_54__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10006), .Y(n11090));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_54__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10002), .Y(n11087));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_55__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10015), .Y(n11084));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_55__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10009), .Y(n11081));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_55__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10004), .Y(n11078));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_56__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10018), .Y(n11075));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_56__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10012), .Y(n11072));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_56__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10006), .Y(n11069));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_57__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10021), .Y(n11066));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_57__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10015), .Y(n11063));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_57__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10009), .Y(n11060));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_58__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10024), .Y(n11057));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_58__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10018), .Y(n11054));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_58__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10012), .Y(n11051));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_59__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10028), .Y(n11048));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_59__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10021), .Y(n11045));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_59__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10015), .Y(n11042));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_60__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10029), .Y(n11039));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_60__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10024), .Y(n11036));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_60__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10018), .Y(n11033));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_61__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10030), .Y(n11030));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_61__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10028), .Y(n11027));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_61__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10021), .Y(n11024));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_62__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10031), .Y(n11021));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_62__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10029), .Y(n11018));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_62__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10024), .Y(n11015));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_63__p0_U6(.A(dpath_mulcore_b3[2]), .B(n10032), .Y(n11012));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_63__p1_U6(.A(dpath_mulcore_b4[2]), .B(n10030), .Y(n11009));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I1_63__p2_U6(.A(dpath_mulcore_b5[2]), .B(n10028), .Y(n11006));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_p2_64__U6(.A(dpath_mulcore_b5[2]), .B(n10029), .Y(n11003));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_p1_64__U6(.A(dpath_mulcore_b4[2]), .B(n10031), .Y(n11000));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_p1_65__U6(.A(dpath_mulcore_b4[2]), .B(n10032), .Y(n10997));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_p2_65__U6(.A(dpath_mulcore_b5[2]), .B(n10030), .Y(n10994));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_p2_66__U6(.A(dpath_mulcore_b5[2]), .B(n10031), .Y(n10991));
XOR2X1 mul_dpath_mulcore_ary1_a0_I1_I2_p2_67__U6(.A(dpath_mulcore_b5[2]), .B(n10032), .Y(n10988));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_p1_2__U6(.A(dpath_mulcore_b7[2]), .B(n9855), .Y(n10985));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_p0_0__U6(.A(dpath_mulcore_b6[2]), .B(n9855), .Y(n10983));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_p0_1__U6(.A(dpath_mulcore_b6[2]), .B(n9858), .Y(n10981));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_p0_2__U6(.A(dpath_mulcore_b6[2]), .B(n9861), .Y(n10978));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_p1_3__U6(.A(dpath_mulcore_b7[2]), .B(n9858), .Y(n10975));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I0_p0_3__U6(.A(dpath_mulcore_b6[2]), .B(n9864), .Y(n10972));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_4__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9867), .Y(n10969));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_4__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9861), .Y(n10966));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_5__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9870), .Y(n10963));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_5__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9864), .Y(n10960));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_6__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9873), .Y(n10957));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_6__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9867), .Y(n10954));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_7__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9876), .Y(n10951));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_7__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9870), .Y(n10948));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_8__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9879), .Y(n10945));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_8__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9873), .Y(n10942));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_9__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9882), .Y(n10939));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_9__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9876), .Y(n10936));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_10__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9885), .Y(n10933));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_10__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9879), .Y(n10930));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_11__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9888), .Y(n10927));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_11__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9882), .Y(n10924));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_12__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9891), .Y(n10921));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_12__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9885), .Y(n10918));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_13__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9894), .Y(n10915));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_13__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9888), .Y(n10912));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_14__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9897), .Y(n10909));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_14__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9891), .Y(n10906));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_15__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9900), .Y(n10903));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_15__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9894), .Y(n10900));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_16__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9903), .Y(n10897));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_16__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9897), .Y(n10894));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_17__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9906), .Y(n10891));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_17__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9900), .Y(n10888));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_18__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9909), .Y(n10885));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_18__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9903), .Y(n10882));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_19__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9912), .Y(n10879));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_19__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9906), .Y(n10876));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_20__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9915), .Y(n10873));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_20__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9909), .Y(n10870));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_21__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9918), .Y(n10867));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_21__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9912), .Y(n10864));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_22__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9921), .Y(n10861));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_22__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9915), .Y(n10858));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_23__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9924), .Y(n10855));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_23__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9918), .Y(n10852));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_24__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9927), .Y(n10849));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_24__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9921), .Y(n10846));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_25__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9930), .Y(n10843));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_25__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9924), .Y(n10840));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_26__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9933), .Y(n10837));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_26__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9927), .Y(n10834));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_27__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9936), .Y(n10831));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_27__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9930), .Y(n10828));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_28__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9939), .Y(n10825));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_28__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9933), .Y(n10822));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_29__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9942), .Y(n10819));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_29__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9936), .Y(n10816));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_30__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9945), .Y(n10813));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_30__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9939), .Y(n10810));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_31__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9948), .Y(n10807));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_31__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9942), .Y(n10804));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_32__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9951), .Y(n10801));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_32__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9945), .Y(n10798));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_33__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9954), .Y(n10795));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_33__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9948), .Y(n10792));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_34__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9957), .Y(n10789));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_34__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9951), .Y(n10786));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_35__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9960), .Y(n10783));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_35__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9954), .Y(n10780));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_36__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9963), .Y(n10777));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_36__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9957), .Y(n10774));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_37__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9966), .Y(n10771));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_37__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9960), .Y(n10768));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_38__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9969), .Y(n10765));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_38__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9963), .Y(n10762));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_39__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9972), .Y(n10759));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_39__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9966), .Y(n10756));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_40__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9975), .Y(n10753));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_40__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9969), .Y(n10750));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_41__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9978), .Y(n10747));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_41__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9972), .Y(n10744));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_42__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9981), .Y(n10741));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_42__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9975), .Y(n10738));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_43__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9984), .Y(n10735));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_43__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9978), .Y(n10732));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_44__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9987), .Y(n10729));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_44__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9981), .Y(n10726));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_45__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9990), .Y(n10723));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_45__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9984), .Y(n10720));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_46__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9993), .Y(n10717));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_46__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9987), .Y(n10714));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_47__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9996), .Y(n10711));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_47__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9990), .Y(n10708));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_48__p0_U6(.A(dpath_mulcore_b6[2]), .B(n9998), .Y(n10705));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_48__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9993), .Y(n10702));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_49__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10000), .Y(n10699));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_49__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9996), .Y(n10696));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_50__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10002), .Y(n10693));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_50__p1_U6(.A(dpath_mulcore_b7[2]), .B(n9998), .Y(n10690));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_51__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10004), .Y(n10687));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_51__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10000), .Y(n10684));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_52__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10006), .Y(n10681));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_52__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10002), .Y(n10678));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_53__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10009), .Y(n10675));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_53__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10004), .Y(n10672));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_54__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10012), .Y(n10669));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_54__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10006), .Y(n10666));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_55__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10015), .Y(n10663));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_55__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10009), .Y(n10660));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_56__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10018), .Y(n10657));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_56__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10012), .Y(n10654));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_57__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10021), .Y(n10651));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_57__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10015), .Y(n10648));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_58__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10024), .Y(n10645));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_58__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10018), .Y(n10642));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_59__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10028), .Y(n10639));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_59__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10021), .Y(n10636));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_60__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10029), .Y(n10633));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_60__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10024), .Y(n10630));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_61__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10030), .Y(n10627));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_61__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10028), .Y(n10624));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_62__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10031), .Y(n10621));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_62__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10029), .Y(n10618));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_63__p0_U6(.A(dpath_mulcore_b6[2]), .B(n10032), .Y(n10615));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I1_63__p1_U6(.A(dpath_mulcore_b7[2]), .B(n10030), .Y(n10612));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I2_p1_64__U6(.A(dpath_mulcore_b7[2]), .B(n10031), .Y(n10609));
XOR2X1 mul_dpath_mulcore_ary1_a0_I2_I2_p1_65__U6(.A(dpath_mulcore_b7[2]), .B(n10032), .Y(n10606));
OR2X1 mul_U1(.A(acc_actc3), .B(acc_actc2), .Y(control_n10));
AND2X1 mul_U2(.A(n2964), .B(n4640), .Y(dpath_n850));
AND2X1 mul_U3(.A(n2966), .B(n4642), .Y(dpath_n856));
AND2X1 mul_U4(.A(n2968), .B(n4644), .Y(dpath_n862));
AND2X1 mul_U5(.A(n2970), .B(n4646), .Y(dpath_n868));
AND2X1 mul_U6(.A(n2972), .B(n4648), .Y(dpath_n874));
AND2X1 mul_U7(.A(n2974), .B(n4650), .Y(dpath_n880));
AND2X1 mul_U8(.A(n2976), .B(n4652), .Y(dpath_n886));
AND2X1 mul_U9(.A(n2978), .B(n4654), .Y(dpath_n892));
AND2X1 mul_U10(.A(n2980), .B(n4656), .Y(dpath_n898));
AND2X1 mul_U11(.A(n2982), .B(n4658), .Y(dpath_n904));
AND2X1 mul_U12(.A(n2986), .B(n4662), .Y(dpath_n916));
AND2X1 mul_U13(.A(n2988), .B(n4664), .Y(dpath_n922));
AND2X1 mul_U14(.A(n2990), .B(n4666), .Y(dpath_n928));
AND2X1 mul_U15(.A(n2996), .B(n4672), .Y(dpath_n946));
AND2X1 mul_U16(.A(n2998), .B(n4674), .Y(dpath_n952));
AND2X1 mul_U17(.A(n3000), .B(n4676), .Y(dpath_n958));
AND2X1 mul_U18(.A(n3002), .B(n4678), .Y(dpath_n964));
AND2X1 mul_U19(.A(n3004), .B(n4680), .Y(dpath_n970));
AND2X1 mul_U20(.A(n2879), .B(n4555), .Y(dpath_n654));
AND2X1 mul_U21(.A(n2888), .B(n4564), .Y(dpath_n680));
AND2X1 mul_U22(.A(n2900), .B(n4576), .Y(dpath_n706));
AND2X1 mul_U23(.A(n2912), .B(n4588), .Y(dpath_n732));
AND2X1 mul_U24(.A(n2924), .B(n4600), .Y(dpath_n758));
AND2X1 mul_U25(.A(n2936), .B(n4612), .Y(dpath_n784));
AND2X1 mul_U26(.A(n2948), .B(n4624), .Y(dpath_n810));
AND2X1 mul_U27(.A(n2962), .B(n4638), .Y(dpath_n844));
OR2X1 mul_U28(.A(acc_actc3), .B(acc_actc2), .Y(dpath_n980));
AND2X1 mul_U29(.A(n923), .B(n13097), .Y(dpath_mulcore_ary1_a1_I0_I2_net43));
OR2X1 mul_U30(.A(n7004), .B(dpath_mulcore_b9[0]), .Y(n13097));
AND2X1 mul_U31(.A(n1121), .B(n13685), .Y(dpath_mulcore_ary1_a1_I0_I2_net47));
OR2X1 mul_U32(.A(n9481), .B(dpath_mulcore_b8[0]), .Y(n13685));
AND2X1 mul_U33(.A(n924), .B(n13100), .Y(dpath_mulcore_ary1_a1_I0_I2_net48));
OR2X1 mul_U34(.A(n7005), .B(dpath_mulcore_b9[0]), .Y(n13100));
AND2X1 mul_U35(.A(n928), .B(n13112), .Y(dpath_mulcore_ary1_a1_I0_I1_63__net32));
OR2X1 mul_U36(.A(n7009), .B(dpath_mulcore_b8[0]), .Y(n13112));
AND2X1 mul_U37(.A(n927), .B(n13109), .Y(dpath_mulcore_ary1_a1_I0_I1_63__net046));
OR2X1 mul_U38(.A(n7008), .B(dpath_mulcore_b9[0]), .Y(n13109));
AND2X1 mul_U39(.A(n931), .B(n13121), .Y(dpath_mulcore_ary1_a1_I0_I1_62__net32));
OR2X1 mul_U40(.A(n7012), .B(dpath_mulcore_b8[0]), .Y(n13121));
AND2X1 mul_U41(.A(n930), .B(n13118), .Y(dpath_mulcore_ary1_a1_I0_I1_62__net046));
OR2X1 mul_U42(.A(n7011), .B(dpath_mulcore_b9[0]), .Y(n13118));
AND2X1 mul_U43(.A(n934), .B(n13130), .Y(dpath_mulcore_ary1_a1_I0_I1_61__net32));
OR2X1 mul_U44(.A(n7015), .B(dpath_mulcore_b8[0]), .Y(n13130));
AND2X1 mul_U45(.A(n933), .B(n13127), .Y(dpath_mulcore_ary1_a1_I0_I1_61__net046));
OR2X1 mul_U46(.A(n7014), .B(dpath_mulcore_b9[0]), .Y(n13127));
AND2X1 mul_U47(.A(n937), .B(n13139), .Y(dpath_mulcore_ary1_a1_I0_I1_60__net32));
OR2X1 mul_U48(.A(n7018), .B(dpath_mulcore_b8[0]), .Y(n13139));
AND2X1 mul_U49(.A(n936), .B(n13136), .Y(dpath_mulcore_ary1_a1_I0_I1_60__net046));
OR2X1 mul_U50(.A(n7017), .B(dpath_mulcore_b9[0]), .Y(n13136));
AND2X1 mul_U51(.A(n940), .B(n13148), .Y(dpath_mulcore_ary1_a1_I0_I1_59__net32));
OR2X1 mul_U52(.A(n7021), .B(dpath_mulcore_b8[0]), .Y(n13148));
AND2X1 mul_U53(.A(n939), .B(n13145), .Y(dpath_mulcore_ary1_a1_I0_I1_59__net046));
OR2X1 mul_U54(.A(n7020), .B(dpath_mulcore_b9[0]), .Y(n13145));
AND2X1 mul_U55(.A(n943), .B(n13157), .Y(dpath_mulcore_ary1_a1_I0_I1_58__net32));
OR2X1 mul_U56(.A(n7024), .B(dpath_mulcore_b8[0]), .Y(n13157));
AND2X1 mul_U57(.A(n942), .B(n13154), .Y(dpath_mulcore_ary1_a1_I0_I1_58__net046));
OR2X1 mul_U58(.A(n7023), .B(dpath_mulcore_b9[0]), .Y(n13154));
AND2X1 mul_U59(.A(n946), .B(n13166), .Y(dpath_mulcore_ary1_a1_I0_I1_57__net32));
OR2X1 mul_U60(.A(n7027), .B(dpath_mulcore_b8[0]), .Y(n13166));
AND2X1 mul_U61(.A(n945), .B(n13163), .Y(dpath_mulcore_ary1_a1_I0_I1_57__net046));
OR2X1 mul_U62(.A(n7026), .B(dpath_mulcore_b9[0]), .Y(n13163));
AND2X1 mul_U63(.A(n949), .B(n13175), .Y(dpath_mulcore_ary1_a1_I0_I1_56__net32));
OR2X1 mul_U64(.A(n7030), .B(dpath_mulcore_b8[0]), .Y(n13175));
AND2X1 mul_U65(.A(n948), .B(n13172), .Y(dpath_mulcore_ary1_a1_I0_I1_56__net046));
OR2X1 mul_U66(.A(n7029), .B(dpath_mulcore_b9[0]), .Y(n13172));
AND2X1 mul_U67(.A(n952), .B(n13184), .Y(dpath_mulcore_ary1_a1_I0_I1_55__net32));
OR2X1 mul_U68(.A(n7033), .B(dpath_mulcore_b8[0]), .Y(n13184));
AND2X1 mul_U69(.A(n951), .B(n13181), .Y(dpath_mulcore_ary1_a1_I0_I1_55__net046));
OR2X1 mul_U70(.A(n7032), .B(dpath_mulcore_b9[0]), .Y(n13181));
AND2X1 mul_U71(.A(n955), .B(n13193), .Y(dpath_mulcore_ary1_a1_I0_I1_54__net32));
OR2X1 mul_U72(.A(n7036), .B(dpath_mulcore_b8[0]), .Y(n13193));
AND2X1 mul_U73(.A(n954), .B(n13190), .Y(dpath_mulcore_ary1_a1_I0_I1_54__net046));
OR2X1 mul_U74(.A(n7035), .B(dpath_mulcore_b9[0]), .Y(n13190));
AND2X1 mul_U75(.A(n958), .B(n13202), .Y(dpath_mulcore_ary1_a1_I0_I1_53__net32));
OR2X1 mul_U76(.A(n7039), .B(dpath_mulcore_b8[0]), .Y(n13202));
AND2X1 mul_U77(.A(n957), .B(n13199), .Y(dpath_mulcore_ary1_a1_I0_I1_53__net046));
OR2X1 mul_U78(.A(n7038), .B(dpath_mulcore_b9[0]), .Y(n13199));
AND2X1 mul_U79(.A(n961), .B(n13211), .Y(dpath_mulcore_ary1_a1_I0_I1_52__net32));
OR2X1 mul_U80(.A(n7042), .B(dpath_mulcore_b8[0]), .Y(n13211));
AND2X1 mul_U81(.A(n960), .B(n13208), .Y(dpath_mulcore_ary1_a1_I0_I1_52__net046));
OR2X1 mul_U82(.A(n7041), .B(dpath_mulcore_b9[0]), .Y(n13208));
AND2X1 mul_U83(.A(n964), .B(n13220), .Y(dpath_mulcore_ary1_a1_I0_I1_51__net32));
OR2X1 mul_U84(.A(n7045), .B(dpath_mulcore_b8[0]), .Y(n13220));
AND2X1 mul_U85(.A(n963), .B(n13217), .Y(dpath_mulcore_ary1_a1_I0_I1_51__net046));
OR2X1 mul_U86(.A(n7044), .B(dpath_mulcore_b9[0]), .Y(n13217));
AND2X1 mul_U87(.A(n967), .B(n13229), .Y(dpath_mulcore_ary1_a1_I0_I1_50__net32));
OR2X1 mul_U88(.A(n7048), .B(dpath_mulcore_b8[0]), .Y(n13229));
AND2X1 mul_U89(.A(n966), .B(n13226), .Y(dpath_mulcore_ary1_a1_I0_I1_50__net046));
OR2X1 mul_U90(.A(n7047), .B(dpath_mulcore_b9[0]), .Y(n13226));
AND2X1 mul_U91(.A(n970), .B(n13238), .Y(dpath_mulcore_ary1_a1_I0_I1_49__net32));
OR2X1 mul_U92(.A(n7051), .B(dpath_mulcore_b8[0]), .Y(n13238));
AND2X1 mul_U93(.A(n969), .B(n13235), .Y(dpath_mulcore_ary1_a1_I0_I1_49__net046));
OR2X1 mul_U94(.A(n7050), .B(dpath_mulcore_b9[0]), .Y(n13235));
AND2X1 mul_U95(.A(n973), .B(n13247), .Y(dpath_mulcore_ary1_a1_I0_I1_48__net32));
OR2X1 mul_U96(.A(n7054), .B(dpath_mulcore_b8[0]), .Y(n13247));
AND2X1 mul_U97(.A(n972), .B(n13244), .Y(dpath_mulcore_ary1_a1_I0_I1_48__net046));
OR2X1 mul_U98(.A(n7053), .B(dpath_mulcore_b9[0]), .Y(n13244));
AND2X1 mul_U99(.A(n976), .B(n13256), .Y(dpath_mulcore_ary1_a1_I0_I1_47__net32));
OR2X1 mul_U100(.A(n7057), .B(dpath_mulcore_b8[0]), .Y(n13256));
AND2X1 mul_U101(.A(n975), .B(n13253), .Y(dpath_mulcore_ary1_a1_I0_I1_47__net046));
OR2X1 mul_U102(.A(n7056), .B(dpath_mulcore_b9[0]), .Y(n13253));
AND2X1 mul_U103(.A(n979), .B(n13265), .Y(dpath_mulcore_ary1_a1_I0_I1_46__net32));
OR2X1 mul_U104(.A(n7060), .B(dpath_mulcore_b8[0]), .Y(n13265));
AND2X1 mul_U105(.A(n978), .B(n13262), .Y(dpath_mulcore_ary1_a1_I0_I1_46__net046));
OR2X1 mul_U106(.A(n7059), .B(dpath_mulcore_b9[0]), .Y(n13262));
AND2X1 mul_U107(.A(n982), .B(n13274), .Y(dpath_mulcore_ary1_a1_I0_I1_45__net32));
OR2X1 mul_U108(.A(n7063), .B(dpath_mulcore_b8[0]), .Y(n13274));
AND2X1 mul_U109(.A(n981), .B(n13271), .Y(dpath_mulcore_ary1_a1_I0_I1_45__net046));
OR2X1 mul_U110(.A(n7062), .B(dpath_mulcore_b9[0]), .Y(n13271));
AND2X1 mul_U111(.A(n985), .B(n13283), .Y(dpath_mulcore_ary1_a1_I0_I1_44__net32));
OR2X1 mul_U112(.A(n7066), .B(dpath_mulcore_b8[0]), .Y(n13283));
AND2X1 mul_U113(.A(n984), .B(n13280), .Y(dpath_mulcore_ary1_a1_I0_I1_44__net046));
OR2X1 mul_U114(.A(n7065), .B(dpath_mulcore_b9[0]), .Y(n13280));
AND2X1 mul_U115(.A(n988), .B(n13292), .Y(dpath_mulcore_ary1_a1_I0_I1_43__net32));
OR2X1 mul_U116(.A(n7069), .B(dpath_mulcore_b8[0]), .Y(n13292));
AND2X1 mul_U117(.A(n987), .B(n13289), .Y(dpath_mulcore_ary1_a1_I0_I1_43__net046));
OR2X1 mul_U118(.A(n7068), .B(dpath_mulcore_b9[0]), .Y(n13289));
AND2X1 mul_U119(.A(n991), .B(n13301), .Y(dpath_mulcore_ary1_a1_I0_I1_42__net32));
OR2X1 mul_U120(.A(n7072), .B(dpath_mulcore_b8[0]), .Y(n13301));
AND2X1 mul_U121(.A(n990), .B(n13298), .Y(dpath_mulcore_ary1_a1_I0_I1_42__net046));
OR2X1 mul_U122(.A(n7071), .B(dpath_mulcore_b9[0]), .Y(n13298));
AND2X1 mul_U123(.A(n994), .B(n13310), .Y(dpath_mulcore_ary1_a1_I0_I1_41__net32));
OR2X1 mul_U124(.A(n7075), .B(dpath_mulcore_b8[0]), .Y(n13310));
AND2X1 mul_U125(.A(n993), .B(n13307), .Y(dpath_mulcore_ary1_a1_I0_I1_41__net046));
OR2X1 mul_U126(.A(n7074), .B(dpath_mulcore_b9[0]), .Y(n13307));
AND2X1 mul_U127(.A(n997), .B(n13319), .Y(dpath_mulcore_ary1_a1_I0_I1_40__net32));
OR2X1 mul_U128(.A(n7078), .B(dpath_mulcore_b8[0]), .Y(n13319));
AND2X1 mul_U129(.A(n996), .B(n13316), .Y(dpath_mulcore_ary1_a1_I0_I1_40__net046));
OR2X1 mul_U130(.A(n7077), .B(dpath_mulcore_b9[0]), .Y(n13316));
AND2X1 mul_U131(.A(n1000), .B(n13328), .Y(dpath_mulcore_ary1_a1_I0_I1_39__net32));
OR2X1 mul_U132(.A(n7081), .B(dpath_mulcore_b8[0]), .Y(n13328));
AND2X1 mul_U133(.A(n999), .B(n13325), .Y(dpath_mulcore_ary1_a1_I0_I1_39__net046));
OR2X1 mul_U134(.A(n7080), .B(dpath_mulcore_b9[0]), .Y(n13325));
AND2X1 mul_U135(.A(n1003), .B(n13337), .Y(dpath_mulcore_ary1_a1_I0_I1_38__net32));
OR2X1 mul_U136(.A(n7084), .B(dpath_mulcore_b8[0]), .Y(n13337));
AND2X1 mul_U137(.A(n1002), .B(n13334), .Y(dpath_mulcore_ary1_a1_I0_I1_38__net046));
OR2X1 mul_U138(.A(n7083), .B(dpath_mulcore_b9[0]), .Y(n13334));
AND2X1 mul_U139(.A(n1006), .B(n13346), .Y(dpath_mulcore_ary1_a1_I0_I1_37__net32));
OR2X1 mul_U140(.A(n7087), .B(dpath_mulcore_b8[0]), .Y(n13346));
AND2X1 mul_U141(.A(n1005), .B(n13343), .Y(dpath_mulcore_ary1_a1_I0_I1_37__net046));
OR2X1 mul_U142(.A(n7086), .B(dpath_mulcore_b9[0]), .Y(n13343));
AND2X1 mul_U143(.A(n1009), .B(n13355), .Y(dpath_mulcore_ary1_a1_I0_I1_36__net32));
OR2X1 mul_U144(.A(n7090), .B(dpath_mulcore_b8[0]), .Y(n13355));
AND2X1 mul_U145(.A(n1008), .B(n13352), .Y(dpath_mulcore_ary1_a1_I0_I1_36__net046));
OR2X1 mul_U146(.A(n7089), .B(dpath_mulcore_b9[0]), .Y(n13352));
AND2X1 mul_U147(.A(n1012), .B(n13364), .Y(dpath_mulcore_ary1_a1_I0_I1_35__net32));
OR2X1 mul_U148(.A(n7093), .B(dpath_mulcore_b8[0]), .Y(n13364));
AND2X1 mul_U149(.A(n1011), .B(n13361), .Y(dpath_mulcore_ary1_a1_I0_I1_35__net046));
OR2X1 mul_U150(.A(n7092), .B(dpath_mulcore_b9[0]), .Y(n13361));
AND2X1 mul_U151(.A(n1015), .B(n13373), .Y(dpath_mulcore_ary1_a1_I0_I1_34__net32));
OR2X1 mul_U152(.A(n7096), .B(dpath_mulcore_b8[0]), .Y(n13373));
AND2X1 mul_U153(.A(n1014), .B(n13370), .Y(dpath_mulcore_ary1_a1_I0_I1_34__net046));
OR2X1 mul_U154(.A(n7095), .B(dpath_mulcore_b9[0]), .Y(n13370));
AND2X1 mul_U155(.A(n1018), .B(n13382), .Y(dpath_mulcore_ary1_a1_I0_I1_33__net32));
OR2X1 mul_U156(.A(n7099), .B(dpath_mulcore_b8[0]), .Y(n13382));
AND2X1 mul_U157(.A(n1017), .B(n13379), .Y(dpath_mulcore_ary1_a1_I0_I1_33__net046));
OR2X1 mul_U158(.A(n7098), .B(dpath_mulcore_b9[0]), .Y(n13379));
AND2X1 mul_U159(.A(n1021), .B(n13391), .Y(dpath_mulcore_ary1_a1_I0_I1_32__net32));
OR2X1 mul_U160(.A(n7102), .B(dpath_mulcore_b8[0]), .Y(n13391));
AND2X1 mul_U161(.A(n1020), .B(n13388), .Y(dpath_mulcore_ary1_a1_I0_I1_32__net046));
OR2X1 mul_U162(.A(n7101), .B(dpath_mulcore_b9[0]), .Y(n13388));
AND2X1 mul_U163(.A(n1024), .B(n13400), .Y(dpath_mulcore_ary1_a1_I0_I1_31__net32));
OR2X1 mul_U164(.A(n7105), .B(dpath_mulcore_b8[0]), .Y(n13400));
AND2X1 mul_U165(.A(n1023), .B(n13397), .Y(dpath_mulcore_ary1_a1_I0_I1_31__net046));
OR2X1 mul_U166(.A(n7104), .B(dpath_mulcore_b9[0]), .Y(n13397));
AND2X1 mul_U167(.A(n1027), .B(n13409), .Y(dpath_mulcore_ary1_a1_I0_I1_30__net32));
OR2X1 mul_U168(.A(n7108), .B(dpath_mulcore_b8[0]), .Y(n13409));
AND2X1 mul_U169(.A(n1026), .B(n13406), .Y(dpath_mulcore_ary1_a1_I0_I1_30__net046));
OR2X1 mul_U170(.A(n7107), .B(dpath_mulcore_b9[0]), .Y(n13406));
AND2X1 mul_U171(.A(n1030), .B(n13418), .Y(dpath_mulcore_ary1_a1_I0_I1_29__net32));
OR2X1 mul_U172(.A(n7111), .B(dpath_mulcore_b8[0]), .Y(n13418));
AND2X1 mul_U173(.A(n1029), .B(n13415), .Y(dpath_mulcore_ary1_a1_I0_I1_29__net046));
OR2X1 mul_U174(.A(n7110), .B(dpath_mulcore_b9[0]), .Y(n13415));
AND2X1 mul_U175(.A(n1033), .B(n13427), .Y(dpath_mulcore_ary1_a1_I0_I1_28__net32));
OR2X1 mul_U176(.A(n7114), .B(dpath_mulcore_b8[0]), .Y(n13427));
AND2X1 mul_U177(.A(n1032), .B(n13424), .Y(dpath_mulcore_ary1_a1_I0_I1_28__net046));
OR2X1 mul_U178(.A(n7113), .B(dpath_mulcore_b9[0]), .Y(n13424));
AND2X1 mul_U179(.A(n1036), .B(n13436), .Y(dpath_mulcore_ary1_a1_I0_I1_27__net32));
OR2X1 mul_U180(.A(n7117), .B(dpath_mulcore_b8[0]), .Y(n13436));
AND2X1 mul_U181(.A(n1035), .B(n13433), .Y(dpath_mulcore_ary1_a1_I0_I1_27__net046));
OR2X1 mul_U182(.A(n7116), .B(dpath_mulcore_b9[0]), .Y(n13433));
AND2X1 mul_U183(.A(n1039), .B(n13445), .Y(dpath_mulcore_ary1_a1_I0_I1_26__net32));
OR2X1 mul_U184(.A(n7120), .B(dpath_mulcore_b8[0]), .Y(n13445));
AND2X1 mul_U185(.A(n1038), .B(n13442), .Y(dpath_mulcore_ary1_a1_I0_I1_26__net046));
OR2X1 mul_U186(.A(n7119), .B(dpath_mulcore_b9[0]), .Y(n13442));
AND2X1 mul_U187(.A(n1042), .B(n13454), .Y(dpath_mulcore_ary1_a1_I0_I1_25__net32));
OR2X1 mul_U188(.A(n7123), .B(dpath_mulcore_b8[0]), .Y(n13454));
AND2X1 mul_U189(.A(n1041), .B(n13451), .Y(dpath_mulcore_ary1_a1_I0_I1_25__net046));
OR2X1 mul_U190(.A(n7122), .B(dpath_mulcore_b9[0]), .Y(n13451));
AND2X1 mul_U191(.A(n1045), .B(n13463), .Y(dpath_mulcore_ary1_a1_I0_I1_24__net32));
OR2X1 mul_U192(.A(n7126), .B(dpath_mulcore_b8[0]), .Y(n13463));
AND2X1 mul_U193(.A(n1044), .B(n13460), .Y(dpath_mulcore_ary1_a1_I0_I1_24__net046));
OR2X1 mul_U194(.A(n7125), .B(dpath_mulcore_b9[0]), .Y(n13460));
AND2X1 mul_U195(.A(n1048), .B(n13472), .Y(dpath_mulcore_ary1_a1_I0_I1_23__net32));
OR2X1 mul_U196(.A(n7129), .B(dpath_mulcore_b8[0]), .Y(n13472));
AND2X1 mul_U197(.A(n1047), .B(n13469), .Y(dpath_mulcore_ary1_a1_I0_I1_23__net046));
OR2X1 mul_U198(.A(n7128), .B(dpath_mulcore_b9[0]), .Y(n13469));
AND2X1 mul_U199(.A(n1051), .B(n13481), .Y(dpath_mulcore_ary1_a1_I0_I1_22__net32));
OR2X1 mul_U200(.A(n7132), .B(dpath_mulcore_b8[0]), .Y(n13481));
AND2X1 mul_U201(.A(n1050), .B(n13478), .Y(dpath_mulcore_ary1_a1_I0_I1_22__net046));
OR2X1 mul_U202(.A(n7131), .B(dpath_mulcore_b9[0]), .Y(n13478));
AND2X1 mul_U203(.A(n1054), .B(n13490), .Y(dpath_mulcore_ary1_a1_I0_I1_21__net32));
OR2X1 mul_U204(.A(n7135), .B(dpath_mulcore_b8[0]), .Y(n13490));
AND2X1 mul_U205(.A(n1053), .B(n13487), .Y(dpath_mulcore_ary1_a1_I0_I1_21__net046));
OR2X1 mul_U206(.A(n7134), .B(dpath_mulcore_b9[0]), .Y(n13487));
AND2X1 mul_U207(.A(n1057), .B(n13499), .Y(dpath_mulcore_ary1_a1_I0_I1_20__net32));
OR2X1 mul_U208(.A(n7138), .B(dpath_mulcore_b8[0]), .Y(n13499));
AND2X1 mul_U209(.A(n1056), .B(n13496), .Y(dpath_mulcore_ary1_a1_I0_I1_20__net046));
OR2X1 mul_U210(.A(n7137), .B(dpath_mulcore_b9[0]), .Y(n13496));
AND2X1 mul_U211(.A(n1060), .B(n13508), .Y(dpath_mulcore_ary1_a1_I0_I1_19__net32));
OR2X1 mul_U212(.A(n7141), .B(dpath_mulcore_b8[0]), .Y(n13508));
AND2X1 mul_U213(.A(n1059), .B(n13505), .Y(dpath_mulcore_ary1_a1_I0_I1_19__net046));
OR2X1 mul_U214(.A(n7140), .B(dpath_mulcore_b9[0]), .Y(n13505));
AND2X1 mul_U215(.A(n1063), .B(n13517), .Y(dpath_mulcore_ary1_a1_I0_I1_18__net32));
OR2X1 mul_U216(.A(n7144), .B(dpath_mulcore_b8[0]), .Y(n13517));
AND2X1 mul_U217(.A(n1062), .B(n13514), .Y(dpath_mulcore_ary1_a1_I0_I1_18__net046));
OR2X1 mul_U218(.A(n7143), .B(dpath_mulcore_b9[0]), .Y(n13514));
AND2X1 mul_U219(.A(n1066), .B(n13526), .Y(dpath_mulcore_ary1_a1_I0_I1_17__net32));
OR2X1 mul_U220(.A(n7147), .B(dpath_mulcore_b8[0]), .Y(n13526));
AND2X1 mul_U221(.A(n1065), .B(n13523), .Y(dpath_mulcore_ary1_a1_I0_I1_17__net046));
OR2X1 mul_U222(.A(n7146), .B(dpath_mulcore_b9[0]), .Y(n13523));
AND2X1 mul_U223(.A(n1069), .B(n13535), .Y(dpath_mulcore_ary1_a1_I0_I1_16__net32));
OR2X1 mul_U224(.A(n7150), .B(dpath_mulcore_b8[0]), .Y(n13535));
AND2X1 mul_U225(.A(n1068), .B(n13532), .Y(dpath_mulcore_ary1_a1_I0_I1_16__net046));
OR2X1 mul_U226(.A(n7149), .B(dpath_mulcore_b9[0]), .Y(n13532));
AND2X1 mul_U227(.A(n1072), .B(n13544), .Y(dpath_mulcore_ary1_a1_I0_I1_15__net32));
OR2X1 mul_U228(.A(n7153), .B(dpath_mulcore_b8[0]), .Y(n13544));
AND2X1 mul_U229(.A(n1071), .B(n13541), .Y(dpath_mulcore_ary1_a1_I0_I1_15__net046));
OR2X1 mul_U230(.A(n7152), .B(dpath_mulcore_b9[0]), .Y(n13541));
AND2X1 mul_U231(.A(n1075), .B(n13553), .Y(dpath_mulcore_ary1_a1_I0_I1_14__net32));
OR2X1 mul_U232(.A(n7156), .B(dpath_mulcore_b8[0]), .Y(n13553));
AND2X1 mul_U233(.A(n1074), .B(n13550), .Y(dpath_mulcore_ary1_a1_I0_I1_14__net046));
OR2X1 mul_U234(.A(n7155), .B(dpath_mulcore_b9[0]), .Y(n13550));
AND2X1 mul_U235(.A(n610), .B(n12148), .Y(dpath_mulcore_ary1_a1_I2_I1_62__net32));
OR2X1 mul_U236(.A(n6686), .B(dpath_mulcore_b14[0]), .Y(n12148));
AND2X1 mul_U237(.A(n609), .B(n12145), .Y(dpath_mulcore_ary1_a1_I2_I1_62__net046));
OR2X1 mul_U238(.A(n6685), .B(dpath_mulcore_b15[0]), .Y(n12145));
INVX1 mul_U239(.A(dpath_mulcore_op1_l[58]), .Y(n10024));
AND2X1 mul_U240(.A(n612), .B(n12154), .Y(dpath_mulcore_ary1_a1_I2_I1_61__net32));
OR2X1 mul_U241(.A(n6688), .B(dpath_mulcore_b14[0]), .Y(n12154));
AND2X1 mul_U242(.A(n611), .B(n12151), .Y(dpath_mulcore_ary1_a1_I2_I1_61__net046));
OR2X1 mul_U243(.A(n6687), .B(dpath_mulcore_b15[0]), .Y(n12151));
INVX1 mul_U244(.A(dpath_mulcore_op1_l[57]), .Y(n10021));
AND2X1 mul_U245(.A(n614), .B(n12160), .Y(dpath_mulcore_ary1_a1_I2_I1_60__net32));
OR2X1 mul_U246(.A(n6690), .B(dpath_mulcore_b14[0]), .Y(n12160));
AND2X1 mul_U247(.A(n613), .B(n12157), .Y(dpath_mulcore_ary1_a1_I2_I1_60__net046));
OR2X1 mul_U248(.A(n6689), .B(dpath_mulcore_b15[0]), .Y(n12157));
INVX1 mul_U249(.A(dpath_mulcore_op1_l[56]), .Y(n10018));
AND2X1 mul_U250(.A(n616), .B(n12166), .Y(dpath_mulcore_ary1_a1_I2_I1_59__net32));
OR2X1 mul_U251(.A(n6692), .B(dpath_mulcore_b14[0]), .Y(n12166));
AND2X1 mul_U252(.A(n615), .B(n12163), .Y(dpath_mulcore_ary1_a1_I2_I1_59__net046));
OR2X1 mul_U253(.A(n6691), .B(dpath_mulcore_b15[0]), .Y(n12163));
INVX1 mul_U254(.A(dpath_mulcore_op1_l[55]), .Y(n10015));
AND2X1 mul_U255(.A(n618), .B(n12172), .Y(dpath_mulcore_ary1_a1_I2_I1_58__net32));
OR2X1 mul_U256(.A(n6694), .B(dpath_mulcore_b14[0]), .Y(n12172));
AND2X1 mul_U257(.A(n617), .B(n12169), .Y(dpath_mulcore_ary1_a1_I2_I1_58__net046));
OR2X1 mul_U258(.A(n6693), .B(dpath_mulcore_b15[0]), .Y(n12169));
INVX1 mul_U259(.A(dpath_mulcore_op1_l[54]), .Y(n10012));
AND2X1 mul_U260(.A(n620), .B(n12178), .Y(dpath_mulcore_ary1_a1_I2_I1_57__net32));
OR2X1 mul_U261(.A(n6696), .B(dpath_mulcore_b14[0]), .Y(n12178));
AND2X1 mul_U262(.A(n619), .B(n12175), .Y(dpath_mulcore_ary1_a1_I2_I1_57__net046));
OR2X1 mul_U263(.A(n6695), .B(dpath_mulcore_b15[0]), .Y(n12175));
INVX1 mul_U264(.A(dpath_mulcore_op1_l[53]), .Y(n10009));
AND2X1 mul_U265(.A(n622), .B(n12184), .Y(dpath_mulcore_ary1_a1_I2_I1_56__net32));
OR2X1 mul_U266(.A(n6698), .B(dpath_mulcore_b14[0]), .Y(n12184));
AND2X1 mul_U267(.A(n621), .B(n12181), .Y(dpath_mulcore_ary1_a1_I2_I1_56__net046));
OR2X1 mul_U268(.A(n6697), .B(dpath_mulcore_b15[0]), .Y(n12181));
INVX1 mul_U269(.A(dpath_mulcore_op1_l[52]), .Y(n10006));
AND2X1 mul_U270(.A(n624), .B(n12190), .Y(dpath_mulcore_ary1_a1_I2_I1_55__net32));
OR2X1 mul_U271(.A(n6700), .B(dpath_mulcore_b14[0]), .Y(n12190));
AND2X1 mul_U272(.A(n623), .B(n12187), .Y(dpath_mulcore_ary1_a1_I2_I1_55__net046));
OR2X1 mul_U273(.A(n6699), .B(dpath_mulcore_b15[0]), .Y(n12187));
INVX1 mul_U274(.A(dpath_mulcore_op1_l[51]), .Y(n10004));
AND2X1 mul_U275(.A(n626), .B(n12196), .Y(dpath_mulcore_ary1_a1_I2_I1_54__net32));
OR2X1 mul_U276(.A(n6702), .B(dpath_mulcore_b14[0]), .Y(n12196));
AND2X1 mul_U277(.A(n625), .B(n12193), .Y(dpath_mulcore_ary1_a1_I2_I1_54__net046));
OR2X1 mul_U278(.A(n6701), .B(dpath_mulcore_b15[0]), .Y(n12193));
INVX1 mul_U279(.A(dpath_mulcore_op1_l[50]), .Y(n10002));
AND2X1 mul_U280(.A(n628), .B(n12202), .Y(dpath_mulcore_ary1_a1_I2_I1_53__net32));
OR2X1 mul_U281(.A(n6704), .B(dpath_mulcore_b14[0]), .Y(n12202));
AND2X1 mul_U282(.A(n627), .B(n12199), .Y(dpath_mulcore_ary1_a1_I2_I1_53__net046));
OR2X1 mul_U283(.A(n6703), .B(dpath_mulcore_b15[0]), .Y(n12199));
INVX1 mul_U284(.A(dpath_mulcore_op1_l[49]), .Y(n10000));
AND2X1 mul_U285(.A(n630), .B(n12208), .Y(dpath_mulcore_ary1_a1_I2_I1_52__net32));
OR2X1 mul_U286(.A(n6706), .B(dpath_mulcore_b14[0]), .Y(n12208));
AND2X1 mul_U287(.A(n629), .B(n12205), .Y(dpath_mulcore_ary1_a1_I2_I1_52__net046));
OR2X1 mul_U288(.A(n6705), .B(dpath_mulcore_b15[0]), .Y(n12205));
INVX1 mul_U289(.A(dpath_mulcore_op1_l[48]), .Y(n9998));
AND2X1 mul_U290(.A(n632), .B(n12214), .Y(dpath_mulcore_ary1_a1_I2_I1_51__net32));
OR2X1 mul_U291(.A(n6708), .B(dpath_mulcore_b14[0]), .Y(n12214));
AND2X1 mul_U292(.A(n631), .B(n12211), .Y(dpath_mulcore_ary1_a1_I2_I1_51__net046));
OR2X1 mul_U293(.A(n6707), .B(dpath_mulcore_b15[0]), .Y(n12211));
INVX1 mul_U294(.A(dpath_mulcore_op1_l[47]), .Y(n9996));
AND2X1 mul_U295(.A(n634), .B(n12220), .Y(dpath_mulcore_ary1_a1_I2_I1_50__net32));
OR2X1 mul_U296(.A(n6710), .B(dpath_mulcore_b14[0]), .Y(n12220));
AND2X1 mul_U297(.A(n633), .B(n12217), .Y(dpath_mulcore_ary1_a1_I2_I1_50__net046));
OR2X1 mul_U298(.A(n6709), .B(dpath_mulcore_b15[0]), .Y(n12217));
INVX1 mul_U299(.A(dpath_mulcore_op1_l[46]), .Y(n9993));
AND2X1 mul_U300(.A(n636), .B(n12226), .Y(dpath_mulcore_ary1_a1_I2_I1_49__net32));
OR2X1 mul_U301(.A(n6712), .B(dpath_mulcore_b14[0]), .Y(n12226));
AND2X1 mul_U302(.A(n635), .B(n12223), .Y(dpath_mulcore_ary1_a1_I2_I1_49__net046));
OR2X1 mul_U303(.A(n6711), .B(dpath_mulcore_b15[0]), .Y(n12223));
INVX1 mul_U304(.A(dpath_mulcore_op1_l[45]), .Y(n9990));
AND2X1 mul_U305(.A(n638), .B(n12232), .Y(dpath_mulcore_ary1_a1_I2_I1_48__net32));
OR2X1 mul_U306(.A(n6714), .B(dpath_mulcore_b14[0]), .Y(n12232));
AND2X1 mul_U307(.A(n637), .B(n12229), .Y(dpath_mulcore_ary1_a1_I2_I1_48__net046));
OR2X1 mul_U308(.A(n6713), .B(dpath_mulcore_b15[0]), .Y(n12229));
INVX1 mul_U309(.A(dpath_mulcore_op1_l[44]), .Y(n9987));
AND2X1 mul_U310(.A(n640), .B(n12238), .Y(dpath_mulcore_ary1_a1_I2_I1_47__net32));
OR2X1 mul_U311(.A(n6716), .B(dpath_mulcore_b14[0]), .Y(n12238));
AND2X1 mul_U312(.A(n639), .B(n12235), .Y(dpath_mulcore_ary1_a1_I2_I1_47__net046));
OR2X1 mul_U313(.A(n6715), .B(dpath_mulcore_b15[0]), .Y(n12235));
INVX1 mul_U314(.A(dpath_mulcore_op1_l[43]), .Y(n9984));
AND2X1 mul_U315(.A(n642), .B(n12244), .Y(dpath_mulcore_ary1_a1_I2_I1_46__net32));
OR2X1 mul_U316(.A(n6718), .B(dpath_mulcore_b14[0]), .Y(n12244));
AND2X1 mul_U317(.A(n641), .B(n12241), .Y(dpath_mulcore_ary1_a1_I2_I1_46__net046));
OR2X1 mul_U318(.A(n6717), .B(dpath_mulcore_b15[0]), .Y(n12241));
INVX1 mul_U319(.A(dpath_mulcore_op1_l[42]), .Y(n9981));
AND2X1 mul_U320(.A(n644), .B(n12250), .Y(dpath_mulcore_ary1_a1_I2_I1_45__net32));
OR2X1 mul_U321(.A(n6720), .B(dpath_mulcore_b14[0]), .Y(n12250));
AND2X1 mul_U322(.A(n643), .B(n12247), .Y(dpath_mulcore_ary1_a1_I2_I1_45__net046));
OR2X1 mul_U323(.A(n6719), .B(dpath_mulcore_b15[0]), .Y(n12247));
INVX1 mul_U324(.A(dpath_mulcore_op1_l[41]), .Y(n9978));
AND2X1 mul_U325(.A(n646), .B(n12256), .Y(dpath_mulcore_ary1_a1_I2_I1_44__net32));
OR2X1 mul_U326(.A(n6722), .B(dpath_mulcore_b14[0]), .Y(n12256));
AND2X1 mul_U327(.A(n645), .B(n12253), .Y(dpath_mulcore_ary1_a1_I2_I1_44__net046));
OR2X1 mul_U328(.A(n6721), .B(dpath_mulcore_b15[0]), .Y(n12253));
INVX1 mul_U329(.A(dpath_mulcore_op1_l[40]), .Y(n9975));
AND2X1 mul_U330(.A(n648), .B(n12262), .Y(dpath_mulcore_ary1_a1_I2_I1_43__net32));
OR2X1 mul_U331(.A(n6724), .B(dpath_mulcore_b14[0]), .Y(n12262));
AND2X1 mul_U332(.A(n647), .B(n12259), .Y(dpath_mulcore_ary1_a1_I2_I1_43__net046));
OR2X1 mul_U333(.A(n6723), .B(dpath_mulcore_b15[0]), .Y(n12259));
INVX1 mul_U334(.A(dpath_mulcore_op1_l[39]), .Y(n9972));
AND2X1 mul_U335(.A(n650), .B(n12268), .Y(dpath_mulcore_ary1_a1_I2_I1_42__net32));
OR2X1 mul_U336(.A(n6726), .B(dpath_mulcore_b14[0]), .Y(n12268));
AND2X1 mul_U337(.A(n649), .B(n12265), .Y(dpath_mulcore_ary1_a1_I2_I1_42__net046));
OR2X1 mul_U338(.A(n6725), .B(dpath_mulcore_b15[0]), .Y(n12265));
INVX1 mul_U339(.A(dpath_mulcore_op1_l[38]), .Y(n9969));
AND2X1 mul_U340(.A(n652), .B(n12274), .Y(dpath_mulcore_ary1_a1_I2_I1_41__net32));
OR2X1 mul_U341(.A(n6728), .B(dpath_mulcore_b14[0]), .Y(n12274));
AND2X1 mul_U342(.A(n651), .B(n12271), .Y(dpath_mulcore_ary1_a1_I2_I1_41__net046));
OR2X1 mul_U343(.A(n6727), .B(dpath_mulcore_b15[0]), .Y(n12271));
INVX1 mul_U344(.A(dpath_mulcore_op1_l[37]), .Y(n9966));
AND2X1 mul_U345(.A(n654), .B(n12280), .Y(dpath_mulcore_ary1_a1_I2_I1_40__net32));
OR2X1 mul_U346(.A(n6730), .B(dpath_mulcore_b14[0]), .Y(n12280));
AND2X1 mul_U347(.A(n653), .B(n12277), .Y(dpath_mulcore_ary1_a1_I2_I1_40__net046));
OR2X1 mul_U348(.A(n6729), .B(dpath_mulcore_b15[0]), .Y(n12277));
INVX1 mul_U349(.A(dpath_mulcore_op1_l[36]), .Y(n9963));
AND2X1 mul_U350(.A(n656), .B(n12286), .Y(dpath_mulcore_ary1_a1_I2_I1_39__net32));
OR2X1 mul_U351(.A(n6732), .B(dpath_mulcore_b14[0]), .Y(n12286));
AND2X1 mul_U352(.A(n655), .B(n12283), .Y(dpath_mulcore_ary1_a1_I2_I1_39__net046));
OR2X1 mul_U353(.A(n6731), .B(dpath_mulcore_b15[0]), .Y(n12283));
INVX1 mul_U354(.A(dpath_mulcore_op1_l[35]), .Y(n9960));
AND2X1 mul_U355(.A(n658), .B(n12292), .Y(dpath_mulcore_ary1_a1_I2_I1_38__net32));
OR2X1 mul_U356(.A(n6734), .B(dpath_mulcore_b14[0]), .Y(n12292));
AND2X1 mul_U357(.A(n657), .B(n12289), .Y(dpath_mulcore_ary1_a1_I2_I1_38__net046));
OR2X1 mul_U358(.A(n6733), .B(dpath_mulcore_b15[0]), .Y(n12289));
INVX1 mul_U359(.A(dpath_mulcore_op1_l[34]), .Y(n9957));
AND2X1 mul_U360(.A(n660), .B(n12298), .Y(dpath_mulcore_ary1_a1_I2_I1_37__net32));
OR2X1 mul_U361(.A(n6736), .B(dpath_mulcore_b14[0]), .Y(n12298));
AND2X1 mul_U362(.A(n659), .B(n12295), .Y(dpath_mulcore_ary1_a1_I2_I1_37__net046));
OR2X1 mul_U363(.A(n6735), .B(dpath_mulcore_b15[0]), .Y(n12295));
INVX1 mul_U364(.A(dpath_mulcore_op1_l[33]), .Y(n9954));
AND2X1 mul_U365(.A(n662), .B(n12304), .Y(dpath_mulcore_ary1_a1_I2_I1_36__net32));
OR2X1 mul_U366(.A(n6738), .B(dpath_mulcore_b14[0]), .Y(n12304));
AND2X1 mul_U367(.A(n661), .B(n12301), .Y(dpath_mulcore_ary1_a1_I2_I1_36__net046));
OR2X1 mul_U368(.A(n6737), .B(dpath_mulcore_b15[0]), .Y(n12301));
INVX1 mul_U369(.A(dpath_mulcore_op1_l[32]), .Y(n9951));
AND2X1 mul_U370(.A(n664), .B(n12310), .Y(dpath_mulcore_ary1_a1_I2_I1_35__net32));
OR2X1 mul_U371(.A(n6740), .B(dpath_mulcore_b14[0]), .Y(n12310));
AND2X1 mul_U372(.A(n663), .B(n12307), .Y(dpath_mulcore_ary1_a1_I2_I1_35__net046));
OR2X1 mul_U373(.A(n6739), .B(dpath_mulcore_b15[0]), .Y(n12307));
INVX1 mul_U374(.A(dpath_mulcore_op1_l[31]), .Y(n9948));
AND2X1 mul_U375(.A(n666), .B(n12316), .Y(dpath_mulcore_ary1_a1_I2_I1_34__net32));
OR2X1 mul_U376(.A(n6742), .B(dpath_mulcore_b14[0]), .Y(n12316));
AND2X1 mul_U377(.A(n665), .B(n12313), .Y(dpath_mulcore_ary1_a1_I2_I1_34__net046));
OR2X1 mul_U378(.A(n6741), .B(dpath_mulcore_b15[0]), .Y(n12313));
INVX1 mul_U379(.A(dpath_mulcore_op1_l[30]), .Y(n9945));
AND2X1 mul_U380(.A(n668), .B(n12322), .Y(dpath_mulcore_ary1_a1_I2_I1_33__net32));
OR2X1 mul_U381(.A(n6744), .B(dpath_mulcore_b14[0]), .Y(n12322));
AND2X1 mul_U382(.A(n667), .B(n12319), .Y(dpath_mulcore_ary1_a1_I2_I1_33__net046));
OR2X1 mul_U383(.A(n6743), .B(dpath_mulcore_b15[0]), .Y(n12319));
INVX1 mul_U384(.A(dpath_mulcore_op1_l[29]), .Y(n9942));
AND2X1 mul_U385(.A(n670), .B(n12328), .Y(dpath_mulcore_ary1_a1_I2_I1_32__net32));
OR2X1 mul_U386(.A(n6746), .B(dpath_mulcore_b14[0]), .Y(n12328));
AND2X1 mul_U387(.A(n669), .B(n12325), .Y(dpath_mulcore_ary1_a1_I2_I1_32__net046));
OR2X1 mul_U388(.A(n6745), .B(dpath_mulcore_b15[0]), .Y(n12325));
INVX1 mul_U389(.A(dpath_mulcore_op1_l[28]), .Y(n9939));
AND2X1 mul_U390(.A(n672), .B(n12334), .Y(dpath_mulcore_ary1_a1_I2_I1_31__net32));
OR2X1 mul_U391(.A(n6748), .B(dpath_mulcore_b14[0]), .Y(n12334));
AND2X1 mul_U392(.A(n671), .B(n12331), .Y(dpath_mulcore_ary1_a1_I2_I1_31__net046));
OR2X1 mul_U393(.A(n6747), .B(dpath_mulcore_b15[0]), .Y(n12331));
INVX1 mul_U394(.A(dpath_mulcore_op1_l[27]), .Y(n9936));
AND2X1 mul_U395(.A(n674), .B(n12340), .Y(dpath_mulcore_ary1_a1_I2_I1_30__net32));
OR2X1 mul_U396(.A(n6750), .B(dpath_mulcore_b14[0]), .Y(n12340));
AND2X1 mul_U397(.A(n673), .B(n12337), .Y(dpath_mulcore_ary1_a1_I2_I1_30__net046));
OR2X1 mul_U398(.A(n6749), .B(dpath_mulcore_b15[0]), .Y(n12337));
INVX1 mul_U399(.A(dpath_mulcore_op1_l[26]), .Y(n9933));
AND2X1 mul_U400(.A(n676), .B(n12346), .Y(dpath_mulcore_ary1_a1_I2_I1_29__net32));
OR2X1 mul_U401(.A(n6752), .B(dpath_mulcore_b14[0]), .Y(n12346));
AND2X1 mul_U402(.A(n675), .B(n12343), .Y(dpath_mulcore_ary1_a1_I2_I1_29__net046));
OR2X1 mul_U403(.A(n6751), .B(dpath_mulcore_b15[0]), .Y(n12343));
INVX1 mul_U404(.A(dpath_mulcore_op1_l[25]), .Y(n9930));
AND2X1 mul_U405(.A(n678), .B(n12352), .Y(dpath_mulcore_ary1_a1_I2_I1_28__net32));
OR2X1 mul_U406(.A(n6754), .B(dpath_mulcore_b14[0]), .Y(n12352));
AND2X1 mul_U407(.A(n677), .B(n12349), .Y(dpath_mulcore_ary1_a1_I2_I1_28__net046));
OR2X1 mul_U408(.A(n6753), .B(dpath_mulcore_b15[0]), .Y(n12349));
INVX1 mul_U409(.A(dpath_mulcore_op1_l[24]), .Y(n9927));
AND2X1 mul_U410(.A(n680), .B(n12358), .Y(dpath_mulcore_ary1_a1_I2_I1_27__net32));
OR2X1 mul_U411(.A(n6756), .B(dpath_mulcore_b14[0]), .Y(n12358));
AND2X1 mul_U412(.A(n679), .B(n12355), .Y(dpath_mulcore_ary1_a1_I2_I1_27__net046));
OR2X1 mul_U413(.A(n6755), .B(dpath_mulcore_b15[0]), .Y(n12355));
INVX1 mul_U414(.A(dpath_mulcore_op1_l[23]), .Y(n9924));
AND2X1 mul_U415(.A(n682), .B(n12364), .Y(dpath_mulcore_ary1_a1_I2_I1_26__net32));
OR2X1 mul_U416(.A(n6758), .B(dpath_mulcore_b14[0]), .Y(n12364));
AND2X1 mul_U417(.A(n681), .B(n12361), .Y(dpath_mulcore_ary1_a1_I2_I1_26__net046));
OR2X1 mul_U418(.A(n6757), .B(dpath_mulcore_b15[0]), .Y(n12361));
INVX1 mul_U419(.A(dpath_mulcore_op1_l[22]), .Y(n9921));
AND2X1 mul_U420(.A(n684), .B(n12370), .Y(dpath_mulcore_ary1_a1_I2_I1_25__net32));
OR2X1 mul_U421(.A(n6760), .B(dpath_mulcore_b14[0]), .Y(n12370));
AND2X1 mul_U422(.A(n683), .B(n12367), .Y(dpath_mulcore_ary1_a1_I2_I1_25__net046));
OR2X1 mul_U423(.A(n6759), .B(dpath_mulcore_b15[0]), .Y(n12367));
INVX1 mul_U424(.A(dpath_mulcore_op1_l[21]), .Y(n9918));
AND2X1 mul_U425(.A(n686), .B(n12376), .Y(dpath_mulcore_ary1_a1_I2_I1_24__net32));
OR2X1 mul_U426(.A(n6762), .B(dpath_mulcore_b14[0]), .Y(n12376));
AND2X1 mul_U427(.A(n685), .B(n12373), .Y(dpath_mulcore_ary1_a1_I2_I1_24__net046));
OR2X1 mul_U428(.A(n6761), .B(dpath_mulcore_b15[0]), .Y(n12373));
INVX1 mul_U429(.A(dpath_mulcore_op1_l[20]), .Y(n9915));
AND2X1 mul_U430(.A(n688), .B(n12382), .Y(dpath_mulcore_ary1_a1_I2_I1_23__net32));
OR2X1 mul_U431(.A(n6764), .B(dpath_mulcore_b14[0]), .Y(n12382));
AND2X1 mul_U432(.A(n687), .B(n12379), .Y(dpath_mulcore_ary1_a1_I2_I1_23__net046));
OR2X1 mul_U433(.A(n6763), .B(dpath_mulcore_b15[0]), .Y(n12379));
INVX1 mul_U434(.A(dpath_mulcore_op1_l[19]), .Y(n9912));
AND2X1 mul_U435(.A(n690), .B(n12388), .Y(dpath_mulcore_ary1_a1_I2_I1_22__net32));
OR2X1 mul_U436(.A(n6766), .B(dpath_mulcore_b14[0]), .Y(n12388));
AND2X1 mul_U437(.A(n689), .B(n12385), .Y(dpath_mulcore_ary1_a1_I2_I1_22__net046));
OR2X1 mul_U438(.A(n6765), .B(dpath_mulcore_b15[0]), .Y(n12385));
INVX1 mul_U439(.A(dpath_mulcore_op1_l[18]), .Y(n9909));
AND2X1 mul_U440(.A(n692), .B(n12394), .Y(dpath_mulcore_ary1_a1_I2_I1_21__net32));
OR2X1 mul_U441(.A(n6768), .B(dpath_mulcore_b14[0]), .Y(n12394));
AND2X1 mul_U442(.A(n691), .B(n12391), .Y(dpath_mulcore_ary1_a1_I2_I1_21__net046));
OR2X1 mul_U443(.A(n6767), .B(dpath_mulcore_b15[0]), .Y(n12391));
INVX1 mul_U444(.A(dpath_mulcore_op1_l[17]), .Y(n9906));
AND2X1 mul_U445(.A(n694), .B(n12400), .Y(dpath_mulcore_ary1_a1_I2_I1_20__net32));
OR2X1 mul_U446(.A(n6770), .B(dpath_mulcore_b14[0]), .Y(n12400));
AND2X1 mul_U447(.A(n693), .B(n12397), .Y(dpath_mulcore_ary1_a1_I2_I1_20__net046));
OR2X1 mul_U448(.A(n6769), .B(dpath_mulcore_b15[0]), .Y(n12397));
INVX1 mul_U449(.A(dpath_mulcore_op1_l[16]), .Y(n9903));
AND2X1 mul_U450(.A(n696), .B(n12406), .Y(dpath_mulcore_ary1_a1_I2_I1_19__net32));
OR2X1 mul_U451(.A(n6772), .B(dpath_mulcore_b14[0]), .Y(n12406));
AND2X1 mul_U452(.A(n695), .B(n12403), .Y(dpath_mulcore_ary1_a1_I2_I1_19__net046));
OR2X1 mul_U453(.A(n6771), .B(dpath_mulcore_b15[0]), .Y(n12403));
INVX1 mul_U454(.A(dpath_mulcore_op1_l[15]), .Y(n9900));
AND2X1 mul_U455(.A(n698), .B(n12412), .Y(dpath_mulcore_ary1_a1_I2_I1_18__net32));
OR2X1 mul_U456(.A(n6774), .B(dpath_mulcore_b14[0]), .Y(n12412));
AND2X1 mul_U457(.A(n697), .B(n12409), .Y(dpath_mulcore_ary1_a1_I2_I1_18__net046));
OR2X1 mul_U458(.A(n6773), .B(dpath_mulcore_b15[0]), .Y(n12409));
INVX1 mul_U459(.A(dpath_mulcore_op1_l[14]), .Y(n9897));
AND2X1 mul_U460(.A(n700), .B(n12418), .Y(dpath_mulcore_ary1_a1_I2_I1_17__net32));
OR2X1 mul_U461(.A(n6776), .B(dpath_mulcore_b14[0]), .Y(n12418));
AND2X1 mul_U462(.A(n699), .B(n12415), .Y(dpath_mulcore_ary1_a1_I2_I1_17__net046));
OR2X1 mul_U463(.A(n6775), .B(dpath_mulcore_b15[0]), .Y(n12415));
INVX1 mul_U464(.A(dpath_mulcore_op1_l[13]), .Y(n9894));
AND2X1 mul_U465(.A(n702), .B(n12424), .Y(dpath_mulcore_ary1_a1_I2_I1_16__net32));
OR2X1 mul_U466(.A(n6778), .B(dpath_mulcore_b14[0]), .Y(n12424));
AND2X1 mul_U467(.A(n701), .B(n12421), .Y(dpath_mulcore_ary1_a1_I2_I1_16__net046));
OR2X1 mul_U468(.A(n6777), .B(dpath_mulcore_b15[0]), .Y(n12421));
INVX1 mul_U469(.A(dpath_mulcore_op1_l[12]), .Y(n9891));
AND2X1 mul_U470(.A(n704), .B(n12430), .Y(dpath_mulcore_ary1_a1_I2_I1_15__net32));
OR2X1 mul_U471(.A(n6780), .B(dpath_mulcore_b14[0]), .Y(n12430));
AND2X1 mul_U472(.A(n703), .B(n12427), .Y(dpath_mulcore_ary1_a1_I2_I1_15__net046));
OR2X1 mul_U473(.A(n6779), .B(dpath_mulcore_b15[0]), .Y(n12427));
INVX1 mul_U474(.A(dpath_mulcore_op1_l[11]), .Y(n9888));
AND2X1 mul_U475(.A(n706), .B(n12436), .Y(dpath_mulcore_ary1_a1_I2_I1_14__net32));
OR2X1 mul_U476(.A(n6782), .B(dpath_mulcore_b14[0]), .Y(n12436));
AND2X1 mul_U477(.A(n705), .B(n12433), .Y(dpath_mulcore_ary1_a1_I2_I1_14__net046));
OR2X1 mul_U478(.A(n6781), .B(dpath_mulcore_b15[0]), .Y(n12433));
INVX1 mul_U479(.A(dpath_mulcore_op1_l[10]), .Y(n9885));
AND2X1 mul_U480(.A(n708), .B(n12442), .Y(dpath_mulcore_ary1_a1_I2_I1_13__net32));
OR2X1 mul_U481(.A(n6784), .B(dpath_mulcore_b14[0]), .Y(n12442));
AND2X1 mul_U482(.A(n707), .B(n12439), .Y(dpath_mulcore_ary1_a1_I2_I1_13__net046));
OR2X1 mul_U483(.A(n6783), .B(dpath_mulcore_b15[0]), .Y(n12439));
INVX1 mul_U484(.A(dpath_mulcore_op1_l[9]), .Y(n9882));
AND2X1 mul_U485(.A(n710), .B(n12448), .Y(dpath_mulcore_ary1_a1_I2_I1_12__net32));
OR2X1 mul_U486(.A(n6786), .B(dpath_mulcore_b14[0]), .Y(n12448));
AND2X1 mul_U487(.A(n709), .B(n12445), .Y(dpath_mulcore_ary1_a1_I2_I1_12__net046));
OR2X1 mul_U488(.A(n6785), .B(dpath_mulcore_b15[0]), .Y(n12445));
INVX1 mul_U489(.A(dpath_mulcore_op1_l[8]), .Y(n9879));
AND2X1 mul_U490(.A(n712), .B(n12454), .Y(dpath_mulcore_ary1_a1_I2_I1_11__net32));
OR2X1 mul_U491(.A(n6788), .B(dpath_mulcore_b14[0]), .Y(n12454));
AND2X1 mul_U492(.A(n711), .B(n12451), .Y(dpath_mulcore_ary1_a1_I2_I1_11__net046));
OR2X1 mul_U493(.A(n6787), .B(dpath_mulcore_b15[0]), .Y(n12451));
INVX1 mul_U494(.A(dpath_mulcore_op1_l[7]), .Y(n9876));
AND2X1 mul_U495(.A(n714), .B(n12460), .Y(dpath_mulcore_ary1_a1_I2_I1_10__net32));
OR2X1 mul_U496(.A(n6790), .B(dpath_mulcore_b14[0]), .Y(n12460));
AND2X1 mul_U497(.A(n713), .B(n12457), .Y(dpath_mulcore_ary1_a1_I2_I1_10__net046));
OR2X1 mul_U498(.A(n6789), .B(dpath_mulcore_b15[0]), .Y(n12457));
INVX1 mul_U499(.A(dpath_mulcore_op1_l[6]), .Y(n9873));
AND2X1 mul_U500(.A(n716), .B(n12466), .Y(dpath_mulcore_ary1_a1_I2_I1_9__net32));
OR2X1 mul_U501(.A(n6792), .B(dpath_mulcore_b14[0]), .Y(n12466));
AND2X1 mul_U502(.A(n715), .B(n12463), .Y(dpath_mulcore_ary1_a1_I2_I1_9__net046));
OR2X1 mul_U503(.A(n6791), .B(dpath_mulcore_b15[0]), .Y(n12463));
INVX1 mul_U504(.A(dpath_mulcore_op1_l[5]), .Y(n9870));
AND2X1 mul_U505(.A(n718), .B(n12472), .Y(dpath_mulcore_ary1_a1_I2_I1_8__net32));
OR2X1 mul_U506(.A(n6794), .B(dpath_mulcore_b14[0]), .Y(n12472));
AND2X1 mul_U507(.A(n717), .B(n12469), .Y(dpath_mulcore_ary1_a1_I2_I1_8__net046));
OR2X1 mul_U508(.A(n6793), .B(dpath_mulcore_b15[0]), .Y(n12469));
INVX1 mul_U509(.A(dpath_mulcore_op1_l[4]), .Y(n9867));
AND2X1 mul_U510(.A(n720), .B(n12478), .Y(dpath_mulcore_ary1_a1_I2_I1_7__net32));
OR2X1 mul_U511(.A(n6796), .B(dpath_mulcore_b14[0]), .Y(n12478));
AND2X1 mul_U512(.A(n719), .B(n12475), .Y(dpath_mulcore_ary1_a1_I2_I1_7__net046));
OR2X1 mul_U513(.A(n6795), .B(dpath_mulcore_b15[0]), .Y(n12475));
INVX1 mul_U514(.A(dpath_mulcore_op1_l[3]), .Y(n9864));
AND2X1 mul_U515(.A(n722), .B(n12484), .Y(dpath_mulcore_ary1_a1_I2_I1_6__net32));
OR2X1 mul_U516(.A(n6798), .B(dpath_mulcore_b14[0]), .Y(n12484));
AND2X1 mul_U517(.A(n721), .B(n12481), .Y(dpath_mulcore_ary1_a1_I2_I1_6__net046));
OR2X1 mul_U518(.A(n6797), .B(dpath_mulcore_b15[0]), .Y(n12481));
AND2X1 mul_U519(.A(n724), .B(n12490), .Y(dpath_mulcore_ary1_a1_I2_I1_5__net32));
OR2X1 mul_U520(.A(n6800), .B(dpath_mulcore_b14[0]), .Y(n12490));
AND2X1 mul_U521(.A(n723), .B(n12487), .Y(dpath_mulcore_ary1_a1_I2_I1_5__net046));
OR2X1 mul_U522(.A(n6799), .B(dpath_mulcore_b15[0]), .Y(n12487));
AND2X1 mul_U523(.A(n726), .B(n12496), .Y(dpath_mulcore_ary1_a1_I2_I1_4__net32));
OR2X1 mul_U524(.A(n6802), .B(dpath_mulcore_b14[0]), .Y(n12496));
AND2X1 mul_U525(.A(n725), .B(n12493), .Y(dpath_mulcore_ary1_a1_I2_I1_4__net046));
OR2X1 mul_U526(.A(n6801), .B(dpath_mulcore_b15[0]), .Y(n12493));
AND2X1 mul_U527(.A(n728), .B(n12502), .Y(dpath_mulcore_ary1_a1_I2_I0_p1_3));
OR2X1 mul_U528(.A(n6804), .B(dpath_mulcore_b15[0]), .Y(n12502));
AND2X1 mul_U529(.A(n727), .B(n12499), .Y(dpath_mulcore_ary1_a1_I2_I0_p0_3));
OR2X1 mul_U530(.A(n6803), .B(dpath_mulcore_b14[0]), .Y(n12499));
INVX1 mul_U531(.A(n12512), .Y(n9838));
OR2X1 mul_U532(.A(n6808), .B(dpath_mulcore_b15[0]), .Y(n12512));
AND2X1 mul_U533(.A(n729), .B(n12505), .Y(dpath_mulcore_ary1_a1_I2_I0_p0_2));
OR2X1 mul_U534(.A(n6805), .B(dpath_mulcore_b14[0]), .Y(n12505));
AND2X1 mul_U535(.A(n1093), .B(n13607), .Y(dpath_mulcore_ary1_a1_I0_I1_8__net32));
OR2X1 mul_U536(.A(n7174), .B(dpath_mulcore_b8[0]), .Y(n13607));
AND2X1 mul_U537(.A(n1092), .B(n13604), .Y(dpath_mulcore_ary1_a1_I0_I1_8__net046));
OR2X1 mul_U538(.A(n7173), .B(dpath_mulcore_b9[0]), .Y(n13604));
AND2X1 mul_U539(.A(n2960), .B(n4636), .Y(dpath_n838));
AND2X1 mul_U540(.A(n1998), .B(n4051), .Y(dpath_mulcore_array2_c1[66]));
AND2X1 mul_U541(.A(n2958), .B(n4634), .Y(dpath_n832));
AND2X1 mul_U542(.A(n1990), .B(n4043), .Y(dpath_mulcore_array2_c2[28]));
AND2X1 mul_U543(.A(n2036), .B(n4089), .Y(dpath_mulcore_array2_c1[28]));
OR2X1 mul_U544(.A(n9467), .B(dpath_mulcore_array2_s1[28]), .Y(n17743));
AND2X1 mul_U545(.A(n1991), .B(n4044), .Y(dpath_mulcore_array2_c2[27]));
AND2X1 mul_U546(.A(n2037), .B(n4090), .Y(dpath_mulcore_array2_c1[27]));
OR2X1 mul_U547(.A(n9468), .B(dpath_mulcore_array2_s1[27]), .Y(n17750));
OR2X1 mul_U548(.A(n5906), .B(n6034), .Y(dpath_areg[29]));
AND2X1 mul_U549(.A(n2965), .B(n4641), .Y(dpath_n849));
AND2X1 mul_U550(.A(n1992), .B(n4045), .Y(dpath_mulcore_array2_c2[26]));
AND2X1 mul_U551(.A(n2038), .B(n4091), .Y(dpath_mulcore_array2_c1[26]));
OR2X1 mul_U552(.A(n9469), .B(dpath_mulcore_array2_s1[26]), .Y(n17757));
OR2X1 mul_U553(.A(n5907), .B(n6035), .Y(dpath_areg[28]));
AND2X1 mul_U554(.A(n2967), .B(n4643), .Y(dpath_n855));
AND2X1 mul_U555(.A(n1993), .B(n4046), .Y(dpath_mulcore_array2_c2[25]));
AND2X1 mul_U556(.A(n2039), .B(n4092), .Y(dpath_mulcore_array2_c1[25]));
OR2X1 mul_U557(.A(n9470), .B(dpath_mulcore_array2_s1[25]), .Y(n17764));
OR2X1 mul_U558(.A(n5908), .B(n6036), .Y(dpath_areg[27]));
AND2X1 mul_U559(.A(n2969), .B(n4645), .Y(dpath_n861));
AND2X1 mul_U560(.A(n1994), .B(n4047), .Y(dpath_mulcore_array2_c2[24]));
AND2X1 mul_U561(.A(n2040), .B(n4093), .Y(dpath_mulcore_array2_c1[24]));
OR2X1 mul_U562(.A(n9471), .B(dpath_mulcore_array2_s1[24]), .Y(n17771));
OR2X1 mul_U563(.A(n5909), .B(n6037), .Y(dpath_areg[26]));
AND2X1 mul_U564(.A(n2971), .B(n4647), .Y(dpath_n867));
AND2X1 mul_U565(.A(n1995), .B(n4048), .Y(dpath_mulcore_array2_c2[23]));
AND2X1 mul_U566(.A(n2041), .B(n4094), .Y(dpath_mulcore_array2_c1[23]));
OR2X1 mul_U567(.A(n9472), .B(dpath_mulcore_array2_s1[23]), .Y(n17778));
OR2X1 mul_U568(.A(n5910), .B(n6038), .Y(dpath_areg[25]));
AND2X1 mul_U569(.A(n2973), .B(n4649), .Y(dpath_n873));
AND2X1 mul_U570(.A(n1996), .B(n4049), .Y(dpath_mulcore_array2_c2[22]));
AND2X1 mul_U571(.A(n2042), .B(n4095), .Y(dpath_mulcore_array2_c1[22]));
OR2X1 mul_U572(.A(n9473), .B(dpath_mulcore_array2_s1[22]), .Y(n17785));
OR2X1 mul_U573(.A(n5911), .B(n6039), .Y(dpath_areg[24]));
AND2X1 mul_U574(.A(n2975), .B(n4651), .Y(dpath_n879));
AND2X1 mul_U575(.A(n1997), .B(n4050), .Y(dpath_mulcore_array2_c2[21]));
AND2X1 mul_U576(.A(n2043), .B(n4096), .Y(dpath_mulcore_array2_c1[21]));
OR2X1 mul_U577(.A(n16368), .B(dpath_mulcore_array2_s1[21]), .Y(n17792));
OR2X1 mul_U578(.A(n5912), .B(n6040), .Y(dpath_areg[23]));
AND2X1 mul_U579(.A(n2977), .B(n4653), .Y(dpath_n885));
AND2X1 mul_U580(.A(n2044), .B(n4097), .Y(dpath_mulcore_array2_c1[20]));
OR2X1 mul_U581(.A(n9428), .B(dpath_mulcore_array2_s1[20]), .Y(n17799));
OR2X1 mul_U582(.A(n5913), .B(n6041), .Y(dpath_areg[22]));
AND2X1 mul_U583(.A(n2979), .B(n4655), .Y(dpath_n891));
OR2X1 mul_U584(.A(n5914), .B(n6042), .Y(dpath_areg[21]));
AND2X1 mul_U585(.A(n2981), .B(n4657), .Y(dpath_n897));
OR2X1 mul_U586(.A(n5915), .B(n6043), .Y(dpath_areg[20]));
AND2X1 mul_U587(.A(n2983), .B(n4659), .Y(dpath_n903));
OR2X1 mul_U588(.A(n5917), .B(n6045), .Y(dpath_areg[19]));
AND2X1 mul_U589(.A(n2987), .B(n4663), .Y(dpath_n915));
OR2X1 mul_U590(.A(n5918), .B(n6046), .Y(dpath_areg[18]));
AND2X1 mul_U591(.A(n2989), .B(n4665), .Y(dpath_n921));
OR2X1 mul_U592(.A(n5919), .B(n6047), .Y(dpath_areg[17]));
AND2X1 mul_U593(.A(n2991), .B(n4667), .Y(dpath_n927));
AND2X1 mul_U594(.A(n2994), .B(n4670), .Y(dpath_n940));
AND2X1 mul_U595(.A(n2992), .B(n4668), .Y(dpath_n934));
AND2X1 mul_U596(.A(n1928), .B(n3981), .Y(dpath_mulcore_array2_c1[13]));
OR2X1 mul_U597(.A(n5922), .B(n6050), .Y(dpath_areg[14]));
AND2X1 mul_U598(.A(n2997), .B(n4673), .Y(dpath_n945));
OR2X1 mul_U599(.A(n5923), .B(n6051), .Y(dpath_areg[13]));
AND2X1 mul_U600(.A(n2999), .B(n4675), .Y(dpath_n951));
OR2X1 mul_U601(.A(n5924), .B(n6052), .Y(dpath_areg[12]));
AND2X1 mul_U602(.A(n3001), .B(n4677), .Y(dpath_n957));
OR2X1 mul_U603(.A(n5925), .B(n6053), .Y(dpath_areg[11]));
AND2X1 mul_U604(.A(n3003), .B(n4679), .Y(dpath_n963));
OR2X1 mul_U605(.A(n5926), .B(n6054), .Y(dpath_areg[10]));
AND2X1 mul_U606(.A(n3005), .B(n4681), .Y(dpath_n969));
OR2X1 mul_U607(.A(n5896), .B(n6024), .Y(dpath_areg[9]));
AND2X1 mul_U608(.A(n2880), .B(n4556), .Y(dpath_n653));
OR2X1 mul_U609(.A(n5897), .B(n6025), .Y(dpath_areg[8]));
AND2X1 mul_U610(.A(n2889), .B(n4565), .Y(dpath_n679));
OR2X1 mul_U611(.A(n5898), .B(n6026), .Y(dpath_areg[7]));
AND2X1 mul_U612(.A(n2901), .B(n4577), .Y(dpath_n705));
OR2X1 mul_U613(.A(n5899), .B(n6027), .Y(dpath_areg[6]));
AND2X1 mul_U614(.A(n2913), .B(n4589), .Y(dpath_n731));
OR2X1 mul_U615(.A(n5900), .B(n6028), .Y(dpath_areg[5]));
AND2X1 mul_U616(.A(n2925), .B(n4601), .Y(dpath_n757));
OR2X1 mul_U617(.A(n5901), .B(n6029), .Y(dpath_areg[4]));
AND2X1 mul_U618(.A(n2937), .B(n4613), .Y(dpath_n783));
OR2X1 mul_U619(.A(n5902), .B(n6030), .Y(dpath_areg[3]));
AND2X1 mul_U620(.A(n2949), .B(n4625), .Y(dpath_n809));
OR2X1 mul_U621(.A(n5905), .B(n6033), .Y(dpath_areg[2]));
AND2X1 mul_U622(.A(n2963), .B(n4639), .Y(dpath_n843));
AND2X1 mul_U623(.A(n2984), .B(n4660), .Y(dpath_n910));
AND2X1 mul_U624(.A(n1115), .B(n13673), .Y(dpath_mulcore_ary1_a0_I0_I2_net38));
OR2X1 mul_U625(.A(n9426), .B(dpath_mulcore_b1[0]), .Y(n13673));
AND2X1 mul_U626(.A(n419), .B(n11569), .Y(dpath_mulcore_ary1_a0_I0_I2_net43));
OR2X1 mul_U627(.A(n6492), .B(dpath_mulcore_b1[0]), .Y(n11569));
AND2X1 mul_U628(.A(n1113), .B(n13669), .Y(dpath_mulcore_ary1_a0_I0_I2_net47));
OR2X1 mul_U629(.A(n9217), .B(dpath_mulcore_b0[0]), .Y(n13669));
AND2X1 mul_U630(.A(n420), .B(n11572), .Y(dpath_mulcore_ary1_a0_I0_I2_net48));
OR2X1 mul_U631(.A(n6493), .B(dpath_mulcore_b1[0]), .Y(n11572));
AND2X1 mul_U632(.A(n424), .B(n11584), .Y(dpath_mulcore_ary1_a0_I0_I1_63__net32));
OR2X1 mul_U633(.A(n6497), .B(dpath_mulcore_b0[0]), .Y(n11584));
AND2X1 mul_U634(.A(n423), .B(n11581), .Y(dpath_mulcore_ary1_a0_I0_I1_63__net046));
OR2X1 mul_U635(.A(n6496), .B(dpath_mulcore_b1[0]), .Y(n11581));
AND2X1 mul_U636(.A(n427), .B(n11593), .Y(dpath_mulcore_ary1_a0_I0_I1_62__net32));
OR2X1 mul_U637(.A(n6500), .B(dpath_mulcore_b0[0]), .Y(n11593));
AND2X1 mul_U638(.A(n426), .B(n11590), .Y(dpath_mulcore_ary1_a0_I0_I1_62__net046));
OR2X1 mul_U639(.A(n6499), .B(dpath_mulcore_b1[0]), .Y(n11590));
AND2X1 mul_U640(.A(n430), .B(n11602), .Y(dpath_mulcore_ary1_a0_I0_I1_61__net32));
OR2X1 mul_U641(.A(n6503), .B(dpath_mulcore_b0[0]), .Y(n11602));
AND2X1 mul_U642(.A(n429), .B(n11599), .Y(dpath_mulcore_ary1_a0_I0_I1_61__net046));
OR2X1 mul_U643(.A(n6502), .B(dpath_mulcore_b1[0]), .Y(n11599));
AND2X1 mul_U644(.A(n433), .B(n11611), .Y(dpath_mulcore_ary1_a0_I0_I1_60__net32));
OR2X1 mul_U645(.A(n6506), .B(dpath_mulcore_b0[0]), .Y(n11611));
AND2X1 mul_U646(.A(n432), .B(n11608), .Y(dpath_mulcore_ary1_a0_I0_I1_60__net046));
OR2X1 mul_U647(.A(n6505), .B(dpath_mulcore_b1[0]), .Y(n11608));
AND2X1 mul_U648(.A(n436), .B(n11620), .Y(dpath_mulcore_ary1_a0_I0_I1_59__net32));
OR2X1 mul_U649(.A(n6509), .B(dpath_mulcore_b0[0]), .Y(n11620));
AND2X1 mul_U650(.A(n435), .B(n11617), .Y(dpath_mulcore_ary1_a0_I0_I1_59__net046));
OR2X1 mul_U651(.A(n6508), .B(dpath_mulcore_b1[0]), .Y(n11617));
AND2X1 mul_U652(.A(n439), .B(n11629), .Y(dpath_mulcore_ary1_a0_I0_I1_58__net32));
OR2X1 mul_U653(.A(n6512), .B(dpath_mulcore_b0[0]), .Y(n11629));
AND2X1 mul_U654(.A(n438), .B(n11626), .Y(dpath_mulcore_ary1_a0_I0_I1_58__net046));
OR2X1 mul_U655(.A(n6511), .B(dpath_mulcore_b1[0]), .Y(n11626));
AND2X1 mul_U656(.A(n442), .B(n11638), .Y(dpath_mulcore_ary1_a0_I0_I1_57__net32));
OR2X1 mul_U657(.A(n6515), .B(dpath_mulcore_b0[0]), .Y(n11638));
AND2X1 mul_U658(.A(n441), .B(n11635), .Y(dpath_mulcore_ary1_a0_I0_I1_57__net046));
OR2X1 mul_U659(.A(n6514), .B(dpath_mulcore_b1[0]), .Y(n11635));
AND2X1 mul_U660(.A(n445), .B(n11647), .Y(dpath_mulcore_ary1_a0_I0_I1_56__net32));
OR2X1 mul_U661(.A(n6518), .B(dpath_mulcore_b0[0]), .Y(n11647));
AND2X1 mul_U662(.A(n444), .B(n11644), .Y(dpath_mulcore_ary1_a0_I0_I1_56__net046));
OR2X1 mul_U663(.A(n6517), .B(dpath_mulcore_b1[0]), .Y(n11644));
AND2X1 mul_U664(.A(n448), .B(n11656), .Y(dpath_mulcore_ary1_a0_I0_I1_55__net32));
OR2X1 mul_U665(.A(n6521), .B(dpath_mulcore_b0[0]), .Y(n11656));
AND2X1 mul_U666(.A(n447), .B(n11653), .Y(dpath_mulcore_ary1_a0_I0_I1_55__net046));
OR2X1 mul_U667(.A(n6520), .B(dpath_mulcore_b1[0]), .Y(n11653));
AND2X1 mul_U668(.A(n451), .B(n11665), .Y(dpath_mulcore_ary1_a0_I0_I1_54__net32));
OR2X1 mul_U669(.A(n6524), .B(dpath_mulcore_b0[0]), .Y(n11665));
AND2X1 mul_U670(.A(n450), .B(n11662), .Y(dpath_mulcore_ary1_a0_I0_I1_54__net046));
OR2X1 mul_U671(.A(n6523), .B(dpath_mulcore_b1[0]), .Y(n11662));
AND2X1 mul_U672(.A(n454), .B(n11674), .Y(dpath_mulcore_ary1_a0_I0_I1_53__net32));
OR2X1 mul_U673(.A(n6527), .B(dpath_mulcore_b0[0]), .Y(n11674));
AND2X1 mul_U674(.A(n453), .B(n11671), .Y(dpath_mulcore_ary1_a0_I0_I1_53__net046));
OR2X1 mul_U675(.A(n6526), .B(dpath_mulcore_b1[0]), .Y(n11671));
AND2X1 mul_U676(.A(n457), .B(n11683), .Y(dpath_mulcore_ary1_a0_I0_I1_52__net32));
OR2X1 mul_U677(.A(n6530), .B(dpath_mulcore_b0[0]), .Y(n11683));
AND2X1 mul_U678(.A(n456), .B(n11680), .Y(dpath_mulcore_ary1_a0_I0_I1_52__net046));
OR2X1 mul_U679(.A(n6529), .B(dpath_mulcore_b1[0]), .Y(n11680));
AND2X1 mul_U680(.A(n460), .B(n11692), .Y(dpath_mulcore_ary1_a0_I0_I1_51__net32));
OR2X1 mul_U681(.A(n6533), .B(dpath_mulcore_b0[0]), .Y(n11692));
AND2X1 mul_U682(.A(n459), .B(n11689), .Y(dpath_mulcore_ary1_a0_I0_I1_51__net046));
OR2X1 mul_U683(.A(n6532), .B(dpath_mulcore_b1[0]), .Y(n11689));
AND2X1 mul_U684(.A(n463), .B(n11701), .Y(dpath_mulcore_ary1_a0_I0_I1_50__net32));
OR2X1 mul_U685(.A(n6536), .B(dpath_mulcore_b0[0]), .Y(n11701));
AND2X1 mul_U686(.A(n462), .B(n11698), .Y(dpath_mulcore_ary1_a0_I0_I1_50__net046));
OR2X1 mul_U687(.A(n6535), .B(dpath_mulcore_b1[0]), .Y(n11698));
AND2X1 mul_U688(.A(n466), .B(n11710), .Y(dpath_mulcore_ary1_a0_I0_I1_49__net32));
OR2X1 mul_U689(.A(n6539), .B(dpath_mulcore_b0[0]), .Y(n11710));
AND2X1 mul_U690(.A(n465), .B(n11707), .Y(dpath_mulcore_ary1_a0_I0_I1_49__net046));
OR2X1 mul_U691(.A(n6538), .B(dpath_mulcore_b1[0]), .Y(n11707));
AND2X1 mul_U692(.A(n469), .B(n11719), .Y(dpath_mulcore_ary1_a0_I0_I1_48__net32));
OR2X1 mul_U693(.A(n6542), .B(dpath_mulcore_b0[0]), .Y(n11719));
AND2X1 mul_U694(.A(n468), .B(n11716), .Y(dpath_mulcore_ary1_a0_I0_I1_48__net046));
OR2X1 mul_U695(.A(n6541), .B(dpath_mulcore_b1[0]), .Y(n11716));
AND2X1 mul_U696(.A(n472), .B(n11728), .Y(dpath_mulcore_ary1_a0_I0_I1_47__net32));
OR2X1 mul_U697(.A(n6545), .B(dpath_mulcore_b0[0]), .Y(n11728));
AND2X1 mul_U698(.A(n471), .B(n11725), .Y(dpath_mulcore_ary1_a0_I0_I1_47__net046));
OR2X1 mul_U699(.A(n6544), .B(dpath_mulcore_b1[0]), .Y(n11725));
AND2X1 mul_U700(.A(n475), .B(n11737), .Y(dpath_mulcore_ary1_a0_I0_I1_46__net32));
OR2X1 mul_U701(.A(n6548), .B(dpath_mulcore_b0[0]), .Y(n11737));
AND2X1 mul_U702(.A(n474), .B(n11734), .Y(dpath_mulcore_ary1_a0_I0_I1_46__net046));
OR2X1 mul_U703(.A(n6547), .B(dpath_mulcore_b1[0]), .Y(n11734));
AND2X1 mul_U704(.A(n478), .B(n11746), .Y(dpath_mulcore_ary1_a0_I0_I1_45__net32));
OR2X1 mul_U705(.A(n6551), .B(dpath_mulcore_b0[0]), .Y(n11746));
AND2X1 mul_U706(.A(n477), .B(n11743), .Y(dpath_mulcore_ary1_a0_I0_I1_45__net046));
OR2X1 mul_U707(.A(n6550), .B(dpath_mulcore_b1[0]), .Y(n11743));
AND2X1 mul_U708(.A(n481), .B(n11755), .Y(dpath_mulcore_ary1_a0_I0_I1_44__net32));
OR2X1 mul_U709(.A(n6554), .B(dpath_mulcore_b0[0]), .Y(n11755));
AND2X1 mul_U710(.A(n480), .B(n11752), .Y(dpath_mulcore_ary1_a0_I0_I1_44__net046));
OR2X1 mul_U711(.A(n6553), .B(dpath_mulcore_b1[0]), .Y(n11752));
AND2X1 mul_U712(.A(n484), .B(n11764), .Y(dpath_mulcore_ary1_a0_I0_I1_43__net32));
OR2X1 mul_U713(.A(n6557), .B(dpath_mulcore_b0[0]), .Y(n11764));
AND2X1 mul_U714(.A(n483), .B(n11761), .Y(dpath_mulcore_ary1_a0_I0_I1_43__net046));
OR2X1 mul_U715(.A(n6556), .B(dpath_mulcore_b1[0]), .Y(n11761));
AND2X1 mul_U716(.A(n487), .B(n11773), .Y(dpath_mulcore_ary1_a0_I0_I1_42__net32));
OR2X1 mul_U717(.A(n6560), .B(dpath_mulcore_b0[0]), .Y(n11773));
AND2X1 mul_U718(.A(n486), .B(n11770), .Y(dpath_mulcore_ary1_a0_I0_I1_42__net046));
OR2X1 mul_U719(.A(n6559), .B(dpath_mulcore_b1[0]), .Y(n11770));
AND2X1 mul_U720(.A(n490), .B(n11782), .Y(dpath_mulcore_ary1_a0_I0_I1_41__net32));
OR2X1 mul_U721(.A(n6563), .B(dpath_mulcore_b0[0]), .Y(n11782));
AND2X1 mul_U722(.A(n489), .B(n11779), .Y(dpath_mulcore_ary1_a0_I0_I1_41__net046));
OR2X1 mul_U723(.A(n6562), .B(dpath_mulcore_b1[0]), .Y(n11779));
AND2X1 mul_U724(.A(n493), .B(n11791), .Y(dpath_mulcore_ary1_a0_I0_I1_40__net32));
OR2X1 mul_U725(.A(n6566), .B(dpath_mulcore_b0[0]), .Y(n11791));
AND2X1 mul_U726(.A(n492), .B(n11788), .Y(dpath_mulcore_ary1_a0_I0_I1_40__net046));
OR2X1 mul_U727(.A(n6565), .B(dpath_mulcore_b1[0]), .Y(n11788));
AND2X1 mul_U728(.A(n496), .B(n11800), .Y(dpath_mulcore_ary1_a0_I0_I1_39__net32));
OR2X1 mul_U729(.A(n6569), .B(dpath_mulcore_b0[0]), .Y(n11800));
AND2X1 mul_U730(.A(n495), .B(n11797), .Y(dpath_mulcore_ary1_a0_I0_I1_39__net046));
OR2X1 mul_U731(.A(n6568), .B(dpath_mulcore_b1[0]), .Y(n11797));
AND2X1 mul_U732(.A(n499), .B(n11809), .Y(dpath_mulcore_ary1_a0_I0_I1_38__net32));
OR2X1 mul_U733(.A(n6572), .B(dpath_mulcore_b0[0]), .Y(n11809));
AND2X1 mul_U734(.A(n498), .B(n11806), .Y(dpath_mulcore_ary1_a0_I0_I1_38__net046));
OR2X1 mul_U735(.A(n6571), .B(dpath_mulcore_b1[0]), .Y(n11806));
AND2X1 mul_U736(.A(n502), .B(n11818), .Y(dpath_mulcore_ary1_a0_I0_I1_37__net32));
OR2X1 mul_U737(.A(n6575), .B(dpath_mulcore_b0[0]), .Y(n11818));
AND2X1 mul_U738(.A(n501), .B(n11815), .Y(dpath_mulcore_ary1_a0_I0_I1_37__net046));
OR2X1 mul_U739(.A(n6574), .B(dpath_mulcore_b1[0]), .Y(n11815));
AND2X1 mul_U740(.A(n505), .B(n11827), .Y(dpath_mulcore_ary1_a0_I0_I1_36__net32));
OR2X1 mul_U741(.A(n6578), .B(dpath_mulcore_b0[0]), .Y(n11827));
AND2X1 mul_U742(.A(n504), .B(n11824), .Y(dpath_mulcore_ary1_a0_I0_I1_36__net046));
OR2X1 mul_U743(.A(n6577), .B(dpath_mulcore_b1[0]), .Y(n11824));
AND2X1 mul_U744(.A(n508), .B(n11836), .Y(dpath_mulcore_ary1_a0_I0_I1_35__net32));
OR2X1 mul_U745(.A(n6581), .B(dpath_mulcore_b0[0]), .Y(n11836));
AND2X1 mul_U746(.A(n507), .B(n11833), .Y(dpath_mulcore_ary1_a0_I0_I1_35__net046));
OR2X1 mul_U747(.A(n6580), .B(dpath_mulcore_b1[0]), .Y(n11833));
AND2X1 mul_U748(.A(n511), .B(n11845), .Y(dpath_mulcore_ary1_a0_I0_I1_34__net32));
OR2X1 mul_U749(.A(n6584), .B(dpath_mulcore_b0[0]), .Y(n11845));
AND2X1 mul_U750(.A(n510), .B(n11842), .Y(dpath_mulcore_ary1_a0_I0_I1_34__net046));
OR2X1 mul_U751(.A(n6583), .B(dpath_mulcore_b1[0]), .Y(n11842));
AND2X1 mul_U752(.A(n514), .B(n11854), .Y(dpath_mulcore_ary1_a0_I0_I1_33__net32));
OR2X1 mul_U753(.A(n6587), .B(dpath_mulcore_b0[0]), .Y(n11854));
AND2X1 mul_U754(.A(n513), .B(n11851), .Y(dpath_mulcore_ary1_a0_I0_I1_33__net046));
OR2X1 mul_U755(.A(n6586), .B(dpath_mulcore_b1[0]), .Y(n11851));
AND2X1 mul_U756(.A(n517), .B(n11863), .Y(dpath_mulcore_ary1_a0_I0_I1_32__net32));
OR2X1 mul_U757(.A(n6590), .B(dpath_mulcore_b0[0]), .Y(n11863));
AND2X1 mul_U758(.A(n516), .B(n11860), .Y(dpath_mulcore_ary1_a0_I0_I1_32__net046));
OR2X1 mul_U759(.A(n6589), .B(dpath_mulcore_b1[0]), .Y(n11860));
AND2X1 mul_U760(.A(n520), .B(n11872), .Y(dpath_mulcore_ary1_a0_I0_I1_31__net32));
OR2X1 mul_U761(.A(n6593), .B(dpath_mulcore_b0[0]), .Y(n11872));
AND2X1 mul_U762(.A(n519), .B(n11869), .Y(dpath_mulcore_ary1_a0_I0_I1_31__net046));
OR2X1 mul_U763(.A(n6592), .B(dpath_mulcore_b1[0]), .Y(n11869));
AND2X1 mul_U764(.A(n523), .B(n11881), .Y(dpath_mulcore_ary1_a0_I0_I1_30__net32));
OR2X1 mul_U765(.A(n6596), .B(dpath_mulcore_b0[0]), .Y(n11881));
AND2X1 mul_U766(.A(n522), .B(n11878), .Y(dpath_mulcore_ary1_a0_I0_I1_30__net046));
OR2X1 mul_U767(.A(n6595), .B(dpath_mulcore_b1[0]), .Y(n11878));
AND2X1 mul_U768(.A(n526), .B(n11890), .Y(dpath_mulcore_ary1_a0_I0_I1_29__net32));
OR2X1 mul_U769(.A(n6599), .B(dpath_mulcore_b0[0]), .Y(n11890));
AND2X1 mul_U770(.A(n525), .B(n11887), .Y(dpath_mulcore_ary1_a0_I0_I1_29__net046));
OR2X1 mul_U771(.A(n6598), .B(dpath_mulcore_b1[0]), .Y(n11887));
AND2X1 mul_U772(.A(n529), .B(n11899), .Y(dpath_mulcore_ary1_a0_I0_I1_28__net32));
OR2X1 mul_U773(.A(n6602), .B(dpath_mulcore_b0[0]), .Y(n11899));
AND2X1 mul_U774(.A(n528), .B(n11896), .Y(dpath_mulcore_ary1_a0_I0_I1_28__net046));
OR2X1 mul_U775(.A(n6601), .B(dpath_mulcore_b1[0]), .Y(n11896));
AND2X1 mul_U776(.A(n532), .B(n11908), .Y(dpath_mulcore_ary1_a0_I0_I1_27__net32));
OR2X1 mul_U777(.A(n6605), .B(dpath_mulcore_b0[0]), .Y(n11908));
AND2X1 mul_U778(.A(n531), .B(n11905), .Y(dpath_mulcore_ary1_a0_I0_I1_27__net046));
OR2X1 mul_U779(.A(n6604), .B(dpath_mulcore_b1[0]), .Y(n11905));
AND2X1 mul_U780(.A(n535), .B(n11917), .Y(dpath_mulcore_ary1_a0_I0_I1_26__net32));
OR2X1 mul_U781(.A(n6608), .B(dpath_mulcore_b0[0]), .Y(n11917));
AND2X1 mul_U782(.A(n534), .B(n11914), .Y(dpath_mulcore_ary1_a0_I0_I1_26__net046));
OR2X1 mul_U783(.A(n6607), .B(dpath_mulcore_b1[0]), .Y(n11914));
AND2X1 mul_U784(.A(n538), .B(n11926), .Y(dpath_mulcore_ary1_a0_I0_I1_25__net32));
OR2X1 mul_U785(.A(n6611), .B(dpath_mulcore_b0[0]), .Y(n11926));
AND2X1 mul_U786(.A(n537), .B(n11923), .Y(dpath_mulcore_ary1_a0_I0_I1_25__net046));
OR2X1 mul_U787(.A(n6610), .B(dpath_mulcore_b1[0]), .Y(n11923));
AND2X1 mul_U788(.A(n541), .B(n11935), .Y(dpath_mulcore_ary1_a0_I0_I1_24__net32));
OR2X1 mul_U789(.A(n6614), .B(dpath_mulcore_b0[0]), .Y(n11935));
AND2X1 mul_U790(.A(n540), .B(n11932), .Y(dpath_mulcore_ary1_a0_I0_I1_24__net046));
OR2X1 mul_U791(.A(n6613), .B(dpath_mulcore_b1[0]), .Y(n11932));
AND2X1 mul_U792(.A(n544), .B(n11944), .Y(dpath_mulcore_ary1_a0_I0_I1_23__net32));
OR2X1 mul_U793(.A(n6617), .B(dpath_mulcore_b0[0]), .Y(n11944));
AND2X1 mul_U794(.A(n543), .B(n11941), .Y(dpath_mulcore_ary1_a0_I0_I1_23__net046));
OR2X1 mul_U795(.A(n6616), .B(dpath_mulcore_b1[0]), .Y(n11941));
AND2X1 mul_U796(.A(n547), .B(n11953), .Y(dpath_mulcore_ary1_a0_I0_I1_22__net32));
OR2X1 mul_U797(.A(n6620), .B(dpath_mulcore_b0[0]), .Y(n11953));
AND2X1 mul_U798(.A(n546), .B(n11950), .Y(dpath_mulcore_ary1_a0_I0_I1_22__net046));
OR2X1 mul_U799(.A(n6619), .B(dpath_mulcore_b1[0]), .Y(n11950));
AND2X1 mul_U800(.A(n550), .B(n11962), .Y(dpath_mulcore_ary1_a0_I0_I1_21__net32));
OR2X1 mul_U801(.A(n6623), .B(dpath_mulcore_b0[0]), .Y(n11962));
AND2X1 mul_U802(.A(n549), .B(n11959), .Y(dpath_mulcore_ary1_a0_I0_I1_21__net046));
OR2X1 mul_U803(.A(n6622), .B(dpath_mulcore_b1[0]), .Y(n11959));
AND2X1 mul_U804(.A(n553), .B(n11971), .Y(dpath_mulcore_ary1_a0_I0_I1_20__net32));
OR2X1 mul_U805(.A(n6626), .B(dpath_mulcore_b0[0]), .Y(n11971));
AND2X1 mul_U806(.A(n552), .B(n11968), .Y(dpath_mulcore_ary1_a0_I0_I1_20__net046));
OR2X1 mul_U807(.A(n6625), .B(dpath_mulcore_b1[0]), .Y(n11968));
AND2X1 mul_U808(.A(n556), .B(n11980), .Y(dpath_mulcore_ary1_a0_I0_I1_19__net32));
OR2X1 mul_U809(.A(n6629), .B(dpath_mulcore_b0[0]), .Y(n11980));
AND2X1 mul_U810(.A(n555), .B(n11977), .Y(dpath_mulcore_ary1_a0_I0_I1_19__net046));
OR2X1 mul_U811(.A(n6628), .B(dpath_mulcore_b1[0]), .Y(n11977));
AND2X1 mul_U812(.A(n559), .B(n11989), .Y(dpath_mulcore_ary1_a0_I0_I1_18__net32));
OR2X1 mul_U813(.A(n6632), .B(dpath_mulcore_b0[0]), .Y(n11989));
AND2X1 mul_U814(.A(n558), .B(n11986), .Y(dpath_mulcore_ary1_a0_I0_I1_18__net046));
OR2X1 mul_U815(.A(n6631), .B(dpath_mulcore_b1[0]), .Y(n11986));
AND2X1 mul_U816(.A(n562), .B(n11998), .Y(dpath_mulcore_ary1_a0_I0_I1_17__net32));
OR2X1 mul_U817(.A(n6635), .B(dpath_mulcore_b0[0]), .Y(n11998));
AND2X1 mul_U818(.A(n561), .B(n11995), .Y(dpath_mulcore_ary1_a0_I0_I1_17__net046));
OR2X1 mul_U819(.A(n6634), .B(dpath_mulcore_b1[0]), .Y(n11995));
AND2X1 mul_U820(.A(n565), .B(n12007), .Y(dpath_mulcore_ary1_a0_I0_I1_16__net32));
OR2X1 mul_U821(.A(n6638), .B(dpath_mulcore_b0[0]), .Y(n12007));
AND2X1 mul_U822(.A(n564), .B(n12004), .Y(dpath_mulcore_ary1_a0_I0_I1_16__net046));
OR2X1 mul_U823(.A(n6637), .B(dpath_mulcore_b1[0]), .Y(n12004));
AND2X1 mul_U824(.A(n568), .B(n12016), .Y(dpath_mulcore_ary1_a0_I0_I1_15__net32));
OR2X1 mul_U825(.A(n6641), .B(dpath_mulcore_b0[0]), .Y(n12016));
AND2X1 mul_U826(.A(n567), .B(n12013), .Y(dpath_mulcore_ary1_a0_I0_I1_15__net046));
OR2X1 mul_U827(.A(n6640), .B(dpath_mulcore_b1[0]), .Y(n12013));
AND2X1 mul_U828(.A(n571), .B(n12025), .Y(dpath_mulcore_ary1_a0_I0_I1_14__net32));
OR2X1 mul_U829(.A(n6644), .B(dpath_mulcore_b0[0]), .Y(n12025));
AND2X1 mul_U830(.A(n570), .B(n12022), .Y(dpath_mulcore_ary1_a0_I0_I1_14__net046));
OR2X1 mul_U831(.A(n6643), .B(dpath_mulcore_b1[0]), .Y(n12022));
INVX1 mul_U832(.A(dpath_mulcore_op1_l[2]), .Y(n9861));
AND2X1 mul_U833(.A(n224), .B(n10974), .Y(dpath_mulcore_ary1_a0_I2_I0_p1_3));
OR2X1 mul_U834(.A(n6292), .B(dpath_mulcore_b7[0]), .Y(n10974));
AND2X1 mul_U835(.A(n223), .B(n10971), .Y(dpath_mulcore_ary1_a0_I2_I0_p0_3));
OR2X1 mul_U836(.A(n6291), .B(dpath_mulcore_b6[0]), .Y(n10971));
INVX1 mul_U837(.A(n10984), .Y(n9853));
OR2X1 mul_U838(.A(n6296), .B(dpath_mulcore_b7[0]), .Y(n10984));
AND2X1 mul_U839(.A(n225), .B(n10977), .Y(dpath_mulcore_ary1_a0_I2_I0_p0_2));
OR2X1 mul_U840(.A(n6293), .B(dpath_mulcore_b6[0]), .Y(n10977));
AND2X1 mul_U841(.A(n589), .B(n12079), .Y(dpath_mulcore_ary1_a0_I0_I1_8__net32));
OR2X1 mul_U842(.A(n6662), .B(dpath_mulcore_b0[0]), .Y(n12079));
AND2X1 mul_U843(.A(n588), .B(n12076), .Y(dpath_mulcore_ary1_a0_I0_I1_8__net046));
OR2X1 mul_U844(.A(n6661), .B(dpath_mulcore_b1[0]), .Y(n12076));
INVX1 mul_U845(.A(dpath_mulcore_op1_l[59]), .Y(n10028));
AND2X1 mul_U846(.A(n739), .B(n12539), .Y(dpath_mulcore_ary1_a1_I1_I1_63__net32));
OR2X1 mul_U847(.A(n6817), .B(dpath_mulcore_b11[0]), .Y(n12539));
AND2X1 mul_U848(.A(n738), .B(n12536), .Y(dpath_mulcore_ary1_a1_I1_I1_63__net046));
OR2X1 mul_U849(.A(n6816), .B(dpath_mulcore_b12[0]), .Y(n12536));
AND2X1 mul_U850(.A(n742), .B(n12548), .Y(dpath_mulcore_ary1_a1_I1_I1_62__net32));
OR2X1 mul_U851(.A(n6820), .B(dpath_mulcore_b11[0]), .Y(n12548));
AND2X1 mul_U852(.A(n741), .B(n12545), .Y(dpath_mulcore_ary1_a1_I1_I1_62__net046));
OR2X1 mul_U853(.A(n6819), .B(dpath_mulcore_b12[0]), .Y(n12545));
AND2X1 mul_U854(.A(n920), .B(n13088), .Y(dpath_mulcore_ary1_a1_I0_I2_net078));
OR2X1 mul_U855(.A(n7001), .B(dpath_mulcore_b10[0]), .Y(n13088));
AND2X1 mul_U856(.A(n745), .B(n12557), .Y(dpath_mulcore_ary1_a1_I1_I1_61__net32));
OR2X1 mul_U857(.A(n6823), .B(dpath_mulcore_b11[0]), .Y(n12557));
AND2X1 mul_U858(.A(n744), .B(n12554), .Y(dpath_mulcore_ary1_a1_I1_I1_61__net046));
OR2X1 mul_U859(.A(n6822), .B(dpath_mulcore_b12[0]), .Y(n12554));
OR2X1 mul_U860(.A(n9482), .B(dpath_mulcore_b9[0]), .Y(n13689));
AND2X1 mul_U861(.A(n921), .B(n13091), .Y(dpath_mulcore_ary1_a1_I0_I2_net8));
OR2X1 mul_U862(.A(n7002), .B(dpath_mulcore_b10[0]), .Y(n13091));
AND2X1 mul_U863(.A(n748), .B(n12566), .Y(dpath_mulcore_ary1_a1_I1_I1_60__net32));
OR2X1 mul_U864(.A(n6826), .B(dpath_mulcore_b11[0]), .Y(n12566));
AND2X1 mul_U865(.A(n747), .B(n12563), .Y(dpath_mulcore_ary1_a1_I1_I1_60__net046));
OR2X1 mul_U866(.A(n6825), .B(dpath_mulcore_b12[0]), .Y(n12563));
AND2X1 mul_U867(.A(n922), .B(n13094), .Y(dpath_mulcore_ary1_a1_I0_I2_net15));
OR2X1 mul_U868(.A(n7003), .B(dpath_mulcore_b10[0]), .Y(n13094));
AND2X1 mul_U869(.A(n751), .B(n12575), .Y(dpath_mulcore_ary1_a1_I1_I1_59__net32));
OR2X1 mul_U870(.A(n6829), .B(dpath_mulcore_b11[0]), .Y(n12575));
AND2X1 mul_U871(.A(n750), .B(n12572), .Y(dpath_mulcore_ary1_a1_I1_I1_59__net046));
OR2X1 mul_U872(.A(n6828), .B(dpath_mulcore_b12[0]), .Y(n12572));
AND2X1 mul_U873(.A(n925), .B(n13103), .Y(dpath_mulcore_ary1_a1_I0_I2_net35));
OR2X1 mul_U874(.A(n7006), .B(dpath_mulcore_b10[0]), .Y(n13103));
AND2X1 mul_U875(.A(n754), .B(n12584), .Y(dpath_mulcore_ary1_a1_I1_I1_58__net32));
OR2X1 mul_U876(.A(n6832), .B(dpath_mulcore_b11[0]), .Y(n12584));
AND2X1 mul_U877(.A(n753), .B(n12581), .Y(dpath_mulcore_ary1_a1_I1_I1_58__net046));
OR2X1 mul_U878(.A(n6831), .B(dpath_mulcore_b12[0]), .Y(n12581));
AND2X1 mul_U879(.A(n926), .B(n13106), .Y(dpath_mulcore_ary1_a1_I0_I1_63__net043));
OR2X1 mul_U880(.A(n7007), .B(dpath_mulcore_b10[0]), .Y(n13106));
AND2X1 mul_U881(.A(n757), .B(n12593), .Y(dpath_mulcore_ary1_a1_I1_I1_57__net32));
OR2X1 mul_U882(.A(n6835), .B(dpath_mulcore_b11[0]), .Y(n12593));
AND2X1 mul_U883(.A(n756), .B(n12590), .Y(dpath_mulcore_ary1_a1_I1_I1_57__net046));
OR2X1 mul_U884(.A(n6834), .B(dpath_mulcore_b12[0]), .Y(n12590));
AND2X1 mul_U885(.A(n929), .B(n13115), .Y(dpath_mulcore_ary1_a1_I0_I1_62__net043));
OR2X1 mul_U886(.A(n7010), .B(dpath_mulcore_b10[0]), .Y(n13115));
AND2X1 mul_U887(.A(n760), .B(n12602), .Y(dpath_mulcore_ary1_a1_I1_I1_56__net32));
OR2X1 mul_U888(.A(n6838), .B(dpath_mulcore_b11[0]), .Y(n12602));
AND2X1 mul_U889(.A(n759), .B(n12599), .Y(dpath_mulcore_ary1_a1_I1_I1_56__net046));
OR2X1 mul_U890(.A(n6837), .B(dpath_mulcore_b12[0]), .Y(n12599));
AND2X1 mul_U891(.A(n932), .B(n13124), .Y(dpath_mulcore_ary1_a1_I0_I1_61__net043));
OR2X1 mul_U892(.A(n7013), .B(dpath_mulcore_b10[0]), .Y(n13124));
AND2X1 mul_U893(.A(n763), .B(n12611), .Y(dpath_mulcore_ary1_a1_I1_I1_55__net32));
OR2X1 mul_U894(.A(n6841), .B(dpath_mulcore_b11[0]), .Y(n12611));
AND2X1 mul_U895(.A(n762), .B(n12608), .Y(dpath_mulcore_ary1_a1_I1_I1_55__net046));
OR2X1 mul_U896(.A(n6840), .B(dpath_mulcore_b12[0]), .Y(n12608));
AND2X1 mul_U897(.A(n935), .B(n13133), .Y(dpath_mulcore_ary1_a1_I0_I1_60__net043));
OR2X1 mul_U898(.A(n7016), .B(dpath_mulcore_b10[0]), .Y(n13133));
AND2X1 mul_U899(.A(n766), .B(n12620), .Y(dpath_mulcore_ary1_a1_I1_I1_54__net32));
OR2X1 mul_U900(.A(n6844), .B(dpath_mulcore_b11[0]), .Y(n12620));
AND2X1 mul_U901(.A(n765), .B(n12617), .Y(dpath_mulcore_ary1_a1_I1_I1_54__net046));
OR2X1 mul_U902(.A(n6843), .B(dpath_mulcore_b12[0]), .Y(n12617));
AND2X1 mul_U903(.A(n938), .B(n13142), .Y(dpath_mulcore_ary1_a1_I0_I1_59__net043));
OR2X1 mul_U904(.A(n7019), .B(dpath_mulcore_b10[0]), .Y(n13142));
AND2X1 mul_U905(.A(n769), .B(n12629), .Y(dpath_mulcore_ary1_a1_I1_I1_53__net32));
OR2X1 mul_U906(.A(n6847), .B(dpath_mulcore_b11[0]), .Y(n12629));
AND2X1 mul_U907(.A(n768), .B(n12626), .Y(dpath_mulcore_ary1_a1_I1_I1_53__net046));
OR2X1 mul_U908(.A(n6846), .B(dpath_mulcore_b12[0]), .Y(n12626));
AND2X1 mul_U909(.A(n941), .B(n13151), .Y(dpath_mulcore_ary1_a1_I0_I1_58__net043));
OR2X1 mul_U910(.A(n7022), .B(dpath_mulcore_b10[0]), .Y(n13151));
AND2X1 mul_U911(.A(n772), .B(n12638), .Y(dpath_mulcore_ary1_a1_I1_I1_52__net32));
OR2X1 mul_U912(.A(n6850), .B(dpath_mulcore_b11[0]), .Y(n12638));
AND2X1 mul_U913(.A(n771), .B(n12635), .Y(dpath_mulcore_ary1_a1_I1_I1_52__net046));
OR2X1 mul_U914(.A(n6849), .B(dpath_mulcore_b12[0]), .Y(n12635));
AND2X1 mul_U915(.A(n944), .B(n13160), .Y(dpath_mulcore_ary1_a1_I0_I1_57__net043));
OR2X1 mul_U916(.A(n7025), .B(dpath_mulcore_b10[0]), .Y(n13160));
AND2X1 mul_U917(.A(n775), .B(n12647), .Y(dpath_mulcore_ary1_a1_I1_I1_51__net32));
OR2X1 mul_U918(.A(n6853), .B(dpath_mulcore_b11[0]), .Y(n12647));
AND2X1 mul_U919(.A(n774), .B(n12644), .Y(dpath_mulcore_ary1_a1_I1_I1_51__net046));
OR2X1 mul_U920(.A(n6852), .B(dpath_mulcore_b12[0]), .Y(n12644));
AND2X1 mul_U921(.A(n947), .B(n13169), .Y(dpath_mulcore_ary1_a1_I0_I1_56__net043));
OR2X1 mul_U922(.A(n7028), .B(dpath_mulcore_b10[0]), .Y(n13169));
AND2X1 mul_U923(.A(n778), .B(n12656), .Y(dpath_mulcore_ary1_a1_I1_I1_50__net32));
OR2X1 mul_U924(.A(n6856), .B(dpath_mulcore_b11[0]), .Y(n12656));
AND2X1 mul_U925(.A(n777), .B(n12653), .Y(dpath_mulcore_ary1_a1_I1_I1_50__net046));
OR2X1 mul_U926(.A(n6855), .B(dpath_mulcore_b12[0]), .Y(n12653));
AND2X1 mul_U927(.A(n950), .B(n13178), .Y(dpath_mulcore_ary1_a1_I0_I1_55__net043));
OR2X1 mul_U928(.A(n7031), .B(dpath_mulcore_b10[0]), .Y(n13178));
AND2X1 mul_U929(.A(n781), .B(n12665), .Y(dpath_mulcore_ary1_a1_I1_I1_49__net32));
OR2X1 mul_U930(.A(n6859), .B(dpath_mulcore_b11[0]), .Y(n12665));
AND2X1 mul_U931(.A(n780), .B(n12662), .Y(dpath_mulcore_ary1_a1_I1_I1_49__net046));
OR2X1 mul_U932(.A(n6858), .B(dpath_mulcore_b12[0]), .Y(n12662));
AND2X1 mul_U933(.A(n953), .B(n13187), .Y(dpath_mulcore_ary1_a1_I0_I1_54__net043));
OR2X1 mul_U934(.A(n7034), .B(dpath_mulcore_b10[0]), .Y(n13187));
AND2X1 mul_U935(.A(n784), .B(n12674), .Y(dpath_mulcore_ary1_a1_I1_I1_48__net32));
OR2X1 mul_U936(.A(n6862), .B(dpath_mulcore_b11[0]), .Y(n12674));
AND2X1 mul_U937(.A(n783), .B(n12671), .Y(dpath_mulcore_ary1_a1_I1_I1_48__net046));
OR2X1 mul_U938(.A(n6861), .B(dpath_mulcore_b12[0]), .Y(n12671));
AND2X1 mul_U939(.A(n956), .B(n13196), .Y(dpath_mulcore_ary1_a1_I0_I1_53__net043));
OR2X1 mul_U940(.A(n7037), .B(dpath_mulcore_b10[0]), .Y(n13196));
AND2X1 mul_U941(.A(n787), .B(n12683), .Y(dpath_mulcore_ary1_a1_I1_I1_47__net32));
OR2X1 mul_U942(.A(n6865), .B(dpath_mulcore_b11[0]), .Y(n12683));
AND2X1 mul_U943(.A(n786), .B(n12680), .Y(dpath_mulcore_ary1_a1_I1_I1_47__net046));
OR2X1 mul_U944(.A(n6864), .B(dpath_mulcore_b12[0]), .Y(n12680));
AND2X1 mul_U945(.A(n959), .B(n13205), .Y(dpath_mulcore_ary1_a1_I0_I1_52__net043));
OR2X1 mul_U946(.A(n7040), .B(dpath_mulcore_b10[0]), .Y(n13205));
AND2X1 mul_U947(.A(n790), .B(n12692), .Y(dpath_mulcore_ary1_a1_I1_I1_46__net32));
OR2X1 mul_U948(.A(n6868), .B(dpath_mulcore_b11[0]), .Y(n12692));
AND2X1 mul_U949(.A(n789), .B(n12689), .Y(dpath_mulcore_ary1_a1_I1_I1_46__net046));
OR2X1 mul_U950(.A(n6867), .B(dpath_mulcore_b12[0]), .Y(n12689));
AND2X1 mul_U951(.A(n962), .B(n13214), .Y(dpath_mulcore_ary1_a1_I0_I1_51__net043));
OR2X1 mul_U952(.A(n7043), .B(dpath_mulcore_b10[0]), .Y(n13214));
AND2X1 mul_U953(.A(n793), .B(n12701), .Y(dpath_mulcore_ary1_a1_I1_I1_45__net32));
OR2X1 mul_U954(.A(n6871), .B(dpath_mulcore_b11[0]), .Y(n12701));
AND2X1 mul_U955(.A(n792), .B(n12698), .Y(dpath_mulcore_ary1_a1_I1_I1_45__net046));
OR2X1 mul_U956(.A(n6870), .B(dpath_mulcore_b12[0]), .Y(n12698));
AND2X1 mul_U957(.A(n965), .B(n13223), .Y(dpath_mulcore_ary1_a1_I0_I1_50__net043));
OR2X1 mul_U958(.A(n7046), .B(dpath_mulcore_b10[0]), .Y(n13223));
AND2X1 mul_U959(.A(n796), .B(n12710), .Y(dpath_mulcore_ary1_a1_I1_I1_44__net32));
OR2X1 mul_U960(.A(n6874), .B(dpath_mulcore_b11[0]), .Y(n12710));
AND2X1 mul_U961(.A(n795), .B(n12707), .Y(dpath_mulcore_ary1_a1_I1_I1_44__net046));
OR2X1 mul_U962(.A(n6873), .B(dpath_mulcore_b12[0]), .Y(n12707));
AND2X1 mul_U963(.A(n968), .B(n13232), .Y(dpath_mulcore_ary1_a1_I0_I1_49__net043));
OR2X1 mul_U964(.A(n7049), .B(dpath_mulcore_b10[0]), .Y(n13232));
AND2X1 mul_U965(.A(n799), .B(n12719), .Y(dpath_mulcore_ary1_a1_I1_I1_43__net32));
OR2X1 mul_U966(.A(n6877), .B(dpath_mulcore_b11[0]), .Y(n12719));
AND2X1 mul_U967(.A(n798), .B(n12716), .Y(dpath_mulcore_ary1_a1_I1_I1_43__net046));
OR2X1 mul_U968(.A(n6876), .B(dpath_mulcore_b12[0]), .Y(n12716));
AND2X1 mul_U969(.A(n971), .B(n13241), .Y(dpath_mulcore_ary1_a1_I0_I1_48__net043));
OR2X1 mul_U970(.A(n7052), .B(dpath_mulcore_b10[0]), .Y(n13241));
AND2X1 mul_U971(.A(n802), .B(n12728), .Y(dpath_mulcore_ary1_a1_I1_I1_42__net32));
OR2X1 mul_U972(.A(n6880), .B(dpath_mulcore_b11[0]), .Y(n12728));
AND2X1 mul_U973(.A(n801), .B(n12725), .Y(dpath_mulcore_ary1_a1_I1_I1_42__net046));
OR2X1 mul_U974(.A(n6879), .B(dpath_mulcore_b12[0]), .Y(n12725));
AND2X1 mul_U975(.A(n974), .B(n13250), .Y(dpath_mulcore_ary1_a1_I0_I1_47__net043));
OR2X1 mul_U976(.A(n7055), .B(dpath_mulcore_b10[0]), .Y(n13250));
AND2X1 mul_U977(.A(n805), .B(n12737), .Y(dpath_mulcore_ary1_a1_I1_I1_41__net32));
OR2X1 mul_U978(.A(n6883), .B(dpath_mulcore_b11[0]), .Y(n12737));
AND2X1 mul_U979(.A(n804), .B(n12734), .Y(dpath_mulcore_ary1_a1_I1_I1_41__net046));
OR2X1 mul_U980(.A(n6882), .B(dpath_mulcore_b12[0]), .Y(n12734));
AND2X1 mul_U981(.A(n977), .B(n13259), .Y(dpath_mulcore_ary1_a1_I0_I1_46__net043));
OR2X1 mul_U982(.A(n7058), .B(dpath_mulcore_b10[0]), .Y(n13259));
AND2X1 mul_U983(.A(n808), .B(n12746), .Y(dpath_mulcore_ary1_a1_I1_I1_40__net32));
OR2X1 mul_U984(.A(n6886), .B(dpath_mulcore_b11[0]), .Y(n12746));
AND2X1 mul_U985(.A(n807), .B(n12743), .Y(dpath_mulcore_ary1_a1_I1_I1_40__net046));
OR2X1 mul_U986(.A(n6885), .B(dpath_mulcore_b12[0]), .Y(n12743));
AND2X1 mul_U987(.A(n980), .B(n13268), .Y(dpath_mulcore_ary1_a1_I0_I1_45__net043));
OR2X1 mul_U988(.A(n7061), .B(dpath_mulcore_b10[0]), .Y(n13268));
AND2X1 mul_U989(.A(n811), .B(n12755), .Y(dpath_mulcore_ary1_a1_I1_I1_39__net32));
OR2X1 mul_U990(.A(n6889), .B(dpath_mulcore_b11[0]), .Y(n12755));
AND2X1 mul_U991(.A(n810), .B(n12752), .Y(dpath_mulcore_ary1_a1_I1_I1_39__net046));
OR2X1 mul_U992(.A(n6888), .B(dpath_mulcore_b12[0]), .Y(n12752));
AND2X1 mul_U993(.A(n983), .B(n13277), .Y(dpath_mulcore_ary1_a1_I0_I1_44__net043));
OR2X1 mul_U994(.A(n7064), .B(dpath_mulcore_b10[0]), .Y(n13277));
AND2X1 mul_U995(.A(n814), .B(n12764), .Y(dpath_mulcore_ary1_a1_I1_I1_38__net32));
OR2X1 mul_U996(.A(n6892), .B(dpath_mulcore_b11[0]), .Y(n12764));
AND2X1 mul_U997(.A(n813), .B(n12761), .Y(dpath_mulcore_ary1_a1_I1_I1_38__net046));
OR2X1 mul_U998(.A(n6891), .B(dpath_mulcore_b12[0]), .Y(n12761));
AND2X1 mul_U999(.A(n986), .B(n13286), .Y(dpath_mulcore_ary1_a1_I0_I1_43__net043));
OR2X1 mul_U1000(.A(n7067), .B(dpath_mulcore_b10[0]), .Y(n13286));
AND2X1 mul_U1001(.A(n817), .B(n12773), .Y(dpath_mulcore_ary1_a1_I1_I1_37__net32));
OR2X1 mul_U1002(.A(n6895), .B(dpath_mulcore_b11[0]), .Y(n12773));
AND2X1 mul_U1003(.A(n816), .B(n12770), .Y(dpath_mulcore_ary1_a1_I1_I1_37__net046));
OR2X1 mul_U1004(.A(n6894), .B(dpath_mulcore_b12[0]), .Y(n12770));
AND2X1 mul_U1005(.A(n989), .B(n13295), .Y(dpath_mulcore_ary1_a1_I0_I1_42__net043));
OR2X1 mul_U1006(.A(n7070), .B(dpath_mulcore_b10[0]), .Y(n13295));
AND2X1 mul_U1007(.A(n820), .B(n12782), .Y(dpath_mulcore_ary1_a1_I1_I1_36__net32));
OR2X1 mul_U1008(.A(n6898), .B(dpath_mulcore_b11[0]), .Y(n12782));
AND2X1 mul_U1009(.A(n819), .B(n12779), .Y(dpath_mulcore_ary1_a1_I1_I1_36__net046));
OR2X1 mul_U1010(.A(n6897), .B(dpath_mulcore_b12[0]), .Y(n12779));
AND2X1 mul_U1011(.A(n992), .B(n13304), .Y(dpath_mulcore_ary1_a1_I0_I1_41__net043));
OR2X1 mul_U1012(.A(n7073), .B(dpath_mulcore_b10[0]), .Y(n13304));
AND2X1 mul_U1013(.A(n823), .B(n12791), .Y(dpath_mulcore_ary1_a1_I1_I1_35__net32));
OR2X1 mul_U1014(.A(n6901), .B(dpath_mulcore_b11[0]), .Y(n12791));
AND2X1 mul_U1015(.A(n822), .B(n12788), .Y(dpath_mulcore_ary1_a1_I1_I1_35__net046));
OR2X1 mul_U1016(.A(n6900), .B(dpath_mulcore_b12[0]), .Y(n12788));
AND2X1 mul_U1017(.A(n995), .B(n13313), .Y(dpath_mulcore_ary1_a1_I0_I1_40__net043));
OR2X1 mul_U1018(.A(n7076), .B(dpath_mulcore_b10[0]), .Y(n13313));
AND2X1 mul_U1019(.A(n826), .B(n12800), .Y(dpath_mulcore_ary1_a1_I1_I1_34__net32));
OR2X1 mul_U1020(.A(n6904), .B(dpath_mulcore_b11[0]), .Y(n12800));
AND2X1 mul_U1021(.A(n825), .B(n12797), .Y(dpath_mulcore_ary1_a1_I1_I1_34__net046));
OR2X1 mul_U1022(.A(n6903), .B(dpath_mulcore_b12[0]), .Y(n12797));
AND2X1 mul_U1023(.A(n998), .B(n13322), .Y(dpath_mulcore_ary1_a1_I0_I1_39__net043));
OR2X1 mul_U1024(.A(n7079), .B(dpath_mulcore_b10[0]), .Y(n13322));
AND2X1 mul_U1025(.A(n829), .B(n12809), .Y(dpath_mulcore_ary1_a1_I1_I1_33__net32));
OR2X1 mul_U1026(.A(n6907), .B(dpath_mulcore_b11[0]), .Y(n12809));
AND2X1 mul_U1027(.A(n828), .B(n12806), .Y(dpath_mulcore_ary1_a1_I1_I1_33__net046));
OR2X1 mul_U1028(.A(n6906), .B(dpath_mulcore_b12[0]), .Y(n12806));
AND2X1 mul_U1029(.A(n1001), .B(n13331), .Y(dpath_mulcore_ary1_a1_I0_I1_38__net043));
OR2X1 mul_U1030(.A(n7082), .B(dpath_mulcore_b10[0]), .Y(n13331));
AND2X1 mul_U1031(.A(n832), .B(n12818), .Y(dpath_mulcore_ary1_a1_I1_I1_32__net32));
OR2X1 mul_U1032(.A(n6910), .B(dpath_mulcore_b11[0]), .Y(n12818));
AND2X1 mul_U1033(.A(n831), .B(n12815), .Y(dpath_mulcore_ary1_a1_I1_I1_32__net046));
OR2X1 mul_U1034(.A(n6909), .B(dpath_mulcore_b12[0]), .Y(n12815));
AND2X1 mul_U1035(.A(n1004), .B(n13340), .Y(dpath_mulcore_ary1_a1_I0_I1_37__net043));
OR2X1 mul_U1036(.A(n7085), .B(dpath_mulcore_b10[0]), .Y(n13340));
AND2X1 mul_U1037(.A(n835), .B(n12827), .Y(dpath_mulcore_ary1_a1_I1_I1_31__net32));
OR2X1 mul_U1038(.A(n6913), .B(dpath_mulcore_b11[0]), .Y(n12827));
AND2X1 mul_U1039(.A(n834), .B(n12824), .Y(dpath_mulcore_ary1_a1_I1_I1_31__net046));
OR2X1 mul_U1040(.A(n6912), .B(dpath_mulcore_b12[0]), .Y(n12824));
AND2X1 mul_U1041(.A(n1007), .B(n13349), .Y(dpath_mulcore_ary1_a1_I0_I1_36__net043));
OR2X1 mul_U1042(.A(n7088), .B(dpath_mulcore_b10[0]), .Y(n13349));
AND2X1 mul_U1043(.A(n838), .B(n12836), .Y(dpath_mulcore_ary1_a1_I1_I1_30__net32));
OR2X1 mul_U1044(.A(n6916), .B(dpath_mulcore_b11[0]), .Y(n12836));
AND2X1 mul_U1045(.A(n837), .B(n12833), .Y(dpath_mulcore_ary1_a1_I1_I1_30__net046));
OR2X1 mul_U1046(.A(n6915), .B(dpath_mulcore_b12[0]), .Y(n12833));
AND2X1 mul_U1047(.A(n1010), .B(n13358), .Y(dpath_mulcore_ary1_a1_I0_I1_35__net043));
OR2X1 mul_U1048(.A(n7091), .B(dpath_mulcore_b10[0]), .Y(n13358));
AND2X1 mul_U1049(.A(n841), .B(n12845), .Y(dpath_mulcore_ary1_a1_I1_I1_29__net32));
OR2X1 mul_U1050(.A(n6919), .B(dpath_mulcore_b11[0]), .Y(n12845));
AND2X1 mul_U1051(.A(n840), .B(n12842), .Y(dpath_mulcore_ary1_a1_I1_I1_29__net046));
OR2X1 mul_U1052(.A(n6918), .B(dpath_mulcore_b12[0]), .Y(n12842));
AND2X1 mul_U1053(.A(n1013), .B(n13367), .Y(dpath_mulcore_ary1_a1_I0_I1_34__net043));
OR2X1 mul_U1054(.A(n7094), .B(dpath_mulcore_b10[0]), .Y(n13367));
AND2X1 mul_U1055(.A(n844), .B(n12854), .Y(dpath_mulcore_ary1_a1_I1_I1_28__net32));
OR2X1 mul_U1056(.A(n6922), .B(dpath_mulcore_b11[0]), .Y(n12854));
AND2X1 mul_U1057(.A(n843), .B(n12851), .Y(dpath_mulcore_ary1_a1_I1_I1_28__net046));
OR2X1 mul_U1058(.A(n6921), .B(dpath_mulcore_b12[0]), .Y(n12851));
AND2X1 mul_U1059(.A(n1016), .B(n13376), .Y(dpath_mulcore_ary1_a1_I0_I1_33__net043));
OR2X1 mul_U1060(.A(n7097), .B(dpath_mulcore_b10[0]), .Y(n13376));
AND2X1 mul_U1061(.A(n847), .B(n12863), .Y(dpath_mulcore_ary1_a1_I1_I1_27__net32));
OR2X1 mul_U1062(.A(n6925), .B(dpath_mulcore_b11[0]), .Y(n12863));
AND2X1 mul_U1063(.A(n846), .B(n12860), .Y(dpath_mulcore_ary1_a1_I1_I1_27__net046));
OR2X1 mul_U1064(.A(n6924), .B(dpath_mulcore_b12[0]), .Y(n12860));
AND2X1 mul_U1065(.A(n1019), .B(n13385), .Y(dpath_mulcore_ary1_a1_I0_I1_32__net043));
OR2X1 mul_U1066(.A(n7100), .B(dpath_mulcore_b10[0]), .Y(n13385));
AND2X1 mul_U1067(.A(n850), .B(n12872), .Y(dpath_mulcore_ary1_a1_I1_I1_26__net32));
OR2X1 mul_U1068(.A(n6928), .B(dpath_mulcore_b11[0]), .Y(n12872));
AND2X1 mul_U1069(.A(n849), .B(n12869), .Y(dpath_mulcore_ary1_a1_I1_I1_26__net046));
OR2X1 mul_U1070(.A(n6927), .B(dpath_mulcore_b12[0]), .Y(n12869));
AND2X1 mul_U1071(.A(n1022), .B(n13394), .Y(dpath_mulcore_ary1_a1_I0_I1_31__net043));
OR2X1 mul_U1072(.A(n7103), .B(dpath_mulcore_b10[0]), .Y(n13394));
AND2X1 mul_U1073(.A(n853), .B(n12881), .Y(dpath_mulcore_ary1_a1_I1_I1_25__net32));
OR2X1 mul_U1074(.A(n6931), .B(dpath_mulcore_b11[0]), .Y(n12881));
AND2X1 mul_U1075(.A(n852), .B(n12878), .Y(dpath_mulcore_ary1_a1_I1_I1_25__net046));
OR2X1 mul_U1076(.A(n6930), .B(dpath_mulcore_b12[0]), .Y(n12878));
AND2X1 mul_U1077(.A(n1025), .B(n13403), .Y(dpath_mulcore_ary1_a1_I0_I1_30__net043));
OR2X1 mul_U1078(.A(n7106), .B(dpath_mulcore_b10[0]), .Y(n13403));
AND2X1 mul_U1079(.A(n856), .B(n12890), .Y(dpath_mulcore_ary1_a1_I1_I1_24__net32));
OR2X1 mul_U1080(.A(n6934), .B(dpath_mulcore_b11[0]), .Y(n12890));
AND2X1 mul_U1081(.A(n855), .B(n12887), .Y(dpath_mulcore_ary1_a1_I1_I1_24__net046));
OR2X1 mul_U1082(.A(n6933), .B(dpath_mulcore_b12[0]), .Y(n12887));
AND2X1 mul_U1083(.A(n1028), .B(n13412), .Y(dpath_mulcore_ary1_a1_I0_I1_29__net043));
OR2X1 mul_U1084(.A(n7109), .B(dpath_mulcore_b10[0]), .Y(n13412));
AND2X1 mul_U1085(.A(n859), .B(n12899), .Y(dpath_mulcore_ary1_a1_I1_I1_23__net32));
OR2X1 mul_U1086(.A(n6937), .B(dpath_mulcore_b11[0]), .Y(n12899));
AND2X1 mul_U1087(.A(n858), .B(n12896), .Y(dpath_mulcore_ary1_a1_I1_I1_23__net046));
OR2X1 mul_U1088(.A(n6936), .B(dpath_mulcore_b12[0]), .Y(n12896));
AND2X1 mul_U1089(.A(n1031), .B(n13421), .Y(dpath_mulcore_ary1_a1_I0_I1_28__net043));
OR2X1 mul_U1090(.A(n7112), .B(dpath_mulcore_b10[0]), .Y(n13421));
AND2X1 mul_U1091(.A(n862), .B(n12908), .Y(dpath_mulcore_ary1_a1_I1_I1_22__net32));
OR2X1 mul_U1092(.A(n6940), .B(dpath_mulcore_b11[0]), .Y(n12908));
AND2X1 mul_U1093(.A(n861), .B(n12905), .Y(dpath_mulcore_ary1_a1_I1_I1_22__net046));
OR2X1 mul_U1094(.A(n6939), .B(dpath_mulcore_b12[0]), .Y(n12905));
AND2X1 mul_U1095(.A(n1034), .B(n13430), .Y(dpath_mulcore_ary1_a1_I0_I1_27__net043));
OR2X1 mul_U1096(.A(n7115), .B(dpath_mulcore_b10[0]), .Y(n13430));
AND2X1 mul_U1097(.A(n865), .B(n12917), .Y(dpath_mulcore_ary1_a1_I1_I1_21__net32));
OR2X1 mul_U1098(.A(n6943), .B(dpath_mulcore_b11[0]), .Y(n12917));
AND2X1 mul_U1099(.A(n864), .B(n12914), .Y(dpath_mulcore_ary1_a1_I1_I1_21__net046));
OR2X1 mul_U1100(.A(n6942), .B(dpath_mulcore_b12[0]), .Y(n12914));
AND2X1 mul_U1101(.A(n1037), .B(n13439), .Y(dpath_mulcore_ary1_a1_I0_I1_26__net043));
OR2X1 mul_U1102(.A(n7118), .B(dpath_mulcore_b10[0]), .Y(n13439));
AND2X1 mul_U1103(.A(n868), .B(n12926), .Y(dpath_mulcore_ary1_a1_I1_I1_20__net32));
OR2X1 mul_U1104(.A(n6946), .B(dpath_mulcore_b11[0]), .Y(n12926));
AND2X1 mul_U1105(.A(n867), .B(n12923), .Y(dpath_mulcore_ary1_a1_I1_I1_20__net046));
OR2X1 mul_U1106(.A(n6945), .B(dpath_mulcore_b12[0]), .Y(n12923));
AND2X1 mul_U1107(.A(n1040), .B(n13448), .Y(dpath_mulcore_ary1_a1_I0_I1_25__net043));
OR2X1 mul_U1108(.A(n7121), .B(dpath_mulcore_b10[0]), .Y(n13448));
AND2X1 mul_U1109(.A(n871), .B(n12935), .Y(dpath_mulcore_ary1_a1_I1_I1_19__net32));
OR2X1 mul_U1110(.A(n6949), .B(dpath_mulcore_b11[0]), .Y(n12935));
AND2X1 mul_U1111(.A(n870), .B(n12932), .Y(dpath_mulcore_ary1_a1_I1_I1_19__net046));
OR2X1 mul_U1112(.A(n6948), .B(dpath_mulcore_b12[0]), .Y(n12932));
AND2X1 mul_U1113(.A(n1043), .B(n13457), .Y(dpath_mulcore_ary1_a1_I0_I1_24__net043));
OR2X1 mul_U1114(.A(n7124), .B(dpath_mulcore_b10[0]), .Y(n13457));
AND2X1 mul_U1115(.A(n874), .B(n12944), .Y(dpath_mulcore_ary1_a1_I1_I1_18__net32));
OR2X1 mul_U1116(.A(n6952), .B(dpath_mulcore_b11[0]), .Y(n12944));
AND2X1 mul_U1117(.A(n873), .B(n12941), .Y(dpath_mulcore_ary1_a1_I1_I1_18__net046));
OR2X1 mul_U1118(.A(n6951), .B(dpath_mulcore_b12[0]), .Y(n12941));
AND2X1 mul_U1119(.A(n1046), .B(n13466), .Y(dpath_mulcore_ary1_a1_I0_I1_23__net043));
OR2X1 mul_U1120(.A(n7127), .B(dpath_mulcore_b10[0]), .Y(n13466));
AND2X1 mul_U1121(.A(n877), .B(n12953), .Y(dpath_mulcore_ary1_a1_I1_I1_17__net32));
OR2X1 mul_U1122(.A(n6955), .B(dpath_mulcore_b11[0]), .Y(n12953));
AND2X1 mul_U1123(.A(n876), .B(n12950), .Y(dpath_mulcore_ary1_a1_I1_I1_17__net046));
OR2X1 mul_U1124(.A(n6954), .B(dpath_mulcore_b12[0]), .Y(n12950));
AND2X1 mul_U1125(.A(n1049), .B(n13475), .Y(dpath_mulcore_ary1_a1_I0_I1_22__net043));
OR2X1 mul_U1126(.A(n7130), .B(dpath_mulcore_b10[0]), .Y(n13475));
AND2X1 mul_U1127(.A(n880), .B(n12962), .Y(dpath_mulcore_ary1_a1_I1_I1_16__net32));
OR2X1 mul_U1128(.A(n6958), .B(dpath_mulcore_b11[0]), .Y(n12962));
AND2X1 mul_U1129(.A(n879), .B(n12959), .Y(dpath_mulcore_ary1_a1_I1_I1_16__net046));
OR2X1 mul_U1130(.A(n6957), .B(dpath_mulcore_b12[0]), .Y(n12959));
AND2X1 mul_U1131(.A(n1052), .B(n13484), .Y(dpath_mulcore_ary1_a1_I0_I1_21__net043));
OR2X1 mul_U1132(.A(n7133), .B(dpath_mulcore_b10[0]), .Y(n13484));
AND2X1 mul_U1133(.A(n883), .B(n12971), .Y(dpath_mulcore_ary1_a1_I1_I1_15__net32));
OR2X1 mul_U1134(.A(n6961), .B(dpath_mulcore_b11[0]), .Y(n12971));
AND2X1 mul_U1135(.A(n882), .B(n12968), .Y(dpath_mulcore_ary1_a1_I1_I1_15__net046));
OR2X1 mul_U1136(.A(n6960), .B(dpath_mulcore_b12[0]), .Y(n12968));
AND2X1 mul_U1137(.A(n1055), .B(n13493), .Y(dpath_mulcore_ary1_a1_I0_I1_20__net043));
OR2X1 mul_U1138(.A(n7136), .B(dpath_mulcore_b10[0]), .Y(n13493));
AND2X1 mul_U1139(.A(n886), .B(n12980), .Y(dpath_mulcore_ary1_a1_I1_I1_14__net32));
OR2X1 mul_U1140(.A(n6964), .B(dpath_mulcore_b11[0]), .Y(n12980));
AND2X1 mul_U1141(.A(n885), .B(n12977), .Y(dpath_mulcore_ary1_a1_I1_I1_14__net046));
OR2X1 mul_U1142(.A(n6963), .B(dpath_mulcore_b12[0]), .Y(n12977));
AND2X1 mul_U1143(.A(n1058), .B(n13502), .Y(dpath_mulcore_ary1_a1_I0_I1_19__net043));
OR2X1 mul_U1144(.A(n7139), .B(dpath_mulcore_b10[0]), .Y(n13502));
AND2X1 mul_U1145(.A(n889), .B(n12989), .Y(dpath_mulcore_ary1_a1_I1_I1_13__net32));
OR2X1 mul_U1146(.A(n6967), .B(dpath_mulcore_b11[0]), .Y(n12989));
AND2X1 mul_U1147(.A(n888), .B(n12986), .Y(dpath_mulcore_ary1_a1_I1_I1_13__net046));
OR2X1 mul_U1148(.A(n6966), .B(dpath_mulcore_b12[0]), .Y(n12986));
AND2X1 mul_U1149(.A(n1061), .B(n13511), .Y(dpath_mulcore_ary1_a1_I0_I1_18__net043));
OR2X1 mul_U1150(.A(n7142), .B(dpath_mulcore_b10[0]), .Y(n13511));
AND2X1 mul_U1151(.A(n892), .B(n12998), .Y(dpath_mulcore_ary1_a1_I1_I1_12__net32));
OR2X1 mul_U1152(.A(n6970), .B(dpath_mulcore_b11[0]), .Y(n12998));
AND2X1 mul_U1153(.A(n891), .B(n12995), .Y(dpath_mulcore_ary1_a1_I1_I1_12__net046));
OR2X1 mul_U1154(.A(n6969), .B(dpath_mulcore_b12[0]), .Y(n12995));
AND2X1 mul_U1155(.A(n1064), .B(n13520), .Y(dpath_mulcore_ary1_a1_I0_I1_17__net043));
OR2X1 mul_U1156(.A(n7145), .B(dpath_mulcore_b10[0]), .Y(n13520));
AND2X1 mul_U1157(.A(n895), .B(n13007), .Y(dpath_mulcore_ary1_a1_I1_I1_11__net32));
OR2X1 mul_U1158(.A(n6973), .B(dpath_mulcore_b11[0]), .Y(n13007));
AND2X1 mul_U1159(.A(n894), .B(n13004), .Y(dpath_mulcore_ary1_a1_I1_I1_11__net046));
OR2X1 mul_U1160(.A(n6972), .B(dpath_mulcore_b12[0]), .Y(n13004));
AND2X1 mul_U1161(.A(n1067), .B(n13529), .Y(dpath_mulcore_ary1_a1_I0_I1_16__net043));
OR2X1 mul_U1162(.A(n7148), .B(dpath_mulcore_b10[0]), .Y(n13529));
AND2X1 mul_U1163(.A(n898), .B(n13016), .Y(dpath_mulcore_ary1_a1_I1_I1_10__net32));
OR2X1 mul_U1164(.A(n6976), .B(dpath_mulcore_b11[0]), .Y(n13016));
AND2X1 mul_U1165(.A(n897), .B(n13013), .Y(dpath_mulcore_ary1_a1_I1_I1_10__net046));
OR2X1 mul_U1166(.A(n6975), .B(dpath_mulcore_b12[0]), .Y(n13013));
AND2X1 mul_U1167(.A(n1070), .B(n13538), .Y(dpath_mulcore_ary1_a1_I0_I1_15__net043));
OR2X1 mul_U1168(.A(n7151), .B(dpath_mulcore_b10[0]), .Y(n13538));
AND2X1 mul_U1169(.A(n901), .B(n13025), .Y(dpath_mulcore_ary1_a1_I1_I1_9__net32));
OR2X1 mul_U1170(.A(n6979), .B(dpath_mulcore_b11[0]), .Y(n13025));
AND2X1 mul_U1171(.A(n900), .B(n13022), .Y(dpath_mulcore_ary1_a1_I1_I1_9__net046));
OR2X1 mul_U1172(.A(n6978), .B(dpath_mulcore_b12[0]), .Y(n13022));
AND2X1 mul_U1173(.A(n1073), .B(n13547), .Y(dpath_mulcore_ary1_a1_I0_I1_14__net043));
OR2X1 mul_U1174(.A(n7154), .B(dpath_mulcore_b10[0]), .Y(n13547));
AND2X1 mul_U1175(.A(n904), .B(n13034), .Y(dpath_mulcore_ary1_a1_I1_I1_8__net32));
OR2X1 mul_U1176(.A(n6982), .B(dpath_mulcore_b11[0]), .Y(n13034));
AND2X1 mul_U1177(.A(n903), .B(n13031), .Y(dpath_mulcore_ary1_a1_I1_I1_8__net046));
OR2X1 mul_U1178(.A(n6981), .B(dpath_mulcore_b12[0]), .Y(n13031));
AND2X1 mul_U1179(.A(n907), .B(n13043), .Y(dpath_mulcore_ary1_a1_I1_I1_7__net32));
OR2X1 mul_U1180(.A(n6985), .B(dpath_mulcore_b11[0]), .Y(n13043));
AND2X1 mul_U1181(.A(n906), .B(n13040), .Y(dpath_mulcore_ary1_a1_I1_I1_7__net046));
OR2X1 mul_U1182(.A(n6984), .B(dpath_mulcore_b12[0]), .Y(n13040));
AND2X1 mul_U1183(.A(n1078), .B(n13562), .Y(dpath_mulcore_ary1_a1_I0_I1_13__net32));
OR2X1 mul_U1184(.A(n7159), .B(dpath_mulcore_b8[0]), .Y(n13562));
AND2X1 mul_U1185(.A(n1077), .B(n13559), .Y(dpath_mulcore_ary1_a1_I0_I1_13__net046));
OR2X1 mul_U1186(.A(n7158), .B(dpath_mulcore_b9[0]), .Y(n13559));
AND2X1 mul_U1187(.A(n910), .B(n13052), .Y(dpath_mulcore_ary1_a1_I1_I1_6__net32));
OR2X1 mul_U1188(.A(n6988), .B(dpath_mulcore_b11[0]), .Y(n13052));
AND2X1 mul_U1189(.A(n909), .B(n13049), .Y(dpath_mulcore_ary1_a1_I1_I1_6__net046));
OR2X1 mul_U1190(.A(n6987), .B(dpath_mulcore_b12[0]), .Y(n13049));
AND2X1 mul_U1191(.A(n1081), .B(n13571), .Y(dpath_mulcore_ary1_a1_I0_I1_12__net32));
OR2X1 mul_U1192(.A(n7162), .B(dpath_mulcore_b8[0]), .Y(n13571));
AND2X1 mul_U1193(.A(n1080), .B(n13568), .Y(dpath_mulcore_ary1_a1_I0_I1_12__net046));
OR2X1 mul_U1194(.A(n7161), .B(dpath_mulcore_b9[0]), .Y(n13568));
AND2X1 mul_U1195(.A(n913), .B(n13061), .Y(dpath_mulcore_ary1_a1_I1_I1_5__net32));
OR2X1 mul_U1196(.A(n6991), .B(dpath_mulcore_b11[0]), .Y(n13061));
AND2X1 mul_U1197(.A(n912), .B(n13058), .Y(dpath_mulcore_ary1_a1_I1_I1_5__net046));
OR2X1 mul_U1198(.A(n6990), .B(dpath_mulcore_b12[0]), .Y(n13058));
OR2X1 mul_U1199(.A(n9751), .B(n5937), .Y(dpath_mulcore_ary1_a1_I2_I0_b1n_1));
OR2X1 mul_U1200(.A(n9751), .B(n5936), .Y(dpath_mulcore_ary1_a1_I2_I0_b1n_0));
AND2X1 mul_U1201(.A(n905), .B(n13037), .Y(dpath_mulcore_ary1_a1_I1_I1_7__net043));
OR2X1 mul_U1202(.A(n6983), .B(dpath_mulcore_b13[0]), .Y(n13037));
AND2X1 mul_U1203(.A(n730), .B(n12508), .Y(dpath_mulcore_ary1_a1_I2_I0_p0_1));
OR2X1 mul_U1204(.A(n6806), .B(dpath_mulcore_b14[0]), .Y(n12508));
OR2X1 mul_U1205(.A(n13712), .B(n5939), .Y(dpath_mulcore_ary1_a1_I2_I0_b0n));
AND2X1 mul_U1206(.A(n7404), .B(n9839), .Y(n13712));
AND2X1 mul_U1207(.A(n908), .B(n13046), .Y(dpath_mulcore_ary1_a1_I1_I1_6__net043));
OR2X1 mul_U1208(.A(n6986), .B(dpath_mulcore_b13[0]), .Y(n13046));
INVX1 mul_U1209(.A(n12510), .Y(n9839));
OR2X1 mul_U1210(.A(n6807), .B(dpath_mulcore_b14[0]), .Y(n12510));
OR2X1 mul_U1211(.A(n9749), .B(n5938), .Y(dpath_mulcore_ary1_a1_I2_I0_b0n_0));
AND2X1 mul_U1212(.A(n1084), .B(n13580), .Y(dpath_mulcore_ary1_a1_I0_I1_11__net32));
OR2X1 mul_U1213(.A(n7165), .B(dpath_mulcore_b8[0]), .Y(n13580));
AND2X1 mul_U1214(.A(n1083), .B(n13577), .Y(dpath_mulcore_ary1_a1_I0_I1_11__net046));
OR2X1 mul_U1215(.A(n7164), .B(dpath_mulcore_b9[0]), .Y(n13577));
AND2X1 mul_U1216(.A(n911), .B(n13055), .Y(dpath_mulcore_ary1_a1_I1_I1_5__net043));
OR2X1 mul_U1217(.A(n6989), .B(dpath_mulcore_b13[0]), .Y(n13055));
AND2X1 mul_U1218(.A(n915), .B(n13069), .Y(dpath_mulcore_ary1_a1_I1_I1_4__net32));
OR2X1 mul_U1219(.A(n6994), .B(dpath_mulcore_b11[0]), .Y(n13069));
AND2X1 mul_U1220(.A(n914), .B(n13066), .Y(dpath_mulcore_ary1_a1_I1_I1_4__net046));
OR2X1 mul_U1221(.A(n6993), .B(dpath_mulcore_b12[0]), .Y(n13066));
AND2X1 mul_U1222(.A(n1087), .B(n13589), .Y(dpath_mulcore_ary1_a1_I0_I1_10__net32));
OR2X1 mul_U1223(.A(n7168), .B(dpath_mulcore_b8[0]), .Y(n13589));
AND2X1 mul_U1224(.A(n1086), .B(n13586), .Y(dpath_mulcore_ary1_a1_I0_I1_10__net046));
OR2X1 mul_U1225(.A(n7167), .B(dpath_mulcore_b9[0]), .Y(n13586));
AND2X1 mul_U1226(.A(n1090), .B(n13598), .Y(dpath_mulcore_ary1_a1_I0_I1_9__net32));
OR2X1 mul_U1227(.A(n7171), .B(dpath_mulcore_b8[0]), .Y(n13598));
AND2X1 mul_U1228(.A(n1089), .B(n13595), .Y(dpath_mulcore_ary1_a1_I0_I1_9__net046));
OR2X1 mul_U1229(.A(n7170), .B(dpath_mulcore_b9[0]), .Y(n13595));
AND2X1 mul_U1230(.A(n1088), .B(n13592), .Y(dpath_mulcore_ary1_a1_I0_I1_9__net043));
OR2X1 mul_U1231(.A(n7169), .B(dpath_mulcore_b10[0]), .Y(n13592));
AND2X1 mul_U1232(.A(n1091), .B(n13601), .Y(dpath_mulcore_ary1_a1_I0_I1_8__net043));
OR2X1 mul_U1233(.A(n7172), .B(dpath_mulcore_b10[0]), .Y(n13601));
AND2X1 mul_U1234(.A(n1096), .B(n13616), .Y(dpath_mulcore_ary1_a1_I0_I1_7__net32));
OR2X1 mul_U1235(.A(n7177), .B(dpath_mulcore_b8[0]), .Y(n13616));
AND2X1 mul_U1236(.A(n1095), .B(n13613), .Y(dpath_mulcore_ary1_a1_I0_I1_7__net046));
OR2X1 mul_U1237(.A(n7176), .B(dpath_mulcore_b9[0]), .Y(n13613));
AND2X1 mul_U1238(.A(n1099), .B(n13625), .Y(dpath_mulcore_ary1_a1_I0_I1_6__net32));
OR2X1 mul_U1239(.A(n7180), .B(dpath_mulcore_b8[0]), .Y(n13625));
AND2X1 mul_U1240(.A(n1098), .B(n13622), .Y(dpath_mulcore_ary1_a1_I0_I1_6__net046));
OR2X1 mul_U1241(.A(n7179), .B(dpath_mulcore_b9[0]), .Y(n13622));
AND2X1 mul_U1242(.A(n1102), .B(n13634), .Y(dpath_mulcore_ary1_a1_I0_I1_5__net32));
OR2X1 mul_U1243(.A(n7183), .B(dpath_mulcore_b8[0]), .Y(n13634));
AND2X1 mul_U1244(.A(n1101), .B(n13631), .Y(dpath_mulcore_ary1_a1_I0_I1_5__net046));
OR2X1 mul_U1245(.A(n7182), .B(dpath_mulcore_b9[0]), .Y(n13631));
AND2X1 mul_U1246(.A(n1104), .B(n13642), .Y(dpath_mulcore_ary1_a1_I0_I1_4__net32));
OR2X1 mul_U1247(.A(n7186), .B(dpath_mulcore_b8[0]), .Y(n13642));
AND2X1 mul_U1248(.A(n1103), .B(n13639), .Y(dpath_mulcore_ary1_a1_I0_I1_4__net046));
OR2X1 mul_U1249(.A(n7185), .B(dpath_mulcore_b9[0]), .Y(n13639));
OR2X1 mul_U1250(.A(n5904), .B(n6032), .Y(dpath_areg[30]));
AND2X1 mul_U1251(.A(n2961), .B(n4637), .Y(dpath_n837));
AND2X1 mul_U1252(.A(n2882), .B(n4558), .Y(dpath_areg[95]));
AND2X1 mul_U1253(.A(n2883), .B(n4559), .Y(dpath_areg[94]));
AND2X1 mul_U1254(.A(n2884), .B(n4560), .Y(dpath_areg[93]));
AND2X1 mul_U1255(.A(n2885), .B(n4561), .Y(dpath_areg[92]));
AND2X1 mul_U1256(.A(n2886), .B(n4562), .Y(dpath_areg[91]));
AND2X1 mul_U1257(.A(n2887), .B(n4563), .Y(dpath_areg[90]));
AND2X1 mul_U1258(.A(n2890), .B(n4566), .Y(dpath_areg[89]));
AND2X1 mul_U1259(.A(n2891), .B(n4567), .Y(dpath_areg[88]));
AND2X1 mul_U1260(.A(n2892), .B(n4568), .Y(dpath_areg[87]));
AND2X1 mul_U1261(.A(n2893), .B(n4569), .Y(dpath_areg[86]));
AND2X1 mul_U1262(.A(n2894), .B(n4570), .Y(dpath_areg[85]));
AND2X1 mul_U1263(.A(n2895), .B(n4571), .Y(dpath_areg[84]));
AND2X1 mul_U1264(.A(n2896), .B(n4572), .Y(dpath_areg[83]));
AND2X1 mul_U1265(.A(n2897), .B(n4573), .Y(dpath_areg[82]));
AND2X1 mul_U1266(.A(n1899), .B(n3952), .Y(dpath_mulcore_array2_c1[79]));
AND2X1 mul_U1267(.A(n2898), .B(n4574), .Y(dpath_areg[81]));
AND2X1 mul_U1268(.A(n1900), .B(n3953), .Y(dpath_mulcore_array2_c1[78]));
AND2X1 mul_U1269(.A(n2899), .B(n4575), .Y(dpath_areg[80]));
AND2X1 mul_U1270(.A(n1901), .B(n3954), .Y(dpath_mulcore_array2_c1[77]));
AND2X1 mul_U1271(.A(n2902), .B(n4578), .Y(dpath_areg[79]));
AND2X1 mul_U1272(.A(n1902), .B(n3955), .Y(dpath_mulcore_array2_c1[76]));
AND2X1 mul_U1273(.A(n2903), .B(n4579), .Y(dpath_areg[78]));
AND2X1 mul_U1274(.A(n1903), .B(n3956), .Y(dpath_mulcore_array2_c1[75]));
AND2X1 mul_U1275(.A(n2904), .B(n4580), .Y(dpath_areg[77]));
AND2X1 mul_U1276(.A(n1904), .B(n3957), .Y(dpath_mulcore_array2_c1[74]));
AND2X1 mul_U1277(.A(n2905), .B(n4581), .Y(dpath_areg[76]));
AND2X1 mul_U1278(.A(n1905), .B(n3958), .Y(dpath_mulcore_array2_c1[73]));
AND2X1 mul_U1279(.A(n2906), .B(n4582), .Y(dpath_areg[75]));
AND2X1 mul_U1280(.A(n1906), .B(n3959), .Y(dpath_mulcore_array2_c1[72]));
AND2X1 mul_U1281(.A(n2907), .B(n4583), .Y(dpath_areg[74]));
AND2X1 mul_U1282(.A(n1907), .B(n3960), .Y(dpath_mulcore_array2_c1[71]));
AND2X1 mul_U1283(.A(n2908), .B(n4584), .Y(dpath_areg[73]));
AND2X1 mul_U1284(.A(n1908), .B(n3961), .Y(dpath_mulcore_array2_c1[70]));
AND2X1 mul_U1285(.A(n2909), .B(n4585), .Y(dpath_areg[72]));
AND2X1 mul_U1286(.A(n1909), .B(n3962), .Y(dpath_mulcore_array2_c1[69]));
AND2X1 mul_U1287(.A(n2910), .B(n4586), .Y(dpath_areg[71]));
AND2X1 mul_U1288(.A(n1910), .B(n3963), .Y(dpath_mulcore_array2_c1[68]));
AND2X1 mul_U1289(.A(n2911), .B(n4587), .Y(dpath_areg[70]));
AND2X1 mul_U1290(.A(n2914), .B(n4590), .Y(dpath_areg[69]));
AND2X1 mul_U1291(.A(n1952), .B(n4005), .Y(dpath_mulcore_array2_c2[66]));
OR2X1 mul_U1292(.A(n9429), .B(dpath_mulcore_array2_s1[66]), .Y(n17477));
AND2X1 mul_U1293(.A(n2915), .B(n4591), .Y(dpath_areg[68]));
AND2X1 mul_U1294(.A(n1953), .B(n4006), .Y(dpath_mulcore_array2_c2[65]));
AND2X1 mul_U1295(.A(n1999), .B(n4052), .Y(dpath_mulcore_array2_c1[65]));
OR2X1 mul_U1296(.A(n9430), .B(dpath_mulcore_array2_s1[65]), .Y(n17484));
AND2X1 mul_U1297(.A(n2916), .B(n4592), .Y(dpath_areg[67]));
AND2X1 mul_U1298(.A(n1954), .B(n4007), .Y(dpath_mulcore_array2_c2[64]));
AND2X1 mul_U1299(.A(n2000), .B(n4053), .Y(dpath_mulcore_array2_c1[64]));
OR2X1 mul_U1300(.A(n9431), .B(dpath_mulcore_array2_s1[64]), .Y(n17491));
AND2X1 mul_U1301(.A(n2917), .B(n4593), .Y(dpath_areg[66]));
AND2X1 mul_U1302(.A(n1955), .B(n4008), .Y(dpath_mulcore_array2_c2[63]));
AND2X1 mul_U1303(.A(n2001), .B(n4054), .Y(dpath_mulcore_array2_c1[63]));
OR2X1 mul_U1304(.A(n9432), .B(dpath_mulcore_array2_s1[63]), .Y(n17498));
AND2X1 mul_U1305(.A(n2918), .B(n4594), .Y(dpath_areg[65]));
AND2X1 mul_U1306(.A(n1956), .B(n4009), .Y(dpath_mulcore_array2_c2[62]));
AND2X1 mul_U1307(.A(n2002), .B(n4055), .Y(dpath_mulcore_array2_c1[62]));
OR2X1 mul_U1308(.A(n9433), .B(dpath_mulcore_array2_s1[62]), .Y(n17505));
AND2X1 mul_U1309(.A(n2919), .B(n4595), .Y(dpath_areg[64]));
AND2X1 mul_U1310(.A(n1957), .B(n4010), .Y(dpath_mulcore_array2_c2[61]));
AND2X1 mul_U1311(.A(n2003), .B(n4056), .Y(dpath_mulcore_array2_c1[61]));
OR2X1 mul_U1312(.A(n9434), .B(dpath_mulcore_array2_s1[61]), .Y(n17512));
AND2X1 mul_U1313(.A(n2920), .B(n4596), .Y(dpath_areg[63]));
AND2X1 mul_U1314(.A(n1958), .B(n4011), .Y(dpath_mulcore_array2_c2[60]));
AND2X1 mul_U1315(.A(n2004), .B(n4057), .Y(dpath_mulcore_array2_c1[60]));
OR2X1 mul_U1316(.A(n9435), .B(dpath_mulcore_array2_s1[60]), .Y(n17519));
AND2X1 mul_U1317(.A(n2921), .B(n4597), .Y(dpath_areg[62]));
AND2X1 mul_U1318(.A(n1959), .B(n4012), .Y(dpath_mulcore_array2_c2[59]));
AND2X1 mul_U1319(.A(n2005), .B(n4058), .Y(dpath_mulcore_array2_c1[59]));
OR2X1 mul_U1320(.A(n9436), .B(dpath_mulcore_array2_s1[59]), .Y(n17526));
AND2X1 mul_U1321(.A(n2922), .B(n4598), .Y(dpath_areg[61]));
AND2X1 mul_U1322(.A(n1960), .B(n4013), .Y(dpath_mulcore_array2_c2[58]));
AND2X1 mul_U1323(.A(n2006), .B(n4059), .Y(dpath_mulcore_array2_c1[58]));
OR2X1 mul_U1324(.A(n9437), .B(dpath_mulcore_array2_s1[58]), .Y(n17533));
AND2X1 mul_U1325(.A(n2923), .B(n4599), .Y(dpath_areg[60]));
AND2X1 mul_U1326(.A(n1961), .B(n4014), .Y(dpath_mulcore_array2_c2[57]));
AND2X1 mul_U1327(.A(n2007), .B(n4060), .Y(dpath_mulcore_array2_c1[57]));
OR2X1 mul_U1328(.A(n9438), .B(dpath_mulcore_array2_s1[57]), .Y(n17540));
AND2X1 mul_U1329(.A(n2926), .B(n4602), .Y(dpath_areg[59]));
AND2X1 mul_U1330(.A(n1962), .B(n4015), .Y(dpath_mulcore_array2_c2[56]));
AND2X1 mul_U1331(.A(n2008), .B(n4061), .Y(dpath_mulcore_array2_c1[56]));
OR2X1 mul_U1332(.A(n9439), .B(dpath_mulcore_array2_s1[56]), .Y(n17547));
AND2X1 mul_U1333(.A(n2927), .B(n4603), .Y(dpath_areg[58]));
AND2X1 mul_U1334(.A(n1963), .B(n4016), .Y(dpath_mulcore_array2_c2[55]));
AND2X1 mul_U1335(.A(n2009), .B(n4062), .Y(dpath_mulcore_array2_c1[55]));
OR2X1 mul_U1336(.A(n9440), .B(dpath_mulcore_array2_s1[55]), .Y(n17554));
AND2X1 mul_U1337(.A(n2928), .B(n4604), .Y(dpath_areg[57]));
AND2X1 mul_U1338(.A(n1964), .B(n4017), .Y(dpath_mulcore_array2_c2[54]));
AND2X1 mul_U1339(.A(n2010), .B(n4063), .Y(dpath_mulcore_array2_c1[54]));
OR2X1 mul_U1340(.A(n9441), .B(dpath_mulcore_array2_s1[54]), .Y(n17561));
AND2X1 mul_U1341(.A(n2929), .B(n4605), .Y(dpath_areg[56]));
AND2X1 mul_U1342(.A(n1965), .B(n4018), .Y(dpath_mulcore_array2_c2[53]));
AND2X1 mul_U1343(.A(n2011), .B(n4064), .Y(dpath_mulcore_array2_c1[53]));
OR2X1 mul_U1344(.A(n9442), .B(dpath_mulcore_array2_s1[53]), .Y(n17568));
AND2X1 mul_U1345(.A(n2930), .B(n4606), .Y(dpath_areg[55]));
AND2X1 mul_U1346(.A(n1966), .B(n4019), .Y(dpath_mulcore_array2_c2[52]));
AND2X1 mul_U1347(.A(n2012), .B(n4065), .Y(dpath_mulcore_array2_c1[52]));
OR2X1 mul_U1348(.A(n9443), .B(dpath_mulcore_array2_s1[52]), .Y(n17575));
AND2X1 mul_U1349(.A(n2931), .B(n4607), .Y(dpath_areg[54]));
AND2X1 mul_U1350(.A(n1967), .B(n4020), .Y(dpath_mulcore_array2_c2[51]));
AND2X1 mul_U1351(.A(n2013), .B(n4066), .Y(dpath_mulcore_array2_c1[51]));
OR2X1 mul_U1352(.A(n9444), .B(dpath_mulcore_array2_s1[51]), .Y(n17582));
AND2X1 mul_U1353(.A(n2932), .B(n4608), .Y(dpath_areg[53]));
AND2X1 mul_U1354(.A(n1968), .B(n4021), .Y(dpath_mulcore_array2_c2[50]));
AND2X1 mul_U1355(.A(n2014), .B(n4067), .Y(dpath_mulcore_array2_c1[50]));
OR2X1 mul_U1356(.A(n9445), .B(dpath_mulcore_array2_s1[50]), .Y(n17589));
AND2X1 mul_U1357(.A(n2933), .B(n4609), .Y(dpath_areg[52]));
AND2X1 mul_U1358(.A(n1969), .B(n4022), .Y(dpath_mulcore_array2_c2[49]));
AND2X1 mul_U1359(.A(n2015), .B(n4068), .Y(dpath_mulcore_array2_c1[49]));
OR2X1 mul_U1360(.A(n9446), .B(dpath_mulcore_array2_s1[49]), .Y(n17596));
AND2X1 mul_U1361(.A(n2934), .B(n4610), .Y(dpath_areg[51]));
AND2X1 mul_U1362(.A(n1970), .B(n4023), .Y(dpath_mulcore_array2_c2[48]));
AND2X1 mul_U1363(.A(n2016), .B(n4069), .Y(dpath_mulcore_array2_c1[48]));
OR2X1 mul_U1364(.A(n9447), .B(dpath_mulcore_array2_s1[48]), .Y(n17603));
AND2X1 mul_U1365(.A(n2935), .B(n4611), .Y(dpath_areg[50]));
AND2X1 mul_U1366(.A(n1971), .B(n4024), .Y(dpath_mulcore_array2_c2[47]));
AND2X1 mul_U1367(.A(n2017), .B(n4070), .Y(dpath_mulcore_array2_c1[47]));
OR2X1 mul_U1368(.A(n9448), .B(dpath_mulcore_array2_s1[47]), .Y(n17610));
AND2X1 mul_U1369(.A(n2938), .B(n4614), .Y(dpath_areg[49]));
AND2X1 mul_U1370(.A(n1972), .B(n4025), .Y(dpath_mulcore_array2_c2[46]));
AND2X1 mul_U1371(.A(n2018), .B(n4071), .Y(dpath_mulcore_array2_c1[46]));
OR2X1 mul_U1372(.A(n9449), .B(dpath_mulcore_array2_s1[46]), .Y(n17617));
AND2X1 mul_U1373(.A(n2939), .B(n4615), .Y(dpath_areg[48]));
AND2X1 mul_U1374(.A(n1973), .B(n4026), .Y(dpath_mulcore_array2_c2[45]));
AND2X1 mul_U1375(.A(n2019), .B(n4072), .Y(dpath_mulcore_array2_c1[45]));
OR2X1 mul_U1376(.A(n9450), .B(dpath_mulcore_array2_s1[45]), .Y(n17624));
AND2X1 mul_U1377(.A(n2940), .B(n4616), .Y(dpath_areg[47]));
AND2X1 mul_U1378(.A(n1974), .B(n4027), .Y(dpath_mulcore_array2_c2[44]));
AND2X1 mul_U1379(.A(n2020), .B(n4073), .Y(dpath_mulcore_array2_c1[44]));
OR2X1 mul_U1380(.A(n9451), .B(dpath_mulcore_array2_s1[44]), .Y(n17631));
AND2X1 mul_U1381(.A(n2941), .B(n4617), .Y(dpath_areg[46]));
AND2X1 mul_U1382(.A(n1975), .B(n4028), .Y(dpath_mulcore_array2_c2[43]));
AND2X1 mul_U1383(.A(n2021), .B(n4074), .Y(dpath_mulcore_array2_c1[43]));
OR2X1 mul_U1384(.A(n9452), .B(dpath_mulcore_array2_s1[43]), .Y(n17638));
AND2X1 mul_U1385(.A(n2942), .B(n4618), .Y(dpath_areg[45]));
AND2X1 mul_U1386(.A(n1976), .B(n4029), .Y(dpath_mulcore_array2_c2[42]));
AND2X1 mul_U1387(.A(n2022), .B(n4075), .Y(dpath_mulcore_array2_c1[42]));
OR2X1 mul_U1388(.A(n9453), .B(dpath_mulcore_array2_s1[42]), .Y(n17645));
AND2X1 mul_U1389(.A(n2943), .B(n4619), .Y(dpath_areg[44]));
AND2X1 mul_U1390(.A(n1977), .B(n4030), .Y(dpath_mulcore_array2_c2[41]));
AND2X1 mul_U1391(.A(n2023), .B(n4076), .Y(dpath_mulcore_array2_c1[41]));
OR2X1 mul_U1392(.A(n9454), .B(dpath_mulcore_array2_s1[41]), .Y(n17652));
AND2X1 mul_U1393(.A(n2944), .B(n4620), .Y(dpath_areg[43]));
AND2X1 mul_U1394(.A(n1978), .B(n4031), .Y(dpath_mulcore_array2_c2[40]));
AND2X1 mul_U1395(.A(n2024), .B(n4077), .Y(dpath_mulcore_array2_c1[40]));
OR2X1 mul_U1396(.A(n9455), .B(dpath_mulcore_array2_s1[40]), .Y(n17659));
AND2X1 mul_U1397(.A(n2945), .B(n4621), .Y(dpath_areg[42]));
AND2X1 mul_U1398(.A(n1979), .B(n4032), .Y(dpath_mulcore_array2_c2[39]));
AND2X1 mul_U1399(.A(n2025), .B(n4078), .Y(dpath_mulcore_array2_c1[39]));
OR2X1 mul_U1400(.A(n9456), .B(dpath_mulcore_array2_s1[39]), .Y(n17666));
INVX1 mul_U1401(.A(n9679), .Y(n9717));
AND2X1 mul_U1402(.A(n2946), .B(n4622), .Y(dpath_areg[41]));
AND2X1 mul_U1403(.A(n1980), .B(n4033), .Y(dpath_mulcore_array2_c2[38]));
AND2X1 mul_U1404(.A(n2026), .B(n4079), .Y(dpath_mulcore_array2_c1[38]));
OR2X1 mul_U1405(.A(n9457), .B(dpath_mulcore_array2_s1[38]), .Y(n17673));
AND2X1 mul_U1406(.A(n2947), .B(n4623), .Y(dpath_areg[40]));
AND2X1 mul_U1407(.A(n1981), .B(n4034), .Y(dpath_mulcore_array2_c2[37]));
AND2X1 mul_U1408(.A(n2027), .B(n4080), .Y(dpath_mulcore_array2_c1[37]));
OR2X1 mul_U1409(.A(n9458), .B(dpath_mulcore_array2_s1[37]), .Y(n17680));
AND2X1 mul_U1410(.A(n2950), .B(n4626), .Y(dpath_areg[39]));
AND2X1 mul_U1411(.A(n1982), .B(n4035), .Y(dpath_mulcore_array2_c2[36]));
AND2X1 mul_U1412(.A(n2028), .B(n4081), .Y(dpath_mulcore_array2_c1[36]));
OR2X1 mul_U1413(.A(n9459), .B(dpath_mulcore_array2_s1[36]), .Y(n17687));
AND2X1 mul_U1414(.A(n2951), .B(n4627), .Y(dpath_areg[38]));
AND2X1 mul_U1415(.A(n1983), .B(n4036), .Y(dpath_mulcore_array2_c2[35]));
AND2X1 mul_U1416(.A(n2029), .B(n4082), .Y(dpath_mulcore_array2_c1[35]));
OR2X1 mul_U1417(.A(n9460), .B(dpath_mulcore_array2_s1[35]), .Y(n17694));
AND2X1 mul_U1418(.A(n2952), .B(n4628), .Y(dpath_areg[37]));
AND2X1 mul_U1419(.A(n1984), .B(n4037), .Y(dpath_mulcore_array2_c2[34]));
AND2X1 mul_U1420(.A(n2030), .B(n4083), .Y(dpath_mulcore_array2_c1[34]));
OR2X1 mul_U1421(.A(n9461), .B(dpath_mulcore_array2_s1[34]), .Y(n17701));
AND2X1 mul_U1422(.A(n2953), .B(n4629), .Y(dpath_areg[36]));
AND2X1 mul_U1423(.A(n1985), .B(n4038), .Y(dpath_mulcore_array2_c2[33]));
AND2X1 mul_U1424(.A(n2031), .B(n4084), .Y(dpath_mulcore_array2_c1[33]));
OR2X1 mul_U1425(.A(n9462), .B(dpath_mulcore_array2_s1[33]), .Y(n17708));
AND2X1 mul_U1426(.A(n2954), .B(n4630), .Y(dpath_areg[35]));
AND2X1 mul_U1427(.A(n1986), .B(n4039), .Y(dpath_mulcore_array2_c2[32]));
AND2X1 mul_U1428(.A(n2032), .B(n4085), .Y(dpath_mulcore_array2_c1[32]));
OR2X1 mul_U1429(.A(n9463), .B(dpath_mulcore_array2_s1[32]), .Y(n17715));
AND2X1 mul_U1430(.A(n2955), .B(n4631), .Y(dpath_areg[34]));
AND2X1 mul_U1431(.A(n1987), .B(n4040), .Y(dpath_mulcore_array2_c2[31]));
AND2X1 mul_U1432(.A(n2033), .B(n4086), .Y(dpath_mulcore_array2_c1[31]));
OR2X1 mul_U1433(.A(n9464), .B(dpath_mulcore_array2_s1[31]), .Y(n17722));
AND2X1 mul_U1434(.A(n2956), .B(n4632), .Y(dpath_areg[33]));
AND2X1 mul_U1435(.A(n1988), .B(n4041), .Y(dpath_mulcore_array2_c2[30]));
AND2X1 mul_U1436(.A(n2034), .B(n4087), .Y(dpath_mulcore_array2_c1[30]));
OR2X1 mul_U1437(.A(n9465), .B(dpath_mulcore_array2_s1[30]), .Y(n17729));
OR2X1 mul_U1438(.A(n5903), .B(n6031), .Y(dpath_areg[31]));
AND2X1 mul_U1439(.A(n2959), .B(n4635), .Y(dpath_n831));
INVX1 mul_U1440(.A(n9679), .Y(n9716));
AND2X1 mul_U1441(.A(n2957), .B(n4633), .Y(dpath_areg[32]));
AND2X1 mul_U1442(.A(n1989), .B(n4042), .Y(dpath_mulcore_array2_c2[29]));
AND2X1 mul_U1443(.A(n2035), .B(n4088), .Y(dpath_mulcore_array2_c1[29]));
OR2X1 mul_U1444(.A(n9466), .B(dpath_mulcore_array2_s1[29]), .Y(n17736));
AND2X1 mul_U1445(.A(n1888), .B(n3941), .Y(dpath_mulcore_array2_c1[18]));
AND2X1 mul_U1446(.A(n1889), .B(n3942), .Y(dpath_mulcore_array2_c1[17]));
AND2X1 mul_U1447(.A(n1890), .B(n3943), .Y(dpath_mulcore_array2_c1[16]));
AND2X1 mul_U1448(.A(n1929), .B(n3982), .Y(dpath_mulcore_array2_c1[12]));
AND2X1 mul_U1449(.A(n1930), .B(n3983), .Y(dpath_mulcore_array2_c1[11]));
AND2X1 mul_U1450(.A(n1931), .B(n3984), .Y(dpath_mulcore_array2_c1[10]));
AND2X1 mul_U1451(.A(n1932), .B(n3985), .Y(dpath_mulcore_array2_c1[9]));
AND2X1 mul_U1452(.A(n1933), .B(n3986), .Y(dpath_mulcore_array2_c1[8]));
AND2X1 mul_U1453(.A(n1934), .B(n3987), .Y(dpath_mulcore_array2_c1[7]));
AND2X1 mul_U1454(.A(n1935), .B(n3988), .Y(dpath_mulcore_array2_c1[6]));
AND2X1 mul_U1455(.A(n1936), .B(n3989), .Y(dpath_mulcore_array2_c1[5]));
AND2X1 mul_U1456(.A(n1948), .B(n4001), .Y(dpath_mulcore_array2_c1[4]));
AND2X1 mul_U1457(.A(n2395), .B(n4320), .Y(dpath_mulcore_array2_co[28]));
AND2X1 mul_U1458(.A(n2397), .B(n4322), .Y(dpath_mulcore_array2_co[27]));
AND2X1 mul_U1459(.A(n2399), .B(n4324), .Y(dpath_mulcore_array2_co[26]));
AND2X1 mul_U1460(.A(n2401), .B(n4326), .Y(dpath_mulcore_array2_co[25]));
AND2X1 mul_U1461(.A(n2403), .B(n4328), .Y(dpath_mulcore_array2_co[24]));
AND2X1 mul_U1462(.A(n2405), .B(n4330), .Y(dpath_mulcore_array2_co[23]));
AND2X1 mul_U1463(.A(n2407), .B(n4332), .Y(dpath_mulcore_array2_co[22]));
AND2X1 mul_U1464(.A(n2409), .B(n4334), .Y(dpath_mulcore_array2_co[21]));
AND2X1 mul_U1465(.A(n2411), .B(n4336), .Y(dpath_mulcore_array2_co[20]));
AND2X1 mul_U1466(.A(n1893), .B(n3946), .Y(dpath_mulcore_array2_c2[19]));
AND2X1 mul_U1467(.A(n1887), .B(n3940), .Y(dpath_mulcore_array2_c1[19]));
AND2X1 mul_U1468(.A(n1894), .B(n3947), .Y(dpath_mulcore_array2_c2[18]));
AND2X1 mul_U1469(.A(n1895), .B(n3948), .Y(dpath_mulcore_array2_c2[17]));
AND2X1 mul_U1470(.A(n1896), .B(n3949), .Y(dpath_mulcore_array2_c2[16]));
AND2X1 mul_U1471(.A(n1897), .B(n3950), .Y(dpath_mulcore_array2_c2[15]));
AND2X1 mul_U1472(.A(n1927), .B(n3980), .Y(dpath_mulcore_array2_c1[14]));
OR2X1 mul_U1473(.A(n5921), .B(n6049), .Y(dpath_areg[15]));
AND2X1 mul_U1474(.A(n2995), .B(n4671), .Y(dpath_n939));
INVX1 mul_U1475(.A(n9678), .Y(n9714));
OR2X1 mul_U1476(.A(n5920), .B(n6048), .Y(dpath_areg[16]));
AND2X1 mul_U1477(.A(n2993), .B(n4669), .Y(dpath_n933));
INVX1 mul_U1478(.A(n9678), .Y(n9715));
OR2X1 mul_U1479(.A(n5916), .B(n6044), .Y(dpath_areg[1]));
AND2X1 mul_U1480(.A(n2985), .B(n4661), .Y(dpath_n909));
AND2X1 mul_U1481(.A(n235), .B(n11011), .Y(dpath_mulcore_ary1_a0_I1_I1_63__net32));
OR2X1 mul_U1482(.A(n6305), .B(dpath_mulcore_b3[0]), .Y(n11011));
AND2X1 mul_U1483(.A(n234), .B(n11008), .Y(dpath_mulcore_ary1_a0_I1_I1_63__net046));
OR2X1 mul_U1484(.A(n6304), .B(dpath_mulcore_b4[0]), .Y(n11008));
AND2X1 mul_U1485(.A(n238), .B(n11020), .Y(dpath_mulcore_ary1_a0_I1_I1_62__net32));
OR2X1 mul_U1486(.A(n6308), .B(dpath_mulcore_b3[0]), .Y(n11020));
AND2X1 mul_U1487(.A(n237), .B(n11017), .Y(dpath_mulcore_ary1_a0_I1_I1_62__net046));
OR2X1 mul_U1488(.A(n6307), .B(dpath_mulcore_b4[0]), .Y(n11017));
AND2X1 mul_U1489(.A(n416), .B(n11560), .Y(dpath_mulcore_ary1_a0_I0_I2_net078));
OR2X1 mul_U1490(.A(n6489), .B(dpath_mulcore_b2[0]), .Y(n11560));
AND2X1 mul_U1491(.A(n241), .B(n11029), .Y(dpath_mulcore_ary1_a0_I1_I1_61__net32));
OR2X1 mul_U1492(.A(n6311), .B(dpath_mulcore_b3[0]), .Y(n11029));
AND2X1 mul_U1493(.A(n240), .B(n11026), .Y(dpath_mulcore_ary1_a0_I1_I1_61__net046));
OR2X1 mul_U1494(.A(n6310), .B(dpath_mulcore_b4[0]), .Y(n11026));
AND2X1 mul_U1495(.A(n417), .B(n11563), .Y(dpath_mulcore_ary1_a0_I0_I2_net8));
OR2X1 mul_U1496(.A(n6490), .B(dpath_mulcore_b2[0]), .Y(n11563));
AND2X1 mul_U1497(.A(n244), .B(n11038), .Y(dpath_mulcore_ary1_a0_I1_I1_60__net32));
OR2X1 mul_U1498(.A(n6314), .B(dpath_mulcore_b3[0]), .Y(n11038));
AND2X1 mul_U1499(.A(n243), .B(n11035), .Y(dpath_mulcore_ary1_a0_I1_I1_60__net046));
OR2X1 mul_U1500(.A(n6313), .B(dpath_mulcore_b4[0]), .Y(n11035));
AND2X1 mul_U1501(.A(n418), .B(n11566), .Y(dpath_mulcore_ary1_a0_I0_I2_net15));
OR2X1 mul_U1502(.A(n6491), .B(dpath_mulcore_b2[0]), .Y(n11566));
AND2X1 mul_U1503(.A(n247), .B(n11047), .Y(dpath_mulcore_ary1_a0_I1_I1_59__net32));
OR2X1 mul_U1504(.A(n6317), .B(dpath_mulcore_b3[0]), .Y(n11047));
AND2X1 mul_U1505(.A(n246), .B(n11044), .Y(dpath_mulcore_ary1_a0_I1_I1_59__net046));
OR2X1 mul_U1506(.A(n6316), .B(dpath_mulcore_b4[0]), .Y(n11044));
AND2X1 mul_U1507(.A(n421), .B(n11575), .Y(dpath_mulcore_ary1_a0_I0_I2_net35));
OR2X1 mul_U1508(.A(n6494), .B(dpath_mulcore_b2[0]), .Y(n11575));
AND2X1 mul_U1509(.A(n250), .B(n11056), .Y(dpath_mulcore_ary1_a0_I1_I1_58__net32));
OR2X1 mul_U1510(.A(n6320), .B(dpath_mulcore_b3[0]), .Y(n11056));
AND2X1 mul_U1511(.A(n249), .B(n11053), .Y(dpath_mulcore_ary1_a0_I1_I1_58__net046));
OR2X1 mul_U1512(.A(n6319), .B(dpath_mulcore_b4[0]), .Y(n11053));
AND2X1 mul_U1513(.A(n422), .B(n11578), .Y(dpath_mulcore_ary1_a0_I0_I1_63__net043));
OR2X1 mul_U1514(.A(n6495), .B(dpath_mulcore_b2[0]), .Y(n11578));
AND2X1 mul_U1515(.A(n253), .B(n11065), .Y(dpath_mulcore_ary1_a0_I1_I1_57__net32));
OR2X1 mul_U1516(.A(n6323), .B(dpath_mulcore_b3[0]), .Y(n11065));
AND2X1 mul_U1517(.A(n252), .B(n11062), .Y(dpath_mulcore_ary1_a0_I1_I1_57__net046));
OR2X1 mul_U1518(.A(n6322), .B(dpath_mulcore_b4[0]), .Y(n11062));
AND2X1 mul_U1519(.A(n425), .B(n11587), .Y(dpath_mulcore_ary1_a0_I0_I1_62__net043));
OR2X1 mul_U1520(.A(n6498), .B(dpath_mulcore_b2[0]), .Y(n11587));
AND2X1 mul_U1521(.A(n256), .B(n11074), .Y(dpath_mulcore_ary1_a0_I1_I1_56__net32));
OR2X1 mul_U1522(.A(n6326), .B(dpath_mulcore_b3[0]), .Y(n11074));
AND2X1 mul_U1523(.A(n255), .B(n11071), .Y(dpath_mulcore_ary1_a0_I1_I1_56__net046));
OR2X1 mul_U1524(.A(n6325), .B(dpath_mulcore_b4[0]), .Y(n11071));
AND2X1 mul_U1525(.A(n428), .B(n11596), .Y(dpath_mulcore_ary1_a0_I0_I1_61__net043));
OR2X1 mul_U1526(.A(n6501), .B(dpath_mulcore_b2[0]), .Y(n11596));
AND2X1 mul_U1527(.A(n259), .B(n11083), .Y(dpath_mulcore_ary1_a0_I1_I1_55__net32));
OR2X1 mul_U1528(.A(n6329), .B(dpath_mulcore_b3[0]), .Y(n11083));
AND2X1 mul_U1529(.A(n258), .B(n11080), .Y(dpath_mulcore_ary1_a0_I1_I1_55__net046));
OR2X1 mul_U1530(.A(n6328), .B(dpath_mulcore_b4[0]), .Y(n11080));
AND2X1 mul_U1531(.A(n431), .B(n11605), .Y(dpath_mulcore_ary1_a0_I0_I1_60__net043));
OR2X1 mul_U1532(.A(n6504), .B(dpath_mulcore_b2[0]), .Y(n11605));
AND2X1 mul_U1533(.A(n262), .B(n11092), .Y(dpath_mulcore_ary1_a0_I1_I1_54__net32));
OR2X1 mul_U1534(.A(n6332), .B(dpath_mulcore_b3[0]), .Y(n11092));
AND2X1 mul_U1535(.A(n261), .B(n11089), .Y(dpath_mulcore_ary1_a0_I1_I1_54__net046));
OR2X1 mul_U1536(.A(n6331), .B(dpath_mulcore_b4[0]), .Y(n11089));
AND2X1 mul_U1537(.A(n434), .B(n11614), .Y(dpath_mulcore_ary1_a0_I0_I1_59__net043));
OR2X1 mul_U1538(.A(n6507), .B(dpath_mulcore_b2[0]), .Y(n11614));
AND2X1 mul_U1539(.A(n265), .B(n11101), .Y(dpath_mulcore_ary1_a0_I1_I1_53__net32));
OR2X1 mul_U1540(.A(n6335), .B(dpath_mulcore_b3[0]), .Y(n11101));
AND2X1 mul_U1541(.A(n264), .B(n11098), .Y(dpath_mulcore_ary1_a0_I1_I1_53__net046));
OR2X1 mul_U1542(.A(n6334), .B(dpath_mulcore_b4[0]), .Y(n11098));
AND2X1 mul_U1543(.A(n437), .B(n11623), .Y(dpath_mulcore_ary1_a0_I0_I1_58__net043));
OR2X1 mul_U1544(.A(n6510), .B(dpath_mulcore_b2[0]), .Y(n11623));
AND2X1 mul_U1545(.A(n268), .B(n11110), .Y(dpath_mulcore_ary1_a0_I1_I1_52__net32));
OR2X1 mul_U1546(.A(n6338), .B(dpath_mulcore_b3[0]), .Y(n11110));
AND2X1 mul_U1547(.A(n267), .B(n11107), .Y(dpath_mulcore_ary1_a0_I1_I1_52__net046));
OR2X1 mul_U1548(.A(n6337), .B(dpath_mulcore_b4[0]), .Y(n11107));
AND2X1 mul_U1549(.A(n440), .B(n11632), .Y(dpath_mulcore_ary1_a0_I0_I1_57__net043));
OR2X1 mul_U1550(.A(n6513), .B(dpath_mulcore_b2[0]), .Y(n11632));
AND2X1 mul_U1551(.A(n271), .B(n11119), .Y(dpath_mulcore_ary1_a0_I1_I1_51__net32));
OR2X1 mul_U1552(.A(n6341), .B(dpath_mulcore_b3[0]), .Y(n11119));
AND2X1 mul_U1553(.A(n270), .B(n11116), .Y(dpath_mulcore_ary1_a0_I1_I1_51__net046));
OR2X1 mul_U1554(.A(n6340), .B(dpath_mulcore_b4[0]), .Y(n11116));
AND2X1 mul_U1555(.A(n443), .B(n11641), .Y(dpath_mulcore_ary1_a0_I0_I1_56__net043));
OR2X1 mul_U1556(.A(n6516), .B(dpath_mulcore_b2[0]), .Y(n11641));
AND2X1 mul_U1557(.A(n274), .B(n11128), .Y(dpath_mulcore_ary1_a0_I1_I1_50__net32));
OR2X1 mul_U1558(.A(n6344), .B(dpath_mulcore_b3[0]), .Y(n11128));
AND2X1 mul_U1559(.A(n273), .B(n11125), .Y(dpath_mulcore_ary1_a0_I1_I1_50__net046));
OR2X1 mul_U1560(.A(n6343), .B(dpath_mulcore_b4[0]), .Y(n11125));
AND2X1 mul_U1561(.A(n446), .B(n11650), .Y(dpath_mulcore_ary1_a0_I0_I1_55__net043));
OR2X1 mul_U1562(.A(n6519), .B(dpath_mulcore_b2[0]), .Y(n11650));
AND2X1 mul_U1563(.A(n277), .B(n11137), .Y(dpath_mulcore_ary1_a0_I1_I1_49__net32));
OR2X1 mul_U1564(.A(n6347), .B(dpath_mulcore_b3[0]), .Y(n11137));
AND2X1 mul_U1565(.A(n276), .B(n11134), .Y(dpath_mulcore_ary1_a0_I1_I1_49__net046));
OR2X1 mul_U1566(.A(n6346), .B(dpath_mulcore_b4[0]), .Y(n11134));
AND2X1 mul_U1567(.A(n449), .B(n11659), .Y(dpath_mulcore_ary1_a0_I0_I1_54__net043));
OR2X1 mul_U1568(.A(n6522), .B(dpath_mulcore_b2[0]), .Y(n11659));
AND2X1 mul_U1569(.A(n280), .B(n11146), .Y(dpath_mulcore_ary1_a0_I1_I1_48__net32));
OR2X1 mul_U1570(.A(n6350), .B(dpath_mulcore_b3[0]), .Y(n11146));
AND2X1 mul_U1571(.A(n279), .B(n11143), .Y(dpath_mulcore_ary1_a0_I1_I1_48__net046));
OR2X1 mul_U1572(.A(n6349), .B(dpath_mulcore_b4[0]), .Y(n11143));
AND2X1 mul_U1573(.A(n452), .B(n11668), .Y(dpath_mulcore_ary1_a0_I0_I1_53__net043));
OR2X1 mul_U1574(.A(n6525), .B(dpath_mulcore_b2[0]), .Y(n11668));
AND2X1 mul_U1575(.A(n283), .B(n11155), .Y(dpath_mulcore_ary1_a0_I1_I1_47__net32));
OR2X1 mul_U1576(.A(n6353), .B(dpath_mulcore_b3[0]), .Y(n11155));
AND2X1 mul_U1577(.A(n282), .B(n11152), .Y(dpath_mulcore_ary1_a0_I1_I1_47__net046));
OR2X1 mul_U1578(.A(n6352), .B(dpath_mulcore_b4[0]), .Y(n11152));
AND2X1 mul_U1579(.A(n455), .B(n11677), .Y(dpath_mulcore_ary1_a0_I0_I1_52__net043));
OR2X1 mul_U1580(.A(n6528), .B(dpath_mulcore_b2[0]), .Y(n11677));
AND2X1 mul_U1581(.A(n286), .B(n11164), .Y(dpath_mulcore_ary1_a0_I1_I1_46__net32));
OR2X1 mul_U1582(.A(n6356), .B(dpath_mulcore_b3[0]), .Y(n11164));
AND2X1 mul_U1583(.A(n285), .B(n11161), .Y(dpath_mulcore_ary1_a0_I1_I1_46__net046));
OR2X1 mul_U1584(.A(n6355), .B(dpath_mulcore_b4[0]), .Y(n11161));
AND2X1 mul_U1585(.A(n458), .B(n11686), .Y(dpath_mulcore_ary1_a0_I0_I1_51__net043));
OR2X1 mul_U1586(.A(n6531), .B(dpath_mulcore_b2[0]), .Y(n11686));
AND2X1 mul_U1587(.A(n289), .B(n11173), .Y(dpath_mulcore_ary1_a0_I1_I1_45__net32));
OR2X1 mul_U1588(.A(n6359), .B(dpath_mulcore_b3[0]), .Y(n11173));
AND2X1 mul_U1589(.A(n288), .B(n11170), .Y(dpath_mulcore_ary1_a0_I1_I1_45__net046));
OR2X1 mul_U1590(.A(n6358), .B(dpath_mulcore_b4[0]), .Y(n11170));
AND2X1 mul_U1591(.A(n461), .B(n11695), .Y(dpath_mulcore_ary1_a0_I0_I1_50__net043));
OR2X1 mul_U1592(.A(n6534), .B(dpath_mulcore_b2[0]), .Y(n11695));
AND2X1 mul_U1593(.A(n292), .B(n11182), .Y(dpath_mulcore_ary1_a0_I1_I1_44__net32));
OR2X1 mul_U1594(.A(n6362), .B(dpath_mulcore_b3[0]), .Y(n11182));
AND2X1 mul_U1595(.A(n291), .B(n11179), .Y(dpath_mulcore_ary1_a0_I1_I1_44__net046));
OR2X1 mul_U1596(.A(n6361), .B(dpath_mulcore_b4[0]), .Y(n11179));
AND2X1 mul_U1597(.A(n464), .B(n11704), .Y(dpath_mulcore_ary1_a0_I0_I1_49__net043));
OR2X1 mul_U1598(.A(n6537), .B(dpath_mulcore_b2[0]), .Y(n11704));
AND2X1 mul_U1599(.A(n295), .B(n11191), .Y(dpath_mulcore_ary1_a0_I1_I1_43__net32));
OR2X1 mul_U1600(.A(n6365), .B(dpath_mulcore_b3[0]), .Y(n11191));
AND2X1 mul_U1601(.A(n294), .B(n11188), .Y(dpath_mulcore_ary1_a0_I1_I1_43__net046));
OR2X1 mul_U1602(.A(n6364), .B(dpath_mulcore_b4[0]), .Y(n11188));
AND2X1 mul_U1603(.A(n467), .B(n11713), .Y(dpath_mulcore_ary1_a0_I0_I1_48__net043));
OR2X1 mul_U1604(.A(n6540), .B(dpath_mulcore_b2[0]), .Y(n11713));
AND2X1 mul_U1605(.A(n298), .B(n11200), .Y(dpath_mulcore_ary1_a0_I1_I1_42__net32));
OR2X1 mul_U1606(.A(n6368), .B(dpath_mulcore_b3[0]), .Y(n11200));
AND2X1 mul_U1607(.A(n297), .B(n11197), .Y(dpath_mulcore_ary1_a0_I1_I1_42__net046));
OR2X1 mul_U1608(.A(n6367), .B(dpath_mulcore_b4[0]), .Y(n11197));
AND2X1 mul_U1609(.A(n470), .B(n11722), .Y(dpath_mulcore_ary1_a0_I0_I1_47__net043));
OR2X1 mul_U1610(.A(n6543), .B(dpath_mulcore_b2[0]), .Y(n11722));
AND2X1 mul_U1611(.A(n301), .B(n11209), .Y(dpath_mulcore_ary1_a0_I1_I1_41__net32));
OR2X1 mul_U1612(.A(n6371), .B(dpath_mulcore_b3[0]), .Y(n11209));
AND2X1 mul_U1613(.A(n300), .B(n11206), .Y(dpath_mulcore_ary1_a0_I1_I1_41__net046));
OR2X1 mul_U1614(.A(n6370), .B(dpath_mulcore_b4[0]), .Y(n11206));
AND2X1 mul_U1615(.A(n473), .B(n11731), .Y(dpath_mulcore_ary1_a0_I0_I1_46__net043));
OR2X1 mul_U1616(.A(n6546), .B(dpath_mulcore_b2[0]), .Y(n11731));
AND2X1 mul_U1617(.A(n304), .B(n11218), .Y(dpath_mulcore_ary1_a0_I1_I1_40__net32));
OR2X1 mul_U1618(.A(n6374), .B(dpath_mulcore_b3[0]), .Y(n11218));
AND2X1 mul_U1619(.A(n303), .B(n11215), .Y(dpath_mulcore_ary1_a0_I1_I1_40__net046));
OR2X1 mul_U1620(.A(n6373), .B(dpath_mulcore_b4[0]), .Y(n11215));
AND2X1 mul_U1621(.A(n476), .B(n11740), .Y(dpath_mulcore_ary1_a0_I0_I1_45__net043));
OR2X1 mul_U1622(.A(n6549), .B(dpath_mulcore_b2[0]), .Y(n11740));
AND2X1 mul_U1623(.A(n307), .B(n11227), .Y(dpath_mulcore_ary1_a0_I1_I1_39__net32));
OR2X1 mul_U1624(.A(n6377), .B(dpath_mulcore_b3[0]), .Y(n11227));
AND2X1 mul_U1625(.A(n306), .B(n11224), .Y(dpath_mulcore_ary1_a0_I1_I1_39__net046));
OR2X1 mul_U1626(.A(n6376), .B(dpath_mulcore_b4[0]), .Y(n11224));
AND2X1 mul_U1627(.A(n479), .B(n11749), .Y(dpath_mulcore_ary1_a0_I0_I1_44__net043));
OR2X1 mul_U1628(.A(n6552), .B(dpath_mulcore_b2[0]), .Y(n11749));
AND2X1 mul_U1629(.A(n310), .B(n11236), .Y(dpath_mulcore_ary1_a0_I1_I1_38__net32));
OR2X1 mul_U1630(.A(n6380), .B(dpath_mulcore_b3[0]), .Y(n11236));
AND2X1 mul_U1631(.A(n309), .B(n11233), .Y(dpath_mulcore_ary1_a0_I1_I1_38__net046));
OR2X1 mul_U1632(.A(n6379), .B(dpath_mulcore_b4[0]), .Y(n11233));
AND2X1 mul_U1633(.A(n482), .B(n11758), .Y(dpath_mulcore_ary1_a0_I0_I1_43__net043));
OR2X1 mul_U1634(.A(n6555), .B(dpath_mulcore_b2[0]), .Y(n11758));
AND2X1 mul_U1635(.A(n313), .B(n11245), .Y(dpath_mulcore_ary1_a0_I1_I1_37__net32));
OR2X1 mul_U1636(.A(n6383), .B(dpath_mulcore_b3[0]), .Y(n11245));
AND2X1 mul_U1637(.A(n312), .B(n11242), .Y(dpath_mulcore_ary1_a0_I1_I1_37__net046));
OR2X1 mul_U1638(.A(n6382), .B(dpath_mulcore_b4[0]), .Y(n11242));
AND2X1 mul_U1639(.A(n485), .B(n11767), .Y(dpath_mulcore_ary1_a0_I0_I1_42__net043));
OR2X1 mul_U1640(.A(n6558), .B(dpath_mulcore_b2[0]), .Y(n11767));
AND2X1 mul_U1641(.A(n316), .B(n11254), .Y(dpath_mulcore_ary1_a0_I1_I1_36__net32));
OR2X1 mul_U1642(.A(n6386), .B(dpath_mulcore_b3[0]), .Y(n11254));
AND2X1 mul_U1643(.A(n315), .B(n11251), .Y(dpath_mulcore_ary1_a0_I1_I1_36__net046));
OR2X1 mul_U1644(.A(n6385), .B(dpath_mulcore_b4[0]), .Y(n11251));
AND2X1 mul_U1645(.A(n488), .B(n11776), .Y(dpath_mulcore_ary1_a0_I0_I1_41__net043));
OR2X1 mul_U1646(.A(n6561), .B(dpath_mulcore_b2[0]), .Y(n11776));
AND2X1 mul_U1647(.A(n319), .B(n11263), .Y(dpath_mulcore_ary1_a0_I1_I1_35__net32));
OR2X1 mul_U1648(.A(n6389), .B(dpath_mulcore_b3[0]), .Y(n11263));
AND2X1 mul_U1649(.A(n318), .B(n11260), .Y(dpath_mulcore_ary1_a0_I1_I1_35__net046));
OR2X1 mul_U1650(.A(n6388), .B(dpath_mulcore_b4[0]), .Y(n11260));
AND2X1 mul_U1651(.A(n491), .B(n11785), .Y(dpath_mulcore_ary1_a0_I0_I1_40__net043));
OR2X1 mul_U1652(.A(n6564), .B(dpath_mulcore_b2[0]), .Y(n11785));
AND2X1 mul_U1653(.A(n322), .B(n11272), .Y(dpath_mulcore_ary1_a0_I1_I1_34__net32));
OR2X1 mul_U1654(.A(n6392), .B(dpath_mulcore_b3[0]), .Y(n11272));
AND2X1 mul_U1655(.A(n321), .B(n11269), .Y(dpath_mulcore_ary1_a0_I1_I1_34__net046));
OR2X1 mul_U1656(.A(n6391), .B(dpath_mulcore_b4[0]), .Y(n11269));
AND2X1 mul_U1657(.A(n494), .B(n11794), .Y(dpath_mulcore_ary1_a0_I0_I1_39__net043));
OR2X1 mul_U1658(.A(n6567), .B(dpath_mulcore_b2[0]), .Y(n11794));
AND2X1 mul_U1659(.A(n325), .B(n11281), .Y(dpath_mulcore_ary1_a0_I1_I1_33__net32));
OR2X1 mul_U1660(.A(n6395), .B(dpath_mulcore_b3[0]), .Y(n11281));
AND2X1 mul_U1661(.A(n324), .B(n11278), .Y(dpath_mulcore_ary1_a0_I1_I1_33__net046));
OR2X1 mul_U1662(.A(n6394), .B(dpath_mulcore_b4[0]), .Y(n11278));
AND2X1 mul_U1663(.A(n497), .B(n11803), .Y(dpath_mulcore_ary1_a0_I0_I1_38__net043));
OR2X1 mul_U1664(.A(n6570), .B(dpath_mulcore_b2[0]), .Y(n11803));
AND2X1 mul_U1665(.A(n328), .B(n11290), .Y(dpath_mulcore_ary1_a0_I1_I1_32__net32));
OR2X1 mul_U1666(.A(n6398), .B(dpath_mulcore_b3[0]), .Y(n11290));
AND2X1 mul_U1667(.A(n327), .B(n11287), .Y(dpath_mulcore_ary1_a0_I1_I1_32__net046));
OR2X1 mul_U1668(.A(n6397), .B(dpath_mulcore_b4[0]), .Y(n11287));
AND2X1 mul_U1669(.A(n500), .B(n11812), .Y(dpath_mulcore_ary1_a0_I0_I1_37__net043));
OR2X1 mul_U1670(.A(n6573), .B(dpath_mulcore_b2[0]), .Y(n11812));
AND2X1 mul_U1671(.A(n331), .B(n11299), .Y(dpath_mulcore_ary1_a0_I1_I1_31__net32));
OR2X1 mul_U1672(.A(n6401), .B(dpath_mulcore_b3[0]), .Y(n11299));
AND2X1 mul_U1673(.A(n330), .B(n11296), .Y(dpath_mulcore_ary1_a0_I1_I1_31__net046));
OR2X1 mul_U1674(.A(n6400), .B(dpath_mulcore_b4[0]), .Y(n11296));
AND2X1 mul_U1675(.A(n503), .B(n11821), .Y(dpath_mulcore_ary1_a0_I0_I1_36__net043));
OR2X1 mul_U1676(.A(n6576), .B(dpath_mulcore_b2[0]), .Y(n11821));
AND2X1 mul_U1677(.A(n334), .B(n11308), .Y(dpath_mulcore_ary1_a0_I1_I1_30__net32));
OR2X1 mul_U1678(.A(n6404), .B(dpath_mulcore_b3[0]), .Y(n11308));
AND2X1 mul_U1679(.A(n333), .B(n11305), .Y(dpath_mulcore_ary1_a0_I1_I1_30__net046));
OR2X1 mul_U1680(.A(n6403), .B(dpath_mulcore_b4[0]), .Y(n11305));
AND2X1 mul_U1681(.A(n506), .B(n11830), .Y(dpath_mulcore_ary1_a0_I0_I1_35__net043));
OR2X1 mul_U1682(.A(n6579), .B(dpath_mulcore_b2[0]), .Y(n11830));
AND2X1 mul_U1683(.A(n337), .B(n11317), .Y(dpath_mulcore_ary1_a0_I1_I1_29__net32));
OR2X1 mul_U1684(.A(n6407), .B(dpath_mulcore_b3[0]), .Y(n11317));
AND2X1 mul_U1685(.A(n336), .B(n11314), .Y(dpath_mulcore_ary1_a0_I1_I1_29__net046));
OR2X1 mul_U1686(.A(n6406), .B(dpath_mulcore_b4[0]), .Y(n11314));
AND2X1 mul_U1687(.A(n509), .B(n11839), .Y(dpath_mulcore_ary1_a0_I0_I1_34__net043));
OR2X1 mul_U1688(.A(n6582), .B(dpath_mulcore_b2[0]), .Y(n11839));
AND2X1 mul_U1689(.A(n340), .B(n11326), .Y(dpath_mulcore_ary1_a0_I1_I1_28__net32));
OR2X1 mul_U1690(.A(n6410), .B(dpath_mulcore_b3[0]), .Y(n11326));
AND2X1 mul_U1691(.A(n339), .B(n11323), .Y(dpath_mulcore_ary1_a0_I1_I1_28__net046));
OR2X1 mul_U1692(.A(n6409), .B(dpath_mulcore_b4[0]), .Y(n11323));
AND2X1 mul_U1693(.A(n512), .B(n11848), .Y(dpath_mulcore_ary1_a0_I0_I1_33__net043));
OR2X1 mul_U1694(.A(n6585), .B(dpath_mulcore_b2[0]), .Y(n11848));
AND2X1 mul_U1695(.A(n343), .B(n11335), .Y(dpath_mulcore_ary1_a0_I1_I1_27__net32));
OR2X1 mul_U1696(.A(n6413), .B(dpath_mulcore_b3[0]), .Y(n11335));
AND2X1 mul_U1697(.A(n342), .B(n11332), .Y(dpath_mulcore_ary1_a0_I1_I1_27__net046));
OR2X1 mul_U1698(.A(n6412), .B(dpath_mulcore_b4[0]), .Y(n11332));
AND2X1 mul_U1699(.A(n515), .B(n11857), .Y(dpath_mulcore_ary1_a0_I0_I1_32__net043));
OR2X1 mul_U1700(.A(n6588), .B(dpath_mulcore_b2[0]), .Y(n11857));
AND2X1 mul_U1701(.A(n346), .B(n11344), .Y(dpath_mulcore_ary1_a0_I1_I1_26__net32));
OR2X1 mul_U1702(.A(n6416), .B(dpath_mulcore_b3[0]), .Y(n11344));
AND2X1 mul_U1703(.A(n345), .B(n11341), .Y(dpath_mulcore_ary1_a0_I1_I1_26__net046));
OR2X1 mul_U1704(.A(n6415), .B(dpath_mulcore_b4[0]), .Y(n11341));
AND2X1 mul_U1705(.A(n518), .B(n11866), .Y(dpath_mulcore_ary1_a0_I0_I1_31__net043));
OR2X1 mul_U1706(.A(n6591), .B(dpath_mulcore_b2[0]), .Y(n11866));
AND2X1 mul_U1707(.A(n349), .B(n11353), .Y(dpath_mulcore_ary1_a0_I1_I1_25__net32));
OR2X1 mul_U1708(.A(n6419), .B(dpath_mulcore_b3[0]), .Y(n11353));
AND2X1 mul_U1709(.A(n348), .B(n11350), .Y(dpath_mulcore_ary1_a0_I1_I1_25__net046));
OR2X1 mul_U1710(.A(n6418), .B(dpath_mulcore_b4[0]), .Y(n11350));
AND2X1 mul_U1711(.A(n521), .B(n11875), .Y(dpath_mulcore_ary1_a0_I0_I1_30__net043));
OR2X1 mul_U1712(.A(n6594), .B(dpath_mulcore_b2[0]), .Y(n11875));
AND2X1 mul_U1713(.A(n352), .B(n11362), .Y(dpath_mulcore_ary1_a0_I1_I1_24__net32));
OR2X1 mul_U1714(.A(n6422), .B(dpath_mulcore_b3[0]), .Y(n11362));
AND2X1 mul_U1715(.A(n351), .B(n11359), .Y(dpath_mulcore_ary1_a0_I1_I1_24__net046));
OR2X1 mul_U1716(.A(n6421), .B(dpath_mulcore_b4[0]), .Y(n11359));
AND2X1 mul_U1717(.A(n524), .B(n11884), .Y(dpath_mulcore_ary1_a0_I0_I1_29__net043));
OR2X1 mul_U1718(.A(n6597), .B(dpath_mulcore_b2[0]), .Y(n11884));
AND2X1 mul_U1719(.A(n355), .B(n11371), .Y(dpath_mulcore_ary1_a0_I1_I1_23__net32));
OR2X1 mul_U1720(.A(n6425), .B(dpath_mulcore_b3[0]), .Y(n11371));
AND2X1 mul_U1721(.A(n354), .B(n11368), .Y(dpath_mulcore_ary1_a0_I1_I1_23__net046));
OR2X1 mul_U1722(.A(n6424), .B(dpath_mulcore_b4[0]), .Y(n11368));
AND2X1 mul_U1723(.A(n527), .B(n11893), .Y(dpath_mulcore_ary1_a0_I0_I1_28__net043));
OR2X1 mul_U1724(.A(n6600), .B(dpath_mulcore_b2[0]), .Y(n11893));
AND2X1 mul_U1725(.A(n358), .B(n11380), .Y(dpath_mulcore_ary1_a0_I1_I1_22__net32));
OR2X1 mul_U1726(.A(n6428), .B(dpath_mulcore_b3[0]), .Y(n11380));
AND2X1 mul_U1727(.A(n357), .B(n11377), .Y(dpath_mulcore_ary1_a0_I1_I1_22__net046));
OR2X1 mul_U1728(.A(n6427), .B(dpath_mulcore_b4[0]), .Y(n11377));
AND2X1 mul_U1729(.A(n530), .B(n11902), .Y(dpath_mulcore_ary1_a0_I0_I1_27__net043));
OR2X1 mul_U1730(.A(n6603), .B(dpath_mulcore_b2[0]), .Y(n11902));
AND2X1 mul_U1731(.A(n361), .B(n11389), .Y(dpath_mulcore_ary1_a0_I1_I1_21__net32));
OR2X1 mul_U1732(.A(n6431), .B(dpath_mulcore_b3[0]), .Y(n11389));
AND2X1 mul_U1733(.A(n360), .B(n11386), .Y(dpath_mulcore_ary1_a0_I1_I1_21__net046));
OR2X1 mul_U1734(.A(n6430), .B(dpath_mulcore_b4[0]), .Y(n11386));
AND2X1 mul_U1735(.A(n533), .B(n11911), .Y(dpath_mulcore_ary1_a0_I0_I1_26__net043));
OR2X1 mul_U1736(.A(n6606), .B(dpath_mulcore_b2[0]), .Y(n11911));
AND2X1 mul_U1737(.A(n364), .B(n11398), .Y(dpath_mulcore_ary1_a0_I1_I1_20__net32));
OR2X1 mul_U1738(.A(n6434), .B(dpath_mulcore_b3[0]), .Y(n11398));
AND2X1 mul_U1739(.A(n363), .B(n11395), .Y(dpath_mulcore_ary1_a0_I1_I1_20__net046));
OR2X1 mul_U1740(.A(n6433), .B(dpath_mulcore_b4[0]), .Y(n11395));
AND2X1 mul_U1741(.A(n536), .B(n11920), .Y(dpath_mulcore_ary1_a0_I0_I1_25__net043));
OR2X1 mul_U1742(.A(n6609), .B(dpath_mulcore_b2[0]), .Y(n11920));
AND2X1 mul_U1743(.A(n367), .B(n11407), .Y(dpath_mulcore_ary1_a0_I1_I1_19__net32));
OR2X1 mul_U1744(.A(n6437), .B(dpath_mulcore_b3[0]), .Y(n11407));
AND2X1 mul_U1745(.A(n366), .B(n11404), .Y(dpath_mulcore_ary1_a0_I1_I1_19__net046));
OR2X1 mul_U1746(.A(n6436), .B(dpath_mulcore_b4[0]), .Y(n11404));
AND2X1 mul_U1747(.A(n539), .B(n11929), .Y(dpath_mulcore_ary1_a0_I0_I1_24__net043));
OR2X1 mul_U1748(.A(n6612), .B(dpath_mulcore_b2[0]), .Y(n11929));
AND2X1 mul_U1749(.A(n370), .B(n11416), .Y(dpath_mulcore_ary1_a0_I1_I1_18__net32));
OR2X1 mul_U1750(.A(n6440), .B(dpath_mulcore_b3[0]), .Y(n11416));
AND2X1 mul_U1751(.A(n369), .B(n11413), .Y(dpath_mulcore_ary1_a0_I1_I1_18__net046));
OR2X1 mul_U1752(.A(n6439), .B(dpath_mulcore_b4[0]), .Y(n11413));
AND2X1 mul_U1753(.A(n542), .B(n11938), .Y(dpath_mulcore_ary1_a0_I0_I1_23__net043));
OR2X1 mul_U1754(.A(n6615), .B(dpath_mulcore_b2[0]), .Y(n11938));
AND2X1 mul_U1755(.A(n373), .B(n11425), .Y(dpath_mulcore_ary1_a0_I1_I1_17__net32));
OR2X1 mul_U1756(.A(n6443), .B(dpath_mulcore_b3[0]), .Y(n11425));
AND2X1 mul_U1757(.A(n372), .B(n11422), .Y(dpath_mulcore_ary1_a0_I1_I1_17__net046));
OR2X1 mul_U1758(.A(n6442), .B(dpath_mulcore_b4[0]), .Y(n11422));
AND2X1 mul_U1759(.A(n545), .B(n11947), .Y(dpath_mulcore_ary1_a0_I0_I1_22__net043));
OR2X1 mul_U1760(.A(n6618), .B(dpath_mulcore_b2[0]), .Y(n11947));
AND2X1 mul_U1761(.A(n376), .B(n11434), .Y(dpath_mulcore_ary1_a0_I1_I1_16__net32));
OR2X1 mul_U1762(.A(n6446), .B(dpath_mulcore_b3[0]), .Y(n11434));
AND2X1 mul_U1763(.A(n375), .B(n11431), .Y(dpath_mulcore_ary1_a0_I1_I1_16__net046));
OR2X1 mul_U1764(.A(n6445), .B(dpath_mulcore_b4[0]), .Y(n11431));
AND2X1 mul_U1765(.A(n548), .B(n11956), .Y(dpath_mulcore_ary1_a0_I0_I1_21__net043));
OR2X1 mul_U1766(.A(n6621), .B(dpath_mulcore_b2[0]), .Y(n11956));
AND2X1 mul_U1767(.A(n379), .B(n11443), .Y(dpath_mulcore_ary1_a0_I1_I1_15__net32));
OR2X1 mul_U1768(.A(n6449), .B(dpath_mulcore_b3[0]), .Y(n11443));
AND2X1 mul_U1769(.A(n378), .B(n11440), .Y(dpath_mulcore_ary1_a0_I1_I1_15__net046));
OR2X1 mul_U1770(.A(n6448), .B(dpath_mulcore_b4[0]), .Y(n11440));
AND2X1 mul_U1771(.A(n551), .B(n11965), .Y(dpath_mulcore_ary1_a0_I0_I1_20__net043));
OR2X1 mul_U1772(.A(n6624), .B(dpath_mulcore_b2[0]), .Y(n11965));
AND2X1 mul_U1773(.A(n382), .B(n11452), .Y(dpath_mulcore_ary1_a0_I1_I1_14__net32));
OR2X1 mul_U1774(.A(n6452), .B(dpath_mulcore_b3[0]), .Y(n11452));
AND2X1 mul_U1775(.A(n381), .B(n11449), .Y(dpath_mulcore_ary1_a0_I1_I1_14__net046));
OR2X1 mul_U1776(.A(n6451), .B(dpath_mulcore_b4[0]), .Y(n11449));
AND2X1 mul_U1777(.A(n554), .B(n11974), .Y(dpath_mulcore_ary1_a0_I0_I1_19__net043));
OR2X1 mul_U1778(.A(n6627), .B(dpath_mulcore_b2[0]), .Y(n11974));
AND2X1 mul_U1779(.A(n385), .B(n11461), .Y(dpath_mulcore_ary1_a0_I1_I1_13__net32));
OR2X1 mul_U1780(.A(n6455), .B(dpath_mulcore_b3[0]), .Y(n11461));
AND2X1 mul_U1781(.A(n384), .B(n11458), .Y(dpath_mulcore_ary1_a0_I1_I1_13__net046));
OR2X1 mul_U1782(.A(n6454), .B(dpath_mulcore_b4[0]), .Y(n11458));
AND2X1 mul_U1783(.A(n557), .B(n11983), .Y(dpath_mulcore_ary1_a0_I0_I1_18__net043));
OR2X1 mul_U1784(.A(n6630), .B(dpath_mulcore_b2[0]), .Y(n11983));
AND2X1 mul_U1785(.A(n388), .B(n11470), .Y(dpath_mulcore_ary1_a0_I1_I1_12__net32));
OR2X1 mul_U1786(.A(n6458), .B(dpath_mulcore_b3[0]), .Y(n11470));
AND2X1 mul_U1787(.A(n387), .B(n11467), .Y(dpath_mulcore_ary1_a0_I1_I1_12__net046));
OR2X1 mul_U1788(.A(n6457), .B(dpath_mulcore_b4[0]), .Y(n11467));
AND2X1 mul_U1789(.A(n560), .B(n11992), .Y(dpath_mulcore_ary1_a0_I0_I1_17__net043));
OR2X1 mul_U1790(.A(n6633), .B(dpath_mulcore_b2[0]), .Y(n11992));
AND2X1 mul_U1791(.A(n391), .B(n11479), .Y(dpath_mulcore_ary1_a0_I1_I1_11__net32));
OR2X1 mul_U1792(.A(n6461), .B(dpath_mulcore_b3[0]), .Y(n11479));
AND2X1 mul_U1793(.A(n390), .B(n11476), .Y(dpath_mulcore_ary1_a0_I1_I1_11__net046));
OR2X1 mul_U1794(.A(n6460), .B(dpath_mulcore_b4[0]), .Y(n11476));
AND2X1 mul_U1795(.A(n563), .B(n12001), .Y(dpath_mulcore_ary1_a0_I0_I1_16__net043));
OR2X1 mul_U1796(.A(n6636), .B(dpath_mulcore_b2[0]), .Y(n12001));
AND2X1 mul_U1797(.A(n394), .B(n11488), .Y(dpath_mulcore_ary1_a0_I1_I1_10__net32));
OR2X1 mul_U1798(.A(n6464), .B(dpath_mulcore_b3[0]), .Y(n11488));
AND2X1 mul_U1799(.A(n393), .B(n11485), .Y(dpath_mulcore_ary1_a0_I1_I1_10__net046));
OR2X1 mul_U1800(.A(n6463), .B(dpath_mulcore_b4[0]), .Y(n11485));
AND2X1 mul_U1801(.A(n566), .B(n12010), .Y(dpath_mulcore_ary1_a0_I0_I1_15__net043));
OR2X1 mul_U1802(.A(n6639), .B(dpath_mulcore_b2[0]), .Y(n12010));
AND2X1 mul_U1803(.A(n397), .B(n11497), .Y(dpath_mulcore_ary1_a0_I1_I1_9__net32));
OR2X1 mul_U1804(.A(n6467), .B(dpath_mulcore_b3[0]), .Y(n11497));
AND2X1 mul_U1805(.A(n396), .B(n11494), .Y(dpath_mulcore_ary1_a0_I1_I1_9__net046));
OR2X1 mul_U1806(.A(n6466), .B(dpath_mulcore_b4[0]), .Y(n11494));
AND2X1 mul_U1807(.A(n569), .B(n12019), .Y(dpath_mulcore_ary1_a0_I0_I1_14__net043));
OR2X1 mul_U1808(.A(n6642), .B(dpath_mulcore_b2[0]), .Y(n12019));
AND2X1 mul_U1809(.A(n400), .B(n11506), .Y(dpath_mulcore_ary1_a0_I1_I1_8__net32));
OR2X1 mul_U1810(.A(n6470), .B(dpath_mulcore_b3[0]), .Y(n11506));
AND2X1 mul_U1811(.A(n399), .B(n11503), .Y(dpath_mulcore_ary1_a0_I1_I1_8__net046));
OR2X1 mul_U1812(.A(n6469), .B(dpath_mulcore_b4[0]), .Y(n11503));
AND2X1 mul_U1813(.A(n403), .B(n11515), .Y(dpath_mulcore_ary1_a0_I1_I1_7__net32));
OR2X1 mul_U1814(.A(n6473), .B(dpath_mulcore_b3[0]), .Y(n11515));
AND2X1 mul_U1815(.A(n402), .B(n11512), .Y(dpath_mulcore_ary1_a0_I1_I1_7__net046));
OR2X1 mul_U1816(.A(n6472), .B(dpath_mulcore_b4[0]), .Y(n11512));
AND2X1 mul_U1817(.A(n574), .B(n12034), .Y(dpath_mulcore_ary1_a0_I0_I1_13__net32));
OR2X1 mul_U1818(.A(n6647), .B(dpath_mulcore_b0[0]), .Y(n12034));
AND2X1 mul_U1819(.A(n573), .B(n12031), .Y(dpath_mulcore_ary1_a0_I0_I1_13__net046));
OR2X1 mul_U1820(.A(n6646), .B(dpath_mulcore_b1[0]), .Y(n12031));
AND2X1 mul_U1821(.A(n406), .B(n11524), .Y(dpath_mulcore_ary1_a0_I1_I1_6__net32));
OR2X1 mul_U1822(.A(n6476), .B(dpath_mulcore_b3[0]), .Y(n11524));
AND2X1 mul_U1823(.A(n405), .B(n11521), .Y(dpath_mulcore_ary1_a0_I1_I1_6__net046));
OR2X1 mul_U1824(.A(n6475), .B(dpath_mulcore_b4[0]), .Y(n11521));
AND2X1 mul_U1825(.A(n577), .B(n12043), .Y(dpath_mulcore_ary1_a0_I0_I1_12__net32));
OR2X1 mul_U1826(.A(n6650), .B(dpath_mulcore_b0[0]), .Y(n12043));
AND2X1 mul_U1827(.A(n576), .B(n12040), .Y(dpath_mulcore_ary1_a0_I0_I1_12__net046));
OR2X1 mul_U1828(.A(n6649), .B(dpath_mulcore_b1[0]), .Y(n12040));
AND2X1 mul_U1829(.A(n409), .B(n11533), .Y(dpath_mulcore_ary1_a0_I1_I1_5__net32));
OR2X1 mul_U1830(.A(n6479), .B(dpath_mulcore_b3[0]), .Y(n11533));
AND2X1 mul_U1831(.A(n408), .B(n11530), .Y(dpath_mulcore_ary1_a0_I1_I1_5__net046));
OR2X1 mul_U1832(.A(n6478), .B(dpath_mulcore_b4[0]), .Y(n11530));
AND2X1 mul_U1833(.A(n106), .B(n10620), .Y(dpath_mulcore_ary1_a0_I2_I1_62__net32));
OR2X1 mul_U1834(.A(n6174), .B(dpath_mulcore_b6[0]), .Y(n10620));
AND2X1 mul_U1835(.A(n105), .B(n10617), .Y(dpath_mulcore_ary1_a0_I2_I1_62__net046));
OR2X1 mul_U1836(.A(n6173), .B(dpath_mulcore_b7[0]), .Y(n10617));
AND2X1 mul_U1837(.A(n108), .B(n10626), .Y(dpath_mulcore_ary1_a0_I2_I1_61__net32));
OR2X1 mul_U1838(.A(n6176), .B(dpath_mulcore_b6[0]), .Y(n10626));
AND2X1 mul_U1839(.A(n107), .B(n10623), .Y(dpath_mulcore_ary1_a0_I2_I1_61__net046));
OR2X1 mul_U1840(.A(n6175), .B(dpath_mulcore_b7[0]), .Y(n10623));
AND2X1 mul_U1841(.A(n110), .B(n10632), .Y(dpath_mulcore_ary1_a0_I2_I1_60__net32));
OR2X1 mul_U1842(.A(n6178), .B(dpath_mulcore_b6[0]), .Y(n10632));
AND2X1 mul_U1843(.A(n109), .B(n10629), .Y(dpath_mulcore_ary1_a0_I2_I1_60__net046));
OR2X1 mul_U1844(.A(n6177), .B(dpath_mulcore_b7[0]), .Y(n10629));
AND2X1 mul_U1845(.A(n112), .B(n10638), .Y(dpath_mulcore_ary1_a0_I2_I1_59__net32));
OR2X1 mul_U1846(.A(n6180), .B(dpath_mulcore_b6[0]), .Y(n10638));
AND2X1 mul_U1847(.A(n111), .B(n10635), .Y(dpath_mulcore_ary1_a0_I2_I1_59__net046));
OR2X1 mul_U1848(.A(n6179), .B(dpath_mulcore_b7[0]), .Y(n10635));
AND2X1 mul_U1849(.A(n114), .B(n10644), .Y(dpath_mulcore_ary1_a0_I2_I1_58__net32));
OR2X1 mul_U1850(.A(n6182), .B(dpath_mulcore_b6[0]), .Y(n10644));
AND2X1 mul_U1851(.A(n113), .B(n10641), .Y(dpath_mulcore_ary1_a0_I2_I1_58__net046));
OR2X1 mul_U1852(.A(n6181), .B(dpath_mulcore_b7[0]), .Y(n10641));
AND2X1 mul_U1853(.A(n116), .B(n10650), .Y(dpath_mulcore_ary1_a0_I2_I1_57__net32));
OR2X1 mul_U1854(.A(n6184), .B(dpath_mulcore_b6[0]), .Y(n10650));
AND2X1 mul_U1855(.A(n115), .B(n10647), .Y(dpath_mulcore_ary1_a0_I2_I1_57__net046));
OR2X1 mul_U1856(.A(n6183), .B(dpath_mulcore_b7[0]), .Y(n10647));
AND2X1 mul_U1857(.A(n118), .B(n10656), .Y(dpath_mulcore_ary1_a0_I2_I1_56__net32));
OR2X1 mul_U1858(.A(n6186), .B(dpath_mulcore_b6[0]), .Y(n10656));
AND2X1 mul_U1859(.A(n117), .B(n10653), .Y(dpath_mulcore_ary1_a0_I2_I1_56__net046));
OR2X1 mul_U1860(.A(n6185), .B(dpath_mulcore_b7[0]), .Y(n10653));
AND2X1 mul_U1861(.A(n120), .B(n10662), .Y(dpath_mulcore_ary1_a0_I2_I1_55__net32));
OR2X1 mul_U1862(.A(n6188), .B(dpath_mulcore_b6[0]), .Y(n10662));
AND2X1 mul_U1863(.A(n119), .B(n10659), .Y(dpath_mulcore_ary1_a0_I2_I1_55__net046));
OR2X1 mul_U1864(.A(n6187), .B(dpath_mulcore_b7[0]), .Y(n10659));
AND2X1 mul_U1865(.A(n122), .B(n10668), .Y(dpath_mulcore_ary1_a0_I2_I1_54__net32));
OR2X1 mul_U1866(.A(n6190), .B(dpath_mulcore_b6[0]), .Y(n10668));
AND2X1 mul_U1867(.A(n121), .B(n10665), .Y(dpath_mulcore_ary1_a0_I2_I1_54__net046));
OR2X1 mul_U1868(.A(n6189), .B(dpath_mulcore_b7[0]), .Y(n10665));
AND2X1 mul_U1869(.A(n124), .B(n10674), .Y(dpath_mulcore_ary1_a0_I2_I1_53__net32));
OR2X1 mul_U1870(.A(n6192), .B(dpath_mulcore_b6[0]), .Y(n10674));
AND2X1 mul_U1871(.A(n123), .B(n10671), .Y(dpath_mulcore_ary1_a0_I2_I1_53__net046));
OR2X1 mul_U1872(.A(n6191), .B(dpath_mulcore_b7[0]), .Y(n10671));
AND2X1 mul_U1873(.A(n126), .B(n10680), .Y(dpath_mulcore_ary1_a0_I2_I1_52__net32));
OR2X1 mul_U1874(.A(n6194), .B(dpath_mulcore_b6[0]), .Y(n10680));
AND2X1 mul_U1875(.A(n125), .B(n10677), .Y(dpath_mulcore_ary1_a0_I2_I1_52__net046));
OR2X1 mul_U1876(.A(n6193), .B(dpath_mulcore_b7[0]), .Y(n10677));
AND2X1 mul_U1877(.A(n128), .B(n10686), .Y(dpath_mulcore_ary1_a0_I2_I1_51__net32));
OR2X1 mul_U1878(.A(n6196), .B(dpath_mulcore_b6[0]), .Y(n10686));
AND2X1 mul_U1879(.A(n127), .B(n10683), .Y(dpath_mulcore_ary1_a0_I2_I1_51__net046));
OR2X1 mul_U1880(.A(n6195), .B(dpath_mulcore_b7[0]), .Y(n10683));
AND2X1 mul_U1881(.A(n130), .B(n10692), .Y(dpath_mulcore_ary1_a0_I2_I1_50__net32));
OR2X1 mul_U1882(.A(n6198), .B(dpath_mulcore_b6[0]), .Y(n10692));
AND2X1 mul_U1883(.A(n129), .B(n10689), .Y(dpath_mulcore_ary1_a0_I2_I1_50__net046));
OR2X1 mul_U1884(.A(n6197), .B(dpath_mulcore_b7[0]), .Y(n10689));
AND2X1 mul_U1885(.A(n132), .B(n10698), .Y(dpath_mulcore_ary1_a0_I2_I1_49__net32));
OR2X1 mul_U1886(.A(n6200), .B(dpath_mulcore_b6[0]), .Y(n10698));
AND2X1 mul_U1887(.A(n131), .B(n10695), .Y(dpath_mulcore_ary1_a0_I2_I1_49__net046));
OR2X1 mul_U1888(.A(n6199), .B(dpath_mulcore_b7[0]), .Y(n10695));
AND2X1 mul_U1889(.A(n134), .B(n10704), .Y(dpath_mulcore_ary1_a0_I2_I1_48__net32));
OR2X1 mul_U1890(.A(n6202), .B(dpath_mulcore_b6[0]), .Y(n10704));
AND2X1 mul_U1891(.A(n133), .B(n10701), .Y(dpath_mulcore_ary1_a0_I2_I1_48__net046));
OR2X1 mul_U1892(.A(n6201), .B(dpath_mulcore_b7[0]), .Y(n10701));
AND2X1 mul_U1893(.A(n136), .B(n10710), .Y(dpath_mulcore_ary1_a0_I2_I1_47__net32));
OR2X1 mul_U1894(.A(n6204), .B(dpath_mulcore_b6[0]), .Y(n10710));
AND2X1 mul_U1895(.A(n135), .B(n10707), .Y(dpath_mulcore_ary1_a0_I2_I1_47__net046));
OR2X1 mul_U1896(.A(n6203), .B(dpath_mulcore_b7[0]), .Y(n10707));
AND2X1 mul_U1897(.A(n138), .B(n10716), .Y(dpath_mulcore_ary1_a0_I2_I1_46__net32));
OR2X1 mul_U1898(.A(n6206), .B(dpath_mulcore_b6[0]), .Y(n10716));
AND2X1 mul_U1899(.A(n137), .B(n10713), .Y(dpath_mulcore_ary1_a0_I2_I1_46__net046));
OR2X1 mul_U1900(.A(n6205), .B(dpath_mulcore_b7[0]), .Y(n10713));
AND2X1 mul_U1901(.A(n140), .B(n10722), .Y(dpath_mulcore_ary1_a0_I2_I1_45__net32));
OR2X1 mul_U1902(.A(n6208), .B(dpath_mulcore_b6[0]), .Y(n10722));
AND2X1 mul_U1903(.A(n139), .B(n10719), .Y(dpath_mulcore_ary1_a0_I2_I1_45__net046));
OR2X1 mul_U1904(.A(n6207), .B(dpath_mulcore_b7[0]), .Y(n10719));
AND2X1 mul_U1905(.A(n142), .B(n10728), .Y(dpath_mulcore_ary1_a0_I2_I1_44__net32));
OR2X1 mul_U1906(.A(n6210), .B(dpath_mulcore_b6[0]), .Y(n10728));
AND2X1 mul_U1907(.A(n141), .B(n10725), .Y(dpath_mulcore_ary1_a0_I2_I1_44__net046));
OR2X1 mul_U1908(.A(n6209), .B(dpath_mulcore_b7[0]), .Y(n10725));
AND2X1 mul_U1909(.A(n144), .B(n10734), .Y(dpath_mulcore_ary1_a0_I2_I1_43__net32));
OR2X1 mul_U1910(.A(n6212), .B(dpath_mulcore_b6[0]), .Y(n10734));
AND2X1 mul_U1911(.A(n143), .B(n10731), .Y(dpath_mulcore_ary1_a0_I2_I1_43__net046));
OR2X1 mul_U1912(.A(n6211), .B(dpath_mulcore_b7[0]), .Y(n10731));
AND2X1 mul_U1913(.A(n146), .B(n10740), .Y(dpath_mulcore_ary1_a0_I2_I1_42__net32));
OR2X1 mul_U1914(.A(n6214), .B(dpath_mulcore_b6[0]), .Y(n10740));
AND2X1 mul_U1915(.A(n145), .B(n10737), .Y(dpath_mulcore_ary1_a0_I2_I1_42__net046));
OR2X1 mul_U1916(.A(n6213), .B(dpath_mulcore_b7[0]), .Y(n10737));
AND2X1 mul_U1917(.A(n148), .B(n10746), .Y(dpath_mulcore_ary1_a0_I2_I1_41__net32));
OR2X1 mul_U1918(.A(n6216), .B(dpath_mulcore_b6[0]), .Y(n10746));
AND2X1 mul_U1919(.A(n147), .B(n10743), .Y(dpath_mulcore_ary1_a0_I2_I1_41__net046));
OR2X1 mul_U1920(.A(n6215), .B(dpath_mulcore_b7[0]), .Y(n10743));
AND2X1 mul_U1921(.A(n150), .B(n10752), .Y(dpath_mulcore_ary1_a0_I2_I1_40__net32));
OR2X1 mul_U1922(.A(n6218), .B(dpath_mulcore_b6[0]), .Y(n10752));
AND2X1 mul_U1923(.A(n149), .B(n10749), .Y(dpath_mulcore_ary1_a0_I2_I1_40__net046));
OR2X1 mul_U1924(.A(n6217), .B(dpath_mulcore_b7[0]), .Y(n10749));
AND2X1 mul_U1925(.A(n152), .B(n10758), .Y(dpath_mulcore_ary1_a0_I2_I1_39__net32));
OR2X1 mul_U1926(.A(n6220), .B(dpath_mulcore_b6[0]), .Y(n10758));
AND2X1 mul_U1927(.A(n151), .B(n10755), .Y(dpath_mulcore_ary1_a0_I2_I1_39__net046));
OR2X1 mul_U1928(.A(n6219), .B(dpath_mulcore_b7[0]), .Y(n10755));
AND2X1 mul_U1929(.A(n154), .B(n10764), .Y(dpath_mulcore_ary1_a0_I2_I1_38__net32));
OR2X1 mul_U1930(.A(n6222), .B(dpath_mulcore_b6[0]), .Y(n10764));
AND2X1 mul_U1931(.A(n153), .B(n10761), .Y(dpath_mulcore_ary1_a0_I2_I1_38__net046));
OR2X1 mul_U1932(.A(n6221), .B(dpath_mulcore_b7[0]), .Y(n10761));
AND2X1 mul_U1933(.A(n156), .B(n10770), .Y(dpath_mulcore_ary1_a0_I2_I1_37__net32));
OR2X1 mul_U1934(.A(n6224), .B(dpath_mulcore_b6[0]), .Y(n10770));
AND2X1 mul_U1935(.A(n155), .B(n10767), .Y(dpath_mulcore_ary1_a0_I2_I1_37__net046));
OR2X1 mul_U1936(.A(n6223), .B(dpath_mulcore_b7[0]), .Y(n10767));
AND2X1 mul_U1937(.A(n158), .B(n10776), .Y(dpath_mulcore_ary1_a0_I2_I1_36__net32));
OR2X1 mul_U1938(.A(n6226), .B(dpath_mulcore_b6[0]), .Y(n10776));
AND2X1 mul_U1939(.A(n157), .B(n10773), .Y(dpath_mulcore_ary1_a0_I2_I1_36__net046));
OR2X1 mul_U1940(.A(n6225), .B(dpath_mulcore_b7[0]), .Y(n10773));
AND2X1 mul_U1941(.A(n160), .B(n10782), .Y(dpath_mulcore_ary1_a0_I2_I1_35__net32));
OR2X1 mul_U1942(.A(n6228), .B(dpath_mulcore_b6[0]), .Y(n10782));
AND2X1 mul_U1943(.A(n159), .B(n10779), .Y(dpath_mulcore_ary1_a0_I2_I1_35__net046));
OR2X1 mul_U1944(.A(n6227), .B(dpath_mulcore_b7[0]), .Y(n10779));
AND2X1 mul_U1945(.A(n162), .B(n10788), .Y(dpath_mulcore_ary1_a0_I2_I1_34__net32));
OR2X1 mul_U1946(.A(n6230), .B(dpath_mulcore_b6[0]), .Y(n10788));
AND2X1 mul_U1947(.A(n161), .B(n10785), .Y(dpath_mulcore_ary1_a0_I2_I1_34__net046));
OR2X1 mul_U1948(.A(n6229), .B(dpath_mulcore_b7[0]), .Y(n10785));
AND2X1 mul_U1949(.A(n164), .B(n10794), .Y(dpath_mulcore_ary1_a0_I2_I1_33__net32));
OR2X1 mul_U1950(.A(n6232), .B(dpath_mulcore_b6[0]), .Y(n10794));
AND2X1 mul_U1951(.A(n163), .B(n10791), .Y(dpath_mulcore_ary1_a0_I2_I1_33__net046));
OR2X1 mul_U1952(.A(n6231), .B(dpath_mulcore_b7[0]), .Y(n10791));
AND2X1 mul_U1953(.A(n166), .B(n10800), .Y(dpath_mulcore_ary1_a0_I2_I1_32__net32));
OR2X1 mul_U1954(.A(n6234), .B(dpath_mulcore_b6[0]), .Y(n10800));
AND2X1 mul_U1955(.A(n165), .B(n10797), .Y(dpath_mulcore_ary1_a0_I2_I1_32__net046));
OR2X1 mul_U1956(.A(n6233), .B(dpath_mulcore_b7[0]), .Y(n10797));
AND2X1 mul_U1957(.A(n168), .B(n10806), .Y(dpath_mulcore_ary1_a0_I2_I1_31__net32));
OR2X1 mul_U1958(.A(n6236), .B(dpath_mulcore_b6[0]), .Y(n10806));
AND2X1 mul_U1959(.A(n167), .B(n10803), .Y(dpath_mulcore_ary1_a0_I2_I1_31__net046));
OR2X1 mul_U1960(.A(n6235), .B(dpath_mulcore_b7[0]), .Y(n10803));
AND2X1 mul_U1961(.A(n170), .B(n10812), .Y(dpath_mulcore_ary1_a0_I2_I1_30__net32));
OR2X1 mul_U1962(.A(n6238), .B(dpath_mulcore_b6[0]), .Y(n10812));
AND2X1 mul_U1963(.A(n169), .B(n10809), .Y(dpath_mulcore_ary1_a0_I2_I1_30__net046));
OR2X1 mul_U1964(.A(n6237), .B(dpath_mulcore_b7[0]), .Y(n10809));
AND2X1 mul_U1965(.A(n172), .B(n10818), .Y(dpath_mulcore_ary1_a0_I2_I1_29__net32));
OR2X1 mul_U1966(.A(n6240), .B(dpath_mulcore_b6[0]), .Y(n10818));
AND2X1 mul_U1967(.A(n171), .B(n10815), .Y(dpath_mulcore_ary1_a0_I2_I1_29__net046));
OR2X1 mul_U1968(.A(n6239), .B(dpath_mulcore_b7[0]), .Y(n10815));
AND2X1 mul_U1969(.A(n174), .B(n10824), .Y(dpath_mulcore_ary1_a0_I2_I1_28__net32));
OR2X1 mul_U1970(.A(n6242), .B(dpath_mulcore_b6[0]), .Y(n10824));
AND2X1 mul_U1971(.A(n173), .B(n10821), .Y(dpath_mulcore_ary1_a0_I2_I1_28__net046));
OR2X1 mul_U1972(.A(n6241), .B(dpath_mulcore_b7[0]), .Y(n10821));
AND2X1 mul_U1973(.A(n176), .B(n10830), .Y(dpath_mulcore_ary1_a0_I2_I1_27__net32));
OR2X1 mul_U1974(.A(n6244), .B(dpath_mulcore_b6[0]), .Y(n10830));
AND2X1 mul_U1975(.A(n175), .B(n10827), .Y(dpath_mulcore_ary1_a0_I2_I1_27__net046));
OR2X1 mul_U1976(.A(n6243), .B(dpath_mulcore_b7[0]), .Y(n10827));
AND2X1 mul_U1977(.A(n178), .B(n10836), .Y(dpath_mulcore_ary1_a0_I2_I1_26__net32));
OR2X1 mul_U1978(.A(n6246), .B(dpath_mulcore_b6[0]), .Y(n10836));
AND2X1 mul_U1979(.A(n177), .B(n10833), .Y(dpath_mulcore_ary1_a0_I2_I1_26__net046));
OR2X1 mul_U1980(.A(n6245), .B(dpath_mulcore_b7[0]), .Y(n10833));
AND2X1 mul_U1981(.A(n180), .B(n10842), .Y(dpath_mulcore_ary1_a0_I2_I1_25__net32));
OR2X1 mul_U1982(.A(n6248), .B(dpath_mulcore_b6[0]), .Y(n10842));
AND2X1 mul_U1983(.A(n179), .B(n10839), .Y(dpath_mulcore_ary1_a0_I2_I1_25__net046));
OR2X1 mul_U1984(.A(n6247), .B(dpath_mulcore_b7[0]), .Y(n10839));
AND2X1 mul_U1985(.A(n182), .B(n10848), .Y(dpath_mulcore_ary1_a0_I2_I1_24__net32));
OR2X1 mul_U1986(.A(n6250), .B(dpath_mulcore_b6[0]), .Y(n10848));
AND2X1 mul_U1987(.A(n181), .B(n10845), .Y(dpath_mulcore_ary1_a0_I2_I1_24__net046));
OR2X1 mul_U1988(.A(n6249), .B(dpath_mulcore_b7[0]), .Y(n10845));
AND2X1 mul_U1989(.A(n184), .B(n10854), .Y(dpath_mulcore_ary1_a0_I2_I1_23__net32));
OR2X1 mul_U1990(.A(n6252), .B(dpath_mulcore_b6[0]), .Y(n10854));
AND2X1 mul_U1991(.A(n183), .B(n10851), .Y(dpath_mulcore_ary1_a0_I2_I1_23__net046));
OR2X1 mul_U1992(.A(n6251), .B(dpath_mulcore_b7[0]), .Y(n10851));
AND2X1 mul_U1993(.A(n186), .B(n10860), .Y(dpath_mulcore_ary1_a0_I2_I1_22__net32));
OR2X1 mul_U1994(.A(n6254), .B(dpath_mulcore_b6[0]), .Y(n10860));
AND2X1 mul_U1995(.A(n185), .B(n10857), .Y(dpath_mulcore_ary1_a0_I2_I1_22__net046));
OR2X1 mul_U1996(.A(n6253), .B(dpath_mulcore_b7[0]), .Y(n10857));
AND2X1 mul_U1997(.A(n188), .B(n10866), .Y(dpath_mulcore_ary1_a0_I2_I1_21__net32));
OR2X1 mul_U1998(.A(n6256), .B(dpath_mulcore_b6[0]), .Y(n10866));
AND2X1 mul_U1999(.A(n187), .B(n10863), .Y(dpath_mulcore_ary1_a0_I2_I1_21__net046));
OR2X1 mul_U2000(.A(n6255), .B(dpath_mulcore_b7[0]), .Y(n10863));
AND2X1 mul_U2001(.A(n190), .B(n10872), .Y(dpath_mulcore_ary1_a0_I2_I1_20__net32));
OR2X1 mul_U2002(.A(n6258), .B(dpath_mulcore_b6[0]), .Y(n10872));
AND2X1 mul_U2003(.A(n189), .B(n10869), .Y(dpath_mulcore_ary1_a0_I2_I1_20__net046));
OR2X1 mul_U2004(.A(n6257), .B(dpath_mulcore_b7[0]), .Y(n10869));
AND2X1 mul_U2005(.A(n192), .B(n10878), .Y(dpath_mulcore_ary1_a0_I2_I1_19__net32));
OR2X1 mul_U2006(.A(n6260), .B(dpath_mulcore_b6[0]), .Y(n10878));
AND2X1 mul_U2007(.A(n191), .B(n10875), .Y(dpath_mulcore_ary1_a0_I2_I1_19__net046));
OR2X1 mul_U2008(.A(n6259), .B(dpath_mulcore_b7[0]), .Y(n10875));
AND2X1 mul_U2009(.A(n194), .B(n10884), .Y(dpath_mulcore_ary1_a0_I2_I1_18__net32));
OR2X1 mul_U2010(.A(n6262), .B(dpath_mulcore_b6[0]), .Y(n10884));
AND2X1 mul_U2011(.A(n193), .B(n10881), .Y(dpath_mulcore_ary1_a0_I2_I1_18__net046));
OR2X1 mul_U2012(.A(n6261), .B(dpath_mulcore_b7[0]), .Y(n10881));
AND2X1 mul_U2013(.A(n196), .B(n10890), .Y(dpath_mulcore_ary1_a0_I2_I1_17__net32));
OR2X1 mul_U2014(.A(n6264), .B(dpath_mulcore_b6[0]), .Y(n10890));
AND2X1 mul_U2015(.A(n195), .B(n10887), .Y(dpath_mulcore_ary1_a0_I2_I1_17__net046));
OR2X1 mul_U2016(.A(n6263), .B(dpath_mulcore_b7[0]), .Y(n10887));
AND2X1 mul_U2017(.A(n198), .B(n10896), .Y(dpath_mulcore_ary1_a0_I2_I1_16__net32));
OR2X1 mul_U2018(.A(n6266), .B(dpath_mulcore_b6[0]), .Y(n10896));
AND2X1 mul_U2019(.A(n197), .B(n10893), .Y(dpath_mulcore_ary1_a0_I2_I1_16__net046));
OR2X1 mul_U2020(.A(n6265), .B(dpath_mulcore_b7[0]), .Y(n10893));
AND2X1 mul_U2021(.A(n200), .B(n10902), .Y(dpath_mulcore_ary1_a0_I2_I1_15__net32));
OR2X1 mul_U2022(.A(n6268), .B(dpath_mulcore_b6[0]), .Y(n10902));
AND2X1 mul_U2023(.A(n199), .B(n10899), .Y(dpath_mulcore_ary1_a0_I2_I1_15__net046));
OR2X1 mul_U2024(.A(n6267), .B(dpath_mulcore_b7[0]), .Y(n10899));
AND2X1 mul_U2025(.A(n202), .B(n10908), .Y(dpath_mulcore_ary1_a0_I2_I1_14__net32));
OR2X1 mul_U2026(.A(n6270), .B(dpath_mulcore_b6[0]), .Y(n10908));
AND2X1 mul_U2027(.A(n201), .B(n10905), .Y(dpath_mulcore_ary1_a0_I2_I1_14__net046));
OR2X1 mul_U2028(.A(n6269), .B(dpath_mulcore_b7[0]), .Y(n10905));
AND2X1 mul_U2029(.A(n204), .B(n10914), .Y(dpath_mulcore_ary1_a0_I2_I1_13__net32));
OR2X1 mul_U2030(.A(n6272), .B(dpath_mulcore_b6[0]), .Y(n10914));
AND2X1 mul_U2031(.A(n203), .B(n10911), .Y(dpath_mulcore_ary1_a0_I2_I1_13__net046));
OR2X1 mul_U2032(.A(n6271), .B(dpath_mulcore_b7[0]), .Y(n10911));
AND2X1 mul_U2033(.A(n206), .B(n10920), .Y(dpath_mulcore_ary1_a0_I2_I1_12__net32));
OR2X1 mul_U2034(.A(n6274), .B(dpath_mulcore_b6[0]), .Y(n10920));
AND2X1 mul_U2035(.A(n205), .B(n10917), .Y(dpath_mulcore_ary1_a0_I2_I1_12__net046));
OR2X1 mul_U2036(.A(n6273), .B(dpath_mulcore_b7[0]), .Y(n10917));
AND2X1 mul_U2037(.A(n208), .B(n10926), .Y(dpath_mulcore_ary1_a0_I2_I1_11__net32));
OR2X1 mul_U2038(.A(n6276), .B(dpath_mulcore_b6[0]), .Y(n10926));
AND2X1 mul_U2039(.A(n207), .B(n10923), .Y(dpath_mulcore_ary1_a0_I2_I1_11__net046));
OR2X1 mul_U2040(.A(n6275), .B(dpath_mulcore_b7[0]), .Y(n10923));
AND2X1 mul_U2041(.A(n210), .B(n10932), .Y(dpath_mulcore_ary1_a0_I2_I1_10__net32));
OR2X1 mul_U2042(.A(n6278), .B(dpath_mulcore_b6[0]), .Y(n10932));
AND2X1 mul_U2043(.A(n209), .B(n10929), .Y(dpath_mulcore_ary1_a0_I2_I1_10__net046));
OR2X1 mul_U2044(.A(n6277), .B(dpath_mulcore_b7[0]), .Y(n10929));
AND2X1 mul_U2045(.A(n212), .B(n10938), .Y(dpath_mulcore_ary1_a0_I2_I1_9__net32));
OR2X1 mul_U2046(.A(n6280), .B(dpath_mulcore_b6[0]), .Y(n10938));
AND2X1 mul_U2047(.A(n211), .B(n10935), .Y(dpath_mulcore_ary1_a0_I2_I1_9__net046));
OR2X1 mul_U2048(.A(n6279), .B(dpath_mulcore_b7[0]), .Y(n10935));
AND2X1 mul_U2049(.A(n214), .B(n10944), .Y(dpath_mulcore_ary1_a0_I2_I1_8__net32));
OR2X1 mul_U2050(.A(n6282), .B(dpath_mulcore_b6[0]), .Y(n10944));
AND2X1 mul_U2051(.A(n213), .B(n10941), .Y(dpath_mulcore_ary1_a0_I2_I1_8__net046));
OR2X1 mul_U2052(.A(n6281), .B(dpath_mulcore_b7[0]), .Y(n10941));
AND2X1 mul_U2053(.A(n216), .B(n10950), .Y(dpath_mulcore_ary1_a0_I2_I1_7__net32));
OR2X1 mul_U2054(.A(n6284), .B(dpath_mulcore_b6[0]), .Y(n10950));
AND2X1 mul_U2055(.A(n215), .B(n10947), .Y(dpath_mulcore_ary1_a0_I2_I1_7__net046));
OR2X1 mul_U2056(.A(n6283), .B(dpath_mulcore_b7[0]), .Y(n10947));
AND2X1 mul_U2057(.A(n218), .B(n10956), .Y(dpath_mulcore_ary1_a0_I2_I1_6__net32));
OR2X1 mul_U2058(.A(n6286), .B(dpath_mulcore_b6[0]), .Y(n10956));
AND2X1 mul_U2059(.A(n217), .B(n10953), .Y(dpath_mulcore_ary1_a0_I2_I1_6__net046));
OR2X1 mul_U2060(.A(n6285), .B(dpath_mulcore_b7[0]), .Y(n10953));
AND2X1 mul_U2061(.A(n220), .B(n10962), .Y(dpath_mulcore_ary1_a0_I2_I1_5__net32));
OR2X1 mul_U2062(.A(n6288), .B(dpath_mulcore_b6[0]), .Y(n10962));
AND2X1 mul_U2063(.A(n219), .B(n10959), .Y(dpath_mulcore_ary1_a0_I2_I1_5__net046));
OR2X1 mul_U2064(.A(n6287), .B(dpath_mulcore_b7[0]), .Y(n10959));
AND2X1 mul_U2065(.A(n222), .B(n10968), .Y(dpath_mulcore_ary1_a0_I2_I1_4__net32));
OR2X1 mul_U2066(.A(n6290), .B(dpath_mulcore_b6[0]), .Y(n10968));
AND2X1 mul_U2067(.A(n221), .B(n10965), .Y(dpath_mulcore_ary1_a0_I2_I1_4__net046));
OR2X1 mul_U2068(.A(n6289), .B(dpath_mulcore_b7[0]), .Y(n10965));
OR2X1 mul_U2069(.A(n9735), .B(n5956), .Y(dpath_mulcore_ary1_a0_I2_I0_b1n_1));
OR2X1 mul_U2070(.A(n9735), .B(n5957), .Y(dpath_mulcore_ary1_a0_I2_I0_b1n_0));
AND2X1 mul_U2071(.A(n401), .B(n11509), .Y(dpath_mulcore_ary1_a0_I1_I1_7__net043));
OR2X1 mul_U2072(.A(n6471), .B(dpath_mulcore_b5[0]), .Y(n11509));
AND2X1 mul_U2073(.A(n226), .B(n10980), .Y(dpath_mulcore_ary1_a0_I2_I0_p0_1));
OR2X1 mul_U2074(.A(n6294), .B(dpath_mulcore_b6[0]), .Y(n10980));
OR2X1 mul_U2075(.A(dpath_mulcore_ary1_a0_I2_I0_n1), .B(n5954), .Y(dpath_mulcore_ary1_a0_I2_I0_b0n));
AND2X1 mul_U2076(.A(n7416), .B(n9854), .Y(dpath_mulcore_ary1_a0_I2_I0_n1));
AND2X1 mul_U2077(.A(n404), .B(n11518), .Y(dpath_mulcore_ary1_a0_I1_I1_6__net043));
OR2X1 mul_U2078(.A(n6474), .B(dpath_mulcore_b5[0]), .Y(n11518));
INVX1 mul_U2079(.A(n10982), .Y(n9854));
OR2X1 mul_U2080(.A(n6295), .B(dpath_mulcore_b6[0]), .Y(n10982));
OR2X1 mul_U2081(.A(n9733), .B(n5955), .Y(dpath_mulcore_ary1_a0_I2_I0_b0n_0));
AND2X1 mul_U2082(.A(n580), .B(n12052), .Y(dpath_mulcore_ary1_a0_I0_I1_11__net32));
OR2X1 mul_U2083(.A(n6653), .B(dpath_mulcore_b0[0]), .Y(n12052));
AND2X1 mul_U2084(.A(n579), .B(n12049), .Y(dpath_mulcore_ary1_a0_I0_I1_11__net046));
OR2X1 mul_U2085(.A(n6652), .B(dpath_mulcore_b1[0]), .Y(n12049));
AND2X1 mul_U2086(.A(n407), .B(n11527), .Y(dpath_mulcore_ary1_a0_I1_I1_5__net043));
OR2X1 mul_U2087(.A(n6477), .B(dpath_mulcore_b5[0]), .Y(n11527));
AND2X1 mul_U2088(.A(n411), .B(n11541), .Y(dpath_mulcore_ary1_a0_I1_I1_4__net32));
OR2X1 mul_U2089(.A(n6482), .B(dpath_mulcore_b3[0]), .Y(n11541));
AND2X1 mul_U2090(.A(n410), .B(n11538), .Y(dpath_mulcore_ary1_a0_I1_I1_4__net046));
OR2X1 mul_U2091(.A(n6481), .B(dpath_mulcore_b4[0]), .Y(n11538));
AND2X1 mul_U2092(.A(n583), .B(n12061), .Y(dpath_mulcore_ary1_a0_I0_I1_10__net32));
OR2X1 mul_U2093(.A(n6656), .B(dpath_mulcore_b0[0]), .Y(n12061));
AND2X1 mul_U2094(.A(n582), .B(n12058), .Y(dpath_mulcore_ary1_a0_I0_I1_10__net046));
OR2X1 mul_U2095(.A(n6655), .B(dpath_mulcore_b1[0]), .Y(n12058));
AND2X1 mul_U2096(.A(n586), .B(n12070), .Y(dpath_mulcore_ary1_a0_I0_I1_9__net32));
OR2X1 mul_U2097(.A(n6659), .B(dpath_mulcore_b0[0]), .Y(n12070));
AND2X1 mul_U2098(.A(n585), .B(n12067), .Y(dpath_mulcore_ary1_a0_I0_I1_9__net046));
OR2X1 mul_U2099(.A(n6658), .B(dpath_mulcore_b1[0]), .Y(n12067));
AND2X1 mul_U2100(.A(n584), .B(n12064), .Y(dpath_mulcore_ary1_a0_I0_I1_9__net043));
OR2X1 mul_U2101(.A(n6657), .B(dpath_mulcore_b2[0]), .Y(n12064));
AND2X1 mul_U2102(.A(n587), .B(n12073), .Y(dpath_mulcore_ary1_a0_I0_I1_8__net043));
OR2X1 mul_U2103(.A(n6660), .B(dpath_mulcore_b2[0]), .Y(n12073));
AND2X1 mul_U2104(.A(n592), .B(n12088), .Y(dpath_mulcore_ary1_a0_I0_I1_7__net32));
OR2X1 mul_U2105(.A(n6665), .B(dpath_mulcore_b0[0]), .Y(n12088));
AND2X1 mul_U2106(.A(n591), .B(n12085), .Y(dpath_mulcore_ary1_a0_I0_I1_7__net046));
OR2X1 mul_U2107(.A(n6664), .B(dpath_mulcore_b1[0]), .Y(n12085));
AND2X1 mul_U2108(.A(n595), .B(n12097), .Y(dpath_mulcore_ary1_a0_I0_I1_6__net32));
OR2X1 mul_U2109(.A(n6668), .B(dpath_mulcore_b0[0]), .Y(n12097));
AND2X1 mul_U2110(.A(n594), .B(n12094), .Y(dpath_mulcore_ary1_a0_I0_I1_6__net046));
OR2X1 mul_U2111(.A(n6667), .B(dpath_mulcore_b1[0]), .Y(n12094));
AND2X1 mul_U2112(.A(n598), .B(n12106), .Y(dpath_mulcore_ary1_a0_I0_I1_5__net32));
OR2X1 mul_U2113(.A(n6671), .B(dpath_mulcore_b0[0]), .Y(n12106));
AND2X1 mul_U2114(.A(n597), .B(n12103), .Y(dpath_mulcore_ary1_a0_I0_I1_5__net046));
OR2X1 mul_U2115(.A(n6670), .B(dpath_mulcore_b1[0]), .Y(n12103));
AND2X1 mul_U2116(.A(n600), .B(n12114), .Y(dpath_mulcore_ary1_a0_I0_I1_4__net32));
OR2X1 mul_U2117(.A(n6674), .B(dpath_mulcore_b0[0]), .Y(n12114));
AND2X1 mul_U2118(.A(n599), .B(n12111), .Y(dpath_mulcore_ary1_a0_I0_I1_4__net046));
OR2X1 mul_U2119(.A(n6673), .B(dpath_mulcore_b1[0]), .Y(n12111));
AND2X1 mul_U2120(.A(n2833), .B(n4509), .Y(dpath_n387));
AND2X1 mul_U2121(.A(n2789), .B(n4465), .Y(dpath_n255));
AND2X1 mul_U2122(.A(n2757), .B(n4433), .Y(dpath_n159));
AND2X1 mul_U2123(.A(n2753), .B(n4429), .Y(dpath_n147));
AND2X1 mul_U2124(.A(n2875), .B(n4551), .Y(dpath_n513));
AND2X1 mul_U2125(.A(n2871), .B(n4547), .Y(dpath_n501));
AND2X1 mul_U2126(.A(n2867), .B(n4543), .Y(dpath_n489));
AND2X1 mul_U2127(.A(n2863), .B(n4539), .Y(dpath_n477));
AND2X1 mul_U2128(.A(n2859), .B(n4535), .Y(dpath_n465));
AND2X1 mul_U2129(.A(n2853), .B(n4529), .Y(dpath_n447));
AND2X1 mul_U2130(.A(n2849), .B(n4525), .Y(dpath_n435));
AND2X1 mul_U2131(.A(n2845), .B(n4521), .Y(dpath_n423));
AND2X1 mul_U2132(.A(n2841), .B(n4517), .Y(dpath_n411));
AND2X1 mul_U2133(.A(n2837), .B(n4513), .Y(dpath_n399));
AND2X1 mul_U2134(.A(n2831), .B(n4507), .Y(dpath_n381));
INVX1 mul_U2135(.A(dpath_mulcore_op1_l[60]), .Y(n10029));
AND2X1 mul_U2136(.A(n608), .B(n12142), .Y(dpath_mulcore_ary1_a1_I2_I1_63__net32));
OR2X1 mul_U2137(.A(n6684), .B(dpath_mulcore_b14[0]), .Y(n12142));
AND2X1 mul_U2138(.A(n607), .B(n12139), .Y(dpath_mulcore_ary1_a1_I2_I1_63__net046));
OR2X1 mul_U2139(.A(n6683), .B(dpath_mulcore_b15[0]), .Y(n12139));
AND2X1 mul_U2140(.A(n1118), .B(n13679), .Y(dpath_mulcore_ary1_a1_I1_I2_net47));
OR2X1 mul_U2141(.A(n9479), .B(dpath_mulcore_b11[0]), .Y(n13679));
AND2X1 mul_U2142(.A(n735), .B(n12527), .Y(dpath_mulcore_ary1_a1_I1_I2_net48));
OR2X1 mul_U2143(.A(n6813), .B(dpath_mulcore_b12[0]), .Y(n12527));
AND2X1 mul_U2144(.A(n734), .B(n12524), .Y(dpath_mulcore_ary1_a1_I1_I2_net43));
OR2X1 mul_U2145(.A(n6812), .B(dpath_mulcore_b12[0]), .Y(n12524));
AND2X1 mul_U2146(.A(n737), .B(n12533), .Y(dpath_mulcore_ary1_a1_I1_I1_63__net043));
OR2X1 mul_U2147(.A(n6815), .B(dpath_mulcore_b13[0]), .Y(n12533));
OR2X1 mul_U2148(.A(n9427), .B(dpath_mulcore_b10[0]), .Y(n13687));
AND2X1 mul_U2149(.A(n740), .B(n12542), .Y(dpath_mulcore_ary1_a1_I1_I1_62__net043));
OR2X1 mul_U2150(.A(n6818), .B(dpath_mulcore_b13[0]), .Y(n12542));
AND2X1 mul_U2151(.A(dpath_mulcore_ary1_a1_I0_I2_net38), .B(n3507), .Y(dpath_mulcore_ary1_a1_c0[66]));
AND2X1 mul_U2152(.A(n743), .B(n12551), .Y(dpath_mulcore_ary1_a1_I1_I1_61__net043));
OR2X1 mul_U2153(.A(n6821), .B(dpath_mulcore_b13[0]), .Y(n12551));
AND2X1 mul_U2154(.A(n1443), .B(n3506), .Y(dpath_mulcore_ary1_a1_c0[65]));
AND2X1 mul_U2155(.A(n746), .B(n12560), .Y(dpath_mulcore_ary1_a1_I1_I1_60__net043));
OR2X1 mul_U2156(.A(n6824), .B(dpath_mulcore_b13[0]), .Y(n12560));
AND2X1 mul_U2157(.A(n1442), .B(n3505), .Y(dpath_mulcore_ary1_a1_c0[64]));
AND2X1 mul_U2158(.A(n749), .B(n12569), .Y(dpath_mulcore_ary1_a1_I1_I1_59__net043));
OR2X1 mul_U2159(.A(n6827), .B(dpath_mulcore_b13[0]), .Y(n12569));
AND2X1 mul_U2160(.A(n1374), .B(n3435), .Y(dpath_mulcore_ary1_a1_c0[63]));
AND2X1 mul_U2161(.A(n752), .B(n12578), .Y(dpath_mulcore_ary1_a1_I1_I1_58__net043));
OR2X1 mul_U2162(.A(n6830), .B(dpath_mulcore_b13[0]), .Y(n12578));
AND2X1 mul_U2163(.A(n1375), .B(n3436), .Y(dpath_mulcore_ary1_a1_c0[62]));
AND2X1 mul_U2164(.A(n755), .B(n12587), .Y(dpath_mulcore_ary1_a1_I1_I1_57__net043));
OR2X1 mul_U2165(.A(n6833), .B(dpath_mulcore_b13[0]), .Y(n12587));
AND2X1 mul_U2166(.A(n1376), .B(n3437), .Y(dpath_mulcore_ary1_a1_c0[61]));
AND2X1 mul_U2167(.A(n758), .B(n12596), .Y(dpath_mulcore_ary1_a1_I1_I1_56__net043));
OR2X1 mul_U2168(.A(n6836), .B(dpath_mulcore_b13[0]), .Y(n12596));
AND2X1 mul_U2169(.A(n1377), .B(n3438), .Y(dpath_mulcore_ary1_a1_c0[60]));
AND2X1 mul_U2170(.A(n761), .B(n12605), .Y(dpath_mulcore_ary1_a1_I1_I1_55__net043));
OR2X1 mul_U2171(.A(n6839), .B(dpath_mulcore_b13[0]), .Y(n12605));
AND2X1 mul_U2172(.A(n1378), .B(n3439), .Y(dpath_mulcore_ary1_a1_c0[59]));
AND2X1 mul_U2173(.A(n764), .B(n12614), .Y(dpath_mulcore_ary1_a1_I1_I1_54__net043));
OR2X1 mul_U2174(.A(n6842), .B(dpath_mulcore_b13[0]), .Y(n12614));
AND2X1 mul_U2175(.A(n1379), .B(n3440), .Y(dpath_mulcore_ary1_a1_c0[58]));
AND2X1 mul_U2176(.A(n767), .B(n12623), .Y(dpath_mulcore_ary1_a1_I1_I1_53__net043));
OR2X1 mul_U2177(.A(n6845), .B(dpath_mulcore_b13[0]), .Y(n12623));
AND2X1 mul_U2178(.A(n1380), .B(n3441), .Y(dpath_mulcore_ary1_a1_c0[57]));
AND2X1 mul_U2179(.A(n770), .B(n12632), .Y(dpath_mulcore_ary1_a1_I1_I1_52__net043));
OR2X1 mul_U2180(.A(n6848), .B(dpath_mulcore_b13[0]), .Y(n12632));
AND2X1 mul_U2181(.A(n1381), .B(n3442), .Y(dpath_mulcore_ary1_a1_c0[56]));
AND2X1 mul_U2182(.A(n773), .B(n12641), .Y(dpath_mulcore_ary1_a1_I1_I1_51__net043));
OR2X1 mul_U2183(.A(n6851), .B(dpath_mulcore_b13[0]), .Y(n12641));
AND2X1 mul_U2184(.A(n1382), .B(n3443), .Y(dpath_mulcore_ary1_a1_c0[55]));
AND2X1 mul_U2185(.A(n776), .B(n12650), .Y(dpath_mulcore_ary1_a1_I1_I1_50__net043));
OR2X1 mul_U2186(.A(n6854), .B(dpath_mulcore_b13[0]), .Y(n12650));
AND2X1 mul_U2187(.A(n1383), .B(n3444), .Y(dpath_mulcore_ary1_a1_c0[54]));
AND2X1 mul_U2188(.A(n779), .B(n12659), .Y(dpath_mulcore_ary1_a1_I1_I1_49__net043));
OR2X1 mul_U2189(.A(n6857), .B(dpath_mulcore_b13[0]), .Y(n12659));
AND2X1 mul_U2190(.A(n1384), .B(n3445), .Y(dpath_mulcore_ary1_a1_c0[53]));
AND2X1 mul_U2191(.A(n782), .B(n12668), .Y(dpath_mulcore_ary1_a1_I1_I1_48__net043));
OR2X1 mul_U2192(.A(n6860), .B(dpath_mulcore_b13[0]), .Y(n12668));
AND2X1 mul_U2193(.A(n1385), .B(n3446), .Y(dpath_mulcore_ary1_a1_c0[52]));
AND2X1 mul_U2194(.A(n785), .B(n12677), .Y(dpath_mulcore_ary1_a1_I1_I1_47__net043));
OR2X1 mul_U2195(.A(n6863), .B(dpath_mulcore_b13[0]), .Y(n12677));
AND2X1 mul_U2196(.A(n1386), .B(n3447), .Y(dpath_mulcore_ary1_a1_c0[51]));
AND2X1 mul_U2197(.A(n788), .B(n12686), .Y(dpath_mulcore_ary1_a1_I1_I1_46__net043));
OR2X1 mul_U2198(.A(n6866), .B(dpath_mulcore_b13[0]), .Y(n12686));
AND2X1 mul_U2199(.A(n1387), .B(n3448), .Y(dpath_mulcore_ary1_a1_c0[50]));
AND2X1 mul_U2200(.A(n791), .B(n12695), .Y(dpath_mulcore_ary1_a1_I1_I1_45__net043));
OR2X1 mul_U2201(.A(n6869), .B(dpath_mulcore_b13[0]), .Y(n12695));
AND2X1 mul_U2202(.A(n1388), .B(n3449), .Y(dpath_mulcore_ary1_a1_c0[49]));
AND2X1 mul_U2203(.A(n794), .B(n12704), .Y(dpath_mulcore_ary1_a1_I1_I1_44__net043));
OR2X1 mul_U2204(.A(n6872), .B(dpath_mulcore_b13[0]), .Y(n12704));
AND2X1 mul_U2205(.A(n1389), .B(n3450), .Y(dpath_mulcore_ary1_a1_c0[48]));
AND2X1 mul_U2206(.A(n797), .B(n12713), .Y(dpath_mulcore_ary1_a1_I1_I1_43__net043));
OR2X1 mul_U2207(.A(n6875), .B(dpath_mulcore_b13[0]), .Y(n12713));
AND2X1 mul_U2208(.A(n1390), .B(n3451), .Y(dpath_mulcore_ary1_a1_c0[47]));
AND2X1 mul_U2209(.A(n800), .B(n12722), .Y(dpath_mulcore_ary1_a1_I1_I1_42__net043));
OR2X1 mul_U2210(.A(n6878), .B(dpath_mulcore_b13[0]), .Y(n12722));
AND2X1 mul_U2211(.A(n1391), .B(n3452), .Y(dpath_mulcore_ary1_a1_c0[46]));
AND2X1 mul_U2212(.A(n803), .B(n12731), .Y(dpath_mulcore_ary1_a1_I1_I1_41__net043));
OR2X1 mul_U2213(.A(n6881), .B(dpath_mulcore_b13[0]), .Y(n12731));
AND2X1 mul_U2214(.A(n1392), .B(n3453), .Y(dpath_mulcore_ary1_a1_c0[45]));
AND2X1 mul_U2215(.A(n806), .B(n12740), .Y(dpath_mulcore_ary1_a1_I1_I1_40__net043));
OR2X1 mul_U2216(.A(n6884), .B(dpath_mulcore_b13[0]), .Y(n12740));
AND2X1 mul_U2217(.A(n1393), .B(n3454), .Y(dpath_mulcore_ary1_a1_c0[44]));
AND2X1 mul_U2218(.A(n809), .B(n12749), .Y(dpath_mulcore_ary1_a1_I1_I1_39__net043));
OR2X1 mul_U2219(.A(n6887), .B(dpath_mulcore_b13[0]), .Y(n12749));
AND2X1 mul_U2220(.A(n1394), .B(n3455), .Y(dpath_mulcore_ary1_a1_c0[43]));
AND2X1 mul_U2221(.A(n812), .B(n12758), .Y(dpath_mulcore_ary1_a1_I1_I1_38__net043));
OR2X1 mul_U2222(.A(n6890), .B(dpath_mulcore_b13[0]), .Y(n12758));
AND2X1 mul_U2223(.A(n1395), .B(n3456), .Y(dpath_mulcore_ary1_a1_c0[42]));
AND2X1 mul_U2224(.A(n815), .B(n12767), .Y(dpath_mulcore_ary1_a1_I1_I1_37__net043));
OR2X1 mul_U2225(.A(n6893), .B(dpath_mulcore_b13[0]), .Y(n12767));
AND2X1 mul_U2226(.A(n1396), .B(n3457), .Y(dpath_mulcore_ary1_a1_c0[41]));
AND2X1 mul_U2227(.A(n818), .B(n12776), .Y(dpath_mulcore_ary1_a1_I1_I1_36__net043));
OR2X1 mul_U2228(.A(n6896), .B(dpath_mulcore_b13[0]), .Y(n12776));
AND2X1 mul_U2229(.A(n1397), .B(n3458), .Y(dpath_mulcore_ary1_a1_c0[40]));
AND2X1 mul_U2230(.A(n821), .B(n12785), .Y(dpath_mulcore_ary1_a1_I1_I1_35__net043));
OR2X1 mul_U2231(.A(n6899), .B(dpath_mulcore_b13[0]), .Y(n12785));
AND2X1 mul_U2232(.A(n1398), .B(n3459), .Y(dpath_mulcore_ary1_a1_c0[39]));
AND2X1 mul_U2233(.A(n824), .B(n12794), .Y(dpath_mulcore_ary1_a1_I1_I1_34__net043));
OR2X1 mul_U2234(.A(n6902), .B(dpath_mulcore_b13[0]), .Y(n12794));
AND2X1 mul_U2235(.A(n1399), .B(n3460), .Y(dpath_mulcore_ary1_a1_c0[38]));
AND2X1 mul_U2236(.A(n827), .B(n12803), .Y(dpath_mulcore_ary1_a1_I1_I1_33__net043));
OR2X1 mul_U2237(.A(n6905), .B(dpath_mulcore_b13[0]), .Y(n12803));
AND2X1 mul_U2238(.A(n1400), .B(n3461), .Y(dpath_mulcore_ary1_a1_c0[37]));
AND2X1 mul_U2239(.A(n830), .B(n12812), .Y(dpath_mulcore_ary1_a1_I1_I1_32__net043));
OR2X1 mul_U2240(.A(n6908), .B(dpath_mulcore_b13[0]), .Y(n12812));
AND2X1 mul_U2241(.A(n1401), .B(n3462), .Y(dpath_mulcore_ary1_a1_c0[36]));
AND2X1 mul_U2242(.A(n833), .B(n12821), .Y(dpath_mulcore_ary1_a1_I1_I1_31__net043));
OR2X1 mul_U2243(.A(n6911), .B(dpath_mulcore_b13[0]), .Y(n12821));
AND2X1 mul_U2244(.A(n1402), .B(n3463), .Y(dpath_mulcore_ary1_a1_c0[35]));
AND2X1 mul_U2245(.A(n836), .B(n12830), .Y(dpath_mulcore_ary1_a1_I1_I1_30__net043));
OR2X1 mul_U2246(.A(n6914), .B(dpath_mulcore_b13[0]), .Y(n12830));
AND2X1 mul_U2247(.A(n1403), .B(n3464), .Y(dpath_mulcore_ary1_a1_c0[34]));
AND2X1 mul_U2248(.A(n839), .B(n12839), .Y(dpath_mulcore_ary1_a1_I1_I1_29__net043));
OR2X1 mul_U2249(.A(n6917), .B(dpath_mulcore_b13[0]), .Y(n12839));
AND2X1 mul_U2250(.A(n1404), .B(n3465), .Y(dpath_mulcore_ary1_a1_c0[33]));
AND2X1 mul_U2251(.A(n842), .B(n12848), .Y(dpath_mulcore_ary1_a1_I1_I1_28__net043));
OR2X1 mul_U2252(.A(n6920), .B(dpath_mulcore_b13[0]), .Y(n12848));
AND2X1 mul_U2253(.A(n1405), .B(n3466), .Y(dpath_mulcore_ary1_a1_c0[32]));
AND2X1 mul_U2254(.A(n845), .B(n12857), .Y(dpath_mulcore_ary1_a1_I1_I1_27__net043));
OR2X1 mul_U2255(.A(n6923), .B(dpath_mulcore_b13[0]), .Y(n12857));
AND2X1 mul_U2256(.A(n1406), .B(n3467), .Y(dpath_mulcore_ary1_a1_c0[31]));
AND2X1 mul_U2257(.A(n848), .B(n12866), .Y(dpath_mulcore_ary1_a1_I1_I1_26__net043));
OR2X1 mul_U2258(.A(n6926), .B(dpath_mulcore_b13[0]), .Y(n12866));
AND2X1 mul_U2259(.A(n1407), .B(n3468), .Y(dpath_mulcore_ary1_a1_c0[30]));
AND2X1 mul_U2260(.A(n851), .B(n12875), .Y(dpath_mulcore_ary1_a1_I1_I1_25__net043));
OR2X1 mul_U2261(.A(n6929), .B(dpath_mulcore_b13[0]), .Y(n12875));
AND2X1 mul_U2262(.A(n1408), .B(n3469), .Y(dpath_mulcore_ary1_a1_c0[29]));
AND2X1 mul_U2263(.A(n854), .B(n12884), .Y(dpath_mulcore_ary1_a1_I1_I1_24__net043));
OR2X1 mul_U2264(.A(n6932), .B(dpath_mulcore_b13[0]), .Y(n12884));
AND2X1 mul_U2265(.A(n1409), .B(n3470), .Y(dpath_mulcore_ary1_a1_c0[28]));
AND2X1 mul_U2266(.A(n857), .B(n12893), .Y(dpath_mulcore_ary1_a1_I1_I1_23__net043));
OR2X1 mul_U2267(.A(n6935), .B(dpath_mulcore_b13[0]), .Y(n12893));
AND2X1 mul_U2268(.A(n1410), .B(n3471), .Y(dpath_mulcore_ary1_a1_c0[27]));
AND2X1 mul_U2269(.A(n860), .B(n12902), .Y(dpath_mulcore_ary1_a1_I1_I1_22__net043));
OR2X1 mul_U2270(.A(n6938), .B(dpath_mulcore_b13[0]), .Y(n12902));
AND2X1 mul_U2271(.A(n1411), .B(n3472), .Y(dpath_mulcore_ary1_a1_c0[26]));
AND2X1 mul_U2272(.A(n863), .B(n12911), .Y(dpath_mulcore_ary1_a1_I1_I1_21__net043));
OR2X1 mul_U2273(.A(n6941), .B(dpath_mulcore_b13[0]), .Y(n12911));
AND2X1 mul_U2274(.A(n1412), .B(n3473), .Y(dpath_mulcore_ary1_a1_c0[25]));
AND2X1 mul_U2275(.A(n866), .B(n12920), .Y(dpath_mulcore_ary1_a1_I1_I1_20__net043));
OR2X1 mul_U2276(.A(n6944), .B(dpath_mulcore_b13[0]), .Y(n12920));
AND2X1 mul_U2277(.A(n1413), .B(n3474), .Y(dpath_mulcore_ary1_a1_c0[24]));
AND2X1 mul_U2278(.A(n869), .B(n12929), .Y(dpath_mulcore_ary1_a1_I1_I1_19__net043));
OR2X1 mul_U2279(.A(n6947), .B(dpath_mulcore_b13[0]), .Y(n12929));
AND2X1 mul_U2280(.A(n1414), .B(n3475), .Y(dpath_mulcore_ary1_a1_c0[23]));
AND2X1 mul_U2281(.A(n872), .B(n12938), .Y(dpath_mulcore_ary1_a1_I1_I1_18__net043));
OR2X1 mul_U2282(.A(n6950), .B(dpath_mulcore_b13[0]), .Y(n12938));
AND2X1 mul_U2283(.A(n1415), .B(n3476), .Y(dpath_mulcore_ary1_a1_c0[22]));
AND2X1 mul_U2284(.A(n875), .B(n12947), .Y(dpath_mulcore_ary1_a1_I1_I1_17__net043));
OR2X1 mul_U2285(.A(n6953), .B(dpath_mulcore_b13[0]), .Y(n12947));
AND2X1 mul_U2286(.A(n1416), .B(n3477), .Y(dpath_mulcore_ary1_a1_c0[21]));
AND2X1 mul_U2287(.A(n878), .B(n12956), .Y(dpath_mulcore_ary1_a1_I1_I1_16__net043));
OR2X1 mul_U2288(.A(n6956), .B(dpath_mulcore_b13[0]), .Y(n12956));
AND2X1 mul_U2289(.A(n1417), .B(n3478), .Y(dpath_mulcore_ary1_a1_c0[20]));
AND2X1 mul_U2290(.A(n881), .B(n12965), .Y(dpath_mulcore_ary1_a1_I1_I1_15__net043));
OR2X1 mul_U2291(.A(n6959), .B(dpath_mulcore_b13[0]), .Y(n12965));
AND2X1 mul_U2292(.A(n1418), .B(n3479), .Y(dpath_mulcore_ary1_a1_c0[19]));
AND2X1 mul_U2293(.A(n884), .B(n12974), .Y(dpath_mulcore_ary1_a1_I1_I1_14__net043));
OR2X1 mul_U2294(.A(n6962), .B(dpath_mulcore_b13[0]), .Y(n12974));
AND2X1 mul_U2295(.A(n1419), .B(n3480), .Y(dpath_mulcore_ary1_a1_c0[18]));
AND2X1 mul_U2296(.A(n887), .B(n12983), .Y(dpath_mulcore_ary1_a1_I1_I1_13__net043));
OR2X1 mul_U2297(.A(n6965), .B(dpath_mulcore_b13[0]), .Y(n12983));
AND2X1 mul_U2298(.A(n1420), .B(n3481), .Y(dpath_mulcore_ary1_a1_c0[17]));
AND2X1 mul_U2299(.A(n890), .B(n12992), .Y(dpath_mulcore_ary1_a1_I1_I1_12__net043));
OR2X1 mul_U2300(.A(n6968), .B(dpath_mulcore_b13[0]), .Y(n12992));
AND2X1 mul_U2301(.A(n1421), .B(n3482), .Y(dpath_mulcore_ary1_a1_c0[16]));
AND2X1 mul_U2302(.A(n893), .B(n13001), .Y(dpath_mulcore_ary1_a1_I1_I1_11__net043));
OR2X1 mul_U2303(.A(n6971), .B(dpath_mulcore_b13[0]), .Y(n13001));
AND2X1 mul_U2304(.A(n1422), .B(n3483), .Y(dpath_mulcore_ary1_a1_c0[15]));
AND2X1 mul_U2305(.A(n896), .B(n13010), .Y(dpath_mulcore_ary1_a1_I1_I1_10__net043));
OR2X1 mul_U2306(.A(n6974), .B(dpath_mulcore_b13[0]), .Y(n13010));
AND2X1 mul_U2307(.A(n1423), .B(n3484), .Y(dpath_mulcore_ary1_a1_c0[14]));
AND2X1 mul_U2308(.A(n899), .B(n13019), .Y(dpath_mulcore_ary1_a1_I1_I1_9__net043));
OR2X1 mul_U2309(.A(n6977), .B(dpath_mulcore_b13[0]), .Y(n13019));
AND2X1 mul_U2310(.A(n1424), .B(n3485), .Y(dpath_mulcore_ary1_a1_c0[13]));
AND2X1 mul_U2311(.A(n902), .B(n13028), .Y(dpath_mulcore_ary1_a1_I1_I1_8__net043));
OR2X1 mul_U2312(.A(n6980), .B(dpath_mulcore_b13[0]), .Y(n13028));
AND2X1 mul_U2313(.A(n1076), .B(n13556), .Y(dpath_mulcore_ary1_a1_I0_I1_13__net043));
OR2X1 mul_U2314(.A(n7157), .B(dpath_mulcore_b10[0]), .Y(n13556));
AND2X1 mul_U2315(.A(n1079), .B(n13565), .Y(dpath_mulcore_ary1_a1_I0_I1_12__net043));
OR2X1 mul_U2316(.A(n7160), .B(dpath_mulcore_b10[0]), .Y(n13565));
AND2X1 mul_U2317(.A(n917), .B(n13075), .Y(dpath_mulcore_ary1_a1_I1_I0_p1_3));
OR2X1 mul_U2318(.A(n6996), .B(dpath_mulcore_b12[0]), .Y(n13075));
AND2X1 mul_U2319(.A(n916), .B(n13072), .Y(dpath_mulcore_ary1_a1_I1_I0_p0_3));
OR2X1 mul_U2320(.A(n6995), .B(dpath_mulcore_b11[0]), .Y(n13072));
AND2X1 mul_U2321(.A(n1106), .B(n13648), .Y(dpath_mulcore_ary1_a1_I0_I0_p1_3));
OR2X1 mul_U2322(.A(n7188), .B(dpath_mulcore_b9[0]), .Y(n13648));
AND2X1 mul_U2323(.A(n1105), .B(n13645), .Y(dpath_mulcore_ary1_a1_I0_I0_p0_3));
OR2X1 mul_U2324(.A(n7187), .B(dpath_mulcore_b8[0]), .Y(n13645));
INVX1 mul_U2325(.A(dpath_mulcore_op1_l[61]), .Y(n10030));
AND2X1 mul_U2326(.A(n1116), .B(n13675), .Y(dpath_mulcore_ary1_a1_I2_I2_net47));
OR2X1 mul_U2327(.A(n9477), .B(dpath_mulcore_b14[0]), .Y(n13675));
AND2X1 mul_U2328(.A(n606), .B(n12136), .Y(dpath_mulcore_ary1_a1_I2_I2_net48));
OR2X1 mul_U2329(.A(n6682), .B(dpath_mulcore_b15[0]), .Y(n12136));
AND2X1 mul_U2330(.A(n1255), .B(n3316), .Y(dpath_mulcore_ary1_a1_c2[62]));
AND2X1 mul_U2331(.A(n1256), .B(n3317), .Y(dpath_mulcore_ary1_a1_c2[61]));
AND2X1 mul_U2332(.A(n1257), .B(n3318), .Y(dpath_mulcore_ary1_a1_c2[60]));
AND2X1 mul_U2333(.A(n1258), .B(n3319), .Y(dpath_mulcore_ary1_a1_c2[59]));
AND2X1 mul_U2334(.A(n1259), .B(n3320), .Y(dpath_mulcore_ary1_a1_c2[58]));
AND2X1 mul_U2335(.A(n1260), .B(n3321), .Y(dpath_mulcore_ary1_a1_c2[57]));
AND2X1 mul_U2336(.A(n1261), .B(n3322), .Y(dpath_mulcore_ary1_a1_c2[56]));
AND2X1 mul_U2337(.A(n1262), .B(n3323), .Y(dpath_mulcore_ary1_a1_c2[55]));
AND2X1 mul_U2338(.A(n1263), .B(n3324), .Y(dpath_mulcore_ary1_a1_c2[54]));
AND2X1 mul_U2339(.A(n1264), .B(n3325), .Y(dpath_mulcore_ary1_a1_c2[53]));
AND2X1 mul_U2340(.A(n1265), .B(n3326), .Y(dpath_mulcore_ary1_a1_c2[52]));
AND2X1 mul_U2341(.A(n1266), .B(n3327), .Y(dpath_mulcore_ary1_a1_c2[51]));
AND2X1 mul_U2342(.A(n1267), .B(n3328), .Y(dpath_mulcore_ary1_a1_c2[50]));
AND2X1 mul_U2343(.A(n1268), .B(n3329), .Y(dpath_mulcore_ary1_a1_c2[49]));
AND2X1 mul_U2344(.A(n1269), .B(n3330), .Y(dpath_mulcore_ary1_a1_c2[48]));
AND2X1 mul_U2345(.A(n1270), .B(n3331), .Y(dpath_mulcore_ary1_a1_c2[47]));
AND2X1 mul_U2346(.A(n1271), .B(n3332), .Y(dpath_mulcore_ary1_a1_c2[46]));
AND2X1 mul_U2347(.A(n1272), .B(n3333), .Y(dpath_mulcore_ary1_a1_c2[45]));
AND2X1 mul_U2348(.A(n1273), .B(n3334), .Y(dpath_mulcore_ary1_a1_c2[44]));
AND2X1 mul_U2349(.A(n1274), .B(n3335), .Y(dpath_mulcore_ary1_a1_c2[43]));
AND2X1 mul_U2350(.A(n1275), .B(n3336), .Y(dpath_mulcore_ary1_a1_c2[42]));
AND2X1 mul_U2351(.A(n1276), .B(n3337), .Y(dpath_mulcore_ary1_a1_c2[41]));
AND2X1 mul_U2352(.A(n1277), .B(n3338), .Y(dpath_mulcore_ary1_a1_c2[40]));
AND2X1 mul_U2353(.A(n1278), .B(n3339), .Y(dpath_mulcore_ary1_a1_c2[39]));
AND2X1 mul_U2354(.A(n1279), .B(n3340), .Y(dpath_mulcore_ary1_a1_c2[38]));
AND2X1 mul_U2355(.A(n1280), .B(n3341), .Y(dpath_mulcore_ary1_a1_c2[37]));
AND2X1 mul_U2356(.A(n1281), .B(n3342), .Y(dpath_mulcore_ary1_a1_c2[36]));
AND2X1 mul_U2357(.A(n1282), .B(n3343), .Y(dpath_mulcore_ary1_a1_c2[35]));
AND2X1 mul_U2358(.A(n1283), .B(n3344), .Y(dpath_mulcore_ary1_a1_c2[34]));
AND2X1 mul_U2359(.A(n1284), .B(n3345), .Y(dpath_mulcore_ary1_a1_c2[33]));
AND2X1 mul_U2360(.A(n1285), .B(n3346), .Y(dpath_mulcore_ary1_a1_c2[32]));
AND2X1 mul_U2361(.A(n1286), .B(n3347), .Y(dpath_mulcore_ary1_a1_c2[31]));
AND2X1 mul_U2362(.A(n1287), .B(n3348), .Y(dpath_mulcore_ary1_a1_c2[30]));
AND2X1 mul_U2363(.A(n1288), .B(n3349), .Y(dpath_mulcore_ary1_a1_c2[29]));
AND2X1 mul_U2364(.A(n1289), .B(n3350), .Y(dpath_mulcore_ary1_a1_c2[28]));
AND2X1 mul_U2365(.A(n1290), .B(n3351), .Y(dpath_mulcore_ary1_a1_c2[27]));
AND2X1 mul_U2366(.A(n1291), .B(n3352), .Y(dpath_mulcore_ary1_a1_c2[26]));
AND2X1 mul_U2367(.A(n1292), .B(n3353), .Y(dpath_mulcore_ary1_a1_c2[25]));
AND2X1 mul_U2368(.A(n1293), .B(n3354), .Y(dpath_mulcore_ary1_a1_c2[24]));
AND2X1 mul_U2369(.A(n1294), .B(n3355), .Y(dpath_mulcore_ary1_a1_c2[23]));
AND2X1 mul_U2370(.A(n1295), .B(n3356), .Y(dpath_mulcore_ary1_a1_c2[22]));
AND2X1 mul_U2371(.A(n1296), .B(n3357), .Y(dpath_mulcore_ary1_a1_c2[21]));
AND2X1 mul_U2372(.A(n1297), .B(n3358), .Y(dpath_mulcore_ary1_a1_c2[20]));
AND2X1 mul_U2373(.A(n1298), .B(n3359), .Y(dpath_mulcore_ary1_a1_c2[19]));
AND2X1 mul_U2374(.A(n1299), .B(n3360), .Y(dpath_mulcore_ary1_a1_c2[18]));
AND2X1 mul_U2375(.A(n1300), .B(n3361), .Y(dpath_mulcore_ary1_a1_c2[17]));
AND2X1 mul_U2376(.A(n1301), .B(n3362), .Y(dpath_mulcore_ary1_a1_c2[16]));
AND2X1 mul_U2377(.A(n1302), .B(n3363), .Y(dpath_mulcore_ary1_a1_c2[15]));
AND2X1 mul_U2378(.A(n1303), .B(n3364), .Y(dpath_mulcore_ary1_a1_c2[14]));
AND2X1 mul_U2379(.A(n1304), .B(n3365), .Y(dpath_mulcore_ary1_a1_c2[13]));
AND2X1 mul_U2380(.A(n1305), .B(n3366), .Y(dpath_mulcore_ary1_a1_c2[12]));
AND2X1 mul_U2381(.A(n1306), .B(n3367), .Y(dpath_mulcore_ary1_a1_c2[11]));
AND2X1 mul_U2382(.A(n1307), .B(n3368), .Y(dpath_mulcore_ary1_a1_c2[10]));
AND2X1 mul_U2383(.A(n1308), .B(n3369), .Y(dpath_mulcore_ary1_a1_c2[9]));
AND2X1 mul_U2384(.A(n1309), .B(n3370), .Y(dpath_mulcore_ary1_a1_c2[8]));
AND2X1 mul_U2385(.A(n1310), .B(n3371), .Y(dpath_mulcore_ary1_a1_c2[7]));
AND2X1 mul_U2386(.A(n1311), .B(n3372), .Y(dpath_mulcore_ary1_a1_c2[6]));
AND2X1 mul_U2387(.A(n1312), .B(n3373), .Y(dpath_mulcore_ary1_a1_c2[5]));
AND2X1 mul_U2388(.A(n1313), .B(n3374), .Y(dpath_mulcore_ary1_a1_c2[4]));
AND2X1 mul_U2389(.A(n1128), .B(n3189), .Y(dpath_mulcore_ary1_a1_c2[3]));
AND2X1 mul_U2390(.A(n1129), .B(n3190), .Y(dpath_mulcore_ary1_a1_c2[2]));
AND2X1 mul_U2391(.A(n7399), .B(dpath_mulcore_ary1_a1_I2_I0_b0n), .Y(dpath_mulcore_ary1_a1_c2[1]));
INVX1 mul_U2392(.A(n13063), .Y(n9835));
OR2X1 mul_U2393(.A(n6992), .B(dpath_mulcore_b13[0]), .Y(n13063));
AND2X1 mul_U2394(.A(n1082), .B(n13574), .Y(dpath_mulcore_ary1_a1_I0_I1_11__net043));
OR2X1 mul_U2395(.A(n7163), .B(dpath_mulcore_b10[0]), .Y(n13574));
OR2X1 mul_U2396(.A(n9747), .B(n5950), .Y(dpath_mulcore_ary1_a1_b5n[1]));
AND2X1 mul_U2397(.A(n1085), .B(n13583), .Y(dpath_mulcore_ary1_a1_I0_I1_10__net043));
OR2X1 mul_U2398(.A(n7166), .B(dpath_mulcore_b10[0]), .Y(n13583));
AND2X1 mul_U2399(.A(n1429), .B(n3490), .Y(dpath_mulcore_ary1_a1_c0[8]));
OR2X1 mul_U2400(.A(n9745), .B(n5941), .Y(dpath_mulcore_ary1_a1_I1_I0_b1n_1));
AND2X1 mul_U2401(.A(n1430), .B(n3491), .Y(dpath_mulcore_ary1_a1_c0[7]));
AND2X1 mul_U2402(.A(n1094), .B(n13610), .Y(dpath_mulcore_ary1_a1_I0_I1_7__net043));
OR2X1 mul_U2403(.A(n7175), .B(dpath_mulcore_b10[0]), .Y(n13610));
AND2X1 mul_U2404(.A(n1097), .B(n13619), .Y(dpath_mulcore_ary1_a1_I0_I1_6__net043));
OR2X1 mul_U2405(.A(n7178), .B(dpath_mulcore_b10[0]), .Y(n13619));
AND2X1 mul_U2406(.A(n1100), .B(n13628), .Y(dpath_mulcore_ary1_a1_I0_I1_5__net043));
OR2X1 mul_U2407(.A(n7181), .B(dpath_mulcore_b10[0]), .Y(n13628));
INVX1 mul_U2408(.A(n13636), .Y(n9829));
OR2X1 mul_U2409(.A(n7184), .B(dpath_mulcore_b10[0]), .Y(n13636));
AND2X1 mul_U2410(.A(n2877), .B(n4553), .Y(dpath_n519));
AND2X1 mul_U2411(.A(n2881), .B(n4557), .Y(dpath_areg[96]));
AND2X1 mul_U2412(.A(n1898), .B(n3951), .Y(dpath_mulcore_array2_c1[80]));
AND2X1 mul_U2413(.A(n1926), .B(n3979), .Y(dpath_mulcore_array2_c2[67]));
AND2X1 mul_U2414(.A(n2319), .B(n4244), .Y(dpath_mulcore_array2_co[66]));
AND2X1 mul_U2415(.A(n2321), .B(n4246), .Y(dpath_mulcore_array2_co[65]));
AND2X1 mul_U2416(.A(n2323), .B(n4248), .Y(dpath_mulcore_array2_co[64]));
AND2X1 mul_U2417(.A(n2325), .B(n4250), .Y(dpath_mulcore_array2_co[63]));
AND2X1 mul_U2418(.A(n2327), .B(n4252), .Y(dpath_mulcore_array2_co[62]));
AND2X1 mul_U2419(.A(n2329), .B(n4254), .Y(dpath_mulcore_array2_co[61]));
AND2X1 mul_U2420(.A(n2331), .B(n4256), .Y(dpath_mulcore_array2_co[60]));
AND2X1 mul_U2421(.A(n2333), .B(n4258), .Y(dpath_mulcore_array2_co[59]));
AND2X1 mul_U2422(.A(n2335), .B(n4260), .Y(dpath_mulcore_array2_co[58]));
AND2X1 mul_U2423(.A(n2337), .B(n4262), .Y(dpath_mulcore_array2_co[57]));
AND2X1 mul_U2424(.A(n2339), .B(n4264), .Y(dpath_mulcore_array2_co[56]));
AND2X1 mul_U2425(.A(n2341), .B(n4266), .Y(dpath_mulcore_array2_co[55]));
AND2X1 mul_U2426(.A(n2343), .B(n4268), .Y(dpath_mulcore_array2_co[54]));
AND2X1 mul_U2427(.A(n2345), .B(n4270), .Y(dpath_mulcore_array2_co[53]));
AND2X1 mul_U2428(.A(n2347), .B(n4272), .Y(dpath_mulcore_array2_co[52]));
AND2X1 mul_U2429(.A(n2349), .B(n4274), .Y(dpath_mulcore_array2_co[51]));
AND2X1 mul_U2430(.A(n2351), .B(n4276), .Y(dpath_mulcore_array2_co[50]));
AND2X1 mul_U2431(.A(n2353), .B(n4278), .Y(dpath_mulcore_array2_co[49]));
AND2X1 mul_U2432(.A(n2355), .B(n4280), .Y(dpath_mulcore_array2_co[48]));
AND2X1 mul_U2433(.A(n2357), .B(n4282), .Y(dpath_mulcore_array2_co[47]));
AND2X1 mul_U2434(.A(n2359), .B(n4284), .Y(dpath_mulcore_array2_co[46]));
AND2X1 mul_U2435(.A(n2361), .B(n4286), .Y(dpath_mulcore_array2_co[45]));
AND2X1 mul_U2436(.A(n2363), .B(n4288), .Y(dpath_mulcore_array2_co[44]));
AND2X1 mul_U2437(.A(n2365), .B(n4290), .Y(dpath_mulcore_array2_co[43]));
AND2X1 mul_U2438(.A(n2367), .B(n4292), .Y(dpath_mulcore_array2_co[42]));
AND2X1 mul_U2439(.A(n2369), .B(n4294), .Y(dpath_mulcore_array2_co[41]));
AND2X1 mul_U2440(.A(n2371), .B(n4296), .Y(dpath_mulcore_array2_co[40]));
AND2X1 mul_U2441(.A(n2373), .B(n4298), .Y(dpath_mulcore_array2_co[39]));
AND2X1 mul_U2442(.A(n2375), .B(n4300), .Y(dpath_mulcore_array2_co[38]));
AND2X1 mul_U2443(.A(n2377), .B(n4302), .Y(dpath_mulcore_array2_co[37]));
AND2X1 mul_U2444(.A(n2379), .B(n4304), .Y(dpath_mulcore_array2_co[36]));
AND2X1 mul_U2445(.A(n2381), .B(n4306), .Y(dpath_mulcore_array2_co[35]));
AND2X1 mul_U2446(.A(n2383), .B(n4308), .Y(dpath_mulcore_array2_co[34]));
AND2X1 mul_U2447(.A(n2385), .B(n4310), .Y(dpath_mulcore_array2_co[33]));
AND2X1 mul_U2448(.A(n2387), .B(n4312), .Y(dpath_mulcore_array2_co[32]));
AND2X1 mul_U2449(.A(n2389), .B(n4314), .Y(dpath_mulcore_array2_co[31]));
AND2X1 mul_U2450(.A(n2391), .B(n4316), .Y(dpath_mulcore_array2_co[30]));
AND2X1 mul_U2451(.A(n2393), .B(n4318), .Y(dpath_mulcore_array2_co[29]));
INVX1 mul_U2452(.A(dpath_mulcore_array2_sc3_29__z), .Y(n10042));
INVX1 mul_U2453(.A(dpath_mulcore_array2_sc3_28__z), .Y(n10041));
INVX1 mul_U2454(.A(dpath_mulcore_array2_sc3_27__z), .Y(n10040));
INVX1 mul_U2455(.A(dpath_mulcore_array2_sc3_26__z), .Y(n10039));
INVX1 mul_U2456(.A(dpath_mulcore_array2_sc3_25__z), .Y(n10038));
INVX1 mul_U2457(.A(dpath_mulcore_array2_sc3_24__z), .Y(n10037));
INVX1 mul_U2458(.A(dpath_mulcore_array2_sc3_23__z), .Y(n10036));
INVX1 mul_U2459(.A(dpath_mulcore_array2_sc3_22__z), .Y(n10035));
INVX1 mul_U2460(.A(dpath_mulcore_array2_sc3_21__z), .Y(n10034));
AND2X1 mul_U2461(.A(n1949), .B(n4002), .Y(dpath_mulcore_array2_c1[3]));
AND2X1 mul_U2462(.A(n1950), .B(n4003), .Y(dpath_mulcore_array2_c1[2]));
AND2X1 mul_U2463(.A(n1951), .B(n4004), .Y(dpath_mulcore_array2_c1[1]));
AND2X1 mul_U2464(.A(n2062), .B(n4115), .Y(dpath_mulcore_array2_c1[0]));
AND2X1 mul_U2465(.A(n1483), .B(n3547), .Y(dpath_mulcore_array2_ain[29]));
AND2X1 mul_U2466(.A(n1484), .B(n3548), .Y(dpath_mulcore_array2_ain[28]));
AND2X1 mul_U2467(.A(n1485), .B(n3549), .Y(dpath_mulcore_array2_ain[27]));
AND2X1 mul_U2468(.A(n1486), .B(n3550), .Y(dpath_mulcore_array2_ain[26]));
AND2X1 mul_U2469(.A(n1487), .B(n3551), .Y(dpath_mulcore_array2_ain[25]));
AND2X1 mul_U2470(.A(n1488), .B(n3552), .Y(dpath_mulcore_array2_ain[24]));
AND2X1 mul_U2471(.A(n1489), .B(n3553), .Y(dpath_mulcore_array2_ain[23]));
AND2X1 mul_U2472(.A(n1490), .B(n3554), .Y(dpath_mulcore_array2_ain[22]));
AND2X1 mul_U2473(.A(n1491), .B(n3555), .Y(dpath_mulcore_array2_ain[21]));
AND2X1 mul_U2474(.A(n1492), .B(n3556), .Y(dpath_mulcore_array2_ain[20]));
AND2X1 mul_U2475(.A(n1519), .B(n3583), .Y(dpath_mulcore_array2_ain[19]));
AND2X1 mul_U2476(.A(n1520), .B(n3584), .Y(dpath_mulcore_array2_ain[18]));
AND2X1 mul_U2477(.A(n1521), .B(n3585), .Y(dpath_mulcore_array2_ain[17]));
AND2X1 mul_U2478(.A(n1522), .B(n3586), .Y(dpath_mulcore_array2_ain[16]));
AND2X1 mul_U2479(.A(n1937), .B(n3990), .Y(dpath_mulcore_array2_c2[14]));
AND2X1 mul_U2480(.A(n1529), .B(n3593), .Y(dpath_mulcore_array2_ain[14]));
AND2X1 mul_U2481(.A(n1530), .B(n3594), .Y(dpath_mulcore_array2_ain[13]));
AND2X1 mul_U2482(.A(n1531), .B(n3595), .Y(dpath_mulcore_array2_ain[12]));
AND2X1 mul_U2483(.A(n1532), .B(n3596), .Y(dpath_mulcore_array2_ain[11]));
AND2X1 mul_U2484(.A(n1533), .B(n3597), .Y(dpath_mulcore_array2_ain[10]));
AND2X1 mul_U2485(.A(n1534), .B(n3598), .Y(dpath_mulcore_array2_ain[9]));
AND2X1 mul_U2486(.A(n1535), .B(n3599), .Y(dpath_mulcore_array2_ain[8]));
AND2X1 mul_U2487(.A(n1536), .B(n3600), .Y(dpath_mulcore_array2_ain[7]));
AND2X1 mul_U2488(.A(n1537), .B(n3601), .Y(dpath_mulcore_array2_ain[6]));
AND2X1 mul_U2489(.A(n1538), .B(n3602), .Y(dpath_mulcore_array2_ain[5]));
AND2X1 mul_U2490(.A(n1524), .B(n3588), .Y(dpath_mulcore_array2_ain[4]));
AND2X1 mul_U2491(.A(n1525), .B(n3589), .Y(dpath_mulcore_array2_ain[3]));
AND2X1 mul_U2492(.A(n1526), .B(n3590), .Y(dpath_mulcore_array2_ain[2]));
AND2X1 mul_U2493(.A(n1527), .B(n3591), .Y(dpath_mulcore_array2_ain[1]));
AND2X1 mul_U2494(.A(n3006), .B(n4682), .Y(dpath_n976));
AND2X1 mul_U2495(.A(dpath_mulcore_ps[31]), .B(dpath_mulcore_pc[30]), .Y(dpath_mulcore_array2_c1x2));
AND2X1 mul_U2496(.A(n1110), .B(n13663), .Y(dpath_mulcore_ary1_a0_I1_I2_net47));
OR2X1 mul_U2497(.A(n9475), .B(dpath_mulcore_b3[0]), .Y(n13663));
AND2X1 mul_U2498(.A(n231), .B(n10999), .Y(dpath_mulcore_ary1_a0_I1_I2_net48));
OR2X1 mul_U2499(.A(n6301), .B(dpath_mulcore_b4[0]), .Y(n10999));
AND2X1 mul_U2500(.A(n230), .B(n10996), .Y(dpath_mulcore_ary1_a0_I1_I2_net43));
OR2X1 mul_U2501(.A(n6300), .B(dpath_mulcore_b4[0]), .Y(n10996));
AND2X1 mul_U2502(.A(n233), .B(n11005), .Y(dpath_mulcore_ary1_a0_I1_I1_63__net043));
OR2X1 mul_U2503(.A(n6303), .B(dpath_mulcore_b5[0]), .Y(n11005));
OR2X1 mul_U2504(.A(n9425), .B(dpath_mulcore_b2[0]), .Y(n13671));
AND2X1 mul_U2505(.A(n1437), .B(n3498), .Y(dpath_mulcore_ary1_a0_c0[67]));
AND2X1 mul_U2506(.A(n236), .B(n11014), .Y(dpath_mulcore_ary1_a0_I1_I1_62__net043));
OR2X1 mul_U2507(.A(n6306), .B(dpath_mulcore_b5[0]), .Y(n11014));
AND2X1 mul_U2508(.A(n1436), .B(n3497), .Y(dpath_mulcore_ary1_a0_c0[66]));
AND2X1 mul_U2509(.A(n239), .B(n11023), .Y(dpath_mulcore_ary1_a0_I1_I1_61__net043));
OR2X1 mul_U2510(.A(n6309), .B(dpath_mulcore_b5[0]), .Y(n11023));
AND2X1 mul_U2511(.A(n1435), .B(n3496), .Y(dpath_mulcore_ary1_a0_c0[65]));
AND2X1 mul_U2512(.A(n242), .B(n11032), .Y(dpath_mulcore_ary1_a0_I1_I1_60__net043));
OR2X1 mul_U2513(.A(n6312), .B(dpath_mulcore_b5[0]), .Y(n11032));
AND2X1 mul_U2514(.A(n1434), .B(n3495), .Y(dpath_mulcore_ary1_a0_c0[64]));
AND2X1 mul_U2515(.A(n245), .B(n11041), .Y(dpath_mulcore_ary1_a0_I1_I1_59__net043));
OR2X1 mul_U2516(.A(n6315), .B(dpath_mulcore_b5[0]), .Y(n11041));
AND2X1 mul_U2517(.A(n1194), .B(n3255), .Y(dpath_mulcore_ary1_a0_c0[63]));
AND2X1 mul_U2518(.A(n248), .B(n11050), .Y(dpath_mulcore_ary1_a0_I1_I1_58__net043));
OR2X1 mul_U2519(.A(n6318), .B(dpath_mulcore_b5[0]), .Y(n11050));
AND2X1 mul_U2520(.A(n1195), .B(n3256), .Y(dpath_mulcore_ary1_a0_c0[62]));
AND2X1 mul_U2521(.A(n251), .B(n11059), .Y(dpath_mulcore_ary1_a0_I1_I1_57__net043));
OR2X1 mul_U2522(.A(n6321), .B(dpath_mulcore_b5[0]), .Y(n11059));
AND2X1 mul_U2523(.A(n1196), .B(n3257), .Y(dpath_mulcore_ary1_a0_c0[61]));
AND2X1 mul_U2524(.A(n254), .B(n11068), .Y(dpath_mulcore_ary1_a0_I1_I1_56__net043));
OR2X1 mul_U2525(.A(n6324), .B(dpath_mulcore_b5[0]), .Y(n11068));
AND2X1 mul_U2526(.A(n1197), .B(n3258), .Y(dpath_mulcore_ary1_a0_c0[60]));
AND2X1 mul_U2527(.A(n257), .B(n11077), .Y(dpath_mulcore_ary1_a0_I1_I1_55__net043));
OR2X1 mul_U2528(.A(n6327), .B(dpath_mulcore_b5[0]), .Y(n11077));
AND2X1 mul_U2529(.A(n1198), .B(n3259), .Y(dpath_mulcore_ary1_a0_c0[59]));
AND2X1 mul_U2530(.A(n260), .B(n11086), .Y(dpath_mulcore_ary1_a0_I1_I1_54__net043));
OR2X1 mul_U2531(.A(n6330), .B(dpath_mulcore_b5[0]), .Y(n11086));
AND2X1 mul_U2532(.A(n1199), .B(n3260), .Y(dpath_mulcore_ary1_a0_c0[58]));
AND2X1 mul_U2533(.A(n263), .B(n11095), .Y(dpath_mulcore_ary1_a0_I1_I1_53__net043));
OR2X1 mul_U2534(.A(n6333), .B(dpath_mulcore_b5[0]), .Y(n11095));
AND2X1 mul_U2535(.A(n1200), .B(n3261), .Y(dpath_mulcore_ary1_a0_c0[57]));
AND2X1 mul_U2536(.A(n266), .B(n11104), .Y(dpath_mulcore_ary1_a0_I1_I1_52__net043));
OR2X1 mul_U2537(.A(n6336), .B(dpath_mulcore_b5[0]), .Y(n11104));
AND2X1 mul_U2538(.A(n1201), .B(n3262), .Y(dpath_mulcore_ary1_a0_c0[56]));
AND2X1 mul_U2539(.A(n269), .B(n11113), .Y(dpath_mulcore_ary1_a0_I1_I1_51__net043));
OR2X1 mul_U2540(.A(n6339), .B(dpath_mulcore_b5[0]), .Y(n11113));
AND2X1 mul_U2541(.A(n1202), .B(n3263), .Y(dpath_mulcore_ary1_a0_c0[55]));
AND2X1 mul_U2542(.A(n272), .B(n11122), .Y(dpath_mulcore_ary1_a0_I1_I1_50__net043));
OR2X1 mul_U2543(.A(n6342), .B(dpath_mulcore_b5[0]), .Y(n11122));
AND2X1 mul_U2544(.A(n1203), .B(n3264), .Y(dpath_mulcore_ary1_a0_c0[54]));
AND2X1 mul_U2545(.A(n275), .B(n11131), .Y(dpath_mulcore_ary1_a0_I1_I1_49__net043));
OR2X1 mul_U2546(.A(n6345), .B(dpath_mulcore_b5[0]), .Y(n11131));
AND2X1 mul_U2547(.A(n1204), .B(n3265), .Y(dpath_mulcore_ary1_a0_c0[53]));
AND2X1 mul_U2548(.A(n278), .B(n11140), .Y(dpath_mulcore_ary1_a0_I1_I1_48__net043));
OR2X1 mul_U2549(.A(n6348), .B(dpath_mulcore_b5[0]), .Y(n11140));
AND2X1 mul_U2550(.A(n1205), .B(n3266), .Y(dpath_mulcore_ary1_a0_c0[52]));
AND2X1 mul_U2551(.A(n281), .B(n11149), .Y(dpath_mulcore_ary1_a0_I1_I1_47__net043));
OR2X1 mul_U2552(.A(n6351), .B(dpath_mulcore_b5[0]), .Y(n11149));
AND2X1 mul_U2553(.A(n1206), .B(n3267), .Y(dpath_mulcore_ary1_a0_c0[51]));
AND2X1 mul_U2554(.A(n284), .B(n11158), .Y(dpath_mulcore_ary1_a0_I1_I1_46__net043));
OR2X1 mul_U2555(.A(n6354), .B(dpath_mulcore_b5[0]), .Y(n11158));
AND2X1 mul_U2556(.A(n1207), .B(n3268), .Y(dpath_mulcore_ary1_a0_c0[50]));
AND2X1 mul_U2557(.A(n287), .B(n11167), .Y(dpath_mulcore_ary1_a0_I1_I1_45__net043));
OR2X1 mul_U2558(.A(n6357), .B(dpath_mulcore_b5[0]), .Y(n11167));
AND2X1 mul_U2559(.A(n1208), .B(n3269), .Y(dpath_mulcore_ary1_a0_c0[49]));
AND2X1 mul_U2560(.A(n290), .B(n11176), .Y(dpath_mulcore_ary1_a0_I1_I1_44__net043));
OR2X1 mul_U2561(.A(n6360), .B(dpath_mulcore_b5[0]), .Y(n11176));
AND2X1 mul_U2562(.A(n1209), .B(n3270), .Y(dpath_mulcore_ary1_a0_c0[48]));
AND2X1 mul_U2563(.A(n293), .B(n11185), .Y(dpath_mulcore_ary1_a0_I1_I1_43__net043));
OR2X1 mul_U2564(.A(n6363), .B(dpath_mulcore_b5[0]), .Y(n11185));
AND2X1 mul_U2565(.A(n1210), .B(n3271), .Y(dpath_mulcore_ary1_a0_c0[47]));
AND2X1 mul_U2566(.A(n296), .B(n11194), .Y(dpath_mulcore_ary1_a0_I1_I1_42__net043));
OR2X1 mul_U2567(.A(n6366), .B(dpath_mulcore_b5[0]), .Y(n11194));
AND2X1 mul_U2568(.A(n1211), .B(n3272), .Y(dpath_mulcore_ary1_a0_c0[46]));
AND2X1 mul_U2569(.A(n299), .B(n11203), .Y(dpath_mulcore_ary1_a0_I1_I1_41__net043));
OR2X1 mul_U2570(.A(n6369), .B(dpath_mulcore_b5[0]), .Y(n11203));
AND2X1 mul_U2571(.A(n1212), .B(n3273), .Y(dpath_mulcore_ary1_a0_c0[45]));
AND2X1 mul_U2572(.A(n302), .B(n11212), .Y(dpath_mulcore_ary1_a0_I1_I1_40__net043));
OR2X1 mul_U2573(.A(n6372), .B(dpath_mulcore_b5[0]), .Y(n11212));
AND2X1 mul_U2574(.A(n1213), .B(n3274), .Y(dpath_mulcore_ary1_a0_c0[44]));
AND2X1 mul_U2575(.A(n305), .B(n11221), .Y(dpath_mulcore_ary1_a0_I1_I1_39__net043));
OR2X1 mul_U2576(.A(n6375), .B(dpath_mulcore_b5[0]), .Y(n11221));
AND2X1 mul_U2577(.A(n1214), .B(n3275), .Y(dpath_mulcore_ary1_a0_c0[43]));
AND2X1 mul_U2578(.A(n308), .B(n11230), .Y(dpath_mulcore_ary1_a0_I1_I1_38__net043));
OR2X1 mul_U2579(.A(n6378), .B(dpath_mulcore_b5[0]), .Y(n11230));
AND2X1 mul_U2580(.A(n1215), .B(n3276), .Y(dpath_mulcore_ary1_a0_c0[42]));
AND2X1 mul_U2581(.A(n311), .B(n11239), .Y(dpath_mulcore_ary1_a0_I1_I1_37__net043));
OR2X1 mul_U2582(.A(n6381), .B(dpath_mulcore_b5[0]), .Y(n11239));
AND2X1 mul_U2583(.A(n1216), .B(n3277), .Y(dpath_mulcore_ary1_a0_c0[41]));
AND2X1 mul_U2584(.A(n314), .B(n11248), .Y(dpath_mulcore_ary1_a0_I1_I1_36__net043));
OR2X1 mul_U2585(.A(n6384), .B(dpath_mulcore_b5[0]), .Y(n11248));
AND2X1 mul_U2586(.A(n1217), .B(n3278), .Y(dpath_mulcore_ary1_a0_c0[40]));
AND2X1 mul_U2587(.A(n317), .B(n11257), .Y(dpath_mulcore_ary1_a0_I1_I1_35__net043));
OR2X1 mul_U2588(.A(n6387), .B(dpath_mulcore_b5[0]), .Y(n11257));
AND2X1 mul_U2589(.A(n1218), .B(n3279), .Y(dpath_mulcore_ary1_a0_c0[39]));
AND2X1 mul_U2590(.A(n320), .B(n11266), .Y(dpath_mulcore_ary1_a0_I1_I1_34__net043));
OR2X1 mul_U2591(.A(n6390), .B(dpath_mulcore_b5[0]), .Y(n11266));
AND2X1 mul_U2592(.A(n1219), .B(n3280), .Y(dpath_mulcore_ary1_a0_c0[38]));
AND2X1 mul_U2593(.A(n323), .B(n11275), .Y(dpath_mulcore_ary1_a0_I1_I1_33__net043));
OR2X1 mul_U2594(.A(n6393), .B(dpath_mulcore_b5[0]), .Y(n11275));
AND2X1 mul_U2595(.A(n1220), .B(n3281), .Y(dpath_mulcore_ary1_a0_c0[37]));
AND2X1 mul_U2596(.A(n326), .B(n11284), .Y(dpath_mulcore_ary1_a0_I1_I1_32__net043));
OR2X1 mul_U2597(.A(n6396), .B(dpath_mulcore_b5[0]), .Y(n11284));
AND2X1 mul_U2598(.A(n1221), .B(n3282), .Y(dpath_mulcore_ary1_a0_c0[36]));
AND2X1 mul_U2599(.A(n329), .B(n11293), .Y(dpath_mulcore_ary1_a0_I1_I1_31__net043));
OR2X1 mul_U2600(.A(n6399), .B(dpath_mulcore_b5[0]), .Y(n11293));
AND2X1 mul_U2601(.A(n1222), .B(n3283), .Y(dpath_mulcore_ary1_a0_c0[35]));
AND2X1 mul_U2602(.A(n332), .B(n11302), .Y(dpath_mulcore_ary1_a0_I1_I1_30__net043));
OR2X1 mul_U2603(.A(n6402), .B(dpath_mulcore_b5[0]), .Y(n11302));
AND2X1 mul_U2604(.A(n1223), .B(n3284), .Y(dpath_mulcore_ary1_a0_c0[34]));
AND2X1 mul_U2605(.A(n335), .B(n11311), .Y(dpath_mulcore_ary1_a0_I1_I1_29__net043));
OR2X1 mul_U2606(.A(n6405), .B(dpath_mulcore_b5[0]), .Y(n11311));
AND2X1 mul_U2607(.A(n1224), .B(n3285), .Y(dpath_mulcore_ary1_a0_c0[33]));
AND2X1 mul_U2608(.A(n338), .B(n11320), .Y(dpath_mulcore_ary1_a0_I1_I1_28__net043));
OR2X1 mul_U2609(.A(n6408), .B(dpath_mulcore_b5[0]), .Y(n11320));
AND2X1 mul_U2610(.A(n1225), .B(n3286), .Y(dpath_mulcore_ary1_a0_c0[32]));
AND2X1 mul_U2611(.A(n341), .B(n11329), .Y(dpath_mulcore_ary1_a0_I1_I1_27__net043));
OR2X1 mul_U2612(.A(n6411), .B(dpath_mulcore_b5[0]), .Y(n11329));
AND2X1 mul_U2613(.A(n1226), .B(n3287), .Y(dpath_mulcore_ary1_a0_c0[31]));
AND2X1 mul_U2614(.A(n344), .B(n11338), .Y(dpath_mulcore_ary1_a0_I1_I1_26__net043));
OR2X1 mul_U2615(.A(n6414), .B(dpath_mulcore_b5[0]), .Y(n11338));
AND2X1 mul_U2616(.A(n1227), .B(n3288), .Y(dpath_mulcore_ary1_a0_c0[30]));
AND2X1 mul_U2617(.A(n347), .B(n11347), .Y(dpath_mulcore_ary1_a0_I1_I1_25__net043));
OR2X1 mul_U2618(.A(n6417), .B(dpath_mulcore_b5[0]), .Y(n11347));
AND2X1 mul_U2619(.A(n1228), .B(n3289), .Y(dpath_mulcore_ary1_a0_c0[29]));
AND2X1 mul_U2620(.A(n350), .B(n11356), .Y(dpath_mulcore_ary1_a0_I1_I1_24__net043));
OR2X1 mul_U2621(.A(n6420), .B(dpath_mulcore_b5[0]), .Y(n11356));
AND2X1 mul_U2622(.A(n1229), .B(n3290), .Y(dpath_mulcore_ary1_a0_c0[28]));
AND2X1 mul_U2623(.A(n353), .B(n11365), .Y(dpath_mulcore_ary1_a0_I1_I1_23__net043));
OR2X1 mul_U2624(.A(n6423), .B(dpath_mulcore_b5[0]), .Y(n11365));
AND2X1 mul_U2625(.A(n1230), .B(n3291), .Y(dpath_mulcore_ary1_a0_c0[27]));
AND2X1 mul_U2626(.A(n356), .B(n11374), .Y(dpath_mulcore_ary1_a0_I1_I1_22__net043));
OR2X1 mul_U2627(.A(n6426), .B(dpath_mulcore_b5[0]), .Y(n11374));
AND2X1 mul_U2628(.A(n1231), .B(n3292), .Y(dpath_mulcore_ary1_a0_c0[26]));
AND2X1 mul_U2629(.A(n359), .B(n11383), .Y(dpath_mulcore_ary1_a0_I1_I1_21__net043));
OR2X1 mul_U2630(.A(n6429), .B(dpath_mulcore_b5[0]), .Y(n11383));
AND2X1 mul_U2631(.A(n1232), .B(n3293), .Y(dpath_mulcore_ary1_a0_c0[25]));
AND2X1 mul_U2632(.A(n362), .B(n11392), .Y(dpath_mulcore_ary1_a0_I1_I1_20__net043));
OR2X1 mul_U2633(.A(n6432), .B(dpath_mulcore_b5[0]), .Y(n11392));
AND2X1 mul_U2634(.A(n1233), .B(n3294), .Y(dpath_mulcore_ary1_a0_c0[24]));
AND2X1 mul_U2635(.A(n365), .B(n11401), .Y(dpath_mulcore_ary1_a0_I1_I1_19__net043));
OR2X1 mul_U2636(.A(n6435), .B(dpath_mulcore_b5[0]), .Y(n11401));
AND2X1 mul_U2637(.A(n1234), .B(n3295), .Y(dpath_mulcore_ary1_a0_c0[23]));
AND2X1 mul_U2638(.A(n368), .B(n11410), .Y(dpath_mulcore_ary1_a0_I1_I1_18__net043));
OR2X1 mul_U2639(.A(n6438), .B(dpath_mulcore_b5[0]), .Y(n11410));
AND2X1 mul_U2640(.A(n1235), .B(n3296), .Y(dpath_mulcore_ary1_a0_c0[22]));
AND2X1 mul_U2641(.A(n371), .B(n11419), .Y(dpath_mulcore_ary1_a0_I1_I1_17__net043));
OR2X1 mul_U2642(.A(n6441), .B(dpath_mulcore_b5[0]), .Y(n11419));
AND2X1 mul_U2643(.A(n1236), .B(n3297), .Y(dpath_mulcore_ary1_a0_c0[21]));
AND2X1 mul_U2644(.A(n374), .B(n11428), .Y(dpath_mulcore_ary1_a0_I1_I1_16__net043));
OR2X1 mul_U2645(.A(n6444), .B(dpath_mulcore_b5[0]), .Y(n11428));
AND2X1 mul_U2646(.A(n1237), .B(n3298), .Y(dpath_mulcore_ary1_a0_c0[20]));
AND2X1 mul_U2647(.A(n377), .B(n11437), .Y(dpath_mulcore_ary1_a0_I1_I1_15__net043));
OR2X1 mul_U2648(.A(n6447), .B(dpath_mulcore_b5[0]), .Y(n11437));
AND2X1 mul_U2649(.A(n1238), .B(n3299), .Y(dpath_mulcore_ary1_a0_c0[19]));
AND2X1 mul_U2650(.A(n380), .B(n11446), .Y(dpath_mulcore_ary1_a0_I1_I1_14__net043));
OR2X1 mul_U2651(.A(n6450), .B(dpath_mulcore_b5[0]), .Y(n11446));
AND2X1 mul_U2652(.A(n1239), .B(n3300), .Y(dpath_mulcore_ary1_a0_c0[18]));
AND2X1 mul_U2653(.A(n383), .B(n11455), .Y(dpath_mulcore_ary1_a0_I1_I1_13__net043));
OR2X1 mul_U2654(.A(n6453), .B(dpath_mulcore_b5[0]), .Y(n11455));
AND2X1 mul_U2655(.A(n1240), .B(n3301), .Y(dpath_mulcore_ary1_a0_c0[17]));
AND2X1 mul_U2656(.A(n386), .B(n11464), .Y(dpath_mulcore_ary1_a0_I1_I1_12__net043));
OR2X1 mul_U2657(.A(n6456), .B(dpath_mulcore_b5[0]), .Y(n11464));
AND2X1 mul_U2658(.A(n1241), .B(n3302), .Y(dpath_mulcore_ary1_a0_c0[16]));
AND2X1 mul_U2659(.A(n389), .B(n11473), .Y(dpath_mulcore_ary1_a0_I1_I1_11__net043));
OR2X1 mul_U2660(.A(n6459), .B(dpath_mulcore_b5[0]), .Y(n11473));
AND2X1 mul_U2661(.A(n1242), .B(n3303), .Y(dpath_mulcore_ary1_a0_c0[15]));
AND2X1 mul_U2662(.A(n392), .B(n11482), .Y(dpath_mulcore_ary1_a0_I1_I1_10__net043));
OR2X1 mul_U2663(.A(n6462), .B(dpath_mulcore_b5[0]), .Y(n11482));
AND2X1 mul_U2664(.A(n1243), .B(n3304), .Y(dpath_mulcore_ary1_a0_c0[14]));
AND2X1 mul_U2665(.A(n395), .B(n11491), .Y(dpath_mulcore_ary1_a0_I1_I1_9__net043));
OR2X1 mul_U2666(.A(n6465), .B(dpath_mulcore_b5[0]), .Y(n11491));
AND2X1 mul_U2667(.A(n1244), .B(n3305), .Y(dpath_mulcore_ary1_a0_c0[13]));
AND2X1 mul_U2668(.A(n398), .B(n11500), .Y(dpath_mulcore_ary1_a0_I1_I1_8__net043));
OR2X1 mul_U2669(.A(n6468), .B(dpath_mulcore_b5[0]), .Y(n11500));
AND2X1 mul_U2670(.A(n572), .B(n12028), .Y(dpath_mulcore_ary1_a0_I0_I1_13__net043));
OR2X1 mul_U2671(.A(n6645), .B(dpath_mulcore_b2[0]), .Y(n12028));
AND2X1 mul_U2672(.A(n575), .B(n12037), .Y(dpath_mulcore_ary1_a0_I0_I1_12__net043));
OR2X1 mul_U2673(.A(n6648), .B(dpath_mulcore_b2[0]), .Y(n12037));
AND2X1 mul_U2674(.A(n413), .B(n11547), .Y(dpath_mulcore_ary1_a0_I1_I0_p1_3));
OR2X1 mul_U2675(.A(n6484), .B(dpath_mulcore_b4[0]), .Y(n11547));
AND2X1 mul_U2676(.A(n412), .B(n11544), .Y(dpath_mulcore_ary1_a0_I1_I0_p0_3));
OR2X1 mul_U2677(.A(n6483), .B(dpath_mulcore_b3[0]), .Y(n11544));
AND2X1 mul_U2678(.A(n602), .B(n12120), .Y(dpath_mulcore_ary1_a0_I0_I0_p1_3));
OR2X1 mul_U2679(.A(n6676), .B(dpath_mulcore_b1[0]), .Y(n12120));
AND2X1 mul_U2680(.A(n601), .B(n12117), .Y(dpath_mulcore_ary1_a0_I0_I0_p0_3));
OR2X1 mul_U2681(.A(n6675), .B(dpath_mulcore_b0[0]), .Y(n12117));
INVX1 mul_U2682(.A(dpath_mulcore_op1_l[1]), .Y(n9858));
AND2X1 mul_U2683(.A(n2064), .B(n4117), .Y(dpath_mulcore_ary1_a0_c2[3]));
AND2X1 mul_U2684(.A(n2063), .B(n4116), .Y(dpath_mulcore_ary1_a0_c2[2]));
AND2X1 mul_U2685(.A(n7396), .B(dpath_mulcore_ary1_a0_I2_I0_b0n), .Y(dpath_mulcore_ary1_a0_c2[1]));
INVX1 mul_U2686(.A(n11535), .Y(n9848));
OR2X1 mul_U2687(.A(n6480), .B(dpath_mulcore_b5[0]), .Y(n11535));
AND2X1 mul_U2688(.A(n578), .B(n12046), .Y(dpath_mulcore_ary1_a0_I0_I1_11__net043));
OR2X1 mul_U2689(.A(n6651), .B(dpath_mulcore_b2[0]), .Y(n12046));
OR2X1 mul_U2690(.A(n9731), .B(n5958), .Y(dpath_mulcore_ary1_a0_b5n[1]));
AND2X1 mul_U2691(.A(n581), .B(n12055), .Y(dpath_mulcore_ary1_a0_I0_I1_10__net043));
OR2X1 mul_U2692(.A(n6654), .B(dpath_mulcore_b2[0]), .Y(n12055));
AND2X1 mul_U2693(.A(n1249), .B(n3310), .Y(dpath_mulcore_ary1_a0_c0[8]));
OR2X1 mul_U2694(.A(n9729), .B(n5929), .Y(dpath_mulcore_ary1_a0_I1_I0_b1n_1));
AND2X1 mul_U2695(.A(n1250), .B(n3311), .Y(dpath_mulcore_ary1_a0_c0[7]));
AND2X1 mul_U2696(.A(n590), .B(n12082), .Y(dpath_mulcore_ary1_a0_I0_I1_7__net043));
OR2X1 mul_U2697(.A(n6663), .B(dpath_mulcore_b2[0]), .Y(n12082));
AND2X1 mul_U2698(.A(n593), .B(n12091), .Y(dpath_mulcore_ary1_a0_I0_I1_6__net043));
OR2X1 mul_U2699(.A(n6666), .B(dpath_mulcore_b2[0]), .Y(n12091));
AND2X1 mul_U2700(.A(n596), .B(n12100), .Y(dpath_mulcore_ary1_a0_I0_I1_5__net043));
OR2X1 mul_U2701(.A(n6669), .B(dpath_mulcore_b2[0]), .Y(n12100));
INVX1 mul_U2702(.A(n12108), .Y(n9842));
OR2X1 mul_U2703(.A(n6672), .B(dpath_mulcore_b2[0]), .Y(n12108));
AND2X1 mul_U2704(.A(n2811), .B(n4487), .Y(dpath_n321));
OR2X1 mul_U2705(.A(n5873), .B(n6001), .Y(dpath_mul_op2_d[2]));
AND2X1 mul_U2706(.A(n2834), .B(n4510), .Y(dpath_n386));
AND2X1 mul_U2707(.A(n2767), .B(n4443), .Y(dpath_n189));
OR2X1 mul_U2708(.A(n5851), .B(n5979), .Y(dpath_mul_op2_d[4]));
AND2X1 mul_U2709(.A(n2790), .B(n4466), .Y(dpath_n254));
INVX1 mul_U2710(.A(dpath_mulcore_booth_b1_in0[2]), .Y(n9807));
INVX1 mul_U2711(.A(dpath_mul_op2_d[4]), .Y(n9808));
INVX1 mul_U2712(.A(dpath_mulcore_booth_b1_in1[2]), .Y(n10084));
INVX1 mul_U2713(.A(dpath_mulcore_booth_b[36]), .Y(n10085));
AND2X1 mul_U2714(.A(n2755), .B(n4431), .Y(dpath_n153));
OR2X1 mul_U2715(.A(n5835), .B(n5963), .Y(dpath_mul_op2_d[6]));
AND2X1 mul_U2716(.A(n2758), .B(n4434), .Y(dpath_n158));
INVX1 mul_U2717(.A(dpath_mulcore_booth_b2_in0[2]), .Y(n9809));
INVX1 mul_U2718(.A(dpath_mul_op2_d[6]), .Y(n9810));
INVX1 mul_U2719(.A(dpath_mulcore_booth_b2_in1[2]), .Y(n10086));
INVX1 mul_U2720(.A(dpath_mulcore_booth_b[38]), .Y(n10087));
AND2X1 mul_U2721(.A(n2751), .B(n4427), .Y(dpath_n138));
OR2X1 mul_U2722(.A(n5833), .B(n5961), .Y(dpath_mul_op2_d[8]));
AND2X1 mul_U2723(.A(n2754), .B(n4430), .Y(dpath_n146));
INVX1 mul_U2724(.A(dpath_mulcore_booth_b3_in0[2]), .Y(n9811));
INVX1 mul_U2725(.A(dpath_mul_op2_d[8]), .Y(n9812));
INVX1 mul_U2726(.A(dpath_mulcore_booth_b3_in1[2]), .Y(n10088));
INVX1 mul_U2727(.A(dpath_mulcore_booth_b[40]), .Y(n10089));
AND2X1 mul_U2728(.A(n2873), .B(n4549), .Y(dpath_n507));
OR2X1 mul_U2729(.A(n5894), .B(n6022), .Y(dpath_mul_op2_d[10]));
AND2X1 mul_U2730(.A(n2876), .B(n4552), .Y(dpath_n512));
INVX1 mul_U2731(.A(dpath_mulcore_booth_b4_in0[2]), .Y(n9813));
INVX1 mul_U2732(.A(dpath_mul_op2_d[10]), .Y(n9787));
INVX1 mul_U2733(.A(dpath_mulcore_booth_b4_in1[2]), .Y(n10090));
INVX1 mul_U2734(.A(dpath_mulcore_booth_b[42]), .Y(n10091));
AND2X1 mul_U2735(.A(n2869), .B(n4545), .Y(dpath_n495));
OR2X1 mul_U2736(.A(n5892), .B(n6020), .Y(dpath_mul_op2_d[12]));
AND2X1 mul_U2737(.A(n2872), .B(n4548), .Y(dpath_n500));
INVX1 mul_U2738(.A(dpath_mulcore_booth_b5_in0[2]), .Y(n9788));
INVX1 mul_U2739(.A(dpath_mul_op2_d[12]), .Y(n9789));
INVX1 mul_U2740(.A(dpath_mulcore_booth_b5_in1[2]), .Y(n10092));
INVX1 mul_U2741(.A(dpath_mulcore_booth_b[44]), .Y(n10093));
AND2X1 mul_U2742(.A(n2865), .B(n4541), .Y(dpath_n483));
OR2X1 mul_U2743(.A(n5890), .B(n6018), .Y(dpath_mul_op2_d[14]));
AND2X1 mul_U2744(.A(n2868), .B(n4544), .Y(dpath_n488));
INVX1 mul_U2745(.A(dpath_mulcore_booth_b6_in0[2]), .Y(n9790));
INVX1 mul_U2746(.A(dpath_mul_op2_d[14]), .Y(n9791));
INVX1 mul_U2747(.A(dpath_mulcore_booth_b6_in1[2]), .Y(n10094));
INVX1 mul_U2748(.A(dpath_mulcore_booth_b[46]), .Y(n10095));
AND2X1 mul_U2749(.A(n2861), .B(n4537), .Y(dpath_n471));
OR2X1 mul_U2750(.A(n5888), .B(n6016), .Y(dpath_mul_op2_d[16]));
AND2X1 mul_U2751(.A(n2864), .B(n4540), .Y(dpath_n476));
INVX1 mul_U2752(.A(dpath_mulcore_booth_b8_in1[2]), .Y(n10097));
AND2X1 mul_U2753(.A(n2857), .B(n4533), .Y(dpath_n459));
INVX1 mul_U2754(.A(dpath_mulcore_booth_b8_in0[2]), .Y(n9793));
OR2X1 mul_U2755(.A(n5886), .B(n6014), .Y(dpath_mul_op2_d[18]));
AND2X1 mul_U2756(.A(n2860), .B(n4536), .Y(dpath_n464));
AND2X1 mul_U2757(.A(n2851), .B(n4527), .Y(dpath_n441));
OR2X1 mul_U2758(.A(n5883), .B(n6011), .Y(dpath_mul_op2_d[20]));
AND2X1 mul_U2759(.A(n2854), .B(n4530), .Y(dpath_n446));
INVX1 mul_U2760(.A(dpath_mulcore_booth_b9_in0[2]), .Y(n9794));
INVX1 mul_U2761(.A(dpath_mul_op2_d[20]), .Y(n9796));
INVX1 mul_U2762(.A(dpath_mulcore_booth_b9_in1[2]), .Y(n10098));
INVX1 mul_U2763(.A(dpath_mulcore_booth_b[52]), .Y(n10099));
AND2X1 mul_U2764(.A(n2847), .B(n4523), .Y(dpath_n429));
OR2X1 mul_U2765(.A(n5881), .B(n6009), .Y(dpath_mul_op2_d[22]));
AND2X1 mul_U2766(.A(n2850), .B(n4526), .Y(dpath_n434));
INVX1 mul_U2767(.A(dpath_mulcore_booth_b10_in0[2]), .Y(n9797));
INVX1 mul_U2768(.A(dpath_mul_op2_d[22]), .Y(n9798));
INVX1 mul_U2769(.A(dpath_mulcore_booth_b10_in1[2]), .Y(n10100));
INVX1 mul_U2770(.A(dpath_mulcore_booth_b[54]), .Y(n10101));
AND2X1 mul_U2771(.A(n2843), .B(n4519), .Y(dpath_n417));
OR2X1 mul_U2772(.A(n5879), .B(n6007), .Y(dpath_mul_op2_d[24]));
AND2X1 mul_U2773(.A(n2846), .B(n4522), .Y(dpath_n422));
INVX1 mul_U2774(.A(dpath_mulcore_booth_b11_in0[2]), .Y(n9799));
INVX1 mul_U2775(.A(dpath_mul_op2_d[24]), .Y(n9800));
INVX1 mul_U2776(.A(dpath_mulcore_booth_b11_in1[2]), .Y(n10102));
INVX1 mul_U2777(.A(dpath_mulcore_booth_b[56]), .Y(n10103));
AND2X1 mul_U2778(.A(n2839), .B(n4515), .Y(dpath_n405));
OR2X1 mul_U2779(.A(n5877), .B(n6005), .Y(dpath_mul_op2_d[26]));
AND2X1 mul_U2780(.A(n2842), .B(n4518), .Y(dpath_n410));
INVX1 mul_U2781(.A(dpath_mulcore_booth_b12_in0[2]), .Y(n9801));
INVX1 mul_U2782(.A(dpath_mul_op2_d[26]), .Y(n9802));
INVX1 mul_U2783(.A(dpath_mulcore_booth_b12_in1[2]), .Y(n10104));
INVX1 mul_U2784(.A(dpath_mulcore_booth_b[58]), .Y(n10105));
AND2X1 mul_U2785(.A(n2835), .B(n4511), .Y(dpath_n393));
OR2X1 mul_U2786(.A(n5875), .B(n6003), .Y(dpath_mul_op2_d[28]));
AND2X1 mul_U2787(.A(n2838), .B(n4514), .Y(dpath_n398));
INVX1 mul_U2788(.A(dpath_mulcore_booth_b13_in0[2]), .Y(n9803));
INVX1 mul_U2789(.A(dpath_mul_op2_d[28]), .Y(n9804));
INVX1 mul_U2790(.A(dpath_mulcore_booth_b13_in1[2]), .Y(n10106));
INVX1 mul_U2791(.A(dpath_mulcore_booth_b[60]), .Y(n10107));
OR2X1 mul_U2792(.A(n5872), .B(n6000), .Y(dpath_mul_op2_d[30]));
AND2X1 mul_U2793(.A(n2832), .B(n4508), .Y(dpath_n380));
INVX1 mul_U2794(.A(dpath_mulcore_booth_b14_in0[2]), .Y(n9805));
INVX1 mul_U2795(.A(dpath_mul_op2_d[30]), .Y(n9806));
INVX1 mul_U2796(.A(dpath_mulcore_booth_b14_in1[2]), .Y(n10108));
INVX1 mul_U2797(.A(dpath_mulcore_booth_b[62]), .Y(n10109));
AND2X1 mul_U2798(.A(n731), .B(n12515), .Y(dpath_mulcore_ary1_a1_I1_I2_net078));
OR2X1 mul_U2799(.A(n6809), .B(dpath_mulcore_b13[0]), .Y(n12515));
AND2X1 mul_U2800(.A(dpath_mulcore_ary1_a1_I1_I2_net38), .B(n3504), .Y(dpath_mulcore_ary1_a1_c1[66]));
OR2X1 mul_U2801(.A(n9480), .B(dpath_mulcore_b12[0]), .Y(n13683));
AND2X1 mul_U2802(.A(n732), .B(n12518), .Y(dpath_mulcore_ary1_a1_I1_I2_net8));
OR2X1 mul_U2803(.A(n6810), .B(dpath_mulcore_b13[0]), .Y(n12518));
AND2X1 mul_U2804(.A(n1441), .B(n3503), .Y(dpath_mulcore_ary1_a1_c1[65]));
AND2X1 mul_U2805(.A(n736), .B(n12530), .Y(dpath_mulcore_ary1_a1_I1_I2_net35));
OR2X1 mul_U2806(.A(n6814), .B(dpath_mulcore_b13[0]), .Y(n12530));
AND2X1 mul_U2807(.A(n1440), .B(n3502), .Y(dpath_mulcore_ary1_a1_c1[64]));
AND2X1 mul_U2808(.A(n733), .B(n12521), .Y(dpath_mulcore_ary1_a1_I1_I2_net15));
OR2X1 mul_U2809(.A(n6811), .B(dpath_mulcore_b13[0]), .Y(n12521));
AND2X1 mul_U2810(.A(n1314), .B(n3375), .Y(dpath_mulcore_ary1_a1_c1[63]));
AND2X1 mul_U2811(.A(n1315), .B(n3376), .Y(dpath_mulcore_ary1_a1_c1[62]));
AND2X1 mul_U2812(.A(n1316), .B(n3377), .Y(dpath_mulcore_ary1_a1_c1[61]));
AND2X1 mul_U2813(.A(n1317), .B(n3378), .Y(dpath_mulcore_ary1_a1_c1[60]));
AND2X1 mul_U2814(.A(n1318), .B(n3379), .Y(dpath_mulcore_ary1_a1_c1[59]));
AND2X1 mul_U2815(.A(n1319), .B(n3380), .Y(dpath_mulcore_ary1_a1_c1[58]));
AND2X1 mul_U2816(.A(n1320), .B(n3381), .Y(dpath_mulcore_ary1_a1_c1[57]));
AND2X1 mul_U2817(.A(n1321), .B(n3382), .Y(dpath_mulcore_ary1_a1_c1[56]));
AND2X1 mul_U2818(.A(n1322), .B(n3383), .Y(dpath_mulcore_ary1_a1_c1[55]));
AND2X1 mul_U2819(.A(n1323), .B(n3384), .Y(dpath_mulcore_ary1_a1_c1[54]));
AND2X1 mul_U2820(.A(n1324), .B(n3385), .Y(dpath_mulcore_ary1_a1_c1[53]));
AND2X1 mul_U2821(.A(n1325), .B(n3386), .Y(dpath_mulcore_ary1_a1_c1[52]));
AND2X1 mul_U2822(.A(n1326), .B(n3387), .Y(dpath_mulcore_ary1_a1_c1[51]));
AND2X1 mul_U2823(.A(n1327), .B(n3388), .Y(dpath_mulcore_ary1_a1_c1[50]));
AND2X1 mul_U2824(.A(n1328), .B(n3389), .Y(dpath_mulcore_ary1_a1_c1[49]));
AND2X1 mul_U2825(.A(n1329), .B(n3390), .Y(dpath_mulcore_ary1_a1_c1[48]));
AND2X1 mul_U2826(.A(n1330), .B(n3391), .Y(dpath_mulcore_ary1_a1_c1[47]));
AND2X1 mul_U2827(.A(n1331), .B(n3392), .Y(dpath_mulcore_ary1_a1_c1[46]));
AND2X1 mul_U2828(.A(n1332), .B(n3393), .Y(dpath_mulcore_ary1_a1_c1[45]));
AND2X1 mul_U2829(.A(n1333), .B(n3394), .Y(dpath_mulcore_ary1_a1_c1[44]));
AND2X1 mul_U2830(.A(n1334), .B(n3395), .Y(dpath_mulcore_ary1_a1_c1[43]));
AND2X1 mul_U2831(.A(n1335), .B(n3396), .Y(dpath_mulcore_ary1_a1_c1[42]));
AND2X1 mul_U2832(.A(n1336), .B(n3397), .Y(dpath_mulcore_ary1_a1_c1[41]));
AND2X1 mul_U2833(.A(n1337), .B(n3398), .Y(dpath_mulcore_ary1_a1_c1[40]));
AND2X1 mul_U2834(.A(n1338), .B(n3399), .Y(dpath_mulcore_ary1_a1_c1[39]));
AND2X1 mul_U2835(.A(n1339), .B(n3400), .Y(dpath_mulcore_ary1_a1_c1[38]));
AND2X1 mul_U2836(.A(n1340), .B(n3401), .Y(dpath_mulcore_ary1_a1_c1[37]));
AND2X1 mul_U2837(.A(n1341), .B(n3402), .Y(dpath_mulcore_ary1_a1_c1[36]));
AND2X1 mul_U2838(.A(n1342), .B(n3403), .Y(dpath_mulcore_ary1_a1_c1[35]));
AND2X1 mul_U2839(.A(n1343), .B(n3404), .Y(dpath_mulcore_ary1_a1_c1[34]));
AND2X1 mul_U2840(.A(n1344), .B(n3405), .Y(dpath_mulcore_ary1_a1_c1[33]));
AND2X1 mul_U2841(.A(n1345), .B(n3406), .Y(dpath_mulcore_ary1_a1_c1[32]));
AND2X1 mul_U2842(.A(n1346), .B(n3407), .Y(dpath_mulcore_ary1_a1_c1[31]));
AND2X1 mul_U2843(.A(n1347), .B(n3408), .Y(dpath_mulcore_ary1_a1_c1[30]));
AND2X1 mul_U2844(.A(n1348), .B(n3409), .Y(dpath_mulcore_ary1_a1_c1[29]));
AND2X1 mul_U2845(.A(n1349), .B(n3410), .Y(dpath_mulcore_ary1_a1_c1[28]));
AND2X1 mul_U2846(.A(n1350), .B(n3411), .Y(dpath_mulcore_ary1_a1_c1[27]));
AND2X1 mul_U2847(.A(n1351), .B(n3412), .Y(dpath_mulcore_ary1_a1_c1[26]));
AND2X1 mul_U2848(.A(n1352), .B(n3413), .Y(dpath_mulcore_ary1_a1_c1[25]));
AND2X1 mul_U2849(.A(n1353), .B(n3414), .Y(dpath_mulcore_ary1_a1_c1[24]));
AND2X1 mul_U2850(.A(n1354), .B(n3415), .Y(dpath_mulcore_ary1_a1_c1[23]));
AND2X1 mul_U2851(.A(n1355), .B(n3416), .Y(dpath_mulcore_ary1_a1_c1[22]));
AND2X1 mul_U2852(.A(n1356), .B(n3417), .Y(dpath_mulcore_ary1_a1_c1[21]));
AND2X1 mul_U2853(.A(n1357), .B(n3418), .Y(dpath_mulcore_ary1_a1_c1[20]));
AND2X1 mul_U2854(.A(n1358), .B(n3419), .Y(dpath_mulcore_ary1_a1_c1[19]));
AND2X1 mul_U2855(.A(n1359), .B(n3420), .Y(dpath_mulcore_ary1_a1_c1[18]));
AND2X1 mul_U2856(.A(n1360), .B(n3421), .Y(dpath_mulcore_ary1_a1_c1[17]));
AND2X1 mul_U2857(.A(n1361), .B(n3422), .Y(dpath_mulcore_ary1_a1_c1[16]));
AND2X1 mul_U2858(.A(n1362), .B(n3423), .Y(dpath_mulcore_ary1_a1_c1[15]));
AND2X1 mul_U2859(.A(n1363), .B(n3424), .Y(dpath_mulcore_ary1_a1_c1[14]));
AND2X1 mul_U2860(.A(n1364), .B(n3425), .Y(dpath_mulcore_ary1_a1_c1[13]));
AND2X1 mul_U2861(.A(n1365), .B(n3426), .Y(dpath_mulcore_ary1_a1_c1[12]));
AND2X1 mul_U2862(.A(n1366), .B(n3427), .Y(dpath_mulcore_ary1_a1_c1[11]));
AND2X1 mul_U2863(.A(n1367), .B(n3428), .Y(dpath_mulcore_ary1_a1_c1[10]));
AND2X1 mul_U2864(.A(n1368), .B(n3429), .Y(dpath_mulcore_ary1_a1_c1[9]));
AND2X1 mul_U2865(.A(n1369), .B(n3430), .Y(dpath_mulcore_ary1_a1_c1[8]));
AND2X1 mul_U2866(.A(n1370), .B(n3431), .Y(dpath_mulcore_ary1_a1_c1[7]));
AND2X1 mul_U2867(.A(n1425), .B(n3486), .Y(dpath_mulcore_ary1_a1_c0[12]));
AND2X1 mul_U2868(.A(n1371), .B(n3432), .Y(dpath_mulcore_ary1_a1_c1[6]));
AND2X1 mul_U2869(.A(n1426), .B(n3487), .Y(dpath_mulcore_ary1_a1_c0[11]));
AND2X1 mul_U2870(.A(n1372), .B(n3433), .Y(dpath_mulcore_ary1_a1_c1[5]));
OR2X1 mul_U2871(.A(n9745), .B(n5940), .Y(dpath_mulcore_ary1_a1_I1_I0_b1n_0));
INVX1 mul_U2872(.A(n13085), .Y(n9831));
OR2X1 mul_U2873(.A(n7000), .B(dpath_mulcore_b12[0]), .Y(n13085));
AND2X1 mul_U2874(.A(n918), .B(n13078), .Y(dpath_mulcore_ary1_a1_I1_I0_p0_2));
OR2X1 mul_U2875(.A(n6997), .B(dpath_mulcore_b11[0]), .Y(n13078));
OR2X1 mul_U2876(.A(n9739), .B(n5945), .Y(dpath_mulcore_ary1_a1_I0_I0_b1n_1));
INVX1 mul_U2877(.A(n13658), .Y(n9827));
OR2X1 mul_U2878(.A(n7192), .B(dpath_mulcore_b9[0]), .Y(n13658));
AND2X1 mul_U2879(.A(n1107), .B(n13651), .Y(dpath_mulcore_ary1_a1_I0_I0_p0_2));
OR2X1 mul_U2880(.A(n7189), .B(dpath_mulcore_b8[0]), .Y(n13651));
INVX1 mul_U2881(.A(dpath_mulcore_op1_l[62]), .Y(n10031));
AND2X1 mul_U2882(.A(n605), .B(n12133), .Y(dpath_mulcore_ary1_a1_I2_I2_net43));
OR2X1 mul_U2883(.A(n6681), .B(dpath_mulcore_b15[0]), .Y(n12133));
OR2X1 mul_U2884(.A(n9747), .B(n5951), .Y(dpath_mulcore_ary1_a1_b5n[0]));
AND2X1 mul_U2885(.A(n1427), .B(n3488), .Y(dpath_mulcore_ary1_a1_c0[10]));
AND2X1 mul_U2886(.A(n1373), .B(n3434), .Y(dpath_mulcore_ary1_a1_c1[4]));
AND2X1 mul_U2887(.A(n1428), .B(n3489), .Y(dpath_mulcore_ary1_a1_c0[9]));
AND2X1 mul_U2888(.A(n1431), .B(n3492), .Y(dpath_mulcore_ary1_a1_c0[6]));
AND2X1 mul_U2889(.A(n1432), .B(n3493), .Y(dpath_mulcore_ary1_a1_c0[5]));
INVX1 mul_U2890(.A(n13083), .Y(n9832));
OR2X1 mul_U2891(.A(n6999), .B(dpath_mulcore_b11[0]), .Y(n13083));
OR2X1 mul_U2892(.A(n9743), .B(n5942), .Y(dpath_mulcore_ary1_a1_I1_I0_b0n_0));
AND2X1 mul_U2893(.A(n1433), .B(n3494), .Y(dpath_mulcore_ary1_a1_c0[4]));
AND2X1 mul_U2894(.A(n1132), .B(n3193), .Y(dpath_mulcore_ary1_a1_c0[3]));
INVX1 mul_U2895(.A(dpath_mulcore_booth_b0_in0[2]), .Y(n9795));
INVX1 mul_U2896(.A(dpath_mulcore_booth_b0_in1[2]), .Y(n10083));
AND2X1 mul_U2897(.A(n2855), .B(n4531), .Y(dpath_n453));
OR2X1 mul_U2898(.A(n5895), .B(n6023), .Y(dpath_mul_op2_d[0]));
AND2X1 mul_U2899(.A(n2878), .B(n4554), .Y(dpath_n518));
AND2X1 mul_U2900(.A(n1482), .B(n3546), .Y(dpath_mulcore_array2_ain[30]));
AND2X1 mul_U2901(.A(n1493), .B(n3557), .Y(dpath_mulcore_array2_ain[95]));
AND2X1 mul_U2902(.A(n1494), .B(n3558), .Y(dpath_mulcore_array2_ain[94]));
AND2X1 mul_U2903(.A(n1495), .B(n3559), .Y(dpath_mulcore_array2_ain[93]));
AND2X1 mul_U2904(.A(n1496), .B(n3560), .Y(dpath_mulcore_array2_ain[92]));
AND2X1 mul_U2905(.A(n1497), .B(n3561), .Y(dpath_mulcore_array2_ain[91]));
AND2X1 mul_U2906(.A(n1498), .B(n3562), .Y(dpath_mulcore_array2_ain[90]));
AND2X1 mul_U2907(.A(n1499), .B(n3563), .Y(dpath_mulcore_array2_ain[89]));
AND2X1 mul_U2908(.A(n1500), .B(n3564), .Y(dpath_mulcore_array2_ain[88]));
AND2X1 mul_U2909(.A(n1501), .B(n3565), .Y(dpath_mulcore_array2_ain[87]));
AND2X1 mul_U2910(.A(n1502), .B(n3566), .Y(dpath_mulcore_array2_ain[86]));
AND2X1 mul_U2911(.A(n1503), .B(n3567), .Y(dpath_mulcore_array2_ain[85]));
AND2X1 mul_U2912(.A(n1504), .B(n3568), .Y(dpath_mulcore_array2_ain[84]));
AND2X1 mul_U2913(.A(n1528), .B(n3592), .Y(dpath_mulcore_array2_ain[83]));
AND2X1 mul_U2914(.A(n2478), .B(n4404), .Y(dpath_mulcore_array2_ain[82]));
AND2X1 mul_U2915(.A(n2045), .B(n4098), .Y(dpath_mulcore_array2_c2[80]));
AND2X1 mul_U2916(.A(n1506), .B(n3570), .Y(dpath_mulcore_array2_ain[81]));
AND2X1 mul_U2917(.A(n2046), .B(n4099), .Y(dpath_mulcore_array2_c2[79]));
AND2X1 mul_U2918(.A(n1507), .B(n3571), .Y(dpath_mulcore_array2_ain[80]));
AND2X1 mul_U2919(.A(n2047), .B(n4100), .Y(dpath_mulcore_array2_c2[78]));
AND2X1 mul_U2920(.A(n1508), .B(n3572), .Y(dpath_mulcore_array2_ain[79]));
AND2X1 mul_U2921(.A(n2048), .B(n4101), .Y(dpath_mulcore_array2_c2[77]));
AND2X1 mul_U2922(.A(n1509), .B(n3573), .Y(dpath_mulcore_array2_ain[78]));
AND2X1 mul_U2923(.A(n2049), .B(n4102), .Y(dpath_mulcore_array2_c2[76]));
AND2X1 mul_U2924(.A(n1510), .B(n3574), .Y(dpath_mulcore_array2_ain[77]));
AND2X1 mul_U2925(.A(n2050), .B(n4103), .Y(dpath_mulcore_array2_c2[75]));
AND2X1 mul_U2926(.A(n1511), .B(n3575), .Y(dpath_mulcore_array2_ain[76]));
AND2X1 mul_U2927(.A(n2051), .B(n4104), .Y(dpath_mulcore_array2_c2[74]));
AND2X1 mul_U2928(.A(n1512), .B(n3576), .Y(dpath_mulcore_array2_ain[75]));
AND2X1 mul_U2929(.A(n2052), .B(n4105), .Y(dpath_mulcore_array2_c2[73]));
AND2X1 mul_U2930(.A(n1513), .B(n3577), .Y(dpath_mulcore_array2_ain[74]));
AND2X1 mul_U2931(.A(n2053), .B(n4106), .Y(dpath_mulcore_array2_c2[72]));
AND2X1 mul_U2932(.A(n1514), .B(n3578), .Y(dpath_mulcore_array2_ain[73]));
AND2X1 mul_U2933(.A(n2054), .B(n4107), .Y(dpath_mulcore_array2_c2[71]));
AND2X1 mul_U2934(.A(n1515), .B(n3579), .Y(dpath_mulcore_array2_ain[72]));
AND2X1 mul_U2935(.A(n2055), .B(n4108), .Y(dpath_mulcore_array2_c2[70]));
AND2X1 mul_U2936(.A(n1516), .B(n3580), .Y(dpath_mulcore_array2_ain[71]));
AND2X1 mul_U2937(.A(n2056), .B(n4109), .Y(dpath_mulcore_array2_c2[69]));
AND2X1 mul_U2938(.A(n1517), .B(n3581), .Y(dpath_mulcore_array2_ain[70]));
AND2X1 mul_U2939(.A(n2057), .B(n4110), .Y(dpath_mulcore_array2_c2[68]));
AND2X1 mul_U2940(.A(n1518), .B(n3582), .Y(dpath_mulcore_array2_ain[69]));
INVX1 mul_U2941(.A(dpath_mulcore_array2_sc3_68__z), .Y(n10081));
AND2X1 mul_U2942(.A(n1444), .B(n3508), .Y(dpath_mulcore_array2_ain[68]));
INVX1 mul_U2943(.A(dpath_mulcore_array2_sc3_67__z), .Y(n10080));
AND2X1 mul_U2944(.A(n1445), .B(n3509), .Y(dpath_mulcore_array2_ain[67]));
INVX1 mul_U2945(.A(dpath_mulcore_array2_sc3_66__z), .Y(n10079));
AND2X1 mul_U2946(.A(n1446), .B(n3510), .Y(dpath_mulcore_array2_ain[66]));
INVX1 mul_U2947(.A(dpath_mulcore_array2_sc3_65__z), .Y(n10078));
AND2X1 mul_U2948(.A(n1447), .B(n3511), .Y(dpath_mulcore_array2_ain[65]));
INVX1 mul_U2949(.A(dpath_mulcore_array2_sc3_64__z), .Y(n10077));
AND2X1 mul_U2950(.A(n1448), .B(n3512), .Y(dpath_mulcore_array2_ain[64]));
INVX1 mul_U2951(.A(dpath_mulcore_array2_sc3_63__z), .Y(n10076));
AND2X1 mul_U2952(.A(n1449), .B(n3513), .Y(dpath_mulcore_array2_ain[63]));
INVX1 mul_U2953(.A(dpath_mulcore_array2_sc3_62__z), .Y(n10075));
AND2X1 mul_U2954(.A(n1450), .B(n3514), .Y(dpath_mulcore_array2_ain[62]));
INVX1 mul_U2955(.A(dpath_mulcore_array2_sc3_61__z), .Y(n10074));
AND2X1 mul_U2956(.A(n1451), .B(n3515), .Y(dpath_mulcore_array2_ain[61]));
INVX1 mul_U2957(.A(dpath_mulcore_array2_sc3_60__z), .Y(n10073));
AND2X1 mul_U2958(.A(n1452), .B(n3516), .Y(dpath_mulcore_array2_ain[60]));
INVX1 mul_U2959(.A(dpath_mulcore_array2_sc3_59__z), .Y(n10072));
AND2X1 mul_U2960(.A(n1453), .B(n3517), .Y(dpath_mulcore_array2_ain[59]));
INVX1 mul_U2961(.A(dpath_mulcore_array2_sc3_58__z), .Y(n10071));
AND2X1 mul_U2962(.A(n1454), .B(n3518), .Y(dpath_mulcore_array2_ain[58]));
INVX1 mul_U2963(.A(dpath_mulcore_array2_sc3_57__z), .Y(n10070));
AND2X1 mul_U2964(.A(n1455), .B(n3519), .Y(dpath_mulcore_array2_ain[57]));
INVX1 mul_U2965(.A(dpath_mulcore_array2_sc3_56__z), .Y(n10069));
AND2X1 mul_U2966(.A(n1456), .B(n3520), .Y(dpath_mulcore_array2_ain[56]));
INVX1 mul_U2967(.A(dpath_mulcore_array2_sc3_55__z), .Y(n10068));
AND2X1 mul_U2968(.A(n1457), .B(n3521), .Y(dpath_mulcore_array2_ain[55]));
INVX1 mul_U2969(.A(dpath_mulcore_array2_sc3_54__z), .Y(n10067));
AND2X1 mul_U2970(.A(n1458), .B(n3522), .Y(dpath_mulcore_array2_ain[54]));
INVX1 mul_U2971(.A(dpath_mulcore_array2_sc3_53__z), .Y(n10066));
AND2X1 mul_U2972(.A(n1459), .B(n3523), .Y(dpath_mulcore_array2_ain[53]));
INVX1 mul_U2973(.A(dpath_mulcore_array2_sc3_52__z), .Y(n10065));
AND2X1 mul_U2974(.A(n1460), .B(n3524), .Y(dpath_mulcore_array2_ain[52]));
INVX1 mul_U2975(.A(dpath_mulcore_array2_sc3_51__z), .Y(n10064));
AND2X1 mul_U2976(.A(n1461), .B(n3525), .Y(dpath_mulcore_array2_ain[51]));
INVX1 mul_U2977(.A(dpath_mulcore_array2_sc3_50__z), .Y(n10063));
AND2X1 mul_U2978(.A(n1462), .B(n3526), .Y(dpath_mulcore_array2_ain[50]));
INVX1 mul_U2979(.A(dpath_mulcore_array2_sc3_49__z), .Y(n10062));
AND2X1 mul_U2980(.A(n1463), .B(n3527), .Y(dpath_mulcore_array2_ain[49]));
INVX1 mul_U2981(.A(dpath_mulcore_array2_sc3_48__z), .Y(n10061));
AND2X1 mul_U2982(.A(n1464), .B(n3528), .Y(dpath_mulcore_array2_ain[48]));
INVX1 mul_U2983(.A(dpath_mulcore_array2_sc3_47__z), .Y(n10060));
AND2X1 mul_U2984(.A(n1465), .B(n3529), .Y(dpath_mulcore_array2_ain[47]));
INVX1 mul_U2985(.A(dpath_mulcore_array2_sc3_46__z), .Y(n10059));
AND2X1 mul_U2986(.A(n1466), .B(n3530), .Y(dpath_mulcore_array2_ain[46]));
INVX1 mul_U2987(.A(dpath_mulcore_array2_sc3_45__z), .Y(n10058));
AND2X1 mul_U2988(.A(n1467), .B(n3531), .Y(dpath_mulcore_array2_ain[45]));
INVX1 mul_U2989(.A(dpath_mulcore_array2_sc3_44__z), .Y(n10057));
AND2X1 mul_U2990(.A(n1468), .B(n3532), .Y(dpath_mulcore_array2_ain[44]));
INVX1 mul_U2991(.A(dpath_mulcore_array2_sc3_43__z), .Y(n10056));
AND2X1 mul_U2992(.A(n1469), .B(n3533), .Y(dpath_mulcore_array2_ain[43]));
INVX1 mul_U2993(.A(dpath_mulcore_array2_sc3_42__z), .Y(n10055));
AND2X1 mul_U2994(.A(n1470), .B(n3534), .Y(dpath_mulcore_array2_ain[42]));
INVX1 mul_U2995(.A(dpath_mulcore_array2_sc3_41__z), .Y(n10054));
AND2X1 mul_U2996(.A(n1471), .B(n3535), .Y(dpath_mulcore_array2_ain[41]));
INVX1 mul_U2997(.A(dpath_mulcore_array2_sc3_40__z), .Y(n10053));
AND2X1 mul_U2998(.A(n1472), .B(n3536), .Y(dpath_mulcore_array2_ain[40]));
INVX1 mul_U2999(.A(dpath_mulcore_array2_sc3_39__z), .Y(n10052));
AND2X1 mul_U3000(.A(n1473), .B(n3537), .Y(dpath_mulcore_array2_ain[39]));
INVX1 mul_U3001(.A(dpath_mulcore_array2_sc3_38__z), .Y(n10051));
AND2X1 mul_U3002(.A(n1474), .B(n3538), .Y(dpath_mulcore_array2_ain[38]));
INVX1 mul_U3003(.A(dpath_mulcore_array2_sc3_37__z), .Y(n10050));
AND2X1 mul_U3004(.A(n1475), .B(n3539), .Y(dpath_mulcore_array2_ain[37]));
INVX1 mul_U3005(.A(dpath_mulcore_array2_sc3_36__z), .Y(n10049));
AND2X1 mul_U3006(.A(n1476), .B(n3540), .Y(dpath_mulcore_array2_ain[36]));
INVX1 mul_U3007(.A(dpath_mulcore_array2_sc3_35__z), .Y(n10048));
AND2X1 mul_U3008(.A(n1477), .B(n3541), .Y(dpath_mulcore_array2_ain[35]));
INVX1 mul_U3009(.A(dpath_mulcore_array2_sc3_34__z), .Y(n10047));
AND2X1 mul_U3010(.A(n1478), .B(n3542), .Y(dpath_mulcore_array2_ain[34]));
INVX1 mul_U3011(.A(dpath_mulcore_array2_sc3_33__z), .Y(n10046));
AND2X1 mul_U3012(.A(n1479), .B(n3543), .Y(dpath_mulcore_array2_ain[33]));
INVX1 mul_U3013(.A(dpath_mulcore_array2_sc3_32__z), .Y(n10045));
AND2X1 mul_U3014(.A(n1480), .B(n3544), .Y(dpath_mulcore_array2_ain[32]));
INVX1 mul_U3015(.A(dpath_mulcore_array2_sc3_31__z), .Y(n10044));
AND2X1 mul_U3016(.A(n1481), .B(n3545), .Y(dpath_mulcore_array2_ain[31]));
INVX1 mul_U3017(.A(dpath_mulcore_array2_sc3_30__z), .Y(n10043));
AND2X1 mul_U3018(.A(n2394), .B(n4319), .Y(dpath_mulcore_array2_c3[29]));
AND2X1 mul_U3019(.A(n2396), .B(n4321), .Y(dpath_mulcore_array2_c3[28]));
AND2X1 mul_U3020(.A(n2398), .B(n4323), .Y(dpath_mulcore_array2_c3[27]));
AND2X1 mul_U3021(.A(n2400), .B(n4325), .Y(dpath_mulcore_array2_c3[26]));
AND2X1 mul_U3022(.A(n2402), .B(n4327), .Y(dpath_mulcore_array2_c3[25]));
AND2X1 mul_U3023(.A(n2404), .B(n4329), .Y(dpath_mulcore_array2_c3[24]));
AND2X1 mul_U3024(.A(n2406), .B(n4331), .Y(dpath_mulcore_array2_c3[23]));
AND2X1 mul_U3025(.A(n2408), .B(n4333), .Y(dpath_mulcore_array2_c3[22]));
AND2X1 mul_U3026(.A(n2410), .B(n4335), .Y(dpath_mulcore_array2_c3[21]));
INVX1 mul_U3027(.A(dpath_mulcore_array2_sc3_20__z), .Y(n10033));
AND2X1 mul_U3028(.A(n1911), .B(n3964), .Y(dpath_mulcore_array2_c3[19]));
AND2X1 mul_U3029(.A(n1912), .B(n3965), .Y(dpath_mulcore_array2_c3[18]));
AND2X1 mul_U3030(.A(n1913), .B(n3966), .Y(dpath_mulcore_array2_c3[17]));
AND2X1 mul_U3031(.A(n1914), .B(n3967), .Y(dpath_mulcore_array2_c3[16]));
AND2X1 mul_U3032(.A(n1915), .B(n3968), .Y(dpath_mulcore_array2_c3[15]));
AND2X1 mul_U3033(.A(n1938), .B(n3991), .Y(dpath_mulcore_array2_c2[13]));
AND2X1 mul_U3034(.A(n1939), .B(n3992), .Y(dpath_mulcore_array2_c2[12]));
AND2X1 mul_U3035(.A(n1940), .B(n3993), .Y(dpath_mulcore_array2_c2[11]));
AND2X1 mul_U3036(.A(n1941), .B(n3994), .Y(dpath_mulcore_array2_c2[10]));
AND2X1 mul_U3037(.A(n1942), .B(n3995), .Y(dpath_mulcore_array2_c2[9]));
AND2X1 mul_U3038(.A(n1943), .B(n3996), .Y(dpath_mulcore_array2_c2[8]));
AND2X1 mul_U3039(.A(n1944), .B(n3997), .Y(dpath_mulcore_array2_c2[7]));
AND2X1 mul_U3040(.A(n1945), .B(n3998), .Y(dpath_mulcore_array2_c2[6]));
AND2X1 mul_U3041(.A(n1946), .B(n3999), .Y(dpath_mulcore_array2_c2[5]));
AND2X1 mul_U3042(.A(dpath_mulcore_array2_s1[4]), .B(n7210), .Y(dpath_mulcore_array2_c2[4]));
AND2X1 mul_U3043(.A(dpath_mulcore_array2_s1[3]), .B(n7211), .Y(dpath_mulcore_array2_c2[3]));
AND2X1 mul_U3044(.A(dpath_mulcore_array2_s1[2]), .B(n7212), .Y(dpath_mulcore_array2_c2[2]));
AND2X1 mul_U3045(.A(dpath_mulcore_array2_s1[1]), .B(n7226), .Y(dpath_mulcore_array2_c2[1]));
AND2X1 mul_U3046(.A(dpath_mulcore_array2_s1[0]), .B(dpath_mulcore_array2_c1x2), .Y(dpath_mulcore_array2_c2[0]));
AND2X1 mul_U3047(.A(n1523), .B(n3587), .Y(dpath_mulcore_array2_ain[15]));
OR2X1 mul_U3048(.A(n5927), .B(n6055), .Y(dpath_areg[0]));
AND2X1 mul_U3049(.A(n3007), .B(n4683), .Y(dpath_n975));
AND2X1 mul_U3050(.A(n1505), .B(n3569), .Y(dpath_mulcore_array2_ain[0]));
AND2X1 mul_U3051(.A(n104), .B(n10614), .Y(dpath_mulcore_ary1_a0_I2_I1_63__net32));
OR2X1 mul_U3052(.A(n6172), .B(dpath_mulcore_b6[0]), .Y(n10614));
AND2X1 mul_U3053(.A(n103), .B(n10611), .Y(dpath_mulcore_ary1_a0_I2_I1_63__net046));
OR2X1 mul_U3054(.A(n6171), .B(dpath_mulcore_b7[0]), .Y(n10611));
AND2X1 mul_U3055(.A(n227), .B(n10987), .Y(dpath_mulcore_ary1_a0_I1_I2_net078));
OR2X1 mul_U3056(.A(n6297), .B(dpath_mulcore_b5[0]), .Y(n10987));
AND2X1 mul_U3057(.A(dpath_mulcore_ary1_a0_I1_I2_net38), .B(n4118), .Y(dpath_mulcore_ary1_a0_c1[66]));
OR2X1 mul_U3058(.A(n9476), .B(dpath_mulcore_b4[0]), .Y(n13667));
AND2X1 mul_U3059(.A(n228), .B(n10990), .Y(dpath_mulcore_ary1_a0_I1_I2_net8));
OR2X1 mul_U3060(.A(n6298), .B(dpath_mulcore_b5[0]), .Y(n10990));
AND2X1 mul_U3061(.A(n2065), .B(n4119), .Y(dpath_mulcore_ary1_a0_c1[65]));
AND2X1 mul_U3062(.A(n232), .B(n11002), .Y(dpath_mulcore_ary1_a0_I1_I2_net35));
OR2X1 mul_U3063(.A(n6302), .B(dpath_mulcore_b5[0]), .Y(n11002));
AND2X1 mul_U3064(.A(n2066), .B(n4120), .Y(dpath_mulcore_ary1_a0_c1[64]));
AND2X1 mul_U3065(.A(n229), .B(n10993), .Y(dpath_mulcore_ary1_a0_I1_I2_net15));
OR2X1 mul_U3066(.A(n6299), .B(dpath_mulcore_b5[0]), .Y(n10993));
AND2X1 mul_U3067(.A(n1134), .B(n3195), .Y(dpath_mulcore_ary1_a0_c1[63]));
AND2X1 mul_U3068(.A(n1135), .B(n3196), .Y(dpath_mulcore_ary1_a0_c1[62]));
AND2X1 mul_U3069(.A(n1136), .B(n3197), .Y(dpath_mulcore_ary1_a0_c1[61]));
AND2X1 mul_U3070(.A(n1137), .B(n3198), .Y(dpath_mulcore_ary1_a0_c1[60]));
AND2X1 mul_U3071(.A(n1138), .B(n3199), .Y(dpath_mulcore_ary1_a0_c1[59]));
AND2X1 mul_U3072(.A(n1139), .B(n3200), .Y(dpath_mulcore_ary1_a0_c1[58]));
AND2X1 mul_U3073(.A(n1140), .B(n3201), .Y(dpath_mulcore_ary1_a0_c1[57]));
AND2X1 mul_U3074(.A(n1141), .B(n3202), .Y(dpath_mulcore_ary1_a0_c1[56]));
AND2X1 mul_U3075(.A(n1142), .B(n3203), .Y(dpath_mulcore_ary1_a0_c1[55]));
AND2X1 mul_U3076(.A(n1143), .B(n3204), .Y(dpath_mulcore_ary1_a0_c1[54]));
AND2X1 mul_U3077(.A(n1144), .B(n3205), .Y(dpath_mulcore_ary1_a0_c1[53]));
AND2X1 mul_U3078(.A(n1145), .B(n3206), .Y(dpath_mulcore_ary1_a0_c1[52]));
AND2X1 mul_U3079(.A(n1146), .B(n3207), .Y(dpath_mulcore_ary1_a0_c1[51]));
AND2X1 mul_U3080(.A(n1147), .B(n3208), .Y(dpath_mulcore_ary1_a0_c1[50]));
AND2X1 mul_U3081(.A(n1148), .B(n3209), .Y(dpath_mulcore_ary1_a0_c1[49]));
AND2X1 mul_U3082(.A(n1149), .B(n3210), .Y(dpath_mulcore_ary1_a0_c1[48]));
AND2X1 mul_U3083(.A(n1150), .B(n3211), .Y(dpath_mulcore_ary1_a0_c1[47]));
AND2X1 mul_U3084(.A(n1151), .B(n3212), .Y(dpath_mulcore_ary1_a0_c1[46]));
AND2X1 mul_U3085(.A(n1152), .B(n3213), .Y(dpath_mulcore_ary1_a0_c1[45]));
AND2X1 mul_U3086(.A(n1153), .B(n3214), .Y(dpath_mulcore_ary1_a0_c1[44]));
AND2X1 mul_U3087(.A(n1154), .B(n3215), .Y(dpath_mulcore_ary1_a0_c1[43]));
AND2X1 mul_U3088(.A(n1155), .B(n3216), .Y(dpath_mulcore_ary1_a0_c1[42]));
AND2X1 mul_U3089(.A(n1156), .B(n3217), .Y(dpath_mulcore_ary1_a0_c1[41]));
AND2X1 mul_U3090(.A(n1157), .B(n3218), .Y(dpath_mulcore_ary1_a0_c1[40]));
AND2X1 mul_U3091(.A(n1158), .B(n3219), .Y(dpath_mulcore_ary1_a0_c1[39]));
AND2X1 mul_U3092(.A(n1159), .B(n3220), .Y(dpath_mulcore_ary1_a0_c1[38]));
AND2X1 mul_U3093(.A(n1160), .B(n3221), .Y(dpath_mulcore_ary1_a0_c1[37]));
AND2X1 mul_U3094(.A(n1161), .B(n3222), .Y(dpath_mulcore_ary1_a0_c1[36]));
AND2X1 mul_U3095(.A(n1162), .B(n3223), .Y(dpath_mulcore_ary1_a0_c1[35]));
AND2X1 mul_U3096(.A(n1163), .B(n3224), .Y(dpath_mulcore_ary1_a0_c1[34]));
AND2X1 mul_U3097(.A(n1164), .B(n3225), .Y(dpath_mulcore_ary1_a0_c1[33]));
AND2X1 mul_U3098(.A(n1165), .B(n3226), .Y(dpath_mulcore_ary1_a0_c1[32]));
AND2X1 mul_U3099(.A(n1166), .B(n3227), .Y(dpath_mulcore_ary1_a0_c1[31]));
AND2X1 mul_U3100(.A(n1167), .B(n3228), .Y(dpath_mulcore_ary1_a0_c1[30]));
AND2X1 mul_U3101(.A(n1168), .B(n3229), .Y(dpath_mulcore_ary1_a0_c1[29]));
AND2X1 mul_U3102(.A(n1169), .B(n3230), .Y(dpath_mulcore_ary1_a0_c1[28]));
AND2X1 mul_U3103(.A(n1170), .B(n3231), .Y(dpath_mulcore_ary1_a0_c1[27]));
AND2X1 mul_U3104(.A(n1171), .B(n3232), .Y(dpath_mulcore_ary1_a0_c1[26]));
AND2X1 mul_U3105(.A(n1172), .B(n3233), .Y(dpath_mulcore_ary1_a0_c1[25]));
AND2X1 mul_U3106(.A(n1173), .B(n3234), .Y(dpath_mulcore_ary1_a0_c1[24]));
AND2X1 mul_U3107(.A(n1174), .B(n3235), .Y(dpath_mulcore_ary1_a0_c1[23]));
AND2X1 mul_U3108(.A(n1175), .B(n3236), .Y(dpath_mulcore_ary1_a0_c1[22]));
AND2X1 mul_U3109(.A(n1176), .B(n3237), .Y(dpath_mulcore_ary1_a0_c1[21]));
AND2X1 mul_U3110(.A(n1177), .B(n3238), .Y(dpath_mulcore_ary1_a0_c1[20]));
AND2X1 mul_U3111(.A(n1178), .B(n3239), .Y(dpath_mulcore_ary1_a0_c1[19]));
AND2X1 mul_U3112(.A(n1179), .B(n3240), .Y(dpath_mulcore_ary1_a0_c1[18]));
AND2X1 mul_U3113(.A(n1180), .B(n3241), .Y(dpath_mulcore_ary1_a0_c1[17]));
AND2X1 mul_U3114(.A(n1181), .B(n3242), .Y(dpath_mulcore_ary1_a0_c1[16]));
AND2X1 mul_U3115(.A(n1182), .B(n3243), .Y(dpath_mulcore_ary1_a0_c1[15]));
AND2X1 mul_U3116(.A(n1183), .B(n3244), .Y(dpath_mulcore_ary1_a0_c1[14]));
AND2X1 mul_U3117(.A(n1184), .B(n3245), .Y(dpath_mulcore_ary1_a0_c1[13]));
AND2X1 mul_U3118(.A(n1185), .B(n3246), .Y(dpath_mulcore_ary1_a0_c1[12]));
AND2X1 mul_U3119(.A(n1186), .B(n3247), .Y(dpath_mulcore_ary1_a0_c1[11]));
AND2X1 mul_U3120(.A(n1187), .B(n3248), .Y(dpath_mulcore_ary1_a0_c1[10]));
AND2X1 mul_U3121(.A(n1188), .B(n3249), .Y(dpath_mulcore_ary1_a0_c1[9]));
AND2X1 mul_U3122(.A(n1189), .B(n3250), .Y(dpath_mulcore_ary1_a0_c1[8]));
AND2X1 mul_U3123(.A(n1190), .B(n3251), .Y(dpath_mulcore_ary1_a0_c1[7]));
AND2X1 mul_U3124(.A(n1245), .B(n3306), .Y(dpath_mulcore_ary1_a0_c0[12]));
AND2X1 mul_U3125(.A(n1191), .B(n3252), .Y(dpath_mulcore_ary1_a0_c1[6]));
AND2X1 mul_U3126(.A(n1246), .B(n3307), .Y(dpath_mulcore_ary1_a0_c0[11]));
AND2X1 mul_U3127(.A(n1192), .B(n3253), .Y(dpath_mulcore_ary1_a0_c1[5]));
OR2X1 mul_U3128(.A(n9729), .B(n5928), .Y(dpath_mulcore_ary1_a0_I1_I0_b1n_0));
INVX1 mul_U3129(.A(n11557), .Y(n9844));
OR2X1 mul_U3130(.A(n6488), .B(dpath_mulcore_b4[0]), .Y(n11557));
AND2X1 mul_U3131(.A(n414), .B(n11550), .Y(dpath_mulcore_ary1_a0_I1_I0_p0_2));
OR2X1 mul_U3132(.A(n6485), .B(dpath_mulcore_b3[0]), .Y(n11550));
OR2X1 mul_U3133(.A(n9723), .B(n5933), .Y(dpath_mulcore_ary1_a0_I0_I0_b1n_1));
INVX1 mul_U3134(.A(n12130), .Y(n9840));
OR2X1 mul_U3135(.A(n6680), .B(dpath_mulcore_b1[0]), .Y(n12130));
AND2X1 mul_U3136(.A(n603), .B(n12123), .Y(dpath_mulcore_ary1_a0_I0_I0_p0_2));
OR2X1 mul_U3137(.A(n6677), .B(dpath_mulcore_b0[0]), .Y(n12123));
INVX1 mul_U3138(.A(dpath_mulcore_op1_l[0]), .Y(n9855));
INVX1 mul_U3139(.A(dpath_mulcore_op1_l[63]), .Y(n10032));
AND2X1 mul_U3140(.A(n2477), .B(dpath_mulcore_ary1_a0_I2_I2_p0_64__n3), .Y(dpath_mulcore_ary1_a0_I2_I2_net47));
OR2X1 mul_U3141(.A(n9483), .B(dpath_mulcore_b6[0]), .Y(dpath_mulcore_ary1_a0_I2_I2_p0_64__n3));
AND2X1 mul_U3142(.A(n102), .B(n10608), .Y(dpath_mulcore_ary1_a0_I2_I2_net48));
OR2X1 mul_U3143(.A(n6170), .B(dpath_mulcore_b7[0]), .Y(n10608));
OR2X1 mul_U3144(.A(n9731), .B(n5959), .Y(dpath_mulcore_ary1_a0_b5n[0]));
AND2X1 mul_U3145(.A(n1247), .B(n3308), .Y(dpath_mulcore_ary1_a0_c0[10]));
AND2X1 mul_U3146(.A(n1193), .B(n3254), .Y(dpath_mulcore_ary1_a0_c1[4]));
AND2X1 mul_U3147(.A(n1248), .B(n3309), .Y(dpath_mulcore_ary1_a0_c0[9]));
AND2X1 mul_U3148(.A(n1251), .B(n3312), .Y(dpath_mulcore_ary1_a0_c0[6]));
AND2X1 mul_U3149(.A(n1252), .B(n3313), .Y(dpath_mulcore_ary1_a0_c0[5]));
INVX1 mul_U3150(.A(n11555), .Y(n9845));
OR2X1 mul_U3151(.A(n6487), .B(dpath_mulcore_b3[0]), .Y(n11555));
OR2X1 mul_U3152(.A(n9727), .B(n5930), .Y(dpath_mulcore_ary1_a0_I1_I0_b0n_0));
AND2X1 mul_U3153(.A(n1253), .B(n3314), .Y(dpath_mulcore_ary1_a0_c0[4]));
AND2X1 mul_U3154(.A(n1126), .B(n3187), .Y(dpath_mulcore_ary1_a0_c0[3]));
INVX1 mul_U3155(.A(acc_actc2), .Y(n9818));
INVX1 mul_U3156(.A(spu_mul_acc), .Y(n9814));
OR2X1 mul_U3157(.A(n5862), .B(n5990), .Y(dpath_mulcore_booth_b1_in0[2]));
AND2X1 mul_U3158(.A(n2812), .B(n4488), .Y(dpath_n320));
OR2X1 mul_U3159(.A(n9807), .B(dpath_mul_op2_d[2]), .Y(dpath_mulcore_booth_encode0_a_n44));
OR2X1 mul_U3160(.A(n10084), .B(dpath_mulcore_booth_b[34]), .Y(n18040));
AND2X1 mul_U3161(.A(n2469), .B(n4373), .Y(n18039));
AND2X1 mul_U3162(.A(n9807), .B(dpath_mulcore_booth_b0_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n74));
AND2X1 mul_U3163(.A(n10084), .B(dpath_mulcore_booth_b0_in1[2]), .Y(n18070));
OR2X1 mul_U3164(.A(n5840), .B(n5968), .Y(dpath_mulcore_booth_b2_in0[2]));
AND2X1 mul_U3165(.A(n2768), .B(n4444), .Y(dpath_n188));
AND2X1 mul_U3166(.A(n2468), .B(n4372), .Y(n18035));
AND2X1 mul_U3167(.A(n9809), .B(dpath_mul_op2_d[4]), .Y(dpath_mulcore_booth_encode0_a_n70));
AND2X1 mul_U3168(.A(n9808), .B(n9807), .Y(dpath_mulcore_booth_encode0_a_n69));
AND2X1 mul_U3169(.A(n10085), .B(n10084), .Y(n18065));
AND2X1 mul_U3170(.A(n10086), .B(dpath_mulcore_booth_b[36]), .Y(n18066));
OR2X1 mul_U3171(.A(n5834), .B(n5962), .Y(dpath_mulcore_booth_b3_in0[2]));
AND2X1 mul_U3172(.A(n2756), .B(n4432), .Y(dpath_n152));
AND2X1 mul_U3173(.A(n2467), .B(n4370), .Y(n18031));
AND2X1 mul_U3174(.A(n9811), .B(dpath_mul_op2_d[6]), .Y(dpath_mulcore_booth_encode0_a_n66));
AND2X1 mul_U3175(.A(n9810), .B(n9809), .Y(dpath_mulcore_booth_encode0_a_n65));
AND2X1 mul_U3176(.A(n10087), .B(n10086), .Y(n18061));
AND2X1 mul_U3177(.A(n10088), .B(dpath_mulcore_booth_b[38]), .Y(n18062));
OR2X1 mul_U3178(.A(n5832), .B(n5960), .Y(dpath_mulcore_booth_b4_in0[2]));
AND2X1 mul_U3179(.A(n2752), .B(n4428), .Y(dpath_n137));
AND2X1 mul_U3180(.A(n2466), .B(n4368), .Y(n18027));
AND2X1 mul_U3181(.A(n9813), .B(dpath_mul_op2_d[8]), .Y(dpath_mulcore_booth_encode0_a_n62));
AND2X1 mul_U3182(.A(n9812), .B(n9811), .Y(dpath_mulcore_booth_encode0_a_n61));
AND2X1 mul_U3183(.A(n10089), .B(n10088), .Y(n18057));
AND2X1 mul_U3184(.A(n10090), .B(dpath_mulcore_booth_b[40]), .Y(n18058));
OR2X1 mul_U3185(.A(n5893), .B(n6021), .Y(dpath_mulcore_booth_b5_in0[2]));
AND2X1 mul_U3186(.A(n2874), .B(n4550), .Y(dpath_n506));
AND2X1 mul_U3187(.A(n2465), .B(n4366), .Y(n18023));
AND2X1 mul_U3188(.A(n9788), .B(dpath_mul_op2_d[10]), .Y(dpath_mulcore_booth_encode0_a_n58));
AND2X1 mul_U3189(.A(n9787), .B(n9813), .Y(dpath_mulcore_booth_encode0_a_n57));
AND2X1 mul_U3190(.A(n10091), .B(n10090), .Y(n18053));
AND2X1 mul_U3191(.A(n10092), .B(dpath_mulcore_booth_b[42]), .Y(n18054));
OR2X1 mul_U3192(.A(n5891), .B(n6019), .Y(dpath_mulcore_booth_b6_in0[2]));
AND2X1 mul_U3193(.A(n2870), .B(n4546), .Y(dpath_n494));
AND2X1 mul_U3194(.A(n2464), .B(n4364), .Y(n18019));
AND2X1 mul_U3195(.A(n9790), .B(dpath_mul_op2_d[12]), .Y(dpath_mulcore_booth_encode0_a_n54));
AND2X1 mul_U3196(.A(n9789), .B(n9788), .Y(dpath_mulcore_booth_encode0_a_n53));
AND2X1 mul_U3197(.A(n10093), .B(n10092), .Y(n18049));
AND2X1 mul_U3198(.A(n10094), .B(dpath_mulcore_booth_b[44]), .Y(n18050));
OR2X1 mul_U3199(.A(n5889), .B(n6017), .Y(dpath_mulcore_booth_b7_in0[2]));
AND2X1 mul_U3200(.A(n2866), .B(n4542), .Y(dpath_n482));
OR2X1 mul_U3201(.A(n9790), .B(dpath_mulcore_booth_b7_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n21));
AND2X1 mul_U3202(.A(n18017), .B(n4362), .Y(n18015));
OR2X1 mul_U3203(.A(n10094), .B(dpath_mulcore_booth_b7_in1[2]), .Y(n18017));
AND2X1 mul_U3204(.A(n9791), .B(n9790), .Y(dpath_mulcore_booth_encode0_a_n49));
AND2X1 mul_U3205(.A(n10095), .B(n10094), .Y(n18045));
OR2X1 mul_U3206(.A(n5887), .B(n6015), .Y(dpath_mulcore_booth_b8_in0[2]));
AND2X1 mul_U3207(.A(n2862), .B(n4538), .Y(dpath_n470));
OR2X1 mul_U3208(.A(n9793), .B(dpath_mul_op2_d[16]), .Y(n17949));
INVX1 mul_U3209(.A(dpath_mulcore_booth_b7_in0[2]), .Y(n9792));
INVX1 mul_U3210(.A(dpath_mulcore_booth_b7_in1[2]), .Y(n10096));
AND2X1 mul_U3211(.A(n18077), .B(n4382), .Y(n18075));
OR2X1 mul_U3212(.A(n10097), .B(dpath_mulcore_booth_b[48]), .Y(n18077));
AND2X1 mul_U3213(.A(n9793), .B(dpath_mulcore_booth_b7_in0[2]), .Y(n18009));
AND2X1 mul_U3214(.A(n10097), .B(dpath_mulcore_booth_b7_in1[2]), .Y(n18137));
OR2X1 mul_U3215(.A(n5885), .B(n6013), .Y(dpath_mulcore_booth_b9_in0[2]));
AND2X1 mul_U3216(.A(n2858), .B(n4534), .Y(dpath_n458));
OR2X1 mul_U3217(.A(n9794), .B(dpath_mul_op2_d[18]), .Y(n17976));
OR2X1 mul_U3218(.A(n10098), .B(dpath_mulcore_booth_b[50]), .Y(n18104));
AND2X1 mul_U3219(.A(n2476), .B(n4395), .Y(n18103));
AND2X1 mul_U3220(.A(n9794), .B(dpath_mulcore_booth_b8_in0[2]), .Y(n18006));
AND2X1 mul_U3221(.A(n10098), .B(dpath_mulcore_booth_b8_in1[2]), .Y(n18134));
OR2X1 mul_U3222(.A(n5882), .B(n6010), .Y(dpath_mulcore_booth_b10_in0[2]));
AND2X1 mul_U3223(.A(n2852), .B(n4528), .Y(dpath_n440));
AND2X1 mul_U3224(.A(n2475), .B(n4394), .Y(n18099));
AND2X1 mul_U3225(.A(n9797), .B(dpath_mul_op2_d[20]), .Y(n18002));
AND2X1 mul_U3226(.A(n9796), .B(n9794), .Y(n18001));
AND2X1 mul_U3227(.A(n10099), .B(n10098), .Y(n18129));
AND2X1 mul_U3228(.A(n10100), .B(dpath_mulcore_booth_b[52]), .Y(n18130));
OR2X1 mul_U3229(.A(n5880), .B(n6008), .Y(dpath_mulcore_booth_b11_in0[2]));
AND2X1 mul_U3230(.A(n2848), .B(n4524), .Y(dpath_n428));
AND2X1 mul_U3231(.A(n2474), .B(n4392), .Y(n18095));
AND2X1 mul_U3232(.A(n9799), .B(dpath_mul_op2_d[22]), .Y(n17998));
AND2X1 mul_U3233(.A(n9798), .B(n9797), .Y(n17997));
AND2X1 mul_U3234(.A(n10101), .B(n10100), .Y(n18125));
AND2X1 mul_U3235(.A(n10102), .B(dpath_mulcore_booth_b[54]), .Y(n18126));
OR2X1 mul_U3236(.A(n5878), .B(n6006), .Y(dpath_mulcore_booth_b12_in0[2]));
AND2X1 mul_U3237(.A(n2844), .B(n4520), .Y(dpath_n416));
AND2X1 mul_U3238(.A(n2473), .B(n4390), .Y(n18091));
AND2X1 mul_U3239(.A(n9801), .B(dpath_mul_op2_d[24]), .Y(n17994));
AND2X1 mul_U3240(.A(n9800), .B(n9799), .Y(n17993));
AND2X1 mul_U3241(.A(n10103), .B(n10102), .Y(n18121));
AND2X1 mul_U3242(.A(n10104), .B(dpath_mulcore_booth_b[56]), .Y(n18122));
OR2X1 mul_U3243(.A(n5876), .B(n6004), .Y(dpath_mulcore_booth_b13_in0[2]));
AND2X1 mul_U3244(.A(n2840), .B(n4516), .Y(dpath_n404));
AND2X1 mul_U3245(.A(n2472), .B(n4388), .Y(n18087));
AND2X1 mul_U3246(.A(n9803), .B(dpath_mul_op2_d[26]), .Y(n17990));
AND2X1 mul_U3247(.A(n9802), .B(n9801), .Y(n17989));
AND2X1 mul_U3248(.A(n10105), .B(n10104), .Y(n18117));
AND2X1 mul_U3249(.A(n10106), .B(dpath_mulcore_booth_b[58]), .Y(n18118));
OR2X1 mul_U3250(.A(n5874), .B(n6002), .Y(dpath_mulcore_booth_b14_in0[2]));
AND2X1 mul_U3251(.A(n2836), .B(n4512), .Y(dpath_n392));
AND2X1 mul_U3252(.A(n2471), .B(n4386), .Y(n18083));
AND2X1 mul_U3253(.A(n9805), .B(dpath_mul_op2_d[28]), .Y(n17986));
AND2X1 mul_U3254(.A(n9804), .B(n9803), .Y(n17985));
AND2X1 mul_U3255(.A(n10107), .B(n10106), .Y(n18113));
AND2X1 mul_U3256(.A(n10108), .B(dpath_mulcore_booth_b[60]), .Y(n18114));
OR2X1 mul_U3257(.A(n9805), .B(dpath_mulcore_booth_b15_in0[2]), .Y(n17953));
AND2X1 mul_U3258(.A(n18081), .B(n4384), .Y(n18079));
OR2X1 mul_U3259(.A(n10108), .B(dpath_mulcore_booth_b15_in1[2]), .Y(n18081));
AND2X1 mul_U3260(.A(n9806), .B(n9805), .Y(n17981));
AND2X1 mul_U3261(.A(n10109), .B(n10108), .Y(n18109));
AND2X1 mul_U3262(.A(n1254), .B(n3315), .Y(dpath_mulcore_ary1_a1_c2[63]));
OR2X1 mul_U3263(.A(n9485), .B(dpath_mulcore_b13[0]), .Y(n13681));
OR2X1 mul_U3264(.A(dpath_mulcore_ary1_a1_s_2[71]), .B(dpath_mulcore_ary1_a1_s1[64]), .Y(n17027));
OR2X1 mul_U3265(.A(dpath_mulcore_ary1_a1_s_2[70]), .B(n9369), .Y(n17052));
INVX1 mul_U3266(.A(dpath_mulcore_ary1_a1_s1[64]), .Y(n10025));
AND2X1 mul_U3267(.A(n1746), .B(n3800), .Y(dpath_mulcore_ary1_a1_c_1[69]));
OR2X1 mul_U3268(.A(dpath_mulcore_ary1_a1_s_2[69]), .B(n9370), .Y(n17059));
AND2X1 mul_U3269(.A(n1747), .B(n3801), .Y(dpath_mulcore_ary1_a1_c_1[68]));
OR2X1 mul_U3270(.A(dpath_mulcore_ary1_a1_s_2[68]), .B(n9371), .Y(n17066));
AND2X1 mul_U3271(.A(n1748), .B(n3802), .Y(dpath_mulcore_ary1_a1_c_1[67]));
OR2X1 mul_U3272(.A(dpath_mulcore_ary1_a1_s_2[67]), .B(n9372), .Y(n17073));
AND2X1 mul_U3273(.A(n1749), .B(n3803), .Y(dpath_mulcore_ary1_a1_c_1[66]));
OR2X1 mul_U3274(.A(dpath_mulcore_ary1_a1_s_2[66]), .B(n9373), .Y(n17080));
AND2X1 mul_U3275(.A(n1750), .B(n3804), .Y(dpath_mulcore_ary1_a1_c_1[65]));
OR2X1 mul_U3276(.A(dpath_mulcore_ary1_a1_s_2[65]), .B(n9374), .Y(n17087));
AND2X1 mul_U3277(.A(n1751), .B(n3805), .Y(dpath_mulcore_ary1_a1_c_1[64]));
OR2X1 mul_U3278(.A(dpath_mulcore_ary1_a1_s_2[64]), .B(n9375), .Y(n17094));
AND2X1 mul_U3279(.A(n1752), .B(n3806), .Y(dpath_mulcore_ary1_a1_c_1[63]));
OR2X1 mul_U3280(.A(dpath_mulcore_ary1_a1_s_2[63]), .B(n9376), .Y(n17101));
AND2X1 mul_U3281(.A(n1753), .B(n3807), .Y(dpath_mulcore_ary1_a1_c_1[62]));
OR2X1 mul_U3282(.A(dpath_mulcore_ary1_a1_s_2[62]), .B(n9377), .Y(n17108));
AND2X1 mul_U3283(.A(n1754), .B(n3808), .Y(dpath_mulcore_ary1_a1_c_1[61]));
OR2X1 mul_U3284(.A(dpath_mulcore_ary1_a1_s_2[61]), .B(n9378), .Y(n17115));
AND2X1 mul_U3285(.A(n1755), .B(n3809), .Y(dpath_mulcore_ary1_a1_c_1[60]));
OR2X1 mul_U3286(.A(dpath_mulcore_ary1_a1_s_2[60]), .B(n9379), .Y(n17122));
AND2X1 mul_U3287(.A(n1756), .B(n3810), .Y(dpath_mulcore_ary1_a1_c_1[59]));
OR2X1 mul_U3288(.A(dpath_mulcore_ary1_a1_s_2[59]), .B(n9380), .Y(n17129));
AND2X1 mul_U3289(.A(n1757), .B(n3811), .Y(dpath_mulcore_ary1_a1_c_1[58]));
OR2X1 mul_U3290(.A(dpath_mulcore_ary1_a1_s_2[58]), .B(n9381), .Y(n17136));
AND2X1 mul_U3291(.A(n1758), .B(n3812), .Y(dpath_mulcore_ary1_a1_c_1[57]));
OR2X1 mul_U3292(.A(dpath_mulcore_ary1_a1_s_2[57]), .B(n9382), .Y(n17143));
AND2X1 mul_U3293(.A(n1759), .B(n3813), .Y(dpath_mulcore_ary1_a1_c_1[56]));
OR2X1 mul_U3294(.A(dpath_mulcore_ary1_a1_s_2[56]), .B(n9383), .Y(n17150));
AND2X1 mul_U3295(.A(n1760), .B(n3814), .Y(dpath_mulcore_ary1_a1_c_1[55]));
OR2X1 mul_U3296(.A(dpath_mulcore_ary1_a1_s_2[55]), .B(n9384), .Y(n17157));
AND2X1 mul_U3297(.A(n1761), .B(n3815), .Y(dpath_mulcore_ary1_a1_c_1[54]));
OR2X1 mul_U3298(.A(dpath_mulcore_ary1_a1_s_2[54]), .B(n9385), .Y(n17164));
AND2X1 mul_U3299(.A(n1762), .B(n3816), .Y(dpath_mulcore_ary1_a1_c_1[53]));
OR2X1 mul_U3300(.A(dpath_mulcore_ary1_a1_s_2[53]), .B(n9386), .Y(n17171));
AND2X1 mul_U3301(.A(n1763), .B(n3817), .Y(dpath_mulcore_ary1_a1_c_1[52]));
OR2X1 mul_U3302(.A(dpath_mulcore_ary1_a1_s_2[52]), .B(n9387), .Y(n17178));
AND2X1 mul_U3303(.A(n1764), .B(n3818), .Y(dpath_mulcore_ary1_a1_c_1[51]));
OR2X1 mul_U3304(.A(dpath_mulcore_ary1_a1_s_2[51]), .B(n9388), .Y(n17185));
AND2X1 mul_U3305(.A(n1765), .B(n3819), .Y(dpath_mulcore_ary1_a1_c_1[50]));
OR2X1 mul_U3306(.A(dpath_mulcore_ary1_a1_s_2[50]), .B(n9389), .Y(n17192));
AND2X1 mul_U3307(.A(n1766), .B(n3820), .Y(dpath_mulcore_ary1_a1_c_1[49]));
OR2X1 mul_U3308(.A(dpath_mulcore_ary1_a1_s_2[49]), .B(n9390), .Y(n17199));
AND2X1 mul_U3309(.A(n1767), .B(n3821), .Y(dpath_mulcore_ary1_a1_c_1[48]));
OR2X1 mul_U3310(.A(dpath_mulcore_ary1_a1_s_2[48]), .B(n9391), .Y(n17206));
AND2X1 mul_U3311(.A(n1768), .B(n3822), .Y(dpath_mulcore_ary1_a1_c_1[47]));
OR2X1 mul_U3312(.A(dpath_mulcore_ary1_a1_s_2[47]), .B(n9392), .Y(n17213));
AND2X1 mul_U3313(.A(n1769), .B(n3823), .Y(dpath_mulcore_ary1_a1_c_1[46]));
OR2X1 mul_U3314(.A(dpath_mulcore_ary1_a1_s_2[46]), .B(n9393), .Y(n17220));
AND2X1 mul_U3315(.A(n1770), .B(n3824), .Y(dpath_mulcore_ary1_a1_c_1[45]));
OR2X1 mul_U3316(.A(dpath_mulcore_ary1_a1_s_2[45]), .B(n9394), .Y(n17227));
AND2X1 mul_U3317(.A(n1771), .B(n3825), .Y(dpath_mulcore_ary1_a1_c_1[44]));
OR2X1 mul_U3318(.A(dpath_mulcore_ary1_a1_s_2[44]), .B(n9395), .Y(n17234));
AND2X1 mul_U3319(.A(n1772), .B(n3826), .Y(dpath_mulcore_ary1_a1_c_1[43]));
OR2X1 mul_U3320(.A(dpath_mulcore_ary1_a1_s_2[43]), .B(n9396), .Y(n17241));
AND2X1 mul_U3321(.A(n1773), .B(n3827), .Y(dpath_mulcore_ary1_a1_c_1[42]));
OR2X1 mul_U3322(.A(dpath_mulcore_ary1_a1_s_2[42]), .B(n9397), .Y(n17248));
AND2X1 mul_U3323(.A(n1774), .B(n3828), .Y(dpath_mulcore_ary1_a1_c_1[41]));
OR2X1 mul_U3324(.A(dpath_mulcore_ary1_a1_s_2[41]), .B(n9398), .Y(n17255));
AND2X1 mul_U3325(.A(n1775), .B(n3829), .Y(dpath_mulcore_ary1_a1_c_1[40]));
OR2X1 mul_U3326(.A(dpath_mulcore_ary1_a1_s_2[40]), .B(n9399), .Y(n17262));
AND2X1 mul_U3327(.A(n1776), .B(n3830), .Y(dpath_mulcore_ary1_a1_c_1[39]));
OR2X1 mul_U3328(.A(dpath_mulcore_ary1_a1_s_2[39]), .B(n9400), .Y(n17269));
AND2X1 mul_U3329(.A(n1777), .B(n3831), .Y(dpath_mulcore_ary1_a1_c_1[38]));
OR2X1 mul_U3330(.A(dpath_mulcore_ary1_a1_s_2[38]), .B(n9401), .Y(n17276));
AND2X1 mul_U3331(.A(n1778), .B(n3832), .Y(dpath_mulcore_ary1_a1_c_1[37]));
OR2X1 mul_U3332(.A(dpath_mulcore_ary1_a1_s_2[37]), .B(n9402), .Y(n17283));
AND2X1 mul_U3333(.A(n1779), .B(n3833), .Y(dpath_mulcore_ary1_a1_c_1[36]));
OR2X1 mul_U3334(.A(dpath_mulcore_ary1_a1_s_2[36]), .B(n9403), .Y(n17290));
AND2X1 mul_U3335(.A(n1780), .B(n3834), .Y(dpath_mulcore_ary1_a1_c_1[35]));
OR2X1 mul_U3336(.A(dpath_mulcore_ary1_a1_s_2[35]), .B(n9404), .Y(n17297));
AND2X1 mul_U3337(.A(n1781), .B(n3835), .Y(dpath_mulcore_ary1_a1_c_1[34]));
OR2X1 mul_U3338(.A(dpath_mulcore_ary1_a1_s_2[34]), .B(n9405), .Y(n17304));
AND2X1 mul_U3339(.A(n1782), .B(n3836), .Y(dpath_mulcore_ary1_a1_c_1[33]));
OR2X1 mul_U3340(.A(dpath_mulcore_ary1_a1_s_2[33]), .B(n9406), .Y(n17311));
AND2X1 mul_U3341(.A(n1783), .B(n3837), .Y(dpath_mulcore_ary1_a1_c_1[32]));
OR2X1 mul_U3342(.A(dpath_mulcore_ary1_a1_s_2[32]), .B(n9407), .Y(n17318));
AND2X1 mul_U3343(.A(n1784), .B(n3838), .Y(dpath_mulcore_ary1_a1_c_1[31]));
OR2X1 mul_U3344(.A(dpath_mulcore_ary1_a1_s_2[31]), .B(n9408), .Y(n17325));
AND2X1 mul_U3345(.A(n1785), .B(n3839), .Y(dpath_mulcore_ary1_a1_c_1[30]));
OR2X1 mul_U3346(.A(dpath_mulcore_ary1_a1_s_2[30]), .B(n9409), .Y(n17332));
AND2X1 mul_U3347(.A(n1786), .B(n3840), .Y(dpath_mulcore_ary1_a1_c_1[29]));
OR2X1 mul_U3348(.A(dpath_mulcore_ary1_a1_s_2[29]), .B(n9410), .Y(n17339));
AND2X1 mul_U3349(.A(n1787), .B(n3841), .Y(dpath_mulcore_ary1_a1_c_1[28]));
OR2X1 mul_U3350(.A(dpath_mulcore_ary1_a1_s_2[28]), .B(n9411), .Y(n17346));
AND2X1 mul_U3351(.A(n1788), .B(n3842), .Y(dpath_mulcore_ary1_a1_c_1[27]));
OR2X1 mul_U3352(.A(dpath_mulcore_ary1_a1_s_2[27]), .B(n9412), .Y(n17353));
AND2X1 mul_U3353(.A(n1789), .B(n3843), .Y(dpath_mulcore_ary1_a1_c_1[26]));
OR2X1 mul_U3354(.A(dpath_mulcore_ary1_a1_s_2[26]), .B(n9413), .Y(n17360));
AND2X1 mul_U3355(.A(n1790), .B(n3844), .Y(dpath_mulcore_ary1_a1_c_1[25]));
OR2X1 mul_U3356(.A(dpath_mulcore_ary1_a1_s_2[25]), .B(n9414), .Y(n17367));
AND2X1 mul_U3357(.A(n1791), .B(n3845), .Y(dpath_mulcore_ary1_a1_c_1[24]));
OR2X1 mul_U3358(.A(dpath_mulcore_ary1_a1_s_2[24]), .B(n9415), .Y(n17374));
AND2X1 mul_U3359(.A(n1792), .B(n3846), .Y(dpath_mulcore_ary1_a1_c_1[23]));
OR2X1 mul_U3360(.A(dpath_mulcore_ary1_a1_s_2[23]), .B(n9416), .Y(n17381));
AND2X1 mul_U3361(.A(n1793), .B(n3847), .Y(dpath_mulcore_ary1_a1_c_1[22]));
OR2X1 mul_U3362(.A(dpath_mulcore_ary1_a1_s_2[22]), .B(n9417), .Y(n17388));
AND2X1 mul_U3363(.A(n1794), .B(n3848), .Y(dpath_mulcore_ary1_a1_c_1[21]));
OR2X1 mul_U3364(.A(dpath_mulcore_ary1_a1_s_2[21]), .B(n9418), .Y(n17395));
AND2X1 mul_U3365(.A(n1795), .B(n3849), .Y(dpath_mulcore_ary1_a1_c_1[20]));
OR2X1 mul_U3366(.A(dpath_mulcore_ary1_a1_s_2[20]), .B(n9419), .Y(n17402));
AND2X1 mul_U3367(.A(n1796), .B(n3850), .Y(dpath_mulcore_ary1_a1_c_1[19]));
OR2X1 mul_U3368(.A(dpath_mulcore_ary1_a1_s_2[19]), .B(n9420), .Y(n17409));
AND2X1 mul_U3369(.A(n1797), .B(n3851), .Y(dpath_mulcore_ary1_a1_c_1[18]));
OR2X1 mul_U3370(.A(dpath_mulcore_ary1_a1_s_2[18]), .B(n9421), .Y(n17416));
AND2X1 mul_U3371(.A(n1798), .B(n3852), .Y(dpath_mulcore_ary1_a1_c_1[17]));
OR2X1 mul_U3372(.A(dpath_mulcore_ary1_a1_s_2[17]), .B(n9422), .Y(n17423));
AND2X1 mul_U3373(.A(n1799), .B(n3853), .Y(dpath_mulcore_ary1_a1_c_1[16]));
OR2X1 mul_U3374(.A(dpath_mulcore_ary1_a1_s_2[16]), .B(n9423), .Y(n17430));
AND2X1 mul_U3375(.A(n1800), .B(n3854), .Y(dpath_mulcore_ary1_a1_c_1[15]));
OR2X1 mul_U3376(.A(dpath_mulcore_ary1_a1_s_2[15]), .B(n9424), .Y(n17437));
AND2X1 mul_U3377(.A(n1801), .B(n3855), .Y(dpath_mulcore_ary1_a1_c_1[14]));
OR2X1 mul_U3378(.A(dpath_mulcore_ary1_a1_s_2[14]), .B(dpath_mulcore_ary1_a1_c_1[13]), .Y(n17444));
AND2X1 mul_U3379(.A(dpath_mulcore_ary1_a1_s0[13]), .B(n7204), .Y(dpath_mulcore_ary1_a1_c_1[13]));
OR2X1 mul_U3380(.A(dpath_mulcore_ary1_a1_s_2[13]), .B(dpath_mulcore_ary1_a1_c_1[12]), .Y(n17451));
AND2X1 mul_U3381(.A(dpath_mulcore_ary1_a1_s0[12]), .B(n7205), .Y(dpath_mulcore_ary1_a1_c_1[12]));
OR2X1 mul_U3382(.A(dpath_mulcore_ary1_a1_s_2[12]), .B(dpath_mulcore_ary1_a1_c_1[11]), .Y(n17458));
AND2X1 mul_U3383(.A(dpath_mulcore_ary1_a1_s0[11]), .B(n7206), .Y(dpath_mulcore_ary1_a1_c_1[11]));
OR2X1 mul_U3384(.A(dpath_mulcore_ary1_a1_s_2[11]), .B(dpath_mulcore_ary1_a1_c_1[10]), .Y(n17465));
AND2X1 mul_U3385(.A(n1130), .B(n3191), .Y(dpath_mulcore_ary1_a1_c1[3]));
AND2X1 mul_U3386(.A(n919), .B(n13081), .Y(dpath_mulcore_ary1_a1_I1_I0_p0_1));
OR2X1 mul_U3387(.A(n6998), .B(dpath_mulcore_b11[0]), .Y(n13081));
OR2X1 mul_U3388(.A(n13723), .B(n5943), .Y(dpath_mulcore_ary1_a1_I1_I0_b0n));
AND2X1 mul_U3389(.A(n7405), .B(n9832), .Y(n13723));
AND2X1 mul_U3390(.A(n1133), .B(n3194), .Y(dpath_mulcore_ary1_a1_c0[2]));
OR2X1 mul_U3391(.A(n9739), .B(n5944), .Y(dpath_mulcore_ary1_a1_I0_I0_b1n_0));
OR2X1 mul_U3392(.A(n9478), .B(dpath_mulcore_b15[0]), .Y(n13677));
AND2X1 mul_U3393(.A(n1438), .B(n3499), .Y(dpath_mulcore_ary1_a1_c2[64]));
AND2X1 mul_U3394(.A(n1742), .B(n3796), .Y(dpath_mulcore_ary1_a1_c_2[75]));
AND2X1 mul_U3395(.A(n1743), .B(n3797), .Y(dpath_mulcore_ary1_a1_c_2[74]));
AND2X1 mul_U3396(.A(n1744), .B(n3798), .Y(dpath_mulcore_ary1_a1_c_2[73]));
AND2X1 mul_U3397(.A(n1745), .B(n3799), .Y(dpath_mulcore_ary1_a1_c_2[72]));
AND2X1 mul_U3398(.A(n1741), .B(n3795), .Y(dpath_mulcore_ary1_a1_c_2[71]));
AND2X1 mul_U3399(.A(n1672), .B(n3731), .Y(dpath_mulcore_ary1_a1_c_2[70]));
AND2X1 mul_U3400(.A(n1673), .B(n3732), .Y(dpath_mulcore_ary1_a1_c_2[69]));
AND2X1 mul_U3401(.A(n1674), .B(n3733), .Y(dpath_mulcore_ary1_a1_c_2[68]));
AND2X1 mul_U3402(.A(n1675), .B(n3734), .Y(dpath_mulcore_ary1_a1_c_2[67]));
AND2X1 mul_U3403(.A(n1676), .B(n3735), .Y(dpath_mulcore_ary1_a1_c_2[66]));
AND2X1 mul_U3404(.A(n1677), .B(n3736), .Y(dpath_mulcore_ary1_a1_c_2[65]));
AND2X1 mul_U3405(.A(n1678), .B(n3737), .Y(dpath_mulcore_ary1_a1_c_2[64]));
AND2X1 mul_U3406(.A(n1679), .B(n3738), .Y(dpath_mulcore_ary1_a1_c_2[63]));
AND2X1 mul_U3407(.A(n1680), .B(n3739), .Y(dpath_mulcore_ary1_a1_c_2[62]));
AND2X1 mul_U3408(.A(n1681), .B(n3740), .Y(dpath_mulcore_ary1_a1_c_2[61]));
AND2X1 mul_U3409(.A(n1682), .B(n3741), .Y(dpath_mulcore_ary1_a1_c_2[60]));
AND2X1 mul_U3410(.A(n1683), .B(n3742), .Y(dpath_mulcore_ary1_a1_c_2[59]));
AND2X1 mul_U3411(.A(n1684), .B(n3743), .Y(dpath_mulcore_ary1_a1_c_2[58]));
AND2X1 mul_U3412(.A(n1685), .B(n3744), .Y(dpath_mulcore_ary1_a1_c_2[57]));
AND2X1 mul_U3413(.A(n1686), .B(n3745), .Y(dpath_mulcore_ary1_a1_c_2[56]));
AND2X1 mul_U3414(.A(n1687), .B(n3746), .Y(dpath_mulcore_ary1_a1_c_2[55]));
AND2X1 mul_U3415(.A(n1688), .B(n3747), .Y(dpath_mulcore_ary1_a1_c_2[54]));
AND2X1 mul_U3416(.A(n1689), .B(n3748), .Y(dpath_mulcore_ary1_a1_c_2[53]));
AND2X1 mul_U3417(.A(n1690), .B(n3749), .Y(dpath_mulcore_ary1_a1_c_2[52]));
AND2X1 mul_U3418(.A(n1691), .B(n3750), .Y(dpath_mulcore_ary1_a1_c_2[51]));
AND2X1 mul_U3419(.A(n1692), .B(n3751), .Y(dpath_mulcore_ary1_a1_c_2[50]));
AND2X1 mul_U3420(.A(n1693), .B(n3752), .Y(dpath_mulcore_ary1_a1_c_2[49]));
AND2X1 mul_U3421(.A(n1694), .B(n3753), .Y(dpath_mulcore_ary1_a1_c_2[48]));
AND2X1 mul_U3422(.A(n1695), .B(n3754), .Y(dpath_mulcore_ary1_a1_c_2[47]));
AND2X1 mul_U3423(.A(n1696), .B(n3755), .Y(dpath_mulcore_ary1_a1_c_2[46]));
AND2X1 mul_U3424(.A(n1697), .B(n3756), .Y(dpath_mulcore_ary1_a1_c_2[45]));
AND2X1 mul_U3425(.A(n1698), .B(n3757), .Y(dpath_mulcore_ary1_a1_c_2[44]));
AND2X1 mul_U3426(.A(n1699), .B(n3758), .Y(dpath_mulcore_ary1_a1_c_2[43]));
AND2X1 mul_U3427(.A(n1700), .B(n3759), .Y(dpath_mulcore_ary1_a1_c_2[42]));
AND2X1 mul_U3428(.A(n1701), .B(n3760), .Y(dpath_mulcore_ary1_a1_c_2[41]));
AND2X1 mul_U3429(.A(n1702), .B(n3761), .Y(dpath_mulcore_ary1_a1_c_2[40]));
AND2X1 mul_U3430(.A(n1703), .B(n3762), .Y(dpath_mulcore_ary1_a1_c_2[39]));
AND2X1 mul_U3431(.A(n1704), .B(n3763), .Y(dpath_mulcore_ary1_a1_c_2[38]));
AND2X1 mul_U3432(.A(n1705), .B(n3764), .Y(dpath_mulcore_ary1_a1_c_2[37]));
AND2X1 mul_U3433(.A(n1706), .B(n3765), .Y(dpath_mulcore_ary1_a1_c_2[36]));
AND2X1 mul_U3434(.A(n1707), .B(n3766), .Y(dpath_mulcore_ary1_a1_c_2[35]));
AND2X1 mul_U3435(.A(n1708), .B(n3767), .Y(dpath_mulcore_ary1_a1_c_2[34]));
AND2X1 mul_U3436(.A(n1709), .B(n3768), .Y(dpath_mulcore_ary1_a1_c_2[33]));
AND2X1 mul_U3437(.A(n1710), .B(n3769), .Y(dpath_mulcore_ary1_a1_c_2[32]));
AND2X1 mul_U3438(.A(n1711), .B(n3770), .Y(dpath_mulcore_ary1_a1_c_2[31]));
AND2X1 mul_U3439(.A(n1712), .B(n3771), .Y(dpath_mulcore_ary1_a1_c_2[30]));
AND2X1 mul_U3440(.A(n1713), .B(n3772), .Y(dpath_mulcore_ary1_a1_c_2[29]));
AND2X1 mul_U3441(.A(n1714), .B(n3773), .Y(dpath_mulcore_ary1_a1_c_2[28]));
AND2X1 mul_U3442(.A(n1715), .B(n3774), .Y(dpath_mulcore_ary1_a1_c_2[27]));
AND2X1 mul_U3443(.A(n1716), .B(n3775), .Y(dpath_mulcore_ary1_a1_c_2[26]));
AND2X1 mul_U3444(.A(n1717), .B(n3776), .Y(dpath_mulcore_ary1_a1_c_2[25]));
AND2X1 mul_U3445(.A(n1718), .B(n3777), .Y(dpath_mulcore_ary1_a1_c_2[24]));
AND2X1 mul_U3446(.A(n1719), .B(n3778), .Y(dpath_mulcore_ary1_a1_c_2[23]));
AND2X1 mul_U3447(.A(n1720), .B(n3779), .Y(dpath_mulcore_ary1_a1_c_2[22]));
AND2X1 mul_U3448(.A(n1721), .B(n3780), .Y(dpath_mulcore_ary1_a1_c_2[21]));
AND2X1 mul_U3449(.A(n1722), .B(n3781), .Y(dpath_mulcore_ary1_a1_c_2[20]));
AND2X1 mul_U3450(.A(n1723), .B(n3782), .Y(dpath_mulcore_ary1_a1_c_2[19]));
AND2X1 mul_U3451(.A(n1724), .B(n3783), .Y(dpath_mulcore_ary1_a1_c_2[18]));
AND2X1 mul_U3452(.A(n1725), .B(n3784), .Y(dpath_mulcore_ary1_a1_c_2[17]));
AND2X1 mul_U3453(.A(n1726), .B(n3785), .Y(dpath_mulcore_ary1_a1_c_2[16]));
AND2X1 mul_U3454(.A(n1727), .B(n3786), .Y(dpath_mulcore_ary1_a1_c_2[15]));
AND2X1 mul_U3455(.A(n1728), .B(n3787), .Y(dpath_mulcore_ary1_a1_c_2[14]));
AND2X1 mul_U3456(.A(n1729), .B(n3788), .Y(dpath_mulcore_ary1_a1_c_2[13]));
AND2X1 mul_U3457(.A(n1730), .B(n3789), .Y(dpath_mulcore_ary1_a1_c_2[12]));
AND2X1 mul_U3458(.A(n1731), .B(n3790), .Y(dpath_mulcore_ary1_a1_c_2[11]));
AND2X1 mul_U3459(.A(dpath_mulcore_ary1_a1_s0[10]), .B(n7207), .Y(dpath_mulcore_ary1_a1_c_1[10]));
AND2X1 mul_U3460(.A(n1735), .B(n3792), .Y(dpath_mulcore_ary1_a1_c_1[9]));
AND2X1 mul_U3461(.A(n1736), .B(n3793), .Y(dpath_mulcore_ary1_a1_c_1[8]));
AND2X1 mul_U3462(.A(n1802), .B(n3856), .Y(dpath_mulcore_ary1_a1_c_1[7]));
OR2X1 mul_U3463(.A(n9741), .B(n5952), .Y(dpath_mulcore_ary1_a1_b2n[1]));
OR2X1 mul_U3464(.A(n9741), .B(n5953), .Y(dpath_mulcore_ary1_a1_b2n[0]));
INVX1 mul_U3465(.A(n9497), .Y(n9579));
AND2X1 mul_U3466(.A(n2829), .B(n4505), .Y(dpath_n375));
OR2X1 mul_U3467(.A(n10083), .B(dpath_mulcore_booth_b[32]), .Y(n18013));
INVX1 mul_U3468(.A(dpath_mulcore_booth_b[31]), .Y(n10082));
OR2X1 mul_U3469(.A(n9795), .B(dpath_mul_op2_d[0]), .Y(dpath_mulcore_booth_encode0_a_n17));
AND2X1 mul_U3470(.A(n10083), .B(dpath_mulcore_booth_b[31]), .Y(n18073));
OR2X1 mul_U3471(.A(n5884), .B(n6012), .Y(dpath_mulcore_booth_b0_in0[2]));
AND2X1 mul_U3472(.A(n2856), .B(n4532), .Y(dpath_n452));
INVX1 mul_U3473(.A(dpath_mul_op2_d[0]), .Y(n9786));
OR2X1 mul_U3474(.A(n9311), .B(dpath_mulcore_addin_sum[96]), .Y(n10578));
OR2X1 mul_U3475(.A(n9310), .B(dpath_mulcore_addin_sum[95]), .Y(n10573));
OR2X1 mul_U3476(.A(n9309), .B(dpath_mulcore_addin_sum[94]), .Y(n10568));
OR2X1 mul_U3477(.A(n9308), .B(dpath_mulcore_addin_sum[93]), .Y(n10563));
OR2X1 mul_U3478(.A(n9307), .B(dpath_mulcore_addin_sum[92]), .Y(n10558));
OR2X1 mul_U3479(.A(n9306), .B(dpath_mulcore_addin_sum[91]), .Y(n10553));
OR2X1 mul_U3480(.A(n9305), .B(dpath_mulcore_addin_sum[90]), .Y(n10546));
OR2X1 mul_U3481(.A(n9304), .B(dpath_mulcore_addin_sum[89]), .Y(n10541));
OR2X1 mul_U3482(.A(n9303), .B(dpath_mulcore_addin_sum[88]), .Y(n10536));
OR2X1 mul_U3483(.A(n9302), .B(dpath_mulcore_addin_sum[87]), .Y(n10531));
OR2X1 mul_U3484(.A(n9301), .B(dpath_mulcore_addin_sum[86]), .Y(n10526));
OR2X1 mul_U3485(.A(n9300), .B(dpath_mulcore_addin_sum[85]), .Y(n10521));
OR2X1 mul_U3486(.A(n9299), .B(dpath_mulcore_addin_sum[84]), .Y(n10516));
OR2X1 mul_U3487(.A(n9298), .B(dpath_mulcore_addin_sum[83]), .Y(n10511));
OR2X1 mul_U3488(.A(n9297), .B(dpath_mulcore_addin_sum[82]), .Y(n10506));
OR2X1 mul_U3489(.A(n9296), .B(dpath_mulcore_addin_sum[81]), .Y(n10501));
OR2X1 mul_U3490(.A(n9295), .B(dpath_mulcore_addin_sum[80]), .Y(n10494));
OR2X1 mul_U3491(.A(n9294), .B(dpath_mulcore_addin_sum[79]), .Y(n10489));
OR2X1 mul_U3492(.A(n9293), .B(dpath_mulcore_addin_sum[78]), .Y(n10484));
OR2X1 mul_U3493(.A(n9292), .B(dpath_mulcore_addin_sum[77]), .Y(n10479));
OR2X1 mul_U3494(.A(n9291), .B(dpath_mulcore_addin_sum[76]), .Y(n10474));
OR2X1 mul_U3495(.A(n9290), .B(dpath_mulcore_addin_sum[75]), .Y(n10469));
OR2X1 mul_U3496(.A(n9289), .B(dpath_mulcore_addin_sum[74]), .Y(n10464));
OR2X1 mul_U3497(.A(n9288), .B(dpath_mulcore_addin_sum[73]), .Y(n10459));
OR2X1 mul_U3498(.A(n9287), .B(dpath_mulcore_addin_sum[72]), .Y(n10454));
OR2X1 mul_U3499(.A(n9286), .B(dpath_mulcore_addin_sum[71]), .Y(n10449));
OR2X1 mul_U3500(.A(n9285), .B(dpath_mulcore_addin_sum[70]), .Y(n10442));
OR2X1 mul_U3501(.A(n9284), .B(dpath_mulcore_addin_sum[69]), .Y(n10437));
OR2X1 mul_U3502(.A(n9283), .B(dpath_mulcore_addin_sum[68]), .Y(n10432));
OR2X1 mul_U3503(.A(n9282), .B(dpath_mulcore_addin_sum[67]), .Y(n10427));
OR2X1 mul_U3504(.A(n9281), .B(dpath_mulcore_addin_sum[66]), .Y(n10422));
OR2X1 mul_U3505(.A(n9280), .B(dpath_mulcore_addin_sum[65]), .Y(n10417));
OR2X1 mul_U3506(.A(n9279), .B(dpath_mulcore_addin_sum[64]), .Y(n10412));
OR2X1 mul_U3507(.A(n9278), .B(dpath_mulcore_addin_sum[63]), .Y(n10407));
OR2X1 mul_U3508(.A(n9277), .B(dpath_mulcore_addin_sum[62]), .Y(n10402));
OR2X1 mul_U3509(.A(n9276), .B(dpath_mulcore_addin_sum[61]), .Y(n10397));
OR2X1 mul_U3510(.A(n9275), .B(dpath_mulcore_addin_sum[60]), .Y(n10390));
OR2X1 mul_U3511(.A(n9274), .B(dpath_mulcore_addin_sum[59]), .Y(n10385));
OR2X1 mul_U3512(.A(n9273), .B(dpath_mulcore_addin_sum[58]), .Y(n10380));
OR2X1 mul_U3513(.A(n9272), .B(dpath_mulcore_addin_sum[57]), .Y(n10375));
OR2X1 mul_U3514(.A(n9271), .B(dpath_mulcore_addin_sum[56]), .Y(n10370));
OR2X1 mul_U3515(.A(n9270), .B(dpath_mulcore_addin_sum[55]), .Y(n10365));
OR2X1 mul_U3516(.A(n9269), .B(dpath_mulcore_addin_sum[54]), .Y(n10360));
OR2X1 mul_U3517(.A(n9268), .B(dpath_mulcore_addin_sum[53]), .Y(n10355));
OR2X1 mul_U3518(.A(n9267), .B(dpath_mulcore_addin_sum[52]), .Y(n10350));
OR2X1 mul_U3519(.A(n9266), .B(dpath_mulcore_addin_sum[51]), .Y(n10345));
OR2X1 mul_U3520(.A(n9265), .B(dpath_mulcore_addin_sum[50]), .Y(n10338));
OR2X1 mul_U3521(.A(n9264), .B(dpath_mulcore_addin_sum[49]), .Y(n10333));
OR2X1 mul_U3522(.A(n9263), .B(dpath_mulcore_addin_sum[48]), .Y(n10328));
OR2X1 mul_U3523(.A(n9262), .B(dpath_mulcore_addin_sum[47]), .Y(n10323));
OR2X1 mul_U3524(.A(n9261), .B(dpath_mulcore_addin_sum[46]), .Y(n10318));
OR2X1 mul_U3525(.A(n9260), .B(dpath_mulcore_addin_sum[45]), .Y(n10313));
OR2X1 mul_U3526(.A(n9259), .B(dpath_mulcore_addin_sum[44]), .Y(n10308));
OR2X1 mul_U3527(.A(n9258), .B(dpath_mulcore_addin_sum[43]), .Y(n10303));
OR2X1 mul_U3528(.A(n9257), .B(dpath_mulcore_addin_sum[42]), .Y(n10298));
OR2X1 mul_U3529(.A(n9234), .B(dpath_mulcore_addin_sum[41]), .Y(n10293));
OR2X1 mul_U3530(.A(n9233), .B(dpath_mulcore_addin_sum[40]), .Y(n10290));
OR2X1 mul_U3531(.A(n9232), .B(dpath_mulcore_addin_sum[39]), .Y(n10287));
OR2X1 mul_U3532(.A(n9231), .B(dpath_mulcore_addin_sum[38]), .Y(n10284));
OR2X1 mul_U3533(.A(n9230), .B(dpath_mulcore_addin_sum[37]), .Y(n10281));
OR2X1 mul_U3534(.A(n9229), .B(dpath_mulcore_addin_sum[36]), .Y(n10278));
OR2X1 mul_U3535(.A(n9228), .B(dpath_mulcore_addin_sum[35]), .Y(n10275));
OR2X1 mul_U3536(.A(n9227), .B(dpath_mulcore_addin_sum[34]), .Y(n10272));
OR2X1 mul_U3537(.A(n9226), .B(dpath_mulcore_addin_sum[33]), .Y(n10269));
OR2X1 mul_U3538(.A(dpath_mulcore_addin_cout[31]), .B(dpath_mulcore_addin_sum[32]), .Y(n10266));
OR2X1 mul_U3539(.A(n9256), .B(dpath_mulcore_addin_sum[31]), .Y(n10248));
OR2X1 mul_U3540(.A(n9255), .B(dpath_mulcore_addin_sum[30]), .Y(n10243));
OR2X1 mul_U3541(.A(n9254), .B(dpath_mulcore_addin_sum[29]), .Y(n10238));
OR2X1 mul_U3542(.A(n9253), .B(dpath_mulcore_addin_sum[28]), .Y(n10231));
OR2X1 mul_U3543(.A(n9252), .B(dpath_mulcore_addin_sum[27]), .Y(n10226));
OR2X1 mul_U3544(.A(n9251), .B(dpath_mulcore_addin_sum[26]), .Y(n10221));
OR2X1 mul_U3545(.A(n9250), .B(dpath_mulcore_addin_sum[25]), .Y(n10216));
OR2X1 mul_U3546(.A(n9249), .B(dpath_mulcore_addin_sum[24]), .Y(n10211));
OR2X1 mul_U3547(.A(n9248), .B(dpath_mulcore_addin_sum[23]), .Y(n10206));
OR2X1 mul_U3548(.A(n9247), .B(dpath_mulcore_addin_sum[22]), .Y(n10201));
OR2X1 mul_U3549(.A(n9246), .B(dpath_mulcore_addin_sum[21]), .Y(n10196));
OR2X1 mul_U3550(.A(n9245), .B(dpath_mulcore_addin_sum[20]), .Y(n10191));
OR2X1 mul_U3551(.A(n9244), .B(dpath_mulcore_addin_sum[19]), .Y(n10186));
OR2X1 mul_U3552(.A(n9243), .B(dpath_mulcore_addin_sum[18]), .Y(n10179));
OR2X1 mul_U3553(.A(n9242), .B(dpath_mulcore_addin_sum[17]), .Y(n10174));
OR2X1 mul_U3554(.A(n9241), .B(dpath_mulcore_addin_sum[16]), .Y(n10169));
OR2X1 mul_U3555(.A(n9240), .B(dpath_mulcore_addin_sum[15]), .Y(n10164));
OR2X1 mul_U3556(.A(n9239), .B(dpath_mulcore_addin_sum[14]), .Y(n10159));
OR2X1 mul_U3557(.A(n9238), .B(dpath_mulcore_addin_sum[13]), .Y(n10154));
OR2X1 mul_U3558(.A(n9237), .B(dpath_mulcore_addin_sum[12]), .Y(n10149));
OR2X1 mul_U3559(.A(n9236), .B(dpath_mulcore_addin_sum[11]), .Y(n10144));
OR2X1 mul_U3560(.A(n9235), .B(dpath_mulcore_addin_sum[10]), .Y(n10139));
OR2X1 mul_U3561(.A(n9225), .B(dpath_mulcore_addin_sum[9]), .Y(n10134));
OR2X1 mul_U3562(.A(n9224), .B(dpath_mulcore_addin_sum[8]), .Y(n10131));
OR2X1 mul_U3563(.A(n9223), .B(dpath_mulcore_addin_sum[7]), .Y(n10128));
OR2X1 mul_U3564(.A(n9222), .B(dpath_mulcore_addin_sum[6]), .Y(n10125));
OR2X1 mul_U3565(.A(n9221), .B(dpath_mulcore_addin_sum[5]), .Y(n10122));
OR2X1 mul_U3566(.A(n9220), .B(dpath_mulcore_addin_sum[4]), .Y(n10119));
OR2X1 mul_U3567(.A(n9219), .B(dpath_mulcore_addin_sum[3]), .Y(n10116));
OR2X1 mul_U3568(.A(n9218), .B(dpath_mulcore_addin_sum[2]), .Y(n10113));
OR2X1 mul_U3569(.A(dpath_mulcore_addin_sum[1]), .B(n10184), .Y(n10110));
INVX1 mul_U3570(.A(n9498), .Y(n9580));
AND2X1 mul_U3571(.A(dpath_mulcore_a1s[80]), .B(dpath_mulcore_a1c[79]), .Y(dpath_mulcore_array2_c2[96]));
AND2X1 mul_U3572(.A(dpath_mulcore_a1s[79]), .B(dpath_mulcore_a1c[78]), .Y(dpath_mulcore_array2_c2[95]));
AND2X1 mul_U3573(.A(dpath_mulcore_a1s[78]), .B(dpath_mulcore_a1c[77]), .Y(dpath_mulcore_array2_c2[94]));
AND2X1 mul_U3574(.A(dpath_mulcore_a1s[77]), .B(dpath_mulcore_a1c[76]), .Y(dpath_mulcore_array2_c2[93]));
AND2X1 mul_U3575(.A(dpath_mulcore_a1s[76]), .B(dpath_mulcore_a1c[75]), .Y(dpath_mulcore_array2_c2[92]));
AND2X1 mul_U3576(.A(dpath_mulcore_a1s[75]), .B(dpath_mulcore_a1c[74]), .Y(dpath_mulcore_array2_c2[91]));
AND2X1 mul_U3577(.A(dpath_mulcore_a1s[74]), .B(dpath_mulcore_a1c[73]), .Y(dpath_mulcore_array2_c2[90]));
AND2X1 mul_U3578(.A(dpath_mulcore_a1s[73]), .B(dpath_mulcore_a1c[72]), .Y(dpath_mulcore_array2_c2[89]));
AND2X1 mul_U3579(.A(dpath_mulcore_a1s[72]), .B(dpath_mulcore_a1c[71]), .Y(dpath_mulcore_array2_c2[88]));
AND2X1 mul_U3580(.A(dpath_mulcore_a1s[71]), .B(dpath_mulcore_a1c[70]), .Y(dpath_mulcore_array2_c2[87]));
AND2X1 mul_U3581(.A(dpath_mulcore_a1s[70]), .B(dpath_mulcore_a1c[69]), .Y(dpath_mulcore_array2_c2[86]));
AND2X1 mul_U3582(.A(dpath_mulcore_a1s[69]), .B(dpath_mulcore_a1c[68]), .Y(dpath_mulcore_array2_c2[85]));
AND2X1 mul_U3583(.A(dpath_mulcore_a1s[68]), .B(dpath_mulcore_a1c[67]), .Y(dpath_mulcore_array2_c2[84]));
AND2X1 mul_U3584(.A(n1892), .B(n3945), .Y(dpath_mulcore_array2_c2[83]));
AND2X1 mul_U3585(.A(n1947), .B(n4000), .Y(dpath_mulcore_array2_c2[82]));
AND2X1 mul_U3586(.A(dpath_mulcore_array2_s2[81]), .B(n7213), .Y(dpath_mulcore_array2_c3[81]));
AND2X1 mul_U3587(.A(dpath_mulcore_array2_s2[80]), .B(n7214), .Y(dpath_mulcore_array2_c3[80]));
AND2X1 mul_U3588(.A(dpath_mulcore_array2_s2[79]), .B(n7215), .Y(dpath_mulcore_array2_c3[79]));
AND2X1 mul_U3589(.A(dpath_mulcore_array2_s2[78]), .B(n7216), .Y(dpath_mulcore_array2_c3[78]));
AND2X1 mul_U3590(.A(dpath_mulcore_array2_s2[77]), .B(n7217), .Y(dpath_mulcore_array2_c3[77]));
AND2X1 mul_U3591(.A(dpath_mulcore_array2_s2[76]), .B(n7218), .Y(dpath_mulcore_array2_c3[76]));
AND2X1 mul_U3592(.A(dpath_mulcore_array2_s2[75]), .B(n7219), .Y(dpath_mulcore_array2_c3[75]));
AND2X1 mul_U3593(.A(dpath_mulcore_array2_s2[74]), .B(n7220), .Y(dpath_mulcore_array2_c3[74]));
AND2X1 mul_U3594(.A(dpath_mulcore_array2_s2[73]), .B(n7221), .Y(dpath_mulcore_array2_c3[73]));
AND2X1 mul_U3595(.A(dpath_mulcore_array2_s2[72]), .B(n7222), .Y(dpath_mulcore_array2_c3[72]));
AND2X1 mul_U3596(.A(dpath_mulcore_array2_s2[71]), .B(n7223), .Y(dpath_mulcore_array2_c3[71]));
AND2X1 mul_U3597(.A(dpath_mulcore_array2_s2[70]), .B(n7224), .Y(dpath_mulcore_array2_c3[70]));
AND2X1 mul_U3598(.A(dpath_mulcore_array2_s2[69]), .B(n7225), .Y(dpath_mulcore_array2_c3[69]));
AND2X1 mul_U3599(.A(n2317), .B(n4242), .Y(dpath_mulcore_array2_c3[68]));
AND2X1 mul_U3600(.A(n2318), .B(n4243), .Y(dpath_mulcore_array2_c3[67]));
AND2X1 mul_U3601(.A(n2320), .B(n4245), .Y(dpath_mulcore_array2_c3[66]));
AND2X1 mul_U3602(.A(n2322), .B(n4247), .Y(dpath_mulcore_array2_c3[65]));
AND2X1 mul_U3603(.A(n2324), .B(n4249), .Y(dpath_mulcore_array2_c3[64]));
AND2X1 mul_U3604(.A(n2326), .B(n4251), .Y(dpath_mulcore_array2_c3[63]));
AND2X1 mul_U3605(.A(n2328), .B(n4253), .Y(dpath_mulcore_array2_c3[62]));
AND2X1 mul_U3606(.A(n2330), .B(n4255), .Y(dpath_mulcore_array2_c3[61]));
AND2X1 mul_U3607(.A(n2332), .B(n4257), .Y(dpath_mulcore_array2_c3[60]));
AND2X1 mul_U3608(.A(n2334), .B(n4259), .Y(dpath_mulcore_array2_c3[59]));
AND2X1 mul_U3609(.A(n2336), .B(n4261), .Y(dpath_mulcore_array2_c3[58]));
AND2X1 mul_U3610(.A(n2338), .B(n4263), .Y(dpath_mulcore_array2_c3[57]));
AND2X1 mul_U3611(.A(n2340), .B(n4265), .Y(dpath_mulcore_array2_c3[56]));
AND2X1 mul_U3612(.A(n2342), .B(n4267), .Y(dpath_mulcore_array2_c3[55]));
AND2X1 mul_U3613(.A(n2344), .B(n4269), .Y(dpath_mulcore_array2_c3[54]));
AND2X1 mul_U3614(.A(n2346), .B(n4271), .Y(dpath_mulcore_array2_c3[53]));
AND2X1 mul_U3615(.A(n2348), .B(n4273), .Y(dpath_mulcore_array2_c3[52]));
AND2X1 mul_U3616(.A(n2350), .B(n4275), .Y(dpath_mulcore_array2_c3[51]));
AND2X1 mul_U3617(.A(n2352), .B(n4277), .Y(dpath_mulcore_array2_c3[50]));
AND2X1 mul_U3618(.A(n2354), .B(n4279), .Y(dpath_mulcore_array2_c3[49]));
AND2X1 mul_U3619(.A(n2356), .B(n4281), .Y(dpath_mulcore_array2_c3[48]));
AND2X1 mul_U3620(.A(n2358), .B(n4283), .Y(dpath_mulcore_array2_c3[47]));
AND2X1 mul_U3621(.A(n2360), .B(n4285), .Y(dpath_mulcore_array2_c3[46]));
AND2X1 mul_U3622(.A(n2362), .B(n4287), .Y(dpath_mulcore_array2_c3[45]));
AND2X1 mul_U3623(.A(n2364), .B(n4289), .Y(dpath_mulcore_array2_c3[44]));
AND2X1 mul_U3624(.A(n2366), .B(n4291), .Y(dpath_mulcore_array2_c3[43]));
AND2X1 mul_U3625(.A(n2368), .B(n4293), .Y(dpath_mulcore_array2_c3[42]));
AND2X1 mul_U3626(.A(n2370), .B(n4295), .Y(dpath_mulcore_array2_c3[41]));
AND2X1 mul_U3627(.A(n2372), .B(n4297), .Y(dpath_mulcore_array2_c3[40]));
AND2X1 mul_U3628(.A(n2374), .B(n4299), .Y(dpath_mulcore_array2_c3[39]));
AND2X1 mul_U3629(.A(n2376), .B(n4301), .Y(dpath_mulcore_array2_c3[38]));
AND2X1 mul_U3630(.A(n2378), .B(n4303), .Y(dpath_mulcore_array2_c3[37]));
AND2X1 mul_U3631(.A(n2380), .B(n4305), .Y(dpath_mulcore_array2_c3[36]));
AND2X1 mul_U3632(.A(n2382), .B(n4307), .Y(dpath_mulcore_array2_c3[35]));
AND2X1 mul_U3633(.A(n2384), .B(n4309), .Y(dpath_mulcore_array2_c3[34]));
AND2X1 mul_U3634(.A(n2386), .B(n4311), .Y(dpath_mulcore_array2_c3[33]));
AND2X1 mul_U3635(.A(n2388), .B(n4313), .Y(dpath_mulcore_array2_c3[32]));
AND2X1 mul_U3636(.A(n2390), .B(n4315), .Y(dpath_mulcore_array2_c3[31]));
AND2X1 mul_U3637(.A(n2392), .B(n4317), .Y(dpath_mulcore_array2_c3[30]));
INVX1 mul_U3638(.A(n9496), .Y(n9575));
INVX1 mul_U3639(.A(n9497), .Y(n9578));
INVX1 mul_U3640(.A(n9675), .Y(n9707));
INVX1 mul_U3641(.A(n9676), .Y(n9708));
INVX1 mul_U3642(.A(n9676), .Y(n9709));
INVX1 mul_U3643(.A(n9676), .Y(n9710));
INVX1 mul_U3644(.A(n9677), .Y(n9711));
INVX1 mul_U3645(.A(n9677), .Y(n9712));
INVX1 mul_U3646(.A(n9677), .Y(n9713));
INVX1 mul_U3647(.A(n9696), .Y(n9694));
AND2X1 mul_U3648(.A(n1846), .B(n3900), .Y(dpath_mulcore_pcout[29]));
AND2X1 mul_U3649(.A(n1847), .B(n3901), .Y(dpath_mulcore_pcout[28]));
AND2X1 mul_U3650(.A(n1848), .B(n3902), .Y(dpath_mulcore_pcout[27]));
AND2X1 mul_U3651(.A(n1849), .B(n3903), .Y(dpath_mulcore_pcout[26]));
AND2X1 mul_U3652(.A(n1850), .B(n3904), .Y(dpath_mulcore_pcout[25]));
AND2X1 mul_U3653(.A(n1851), .B(n3905), .Y(dpath_mulcore_pcout[24]));
AND2X1 mul_U3654(.A(n1852), .B(n3906), .Y(dpath_mulcore_pcout[23]));
AND2X1 mul_U3655(.A(n1853), .B(n3907), .Y(dpath_mulcore_pcout[22]));
AND2X1 mul_U3656(.A(n1854), .B(n3908), .Y(dpath_mulcore_pcout[21]));
AND2X1 mul_U3657(.A(n1855), .B(n3909), .Y(dpath_mulcore_pcout[20]));
AND2X1 mul_U3658(.A(n2058), .B(n4111), .Y(dpath_mulcore_pcout[19]));
AND2X1 mul_U3659(.A(n2059), .B(n4112), .Y(dpath_mulcore_pcout[18]));
AND2X1 mul_U3660(.A(n2060), .B(n4113), .Y(dpath_mulcore_pcout[17]));
AND2X1 mul_U3661(.A(n2061), .B(n4114), .Y(dpath_mulcore_pcout[16]));
AND2X1 mul_U3662(.A(n1916), .B(n3969), .Y(dpath_mulcore_pcout[14]));
INVX1 mul_U3663(.A(n9696), .Y(n9695));
AND2X1 mul_U3664(.A(n1917), .B(n3970), .Y(dpath_mulcore_pcout[13]));
AND2X1 mul_U3665(.A(n1918), .B(n3971), .Y(dpath_mulcore_pcout[12]));
AND2X1 mul_U3666(.A(n1919), .B(n3972), .Y(dpath_mulcore_pcout[11]));
AND2X1 mul_U3667(.A(n1920), .B(n3973), .Y(dpath_mulcore_pcout[10]));
AND2X1 mul_U3668(.A(n1921), .B(n3974), .Y(dpath_mulcore_pcout[9]));
AND2X1 mul_U3669(.A(n1922), .B(n3975), .Y(dpath_mulcore_pcout[8]));
INVX1 mul_U3670(.A(n9673), .Y(n9702));
AND2X1 mul_U3671(.A(n1923), .B(n3976), .Y(dpath_mulcore_pcout[7]));
INVX1 mul_U3672(.A(n9699), .Y(n9690));
INVX1 mul_U3673(.A(n9674), .Y(n9703));
AND2X1 mul_U3674(.A(n1924), .B(n3977), .Y(dpath_mulcore_pcout[6]));
INVX1 mul_U3675(.A(n9699), .Y(n9689));
AND2X1 mul_U3676(.A(n1925), .B(n3978), .Y(dpath_mulcore_pcout[5]));
INVX1 mul_U3677(.A(n9698), .Y(n9693));
INVX1 mul_U3678(.A(n9674), .Y(n9704));
AND2X1 mul_U3679(.A(n1882), .B(n3936), .Y(dpath_mulcore_pcout[4]));
INVX1 mul_U3680(.A(n9674), .Y(n9705));
AND2X1 mul_U3681(.A(n1883), .B(n3937), .Y(dpath_mulcore_pcout[3]));
INVX1 mul_U3682(.A(n9700), .Y(n9688));
INVX1 mul_U3683(.A(n9675), .Y(n9706));
AND2X1 mul_U3684(.A(n1884), .B(n3938), .Y(dpath_mulcore_pcout[2]));
INVX1 mul_U3685(.A(n9700), .Y(n9687));
AND2X1 mul_U3686(.A(n1885), .B(n3939), .Y(dpath_mulcore_pcout[1]));
INVX1 mul_U3687(.A(n9701), .Y(n9686));
AND2X1 mul_U3688(.A(n7407), .B(dpath_mulcore_array2_s2[0]), .Y(dpath_mulcore_pcout[0]));
OR2X1 mul_U3689(.A(n9484), .B(dpath_mulcore_b5[0]), .Y(n13665));
OR2X1 mul_U3690(.A(dpath_mulcore_ary1_a0_s_2[71]), .B(dpath_mulcore_ary1_a0_s1[64]), .Y(dpath_mulcore_ary1_a0_sc3_71__n4));
OR2X1 mul_U3691(.A(dpath_mulcore_ary1_a0_s_2[70]), .B(n9313), .Y(n16608));
INVX1 mul_U3692(.A(dpath_mulcore_ary1_a0_s1[64]), .Y(n10026));
AND2X1 mul_U3693(.A(n1612), .B(n3671), .Y(dpath_mulcore_ary1_a0_c_1[69]));
OR2X1 mul_U3694(.A(dpath_mulcore_ary1_a0_s_2[69]), .B(n9314), .Y(n16615));
AND2X1 mul_U3695(.A(n1613), .B(n3672), .Y(dpath_mulcore_ary1_a0_c_1[68]));
OR2X1 mul_U3696(.A(dpath_mulcore_ary1_a0_s_2[68]), .B(n9315), .Y(n16622));
AND2X1 mul_U3697(.A(n1614), .B(n3673), .Y(dpath_mulcore_ary1_a0_c_1[67]));
OR2X1 mul_U3698(.A(dpath_mulcore_ary1_a0_s_2[67]), .B(n9316), .Y(n16629));
AND2X1 mul_U3699(.A(n1615), .B(n3674), .Y(dpath_mulcore_ary1_a0_c_1[66]));
OR2X1 mul_U3700(.A(dpath_mulcore_ary1_a0_s_2[66]), .B(n9317), .Y(n16636));
AND2X1 mul_U3701(.A(n1616), .B(n3675), .Y(dpath_mulcore_ary1_a0_c_1[65]));
OR2X1 mul_U3702(.A(dpath_mulcore_ary1_a0_s_2[65]), .B(n9318), .Y(n16643));
AND2X1 mul_U3703(.A(n1617), .B(n3676), .Y(dpath_mulcore_ary1_a0_c_1[64]));
OR2X1 mul_U3704(.A(dpath_mulcore_ary1_a0_s_2[64]), .B(n9319), .Y(n16650));
AND2X1 mul_U3705(.A(n1618), .B(n3677), .Y(dpath_mulcore_ary1_a0_c_1[63]));
OR2X1 mul_U3706(.A(dpath_mulcore_ary1_a0_s_2[63]), .B(n9320), .Y(n16657));
AND2X1 mul_U3707(.A(n1619), .B(n3678), .Y(dpath_mulcore_ary1_a0_c_1[62]));
OR2X1 mul_U3708(.A(dpath_mulcore_ary1_a0_s_2[62]), .B(n9321), .Y(n16664));
AND2X1 mul_U3709(.A(n1620), .B(n3679), .Y(dpath_mulcore_ary1_a0_c_1[61]));
OR2X1 mul_U3710(.A(dpath_mulcore_ary1_a0_s_2[61]), .B(n9322), .Y(n16671));
AND2X1 mul_U3711(.A(n1621), .B(n3680), .Y(dpath_mulcore_ary1_a0_c_1[60]));
OR2X1 mul_U3712(.A(dpath_mulcore_ary1_a0_s_2[60]), .B(n9323), .Y(n16678));
AND2X1 mul_U3713(.A(n1622), .B(n3681), .Y(dpath_mulcore_ary1_a0_c_1[59]));
OR2X1 mul_U3714(.A(dpath_mulcore_ary1_a0_s_2[59]), .B(n9324), .Y(n16685));
AND2X1 mul_U3715(.A(n1623), .B(n3682), .Y(dpath_mulcore_ary1_a0_c_1[58]));
OR2X1 mul_U3716(.A(dpath_mulcore_ary1_a0_s_2[58]), .B(n9325), .Y(n16692));
AND2X1 mul_U3717(.A(n1624), .B(n3683), .Y(dpath_mulcore_ary1_a0_c_1[57]));
OR2X1 mul_U3718(.A(dpath_mulcore_ary1_a0_s_2[57]), .B(n9326), .Y(n16699));
AND2X1 mul_U3719(.A(n1625), .B(n3684), .Y(dpath_mulcore_ary1_a0_c_1[56]));
OR2X1 mul_U3720(.A(dpath_mulcore_ary1_a0_s_2[56]), .B(n9327), .Y(n16706));
AND2X1 mul_U3721(.A(n1626), .B(n3685), .Y(dpath_mulcore_ary1_a0_c_1[55]));
OR2X1 mul_U3722(.A(dpath_mulcore_ary1_a0_s_2[55]), .B(n9328), .Y(n16713));
AND2X1 mul_U3723(.A(n1627), .B(n3686), .Y(dpath_mulcore_ary1_a0_c_1[54]));
OR2X1 mul_U3724(.A(dpath_mulcore_ary1_a0_s_2[54]), .B(n9329), .Y(n16720));
AND2X1 mul_U3725(.A(n1628), .B(n3687), .Y(dpath_mulcore_ary1_a0_c_1[53]));
OR2X1 mul_U3726(.A(dpath_mulcore_ary1_a0_s_2[53]), .B(n9330), .Y(n16727));
AND2X1 mul_U3727(.A(n1629), .B(n3688), .Y(dpath_mulcore_ary1_a0_c_1[52]));
OR2X1 mul_U3728(.A(dpath_mulcore_ary1_a0_s_2[52]), .B(n9331), .Y(n16734));
AND2X1 mul_U3729(.A(n1630), .B(n3689), .Y(dpath_mulcore_ary1_a0_c_1[51]));
OR2X1 mul_U3730(.A(dpath_mulcore_ary1_a0_s_2[51]), .B(n9332), .Y(n16741));
INVX1 mul_U3731(.A(n9492), .Y(n9565));
AND2X1 mul_U3732(.A(n1631), .B(n3690), .Y(dpath_mulcore_ary1_a0_c_1[50]));
OR2X1 mul_U3733(.A(dpath_mulcore_ary1_a0_s_2[50]), .B(n9333), .Y(n16748));
AND2X1 mul_U3734(.A(n1632), .B(n3691), .Y(dpath_mulcore_ary1_a0_c_1[49]));
OR2X1 mul_U3735(.A(dpath_mulcore_ary1_a0_s_2[49]), .B(n9334), .Y(n16755));
AND2X1 mul_U3736(.A(n1633), .B(n3692), .Y(dpath_mulcore_ary1_a0_c_1[48]));
OR2X1 mul_U3737(.A(dpath_mulcore_ary1_a0_s_2[48]), .B(n9335), .Y(n16762));
AND2X1 mul_U3738(.A(n1634), .B(n3693), .Y(dpath_mulcore_ary1_a0_c_1[47]));
OR2X1 mul_U3739(.A(dpath_mulcore_ary1_a0_s_2[47]), .B(n9336), .Y(n16769));
AND2X1 mul_U3740(.A(n1635), .B(n3694), .Y(dpath_mulcore_ary1_a0_c_1[46]));
OR2X1 mul_U3741(.A(dpath_mulcore_ary1_a0_s_2[46]), .B(n9337), .Y(n16776));
INVX1 mul_U3742(.A(n9499), .Y(n9582));
AND2X1 mul_U3743(.A(n1636), .B(n3695), .Y(dpath_mulcore_ary1_a0_c_1[45]));
OR2X1 mul_U3744(.A(dpath_mulcore_ary1_a0_s_2[45]), .B(n9338), .Y(n16783));
AND2X1 mul_U3745(.A(n1637), .B(n3696), .Y(dpath_mulcore_ary1_a0_c_1[44]));
OR2X1 mul_U3746(.A(dpath_mulcore_ary1_a0_s_2[44]), .B(n9339), .Y(n16790));
AND2X1 mul_U3747(.A(n1638), .B(n3697), .Y(dpath_mulcore_ary1_a0_c_1[43]));
OR2X1 mul_U3748(.A(dpath_mulcore_ary1_a0_s_2[43]), .B(n9340), .Y(n16797));
AND2X1 mul_U3749(.A(n1639), .B(n3698), .Y(dpath_mulcore_ary1_a0_c_1[42]));
OR2X1 mul_U3750(.A(dpath_mulcore_ary1_a0_s_2[42]), .B(n9341), .Y(n16804));
AND2X1 mul_U3751(.A(n1640), .B(n3699), .Y(dpath_mulcore_ary1_a0_c_1[41]));
OR2X1 mul_U3752(.A(dpath_mulcore_ary1_a0_s_2[41]), .B(n9342), .Y(n16811));
AND2X1 mul_U3753(.A(n1641), .B(n3700), .Y(dpath_mulcore_ary1_a0_c_1[40]));
OR2X1 mul_U3754(.A(dpath_mulcore_ary1_a0_s_2[40]), .B(n9343), .Y(n16818));
AND2X1 mul_U3755(.A(n1642), .B(n3701), .Y(dpath_mulcore_ary1_a0_c_1[39]));
OR2X1 mul_U3756(.A(dpath_mulcore_ary1_a0_s_2[39]), .B(n9344), .Y(n16825));
AND2X1 mul_U3757(.A(n1643), .B(n3702), .Y(dpath_mulcore_ary1_a0_c_1[38]));
OR2X1 mul_U3758(.A(dpath_mulcore_ary1_a0_s_2[38]), .B(n9345), .Y(n16832));
AND2X1 mul_U3759(.A(n1644), .B(n3703), .Y(dpath_mulcore_ary1_a0_c_1[37]));
OR2X1 mul_U3760(.A(dpath_mulcore_ary1_a0_s_2[37]), .B(n9346), .Y(n16839));
AND2X1 mul_U3761(.A(n1645), .B(n3704), .Y(dpath_mulcore_ary1_a0_c_1[36]));
OR2X1 mul_U3762(.A(dpath_mulcore_ary1_a0_s_2[36]), .B(n9347), .Y(n16846));
AND2X1 mul_U3763(.A(n1646), .B(n3705), .Y(dpath_mulcore_ary1_a0_c_1[35]));
OR2X1 mul_U3764(.A(dpath_mulcore_ary1_a0_s_2[35]), .B(n9348), .Y(n16853));
AND2X1 mul_U3765(.A(n1647), .B(n3706), .Y(dpath_mulcore_ary1_a0_c_1[34]));
OR2X1 mul_U3766(.A(dpath_mulcore_ary1_a0_s_2[34]), .B(n9349), .Y(n16860));
AND2X1 mul_U3767(.A(n1648), .B(n3707), .Y(dpath_mulcore_ary1_a0_c_1[33]));
OR2X1 mul_U3768(.A(dpath_mulcore_ary1_a0_s_2[33]), .B(n9350), .Y(n16867));
AND2X1 mul_U3769(.A(n1649), .B(n3708), .Y(dpath_mulcore_ary1_a0_c_1[32]));
OR2X1 mul_U3770(.A(dpath_mulcore_ary1_a0_s_2[32]), .B(n9351), .Y(n16874));
AND2X1 mul_U3771(.A(n1650), .B(n3709), .Y(dpath_mulcore_ary1_a0_c_1[31]));
OR2X1 mul_U3772(.A(dpath_mulcore_ary1_a0_s_2[31]), .B(n9352), .Y(n16881));
AND2X1 mul_U3773(.A(n1651), .B(n3710), .Y(dpath_mulcore_ary1_a0_c_1[30]));
OR2X1 mul_U3774(.A(dpath_mulcore_ary1_a0_s_2[30]), .B(n9353), .Y(n16888));
AND2X1 mul_U3775(.A(n1652), .B(n3711), .Y(dpath_mulcore_ary1_a0_c_1[29]));
OR2X1 mul_U3776(.A(dpath_mulcore_ary1_a0_s_2[29]), .B(n9354), .Y(n16895));
AND2X1 mul_U3777(.A(n1653), .B(n3712), .Y(dpath_mulcore_ary1_a0_c_1[28]));
OR2X1 mul_U3778(.A(dpath_mulcore_ary1_a0_s_2[28]), .B(n9355), .Y(n16902));
AND2X1 mul_U3779(.A(n1654), .B(n3713), .Y(dpath_mulcore_ary1_a0_c_1[27]));
OR2X1 mul_U3780(.A(dpath_mulcore_ary1_a0_s_2[27]), .B(n9356), .Y(n16909));
AND2X1 mul_U3781(.A(n1655), .B(n3714), .Y(dpath_mulcore_ary1_a0_c_1[26]));
OR2X1 mul_U3782(.A(dpath_mulcore_ary1_a0_s_2[26]), .B(n9357), .Y(n16916));
AND2X1 mul_U3783(.A(n1656), .B(n3715), .Y(dpath_mulcore_ary1_a0_c_1[25]));
OR2X1 mul_U3784(.A(dpath_mulcore_ary1_a0_s_2[25]), .B(n9358), .Y(n16923));
AND2X1 mul_U3785(.A(n1657), .B(n3716), .Y(dpath_mulcore_ary1_a0_c_1[24]));
OR2X1 mul_U3786(.A(dpath_mulcore_ary1_a0_s_2[24]), .B(n9359), .Y(n16930));
AND2X1 mul_U3787(.A(n1658), .B(n3717), .Y(dpath_mulcore_ary1_a0_c_1[23]));
OR2X1 mul_U3788(.A(dpath_mulcore_ary1_a0_s_2[23]), .B(n9360), .Y(n16937));
AND2X1 mul_U3789(.A(n1659), .B(n3718), .Y(dpath_mulcore_ary1_a0_c_1[22]));
OR2X1 mul_U3790(.A(dpath_mulcore_ary1_a0_s_2[22]), .B(n9361), .Y(n16944));
AND2X1 mul_U3791(.A(n1660), .B(n3719), .Y(dpath_mulcore_ary1_a0_c_1[21]));
OR2X1 mul_U3792(.A(dpath_mulcore_ary1_a0_s_2[21]), .B(n9362), .Y(n16951));
AND2X1 mul_U3793(.A(n1661), .B(n3720), .Y(dpath_mulcore_ary1_a0_c_1[20]));
OR2X1 mul_U3794(.A(dpath_mulcore_ary1_a0_s_2[20]), .B(n9363), .Y(n16958));
AND2X1 mul_U3795(.A(n1662), .B(n3721), .Y(dpath_mulcore_ary1_a0_c_1[19]));
OR2X1 mul_U3796(.A(dpath_mulcore_ary1_a0_s_2[19]), .B(n9364), .Y(n16965));
AND2X1 mul_U3797(.A(n1663), .B(n3722), .Y(dpath_mulcore_ary1_a0_c_1[18]));
OR2X1 mul_U3798(.A(dpath_mulcore_ary1_a0_s_2[18]), .B(n9365), .Y(n16972));
AND2X1 mul_U3799(.A(n1664), .B(n3723), .Y(dpath_mulcore_ary1_a0_c_1[17]));
OR2X1 mul_U3800(.A(dpath_mulcore_ary1_a0_s_2[17]), .B(n9366), .Y(n16979));
AND2X1 mul_U3801(.A(n1665), .B(n3724), .Y(dpath_mulcore_ary1_a0_c_1[16]));
OR2X1 mul_U3802(.A(dpath_mulcore_ary1_a0_s_2[16]), .B(n9367), .Y(n16986));
AND2X1 mul_U3803(.A(n1666), .B(n3725), .Y(dpath_mulcore_ary1_a0_c_1[15]));
OR2X1 mul_U3804(.A(dpath_mulcore_ary1_a0_s_2[15]), .B(n9368), .Y(n16993));
AND2X1 mul_U3805(.A(n1667), .B(n3726), .Y(dpath_mulcore_ary1_a0_c_1[14]));
OR2X1 mul_U3806(.A(dpath_mulcore_ary1_a0_s_2[14]), .B(dpath_mulcore_ary1_a0_c_1[13]), .Y(n17000));
AND2X1 mul_U3807(.A(dpath_mulcore_ary1_a0_s0[13]), .B(n7200), .Y(dpath_mulcore_ary1_a0_c_1[13]));
OR2X1 mul_U3808(.A(dpath_mulcore_ary1_a0_s_2[13]), .B(dpath_mulcore_ary1_a0_c_1[12]), .Y(n17007));
AND2X1 mul_U3809(.A(dpath_mulcore_ary1_a0_s0[12]), .B(n7201), .Y(dpath_mulcore_ary1_a0_c_1[12]));
OR2X1 mul_U3810(.A(dpath_mulcore_ary1_a0_s_2[12]), .B(dpath_mulcore_ary1_a0_c_1[11]), .Y(n17014));
AND2X1 mul_U3811(.A(dpath_mulcore_ary1_a0_s0[11]), .B(n7202), .Y(dpath_mulcore_ary1_a0_c_1[11]));
OR2X1 mul_U3812(.A(dpath_mulcore_ary1_a0_s_2[11]), .B(dpath_mulcore_ary1_a0_c_1[10]), .Y(n17021));
AND2X1 mul_U3813(.A(n1124), .B(n3185), .Y(dpath_mulcore_ary1_a0_c1[3]));
AND2X1 mul_U3814(.A(n415), .B(n11553), .Y(dpath_mulcore_ary1_a0_I1_I0_p0_1));
OR2X1 mul_U3815(.A(n6486), .B(dpath_mulcore_b3[0]), .Y(n11553));
OR2X1 mul_U3816(.A(n13690), .B(n5931), .Y(dpath_mulcore_ary1_a0_I1_I0_b0n));
AND2X1 mul_U3817(.A(n7402), .B(n9845), .Y(n13690));
AND2X1 mul_U3818(.A(n1127), .B(n3188), .Y(dpath_mulcore_ary1_a0_c0[2]));
OR2X1 mul_U3819(.A(n9723), .B(n5932), .Y(dpath_mulcore_ary1_a0_I0_I0_b1n_0));
INVX1 mul_U3820(.A(n9499), .Y(n9581));
INVX1 mul_U3821(.A(n9495), .Y(n9572));
AND2X1 mul_U3822(.A(n101), .B(n10605), .Y(dpath_mulcore_ary1_a0_I2_I2_net43));
OR2X1 mul_U3823(.A(n6169), .B(dpath_mulcore_b7[0]), .Y(n10605));
AND2X1 mul_U3824(.A(n1608), .B(n3667), .Y(dpath_mulcore_ary1_a0_c_2[75]));
AND2X1 mul_U3825(.A(n1609), .B(n3668), .Y(dpath_mulcore_ary1_a0_c_2[74]));
AND2X1 mul_U3826(.A(n1610), .B(n3669), .Y(dpath_mulcore_ary1_a0_c_2[73]));
AND2X1 mul_U3827(.A(n1611), .B(n3670), .Y(dpath_mulcore_ary1_a0_c_2[72]));
AND2X1 mul_U3828(.A(n1607), .B(n3666), .Y(dpath_mulcore_ary1_a0_c_2[71]));
AND2X1 mul_U3829(.A(n2479), .B(n4405), .Y(dpath_mulcore_ary1_a0_c_2[70]));
AND2X1 mul_U3830(.A(n1539), .B(n3603), .Y(dpath_mulcore_ary1_a0_c_2[69]));
AND2X1 mul_U3831(.A(n1540), .B(n3604), .Y(dpath_mulcore_ary1_a0_c_2[68]));
AND2X1 mul_U3832(.A(n1541), .B(n3605), .Y(dpath_mulcore_ary1_a0_c_2[67]));
AND2X1 mul_U3833(.A(n1542), .B(n3606), .Y(dpath_mulcore_ary1_a0_c_2[66]));
AND2X1 mul_U3834(.A(n1543), .B(n3607), .Y(dpath_mulcore_ary1_a0_c_2[65]));
AND2X1 mul_U3835(.A(n1544), .B(n3608), .Y(dpath_mulcore_ary1_a0_c_2[64]));
AND2X1 mul_U3836(.A(n1545), .B(n3609), .Y(dpath_mulcore_ary1_a0_c_2[63]));
AND2X1 mul_U3837(.A(n1546), .B(n3610), .Y(dpath_mulcore_ary1_a0_c_2[62]));
AND2X1 mul_U3838(.A(n1547), .B(n3611), .Y(dpath_mulcore_ary1_a0_c_2[61]));
AND2X1 mul_U3839(.A(n1548), .B(n3612), .Y(dpath_mulcore_ary1_a0_c_2[60]));
AND2X1 mul_U3840(.A(n1549), .B(n3613), .Y(dpath_mulcore_ary1_a0_c_2[59]));
AND2X1 mul_U3841(.A(n1550), .B(n3614), .Y(dpath_mulcore_ary1_a0_c_2[58]));
AND2X1 mul_U3842(.A(n1551), .B(n3615), .Y(dpath_mulcore_ary1_a0_c_2[57]));
AND2X1 mul_U3843(.A(n1552), .B(n3616), .Y(dpath_mulcore_ary1_a0_c_2[56]));
AND2X1 mul_U3844(.A(n1553), .B(n3617), .Y(dpath_mulcore_ary1_a0_c_2[55]));
AND2X1 mul_U3845(.A(n1554), .B(n3618), .Y(dpath_mulcore_ary1_a0_c_2[54]));
AND2X1 mul_U3846(.A(n1555), .B(n3619), .Y(dpath_mulcore_ary1_a0_c_2[53]));
AND2X1 mul_U3847(.A(n1556), .B(n3620), .Y(dpath_mulcore_ary1_a0_c_2[52]));
AND2X1 mul_U3848(.A(n1557), .B(n3621), .Y(dpath_mulcore_ary1_a0_c_2[51]));
AND2X1 mul_U3849(.A(n1558), .B(n3622), .Y(dpath_mulcore_ary1_a0_c_2[50]));
AND2X1 mul_U3850(.A(n1559), .B(n3623), .Y(dpath_mulcore_ary1_a0_c_2[49]));
AND2X1 mul_U3851(.A(n1560), .B(n3624), .Y(dpath_mulcore_ary1_a0_c_2[48]));
AND2X1 mul_U3852(.A(n1561), .B(n3625), .Y(dpath_mulcore_ary1_a0_c_2[47]));
AND2X1 mul_U3853(.A(n1562), .B(n3626), .Y(dpath_mulcore_ary1_a0_c_2[46]));
AND2X1 mul_U3854(.A(n1563), .B(n3627), .Y(dpath_mulcore_ary1_a0_c_2[45]));
AND2X1 mul_U3855(.A(n1564), .B(n3628), .Y(dpath_mulcore_ary1_a0_c_2[44]));
AND2X1 mul_U3856(.A(n1565), .B(n3629), .Y(dpath_mulcore_ary1_a0_c_2[43]));
AND2X1 mul_U3857(.A(n1566), .B(n3630), .Y(dpath_mulcore_ary1_a0_c_2[42]));
AND2X1 mul_U3858(.A(n1567), .B(n3631), .Y(dpath_mulcore_ary1_a0_c_2[41]));
AND2X1 mul_U3859(.A(n1568), .B(n3632), .Y(dpath_mulcore_ary1_a0_c_2[40]));
AND2X1 mul_U3860(.A(n1569), .B(n3633), .Y(dpath_mulcore_ary1_a0_c_2[39]));
AND2X1 mul_U3861(.A(n1570), .B(n3634), .Y(dpath_mulcore_ary1_a0_c_2[38]));
AND2X1 mul_U3862(.A(n1571), .B(n3635), .Y(dpath_mulcore_ary1_a0_c_2[37]));
AND2X1 mul_U3863(.A(n1572), .B(n3636), .Y(dpath_mulcore_ary1_a0_c_2[36]));
AND2X1 mul_U3864(.A(n1573), .B(n3637), .Y(dpath_mulcore_ary1_a0_c_2[35]));
AND2X1 mul_U3865(.A(n1574), .B(n3638), .Y(dpath_mulcore_ary1_a0_c_2[34]));
AND2X1 mul_U3866(.A(n1575), .B(n3639), .Y(dpath_mulcore_ary1_a0_c_2[33]));
AND2X1 mul_U3867(.A(n1576), .B(n3640), .Y(dpath_mulcore_ary1_a0_c_2[32]));
AND2X1 mul_U3868(.A(n1577), .B(n3641), .Y(dpath_mulcore_ary1_a0_c_2[31]));
AND2X1 mul_U3869(.A(n1578), .B(n3642), .Y(dpath_mulcore_ary1_a0_c_2[30]));
AND2X1 mul_U3870(.A(n1579), .B(n3643), .Y(dpath_mulcore_ary1_a0_c_2[29]));
AND2X1 mul_U3871(.A(n1580), .B(n3644), .Y(dpath_mulcore_ary1_a0_c_2[28]));
AND2X1 mul_U3872(.A(n1581), .B(n3645), .Y(dpath_mulcore_ary1_a0_c_2[27]));
AND2X1 mul_U3873(.A(n1582), .B(n3646), .Y(dpath_mulcore_ary1_a0_c_2[26]));
AND2X1 mul_U3874(.A(n1583), .B(n3647), .Y(dpath_mulcore_ary1_a0_c_2[25]));
AND2X1 mul_U3875(.A(n1584), .B(n3648), .Y(dpath_mulcore_ary1_a0_c_2[24]));
AND2X1 mul_U3876(.A(n1585), .B(n3649), .Y(dpath_mulcore_ary1_a0_c_2[23]));
AND2X1 mul_U3877(.A(n1586), .B(n3650), .Y(dpath_mulcore_ary1_a0_c_2[22]));
AND2X1 mul_U3878(.A(n1587), .B(n3651), .Y(dpath_mulcore_ary1_a0_c_2[21]));
AND2X1 mul_U3879(.A(n1588), .B(n3652), .Y(dpath_mulcore_ary1_a0_c_2[20]));
AND2X1 mul_U3880(.A(n1589), .B(n3653), .Y(dpath_mulcore_ary1_a0_c_2[19]));
AND2X1 mul_U3881(.A(n1590), .B(n3654), .Y(dpath_mulcore_ary1_a0_c_2[18]));
AND2X1 mul_U3882(.A(n1591), .B(n3655), .Y(dpath_mulcore_ary1_a0_c_2[17]));
AND2X1 mul_U3883(.A(n1592), .B(n3656), .Y(dpath_mulcore_ary1_a0_c_2[16]));
AND2X1 mul_U3884(.A(n1593), .B(n3657), .Y(dpath_mulcore_ary1_a0_c_2[15]));
AND2X1 mul_U3885(.A(n1594), .B(n3658), .Y(dpath_mulcore_ary1_a0_c_2[14]));
INVX1 mul_U3886(.A(n9493), .Y(n9567));
AND2X1 mul_U3887(.A(n1595), .B(n3659), .Y(dpath_mulcore_ary1_a0_c_2[13]));
AND2X1 mul_U3888(.A(n1596), .B(n3660), .Y(dpath_mulcore_ary1_a0_c_2[12]));
AND2X1 mul_U3889(.A(n1597), .B(n3661), .Y(dpath_mulcore_ary1_a0_c_2[11]));
AND2X1 mul_U3890(.A(dpath_mulcore_ary1_a0_s0[10]), .B(n7203), .Y(dpath_mulcore_ary1_a0_c_1[10]));
INVX1 mul_U3891(.A(n9492), .Y(n9566));
AND2X1 mul_U3892(.A(n1601), .B(n3663), .Y(dpath_mulcore_ary1_a0_c_1[9]));
AND2X1 mul_U3893(.A(n1602), .B(n3664), .Y(dpath_mulcore_ary1_a0_c_1[8]));
AND2X1 mul_U3894(.A(n1668), .B(n3727), .Y(dpath_mulcore_ary1_a0_c_1[7]));
OR2X1 mul_U3895(.A(n9725), .B(n5948), .Y(dpath_mulcore_ary1_a0_b2n[1]));
INVX1 mul_U3896(.A(n9494), .Y(n9570));
OR2X1 mul_U3897(.A(n9725), .B(n5949), .Y(dpath_mulcore_ary1_a0_b2n[0]));
AND2X1 mul_U3898(.A(control_n22), .B(spu_mul_req_vld), .Y(control_n18));
AND2X1 mul_U3899(.A(n3086), .B(n9816), .Y(control_n22));
INVX1 mul_U3900(.A(n9494), .Y(n9571));
INVX1 mul_U3901(.A(control_c1_act), .Y(n9816));
INVX1 mul_U3902(.A(control_favor_e), .Y(n9817));
AND2X1 mul_U3903(.A(n2490), .B(n4419), .Y(dpath_mulcore_booth_encode0_a_n43));
AND2X1 mul_U3904(.A(n5497), .B(n4426), .Y(dpath_mulcore_booth_b1_in0[0]));
AND2X1 mul_U3905(.A(n5440), .B(n4380), .Y(dpath_mulcore_booth_b1_in1[0]));
AND2X1 mul_U3906(.A(dpath_mulcore_booth_encode0_a_n39), .B(n4417), .Y(dpath_mulcore_booth_b2_in0[1]));
AND2X1 mul_U3907(.A(n2489), .B(n4418), .Y(dpath_mulcore_booth_encode0_a_n39));
AND2X1 mul_U3908(.A(n18035), .B(n4371), .Y(dpath_mulcore_booth_b2_in1[1]));
AND2X1 mul_U3909(.A(n5494), .B(n4425), .Y(dpath_mulcore_booth_b2_in0[0]));
AND2X1 mul_U3910(.A(n5437), .B(n4379), .Y(dpath_mulcore_booth_b2_in1[0]));
AND2X1 mul_U3911(.A(dpath_mulcore_booth_encode0_a_n35), .B(n4415), .Y(dpath_mulcore_booth_b3_in0[1]));
AND2X1 mul_U3912(.A(n2488), .B(n4416), .Y(dpath_mulcore_booth_encode0_a_n35));
AND2X1 mul_U3913(.A(n18031), .B(n4369), .Y(dpath_mulcore_booth_b3_in1[1]));
AND2X1 mul_U3914(.A(n5492), .B(n4424), .Y(dpath_mulcore_booth_b3_in0[0]));
AND2X1 mul_U3915(.A(n5435), .B(n4378), .Y(dpath_mulcore_booth_b3_in1[0]));
AND2X1 mul_U3916(.A(dpath_mulcore_booth_encode0_a_n31), .B(n4413), .Y(dpath_mulcore_booth_b4_in0[1]));
AND2X1 mul_U3917(.A(n2487), .B(n4414), .Y(dpath_mulcore_booth_encode0_a_n31));
AND2X1 mul_U3918(.A(n18027), .B(n4367), .Y(dpath_mulcore_booth_b4_in1[1]));
AND2X1 mul_U3919(.A(n5490), .B(n4423), .Y(dpath_mulcore_booth_b4_in0[0]));
AND2X1 mul_U3920(.A(n5433), .B(n4377), .Y(dpath_mulcore_booth_b4_in1[0]));
AND2X1 mul_U3921(.A(dpath_mulcore_booth_encode0_a_n27), .B(n4411), .Y(dpath_mulcore_booth_b5_in0[1]));
AND2X1 mul_U3922(.A(n2486), .B(n4412), .Y(dpath_mulcore_booth_encode0_a_n27));
AND2X1 mul_U3923(.A(n18023), .B(n4365), .Y(dpath_mulcore_booth_b5_in1[1]));
AND2X1 mul_U3924(.A(n5488), .B(n4422), .Y(dpath_mulcore_booth_b5_in0[0]));
AND2X1 mul_U3925(.A(n5431), .B(n4376), .Y(dpath_mulcore_booth_b5_in1[0]));
AND2X1 mul_U3926(.A(dpath_mulcore_booth_encode0_a_n23), .B(n4409), .Y(dpath_mulcore_booth_b6_in0[1]));
AND2X1 mul_U3927(.A(n2485), .B(n4410), .Y(dpath_mulcore_booth_encode0_a_n23));
AND2X1 mul_U3928(.A(n18019), .B(n4363), .Y(dpath_mulcore_booth_b6_in1[1]));
AND2X1 mul_U3929(.A(n5486), .B(n4421), .Y(dpath_mulcore_booth_b6_in0[0]));
AND2X1 mul_U3930(.A(n5429), .B(n4375), .Y(dpath_mulcore_booth_b6_in1[0]));
AND2X1 mul_U3931(.A(dpath_mulcore_booth_encode0_a_n19), .B(n4407), .Y(dpath_mulcore_booth_b7_in0[1]));
AND2X1 mul_U3932(.A(dpath_mulcore_booth_encode0_a_n21), .B(n4408), .Y(dpath_mulcore_booth_encode0_a_n19));
AND2X1 mul_U3933(.A(n18015), .B(n4361), .Y(dpath_mulcore_booth_b7_in1[1]));
AND2X1 mul_U3934(.A(n5483), .B(n4420), .Y(dpath_mulcore_booth_b7_in0[0]));
AND2X1 mul_U3935(.A(n5426), .B(n4374), .Y(dpath_mulcore_booth_b7_in1[0]));
AND2X1 mul_U3936(.A(n17947), .B(n4337), .Y(dpath_mulcore_booth_b8_in0[1]));
AND2X1 mul_U3937(.A(n17949), .B(n4338), .Y(n17947));
AND2X1 mul_U3938(.A(n18075), .B(n4381), .Y(dpath_mulcore_booth_b8_in1[1]));
AND2X1 mul_U3939(.A(n5416), .B(n4359), .Y(dpath_mulcore_booth_b8_in0[0]));
AND2X1 mul_U3940(.A(n5468), .B(n4403), .Y(dpath_mulcore_booth_b8_in1[0]));
AND2X1 mul_U3941(.A(n2462), .B(n4351), .Y(n17975));
AND2X1 mul_U3942(.A(n5414), .B(n4358), .Y(dpath_mulcore_booth_b9_in0[0]));
AND2X1 mul_U3943(.A(n5466), .B(n4402), .Y(dpath_mulcore_booth_b9_in1[0]));
AND2X1 mul_U3944(.A(n17971), .B(n4349), .Y(dpath_mulcore_booth_b10_in0[1]));
AND2X1 mul_U3945(.A(n2461), .B(n4350), .Y(n17971));
AND2X1 mul_U3946(.A(n18099), .B(n4393), .Y(dpath_mulcore_booth_b10_in1[1]));
AND2X1 mul_U3947(.A(n5411), .B(n4357), .Y(dpath_mulcore_booth_b10_in0[0]));
AND2X1 mul_U3948(.A(n5463), .B(n4401), .Y(dpath_mulcore_booth_b10_in1[0]));
AND2X1 mul_U3949(.A(n17967), .B(n4347), .Y(dpath_mulcore_booth_b11_in0[1]));
AND2X1 mul_U3950(.A(n2460), .B(n4348), .Y(n17967));
AND2X1 mul_U3951(.A(n18095), .B(n4391), .Y(dpath_mulcore_booth_b11_in1[1]));
AND2X1 mul_U3952(.A(n5409), .B(n4356), .Y(dpath_mulcore_booth_b11_in0[0]));
AND2X1 mul_U3953(.A(n5461), .B(n4400), .Y(dpath_mulcore_booth_b11_in1[0]));
AND2X1 mul_U3954(.A(n17963), .B(n4345), .Y(dpath_mulcore_booth_b12_in0[1]));
AND2X1 mul_U3955(.A(n2459), .B(n4346), .Y(n17963));
AND2X1 mul_U3956(.A(n18091), .B(n4389), .Y(dpath_mulcore_booth_b12_in1[1]));
AND2X1 mul_U3957(.A(n5407), .B(n4355), .Y(dpath_mulcore_booth_b12_in0[0]));
AND2X1 mul_U3958(.A(n5459), .B(n4399), .Y(dpath_mulcore_booth_b12_in1[0]));
AND2X1 mul_U3959(.A(n17959), .B(n4343), .Y(dpath_mulcore_booth_b13_in0[1]));
AND2X1 mul_U3960(.A(n2458), .B(n4344), .Y(n17959));
AND2X1 mul_U3961(.A(n18087), .B(n4387), .Y(dpath_mulcore_booth_b13_in1[1]));
AND2X1 mul_U3962(.A(n5405), .B(n4354), .Y(dpath_mulcore_booth_b13_in0[0]));
AND2X1 mul_U3963(.A(n5457), .B(n4398), .Y(dpath_mulcore_booth_b13_in1[0]));
AND2X1 mul_U3964(.A(n17955), .B(n4341), .Y(dpath_mulcore_booth_b14_in0[1]));
AND2X1 mul_U3965(.A(n2457), .B(n4342), .Y(n17955));
AND2X1 mul_U3966(.A(n18083), .B(n4385), .Y(dpath_mulcore_booth_b14_in1[1]));
AND2X1 mul_U3967(.A(n5403), .B(n4353), .Y(dpath_mulcore_booth_b14_in0[0]));
AND2X1 mul_U3968(.A(n5455), .B(n4397), .Y(dpath_mulcore_booth_b14_in1[0]));
AND2X1 mul_U3969(.A(n17951), .B(n4339), .Y(dpath_mulcore_booth_b15_in0[1]));
AND2X1 mul_U3970(.A(n17953), .B(n4340), .Y(n17951));
AND2X1 mul_U3971(.A(n18079), .B(n4383), .Y(dpath_mulcore_booth_b15_in1[1]));
AND2X1 mul_U3972(.A(n5400), .B(n4352), .Y(dpath_mulcore_booth_b15_in0[0]));
AND2X1 mul_U3973(.A(n5452), .B(n4396), .Y(dpath_mulcore_booth_b15_in1[0]));
AND2X1 mul_U3974(.A(n1733), .B(n2), .Y(dpath_mulcore_ary1_a1_c_2[76]));
AND2X1 mul_U3975(.A(n2191), .B(n4181), .Y(dpath_mulcore_ary1_a1_co[71]));
AND2X1 mul_U3976(.A(n2198), .B(n4182), .Y(dpath_mulcore_ary1_a1_co[70]));
AND2X1 mul_U3977(.A(n2200), .B(n4183), .Y(dpath_mulcore_ary1_a1_co[69]));
AND2X1 mul_U3978(.A(n2202), .B(n4184), .Y(dpath_mulcore_ary1_a1_co[68]));
AND2X1 mul_U3979(.A(n2204), .B(n4185), .Y(dpath_mulcore_ary1_a1_co[67]));
AND2X1 mul_U3980(.A(n2206), .B(n4186), .Y(dpath_mulcore_ary1_a1_co[66]));
AND2X1 mul_U3981(.A(n2208), .B(n4187), .Y(dpath_mulcore_ary1_a1_co[65]));
AND2X1 mul_U3982(.A(n2210), .B(n4188), .Y(dpath_mulcore_ary1_a1_co[64]));
AND2X1 mul_U3983(.A(n2212), .B(n4189), .Y(dpath_mulcore_ary1_a1_co[63]));
AND2X1 mul_U3984(.A(n2214), .B(n4190), .Y(dpath_mulcore_ary1_a1_co[62]));
AND2X1 mul_U3985(.A(n2216), .B(n4191), .Y(dpath_mulcore_ary1_a1_co[61]));
AND2X1 mul_U3986(.A(n2218), .B(n4192), .Y(dpath_mulcore_ary1_a1_co[60]));
AND2X1 mul_U3987(.A(n2220), .B(n4193), .Y(dpath_mulcore_ary1_a1_co[59]));
AND2X1 mul_U3988(.A(n2222), .B(n4194), .Y(dpath_mulcore_ary1_a1_co[58]));
AND2X1 mul_U3989(.A(n2224), .B(n4195), .Y(dpath_mulcore_ary1_a1_co[57]));
AND2X1 mul_U3990(.A(n2226), .B(n4196), .Y(dpath_mulcore_ary1_a1_co[56]));
AND2X1 mul_U3991(.A(n2228), .B(n4197), .Y(dpath_mulcore_ary1_a1_co[55]));
AND2X1 mul_U3992(.A(n2230), .B(n4198), .Y(dpath_mulcore_ary1_a1_co[54]));
AND2X1 mul_U3993(.A(n2232), .B(n4199), .Y(dpath_mulcore_ary1_a1_co[53]));
AND2X1 mul_U3994(.A(n2234), .B(n4200), .Y(dpath_mulcore_ary1_a1_co[52]));
AND2X1 mul_U3995(.A(n2236), .B(n4201), .Y(dpath_mulcore_ary1_a1_co[51]));
AND2X1 mul_U3996(.A(n2238), .B(n4202), .Y(dpath_mulcore_ary1_a1_co[50]));
AND2X1 mul_U3997(.A(n2240), .B(n4203), .Y(dpath_mulcore_ary1_a1_co[49]));
AND2X1 mul_U3998(.A(n2242), .B(n4204), .Y(dpath_mulcore_ary1_a1_co[48]));
AND2X1 mul_U3999(.A(n2244), .B(n4205), .Y(dpath_mulcore_ary1_a1_co[47]));
AND2X1 mul_U4000(.A(n2246), .B(n4206), .Y(dpath_mulcore_ary1_a1_co[46]));
AND2X1 mul_U4001(.A(n2248), .B(n4207), .Y(dpath_mulcore_ary1_a1_co[45]));
AND2X1 mul_U4002(.A(n2250), .B(n4208), .Y(dpath_mulcore_ary1_a1_co[44]));
AND2X1 mul_U4003(.A(n2252), .B(n4209), .Y(dpath_mulcore_ary1_a1_co[43]));
AND2X1 mul_U4004(.A(n2254), .B(n4210), .Y(dpath_mulcore_ary1_a1_co[42]));
AND2X1 mul_U4005(.A(n2256), .B(n4211), .Y(dpath_mulcore_ary1_a1_co[41]));
AND2X1 mul_U4006(.A(n2258), .B(n4212), .Y(dpath_mulcore_ary1_a1_co[40]));
AND2X1 mul_U4007(.A(n2260), .B(n4213), .Y(dpath_mulcore_ary1_a1_co[39]));
AND2X1 mul_U4008(.A(n2262), .B(n4214), .Y(dpath_mulcore_ary1_a1_co[38]));
AND2X1 mul_U4009(.A(n2264), .B(n4215), .Y(dpath_mulcore_ary1_a1_co[37]));
AND2X1 mul_U4010(.A(n2266), .B(n4216), .Y(dpath_mulcore_ary1_a1_co[36]));
AND2X1 mul_U4011(.A(n2268), .B(n4217), .Y(dpath_mulcore_ary1_a1_co[35]));
AND2X1 mul_U4012(.A(n2270), .B(n4218), .Y(dpath_mulcore_ary1_a1_co[34]));
AND2X1 mul_U4013(.A(n2272), .B(n4219), .Y(dpath_mulcore_ary1_a1_co[33]));
AND2X1 mul_U4014(.A(n2274), .B(n4220), .Y(dpath_mulcore_ary1_a1_co[32]));
AND2X1 mul_U4015(.A(n2276), .B(n4221), .Y(dpath_mulcore_ary1_a1_co[31]));
AND2X1 mul_U4016(.A(n2278), .B(n4222), .Y(dpath_mulcore_ary1_a1_co[30]));
AND2X1 mul_U4017(.A(n2280), .B(n4223), .Y(dpath_mulcore_ary1_a1_co[29]));
AND2X1 mul_U4018(.A(n2282), .B(n4224), .Y(dpath_mulcore_ary1_a1_co[28]));
AND2X1 mul_U4019(.A(n2284), .B(n4225), .Y(dpath_mulcore_ary1_a1_co[27]));
AND2X1 mul_U4020(.A(n2286), .B(n4226), .Y(dpath_mulcore_ary1_a1_co[26]));
AND2X1 mul_U4021(.A(n2288), .B(n4227), .Y(dpath_mulcore_ary1_a1_co[25]));
AND2X1 mul_U4022(.A(n2290), .B(n4228), .Y(dpath_mulcore_ary1_a1_co[24]));
AND2X1 mul_U4023(.A(n2292), .B(n4229), .Y(dpath_mulcore_ary1_a1_co[23]));
AND2X1 mul_U4024(.A(n2294), .B(n4230), .Y(dpath_mulcore_ary1_a1_co[22]));
AND2X1 mul_U4025(.A(n2296), .B(n4231), .Y(dpath_mulcore_ary1_a1_co[21]));
AND2X1 mul_U4026(.A(n2298), .B(n4232), .Y(dpath_mulcore_ary1_a1_co[20]));
AND2X1 mul_U4027(.A(n2300), .B(n4233), .Y(dpath_mulcore_ary1_a1_co[19]));
AND2X1 mul_U4028(.A(n2302), .B(n4234), .Y(dpath_mulcore_ary1_a1_co[18]));
AND2X1 mul_U4029(.A(n2304), .B(n4235), .Y(dpath_mulcore_ary1_a1_co[17]));
AND2X1 mul_U4030(.A(n2306), .B(n4236), .Y(dpath_mulcore_ary1_a1_co[16]));
AND2X1 mul_U4031(.A(n2308), .B(n4237), .Y(dpath_mulcore_ary1_a1_co[15]));
AND2X1 mul_U4032(.A(n2310), .B(n4238), .Y(dpath_mulcore_ary1_a1_co[14]));
AND2X1 mul_U4033(.A(n2312), .B(n4239), .Y(dpath_mulcore_ary1_a1_co[13]));
AND2X1 mul_U4034(.A(n2314), .B(n4240), .Y(dpath_mulcore_ary1_a1_co[12]));
AND2X1 mul_U4035(.A(n2316), .B(n4241), .Y(dpath_mulcore_ary1_a1_co[11]));
AND2X1 mul_U4036(.A(n1131), .B(n3192), .Y(dpath_mulcore_ary1_a1_c1[2]));
AND2X1 mul_U4037(.A(n7400), .B(dpath_mulcore_ary1_a1_I1_I0_b0n), .Y(dpath_mulcore_ary1_a1_c1[1]));
AND2X1 mul_U4038(.A(dpath_mulcore_ary1_a1_s0[2]), .B(dpath_mulcore_ary1_a1_c0[1]), .Y(dpath_mulcore_ary1_a1_c_1[2]));
AND2X1 mul_U4039(.A(n7401), .B(dpath_mulcore_ary1_a1_I0_I0_b0n), .Y(dpath_mulcore_ary1_a1_c0[1]));
AND2X1 mul_U4040(.A(n1108), .B(n13654), .Y(dpath_mulcore_ary1_a1_I0_I0_p0_1));
OR2X1 mul_U4041(.A(n7190), .B(dpath_mulcore_b8[0]), .Y(n13654));
OR2X1 mul_U4042(.A(n13734), .B(n5947), .Y(dpath_mulcore_ary1_a1_I0_I0_b0n));
AND2X1 mul_U4043(.A(n7406), .B(n9828), .Y(n13734));
INVX1 mul_U4044(.A(n13656), .Y(n9828));
OR2X1 mul_U4045(.A(n7191), .B(dpath_mulcore_b8[0]), .Y(n13656));
OR2X1 mul_U4046(.A(n9737), .B(n5946), .Y(dpath_mulcore_ary1_a1_I0_I0_b0n_0));
AND2X1 mul_U4047(.A(dpath_mulcore_ary1_a1_I2_I2_net38), .B(n3501), .Y(dpath_mulcore_ary1_a1_c2[66]));
AND2X1 mul_U4048(.A(n1439), .B(n3500), .Y(dpath_mulcore_ary1_a1_c2[65]));
INVX1 mul_U4049(.A(n9579), .Y(n9519));
INVX1 mul_U4050(.A(dpath_mulcore_ary1_a1_sc3_76__z), .Y(n10022));
INVX1 mul_U4051(.A(dpath_mulcore_ary1_a1_sc3_75__z), .Y(n10019));
INVX1 mul_U4052(.A(dpath_mulcore_ary1_a1_sc3_74__z), .Y(n10016));
INVX1 mul_U4053(.A(dpath_mulcore_ary1_a1_sc3_73__z), .Y(n10013));
INVX1 mul_U4054(.A(dpath_mulcore_ary1_a1_sc3_72__z), .Y(n10010));
INVX1 mul_U4055(.A(dpath_mulcore_ary1_a1_sc3_71__z), .Y(n10007));
INVX1 mul_U4056(.A(dpath_mulcore_ary1_a1_sc3_70__z), .Y(n10005));
INVX1 mul_U4057(.A(dpath_mulcore_ary1_a1_sc3_69__z), .Y(n10003));
INVX1 mul_U4058(.A(dpath_mulcore_ary1_a1_sc3_68__z), .Y(n10001));
INVX1 mul_U4059(.A(dpath_mulcore_ary1_a1_sc3_67__z), .Y(n9999));
INVX1 mul_U4060(.A(dpath_mulcore_ary1_a1_sc3_66__z), .Y(n9997));
INVX1 mul_U4061(.A(dpath_mulcore_ary1_a1_sc3_65__z), .Y(n9994));
INVX1 mul_U4062(.A(dpath_mulcore_ary1_a1_sc3_64__z), .Y(n9991));
INVX1 mul_U4063(.A(dpath_mulcore_ary1_a1_sc3_63__z), .Y(n9988));
INVX1 mul_U4064(.A(dpath_mulcore_ary1_a1_sc3_62__z), .Y(n9985));
INVX1 mul_U4065(.A(dpath_mulcore_ary1_a1_sc3_61__z), .Y(n9982));
INVX1 mul_U4066(.A(dpath_mulcore_ary1_a1_sc3_60__z), .Y(n9979));
INVX1 mul_U4067(.A(dpath_mulcore_ary1_a1_sc3_59__z), .Y(n9976));
INVX1 mul_U4068(.A(dpath_mulcore_ary1_a1_sc3_58__z), .Y(n9973));
INVX1 mul_U4069(.A(dpath_mulcore_ary1_a1_sc3_57__z), .Y(n9970));
INVX1 mul_U4070(.A(dpath_mulcore_ary1_a1_sc3_56__z), .Y(n9967));
INVX1 mul_U4071(.A(dpath_mulcore_ary1_a1_sc3_55__z), .Y(n9964));
INVX1 mul_U4072(.A(dpath_mulcore_ary1_a1_sc3_54__z), .Y(n9961));
INVX1 mul_U4073(.A(dpath_mulcore_ary1_a1_sc3_53__z), .Y(n9958));
INVX1 mul_U4074(.A(dpath_mulcore_ary1_a1_sc3_52__z), .Y(n9955));
INVX1 mul_U4075(.A(dpath_mulcore_ary1_a1_sc3_51__z), .Y(n9952));
INVX1 mul_U4076(.A(dpath_mulcore_ary1_a1_sc3_50__z), .Y(n9949));
INVX1 mul_U4077(.A(dpath_mulcore_ary1_a1_sc3_49__z), .Y(n9946));
INVX1 mul_U4078(.A(dpath_mulcore_ary1_a1_sc3_48__z), .Y(n9943));
INVX1 mul_U4079(.A(dpath_mulcore_ary1_a1_sc3_47__z), .Y(n9940));
INVX1 mul_U4080(.A(dpath_mulcore_ary1_a1_sc3_46__z), .Y(n9937));
INVX1 mul_U4081(.A(dpath_mulcore_ary1_a1_sc3_45__z), .Y(n9934));
INVX1 mul_U4082(.A(dpath_mulcore_ary1_a1_sc3_44__z), .Y(n9931));
INVX1 mul_U4083(.A(dpath_mulcore_ary1_a1_sc3_43__z), .Y(n9928));
INVX1 mul_U4084(.A(dpath_mulcore_ary1_a1_sc3_42__z), .Y(n9925));
INVX1 mul_U4085(.A(dpath_mulcore_ary1_a1_sc3_41__z), .Y(n9922));
INVX1 mul_U4086(.A(dpath_mulcore_ary1_a1_sc3_40__z), .Y(n9919));
INVX1 mul_U4087(.A(dpath_mulcore_ary1_a1_sc3_39__z), .Y(n9916));
INVX1 mul_U4088(.A(dpath_mulcore_ary1_a1_sc3_38__z), .Y(n9913));
INVX1 mul_U4089(.A(dpath_mulcore_ary1_a1_sc3_37__z), .Y(n9910));
INVX1 mul_U4090(.A(dpath_mulcore_ary1_a1_sc3_36__z), .Y(n9907));
INVX1 mul_U4091(.A(dpath_mulcore_ary1_a1_sc3_35__z), .Y(n9904));
INVX1 mul_U4092(.A(dpath_mulcore_ary1_a1_sc3_34__z), .Y(n9901));
INVX1 mul_U4093(.A(dpath_mulcore_ary1_a1_sc3_33__z), .Y(n9898));
INVX1 mul_U4094(.A(dpath_mulcore_ary1_a1_sc3_32__z), .Y(n9895));
INVX1 mul_U4095(.A(dpath_mulcore_ary1_a1_sc3_31__z), .Y(n9892));
INVX1 mul_U4096(.A(dpath_mulcore_ary1_a1_sc3_30__z), .Y(n9889));
INVX1 mul_U4097(.A(dpath_mulcore_ary1_a1_sc3_29__z), .Y(n9886));
INVX1 mul_U4098(.A(dpath_mulcore_ary1_a1_sc3_28__z), .Y(n9883));
INVX1 mul_U4099(.A(dpath_mulcore_ary1_a1_sc3_27__z), .Y(n9880));
INVX1 mul_U4100(.A(dpath_mulcore_ary1_a1_sc3_26__z), .Y(n9877));
INVX1 mul_U4101(.A(dpath_mulcore_ary1_a1_sc3_25__z), .Y(n9874));
INVX1 mul_U4102(.A(dpath_mulcore_ary1_a1_sc3_24__z), .Y(n9871));
INVX1 mul_U4103(.A(dpath_mulcore_ary1_a1_sc3_23__z), .Y(n9868));
INVX1 mul_U4104(.A(dpath_mulcore_ary1_a1_sc3_22__z), .Y(n9865));
INVX1 mul_U4105(.A(dpath_mulcore_ary1_a1_sc3_21__z), .Y(n9862));
INVX1 mul_U4106(.A(dpath_mulcore_ary1_a1_sc3_20__z), .Y(n9859));
INVX1 mul_U4107(.A(dpath_mulcore_ary1_a1_sc3_19__z), .Y(n9856));
INVX1 mul_U4108(.A(dpath_mulcore_ary1_a1_sc3_18__z), .Y(n9826));
INVX1 mul_U4109(.A(dpath_mulcore_ary1_a1_sc3_17__z), .Y(n9824));
INVX1 mul_U4110(.A(dpath_mulcore_ary1_a1_sc3_16__z), .Y(n9825));
INVX1 mul_U4111(.A(dpath_mulcore_ary1_a1_sc3_15__z), .Y(n9836));
INVX1 mul_U4112(.A(dpath_mulcore_ary1_a1_sc3_14__z), .Y(n9837));
INVX1 mul_U4113(.A(dpath_mulcore_ary1_a1_sc3_13__z), .Y(n9833));
INVX1 mul_U4114(.A(dpath_mulcore_ary1_a1_sc3_12__z), .Y(n9834));
AND2X1 mul_U4115(.A(n1732), .B(n3791), .Y(dpath_mulcore_ary1_a1_c_2[10]));
INVX1 mul_U4116(.A(n9575), .Y(n9531));
AND2X1 mul_U4117(.A(n1803), .B(n3857), .Y(dpath_mulcore_ary1_a1_c_1[6]));
AND2X1 mul_U4118(.A(n1804), .B(n3858), .Y(dpath_mulcore_ary1_a1_c_1[5]));
AND2X1 mul_U4119(.A(n1805), .B(n3859), .Y(dpath_mulcore_ary1_a1_c_1[4]));
AND2X1 mul_U4120(.A(n1737), .B(n3794), .Y(dpath_mulcore_ary1_a1_c_1[3]));
INVX1 mul_U4121(.A(n9575), .Y(n9529));
AND2X1 mul_U4122(.A(n2759), .B(n4435), .Y(dpath_n165));
AND2X1 mul_U4123(.A(n2760), .B(n4436), .Y(dpath_n164));
AND2X1 mul_U4124(.A(n2761), .B(n4437), .Y(dpath_n171));
AND2X1 mul_U4125(.A(n2762), .B(n4438), .Y(dpath_n170));
AND2X1 mul_U4126(.A(n2763), .B(n4439), .Y(dpath_n177));
AND2X1 mul_U4127(.A(n2764), .B(n4440), .Y(dpath_n176));
AND2X1 mul_U4128(.A(n2765), .B(n4441), .Y(dpath_n183));
AND2X1 mul_U4129(.A(n2766), .B(n4442), .Y(dpath_n182));
AND2X1 mul_U4130(.A(n2769), .B(n4445), .Y(dpath_n195));
AND2X1 mul_U4131(.A(n2770), .B(n4446), .Y(dpath_n194));
AND2X1 mul_U4132(.A(n2771), .B(n4447), .Y(dpath_n201));
AND2X1 mul_U4133(.A(n2772), .B(n4448), .Y(dpath_n200));
AND2X1 mul_U4134(.A(n2773), .B(n4449), .Y(dpath_n207));
AND2X1 mul_U4135(.A(n2774), .B(n4450), .Y(dpath_n206));
AND2X1 mul_U4136(.A(n2775), .B(n4451), .Y(dpath_n213));
AND2X1 mul_U4137(.A(n2776), .B(n4452), .Y(dpath_n212));
AND2X1 mul_U4138(.A(n2777), .B(n4453), .Y(dpath_n219));
AND2X1 mul_U4139(.A(n2778), .B(n4454), .Y(dpath_n218));
AND2X1 mul_U4140(.A(n2779), .B(n4455), .Y(dpath_n225));
AND2X1 mul_U4141(.A(n2780), .B(n4456), .Y(dpath_n224));
AND2X1 mul_U4142(.A(n2781), .B(n4457), .Y(dpath_n231));
AND2X1 mul_U4143(.A(n2782), .B(n4458), .Y(dpath_n230));
AND2X1 mul_U4144(.A(n2783), .B(n4459), .Y(dpath_n237));
AND2X1 mul_U4145(.A(n2784), .B(n4460), .Y(dpath_n236));
AND2X1 mul_U4146(.A(n2785), .B(n4461), .Y(dpath_n243));
AND2X1 mul_U4147(.A(n2786), .B(n4462), .Y(dpath_n242));
AND2X1 mul_U4148(.A(n2787), .B(n4463), .Y(dpath_n249));
AND2X1 mul_U4149(.A(n2788), .B(n4464), .Y(dpath_n248));
AND2X1 mul_U4150(.A(n2791), .B(n4467), .Y(dpath_n261));
AND2X1 mul_U4151(.A(n2792), .B(n4468), .Y(dpath_n260));
AND2X1 mul_U4152(.A(n2793), .B(n4469), .Y(dpath_n267));
AND2X1 mul_U4153(.A(n2794), .B(n4470), .Y(dpath_n266));
AND2X1 mul_U4154(.A(n2795), .B(n4471), .Y(dpath_n273));
AND2X1 mul_U4155(.A(n2796), .B(n4472), .Y(dpath_n272));
AND2X1 mul_U4156(.A(n2797), .B(n4473), .Y(dpath_n279));
AND2X1 mul_U4157(.A(n2798), .B(n4474), .Y(dpath_n278));
AND2X1 mul_U4158(.A(n2799), .B(n4475), .Y(dpath_n285));
AND2X1 mul_U4159(.A(n2800), .B(n4476), .Y(dpath_n284));
AND2X1 mul_U4160(.A(n2801), .B(n4477), .Y(dpath_n291));
AND2X1 mul_U4161(.A(n2802), .B(n4478), .Y(dpath_n290));
AND2X1 mul_U4162(.A(n2803), .B(n4479), .Y(dpath_n297));
AND2X1 mul_U4163(.A(n2804), .B(n4480), .Y(dpath_n296));
INVX1 mul_U4164(.A(n9577), .Y(n9526));
AND2X1 mul_U4165(.A(n2805), .B(n4481), .Y(dpath_n303));
AND2X1 mul_U4166(.A(n2806), .B(n4482), .Y(dpath_n302));
INVX1 mul_U4167(.A(n9579), .Y(n9520));
AND2X1 mul_U4168(.A(n2807), .B(n4483), .Y(dpath_n309));
AND2X1 mul_U4169(.A(n2808), .B(n4484), .Y(dpath_n308));
INVX1 mul_U4170(.A(n9579), .Y(n9521));
AND2X1 mul_U4171(.A(n2809), .B(n4485), .Y(dpath_n315));
AND2X1 mul_U4172(.A(n2810), .B(n4486), .Y(dpath_n314));
AND2X1 mul_U4173(.A(n2813), .B(n4489), .Y(dpath_n327));
AND2X1 mul_U4174(.A(n2814), .B(n4490), .Y(dpath_n326));
AND2X1 mul_U4175(.A(n2815), .B(n4491), .Y(dpath_n333));
AND2X1 mul_U4176(.A(n2816), .B(n4492), .Y(dpath_n332));
AND2X1 mul_U4177(.A(n2817), .B(n4493), .Y(dpath_n339));
AND2X1 mul_U4178(.A(n2818), .B(n4494), .Y(dpath_n338));
AND2X1 mul_U4179(.A(n2819), .B(n4495), .Y(dpath_n345));
AND2X1 mul_U4180(.A(n2820), .B(n4496), .Y(dpath_n344));
AND2X1 mul_U4181(.A(n2821), .B(n4497), .Y(dpath_n351));
AND2X1 mul_U4182(.A(n2822), .B(n4498), .Y(dpath_n350));
AND2X1 mul_U4183(.A(n2823), .B(n4499), .Y(dpath_n357));
AND2X1 mul_U4184(.A(n2824), .B(n4500), .Y(dpath_n356));
AND2X1 mul_U4185(.A(n2825), .B(n4501), .Y(dpath_n363));
AND2X1 mul_U4186(.A(n2826), .B(n4502), .Y(dpath_n362));
AND2X1 mul_U4187(.A(n2827), .B(n4503), .Y(dpath_n369));
AND2X1 mul_U4188(.A(n2828), .B(n4504), .Y(dpath_n368));
INVX1 mul_U4189(.A(n9577), .Y(n9525));
OR2X1 mul_U4190(.A(n5871), .B(n5999), .Y(dpath_mulcore_booth_b15_in0[2]));
AND2X1 mul_U4191(.A(n2830), .B(n4506), .Y(dpath_n374));
AND2X1 mul_U4192(.A(n2463), .B(c0_act), .Y(dpath_mulcore_booth_out_mux0_n4));
AND2X1 mul_U4193(.A(n18013), .B(n4360), .Y(n18011));
AND2X1 mul_U4194(.A(n2470), .B(c0_act), .Y(dpath_mulcore_booth_out_mux0_n6));
AND2X1 mul_U4195(.A(dpath_acc_reg[129]), .B(n10598), .Y(n10602));
AND2X1 mul_U4196(.A(dpath_mulcore_add_co96), .B(dpath_acc_reg[132]), .Y(n10598));
AND2X1 mul_U4197(.A(n10595), .B(n10594), .Y(n10596));
AND2X1 mul_U4198(.A(dpath_acc_reg[132]), .B(dpath_acc_reg[131]), .Y(n10595));
AND2X1 mul_U4199(.A(n10592), .B(dpath_acc_reg[129]), .Y(n10594));
AND2X1 mul_U4200(.A(dpath_mulcore_add_co96), .B(dpath_acc_reg[130]), .Y(n10592));
AND2X1 mul_U4201(.A(n100), .B(n3183), .Y(n10582));
AND2X1 mul_U4202(.A(n99), .B(n3182), .Y(n10577));
AND2X1 mul_U4203(.A(n98), .B(n3181), .Y(n10572));
AND2X1 mul_U4204(.A(n97), .B(n3180), .Y(n10567));
AND2X1 mul_U4205(.A(n96), .B(n3179), .Y(n10562));
AND2X1 mul_U4206(.A(n95), .B(n3178), .Y(n10557));
AND2X1 mul_U4207(.A(n94), .B(n3177), .Y(n10552));
AND2X1 mul_U4208(.A(n93), .B(n3176), .Y(n10545));
AND2X1 mul_U4209(.A(n92), .B(n3175), .Y(n10540));
AND2X1 mul_U4210(.A(n91), .B(n3174), .Y(n10535));
AND2X1 mul_U4211(.A(n90), .B(n3173), .Y(n10530));
AND2X1 mul_U4212(.A(n89), .B(n3172), .Y(n10525));
AND2X1 mul_U4213(.A(n88), .B(n3171), .Y(n10520));
AND2X1 mul_U4214(.A(n87), .B(n3170), .Y(n10515));
AND2X1 mul_U4215(.A(n86), .B(n3169), .Y(n10510));
AND2X1 mul_U4216(.A(n85), .B(n3168), .Y(n10505));
AND2X1 mul_U4217(.A(n84), .B(n3167), .Y(n10500));
AND2X1 mul_U4218(.A(n83), .B(n3166), .Y(n10493));
AND2X1 mul_U4219(.A(n82), .B(n3165), .Y(n10488));
AND2X1 mul_U4220(.A(n81), .B(n3164), .Y(n10483));
AND2X1 mul_U4221(.A(n80), .B(n3163), .Y(n10478));
AND2X1 mul_U4222(.A(n79), .B(n3162), .Y(n10473));
AND2X1 mul_U4223(.A(n78), .B(n3161), .Y(n10468));
AND2X1 mul_U4224(.A(n77), .B(n3160), .Y(n10463));
AND2X1 mul_U4225(.A(n76), .B(n3159), .Y(n10458));
AND2X1 mul_U4226(.A(n75), .B(n3158), .Y(n10453));
AND2X1 mul_U4227(.A(n74), .B(n3157), .Y(n10448));
AND2X1 mul_U4228(.A(n73), .B(n3156), .Y(n10441));
AND2X1 mul_U4229(.A(n72), .B(n3155), .Y(n10436));
AND2X1 mul_U4230(.A(n71), .B(n3154), .Y(n10431));
AND2X1 mul_U4231(.A(n70), .B(n3153), .Y(n10426));
AND2X1 mul_U4232(.A(n69), .B(n3152), .Y(n10421));
AND2X1 mul_U4233(.A(n68), .B(n3151), .Y(n10416));
AND2X1 mul_U4234(.A(n67), .B(n3150), .Y(n10411));
AND2X1 mul_U4235(.A(n66), .B(n3149), .Y(n10406));
AND2X1 mul_U4236(.A(n65), .B(n3148), .Y(n10401));
AND2X1 mul_U4237(.A(n64), .B(n3147), .Y(n10396));
AND2X1 mul_U4238(.A(n63), .B(n3146), .Y(n10389));
AND2X1 mul_U4239(.A(n62), .B(n3145), .Y(n10384));
AND2X1 mul_U4240(.A(n61), .B(n3144), .Y(n10379));
AND2X1 mul_U4241(.A(n60), .B(n3143), .Y(n10374));
AND2X1 mul_U4242(.A(n59), .B(n3142), .Y(n10369));
AND2X1 mul_U4243(.A(n58), .B(n3141), .Y(n10364));
AND2X1 mul_U4244(.A(n57), .B(n3140), .Y(n10359));
AND2X1 mul_U4245(.A(n56), .B(n3139), .Y(n10354));
AND2X1 mul_U4246(.A(n55), .B(n3138), .Y(n10349));
AND2X1 mul_U4247(.A(n54), .B(n3137), .Y(n10344));
AND2X1 mul_U4248(.A(n53), .B(n3136), .Y(n10337));
AND2X1 mul_U4249(.A(n52), .B(n3135), .Y(n10332));
AND2X1 mul_U4250(.A(n51), .B(n3134), .Y(n10327));
AND2X1 mul_U4251(.A(n50), .B(n3133), .Y(n10322));
AND2X1 mul_U4252(.A(n49), .B(n3132), .Y(n10317));
AND2X1 mul_U4253(.A(n48), .B(n3131), .Y(n10312));
AND2X1 mul_U4254(.A(n47), .B(n3130), .Y(n10307));
AND2X1 mul_U4255(.A(n46), .B(n3129), .Y(n10302));
AND2X1 mul_U4256(.A(n45), .B(n3128), .Y(n10297));
AND2X1 mul_U4257(.A(n44), .B(n3127), .Y(n10590));
AND2X1 mul_U4258(.A(n43), .B(n3126), .Y(n10588));
AND2X1 mul_U4259(.A(n42), .B(n3125), .Y(n10586));
AND2X1 mul_U4260(.A(n41), .B(n3124), .Y(n10584));
AND2X1 mul_U4261(.A(n40), .B(n3123), .Y(n10551));
AND2X1 mul_U4262(.A(n39), .B(n3122), .Y(n10499));
AND2X1 mul_U4263(.A(n38), .B(n3121), .Y(n10447));
AND2X1 mul_U4264(.A(n37), .B(n3120), .Y(n10395));
AND2X1 mul_U4265(.A(n36), .B(n3119), .Y(n10343));
AND2X1 mul_U4266(.A(n35), .B(n3118), .Y(dpath_mulcore_add_co31));
AND2X1 mul_U4267(.A(n34), .B(n3117), .Y(n10247));
AND2X1 mul_U4268(.A(n33), .B(n3116), .Y(n10242));
AND2X1 mul_U4269(.A(n32), .B(n3115), .Y(n10237));
AND2X1 mul_U4270(.A(n31), .B(n3114), .Y(n10230));
AND2X1 mul_U4271(.A(n30), .B(n3113), .Y(n10225));
AND2X1 mul_U4272(.A(n29), .B(n3112), .Y(n10220));
AND2X1 mul_U4273(.A(n28), .B(n3111), .Y(n10215));
AND2X1 mul_U4274(.A(n27), .B(n3110), .Y(n10210));
AND2X1 mul_U4275(.A(n26), .B(n3109), .Y(n10205));
AND2X1 mul_U4276(.A(n25), .B(n3108), .Y(n10200));
AND2X1 mul_U4277(.A(n24), .B(n3107), .Y(n10195));
AND2X1 mul_U4278(.A(n23), .B(n3106), .Y(n10190));
AND2X1 mul_U4279(.A(n22), .B(n3105), .Y(n10185));
AND2X1 mul_U4280(.A(n21), .B(n3104), .Y(n10178));
AND2X1 mul_U4281(.A(n20), .B(n3103), .Y(n10173));
AND2X1 mul_U4282(.A(n19), .B(n3102), .Y(n10168));
AND2X1 mul_U4283(.A(n18), .B(n3101), .Y(n10163));
AND2X1 mul_U4284(.A(n17), .B(n3100), .Y(n10158));
AND2X1 mul_U4285(.A(n16), .B(n3099), .Y(n10153));
AND2X1 mul_U4286(.A(n15), .B(n3098), .Y(n10148));
AND2X1 mul_U4287(.A(n14), .B(n3097), .Y(n10143));
AND2X1 mul_U4288(.A(n13), .B(n3096), .Y(n10138));
AND2X1 mul_U4289(.A(n12), .B(n3095), .Y(n10264));
AND2X1 mul_U4290(.A(n11), .B(n3094), .Y(n10262));
AND2X1 mul_U4291(.A(n10), .B(n3093), .Y(n10260));
AND2X1 mul_U4292(.A(n9), .B(n3092), .Y(n10258));
INVX1 mul_U4293(.A(n9580), .Y(n9515));
AND2X1 mul_U4294(.A(n8), .B(n3091), .Y(n10256));
INVX1 mul_U4295(.A(n9580), .Y(n9516));
AND2X1 mul_U4296(.A(n7), .B(n3090), .Y(n10254));
AND2X1 mul_U4297(.A(n6), .B(n3089), .Y(n10252));
AND2X1 mul_U4298(.A(n5), .B(n3088), .Y(n10236));
AND2X1 mul_U4299(.A(dpath_mulcore_addin_cin), .B(dpath_mulcore_addin_sum[0]), .Y(n10184));
AND2X1 mul_U4300(.A(n1856), .B(n3910), .Y(dpath_mulcore_pcout[96]));
AND2X1 mul_U4301(.A(n1857), .B(n3911), .Y(dpath_mulcore_pcout[95]));
AND2X1 mul_U4302(.A(n1858), .B(n3912), .Y(dpath_mulcore_pcout[94]));
AND2X1 mul_U4303(.A(n1859), .B(n3913), .Y(dpath_mulcore_pcout[93]));
AND2X1 mul_U4304(.A(n1860), .B(n3914), .Y(dpath_mulcore_pcout[92]));
AND2X1 mul_U4305(.A(n1861), .B(n3915), .Y(dpath_mulcore_pcout[91]));
AND2X1 mul_U4306(.A(n1862), .B(n3916), .Y(dpath_mulcore_pcout[90]));
AND2X1 mul_U4307(.A(n1863), .B(n3917), .Y(dpath_mulcore_pcout[89]));
AND2X1 mul_U4308(.A(n1864), .B(n3918), .Y(dpath_mulcore_pcout[88]));
AND2X1 mul_U4309(.A(n1865), .B(n3919), .Y(dpath_mulcore_pcout[87]));
AND2X1 mul_U4310(.A(n1866), .B(n3920), .Y(dpath_mulcore_pcout[86]));
AND2X1 mul_U4311(.A(n1867), .B(n3921), .Y(dpath_mulcore_pcout[85]));
AND2X1 mul_U4312(.A(n1868), .B(n3922), .Y(dpath_mulcore_pcout[84]));
AND2X1 mul_U4313(.A(n1891), .B(n3944), .Y(dpath_mulcore_pcout[83]));
AND2X1 mul_U4314(.A(n1806), .B(n3860), .Y(dpath_mulcore_pcout[82]));
AND2X1 mul_U4315(.A(n1869), .B(n3923), .Y(dpath_mulcore_pcout[81]));
AND2X1 mul_U4316(.A(n1870), .B(n3924), .Y(dpath_mulcore_pcout[80]));
AND2X1 mul_U4317(.A(n1871), .B(n3925), .Y(dpath_mulcore_pcout[79]));
AND2X1 mul_U4318(.A(n1872), .B(n3926), .Y(dpath_mulcore_pcout[78]));
AND2X1 mul_U4319(.A(n1873), .B(n3927), .Y(dpath_mulcore_pcout[77]));
AND2X1 mul_U4320(.A(n1874), .B(n3928), .Y(dpath_mulcore_pcout[76]));
AND2X1 mul_U4321(.A(n1875), .B(n3929), .Y(dpath_mulcore_pcout[75]));
AND2X1 mul_U4322(.A(n1876), .B(n3930), .Y(dpath_mulcore_pcout[74]));
AND2X1 mul_U4323(.A(n1877), .B(n3931), .Y(dpath_mulcore_pcout[73]));
AND2X1 mul_U4324(.A(n1878), .B(n3932), .Y(dpath_mulcore_pcout[72]));
AND2X1 mul_U4325(.A(n1879), .B(n3933), .Y(dpath_mulcore_pcout[71]));
AND2X1 mul_U4326(.A(n1880), .B(n3934), .Y(dpath_mulcore_pcout[70]));
AND2X1 mul_U4327(.A(n1881), .B(n3935), .Y(dpath_mulcore_pcout[69]));
AND2X1 mul_U4328(.A(n1807), .B(n3861), .Y(dpath_mulcore_pcout[68]));
AND2X1 mul_U4329(.A(n1808), .B(n3862), .Y(dpath_mulcore_pcout[67]));
AND2X1 mul_U4330(.A(n1809), .B(n3863), .Y(dpath_mulcore_pcout[66]));
AND2X1 mul_U4331(.A(n1810), .B(n3864), .Y(dpath_mulcore_pcout[65]));
AND2X1 mul_U4332(.A(n1811), .B(n3865), .Y(dpath_mulcore_pcout[64]));
AND2X1 mul_U4333(.A(n1812), .B(n3866), .Y(dpath_mulcore_pcout[63]));
AND2X1 mul_U4334(.A(n1813), .B(n3867), .Y(dpath_mulcore_pcout[62]));
AND2X1 mul_U4335(.A(n1814), .B(n3868), .Y(dpath_mulcore_pcout[61]));
AND2X1 mul_U4336(.A(n1815), .B(n3869), .Y(dpath_mulcore_pcout[60]));
AND2X1 mul_U4337(.A(n1816), .B(n3870), .Y(dpath_mulcore_pcout[59]));
AND2X1 mul_U4338(.A(n1817), .B(n3871), .Y(dpath_mulcore_pcout[58]));
AND2X1 mul_U4339(.A(n1818), .B(n3872), .Y(dpath_mulcore_pcout[57]));
AND2X1 mul_U4340(.A(n1819), .B(n3873), .Y(dpath_mulcore_pcout[56]));
AND2X1 mul_U4341(.A(n1820), .B(n3874), .Y(dpath_mulcore_pcout[55]));
AND2X1 mul_U4342(.A(n1821), .B(n3875), .Y(dpath_mulcore_pcout[54]));
AND2X1 mul_U4343(.A(n1822), .B(n3876), .Y(dpath_mulcore_pcout[53]));
AND2X1 mul_U4344(.A(n1823), .B(n3877), .Y(dpath_mulcore_pcout[52]));
AND2X1 mul_U4345(.A(n1824), .B(n3878), .Y(dpath_mulcore_pcout[51]));
AND2X1 mul_U4346(.A(n1825), .B(n3879), .Y(dpath_mulcore_pcout[50]));
AND2X1 mul_U4347(.A(n1826), .B(n3880), .Y(dpath_mulcore_pcout[49]));
AND2X1 mul_U4348(.A(n1827), .B(n3881), .Y(dpath_mulcore_pcout[48]));
AND2X1 mul_U4349(.A(n1828), .B(n3882), .Y(dpath_mulcore_pcout[47]));
AND2X1 mul_U4350(.A(n1829), .B(n3883), .Y(dpath_mulcore_pcout[46]));
AND2X1 mul_U4351(.A(n1830), .B(n3884), .Y(dpath_mulcore_pcout[45]));
AND2X1 mul_U4352(.A(n1831), .B(n3885), .Y(dpath_mulcore_pcout[44]));
AND2X1 mul_U4353(.A(n1832), .B(n3886), .Y(dpath_mulcore_pcout[43]));
AND2X1 mul_U4354(.A(n1833), .B(n3887), .Y(dpath_mulcore_pcout[42]));
AND2X1 mul_U4355(.A(n1834), .B(n3888), .Y(dpath_mulcore_pcout[41]));
AND2X1 mul_U4356(.A(n1835), .B(n3889), .Y(dpath_mulcore_pcout[40]));
AND2X1 mul_U4357(.A(n1836), .B(n3890), .Y(dpath_mulcore_pcout[39]));
AND2X1 mul_U4358(.A(n1837), .B(n3891), .Y(dpath_mulcore_pcout[38]));
AND2X1 mul_U4359(.A(n1838), .B(n3892), .Y(dpath_mulcore_pcout[37]));
INVX1 mul_U4360(.A(n9580), .Y(n9514));
AND2X1 mul_U4361(.A(n1839), .B(n3893), .Y(dpath_mulcore_pcout[36]));
AND2X1 mul_U4362(.A(n1840), .B(n3894), .Y(dpath_mulcore_pcout[35]));
AND2X1 mul_U4363(.A(n1841), .B(n3895), .Y(dpath_mulcore_pcout[34]));
AND2X1 mul_U4364(.A(n1842), .B(n3896), .Y(dpath_mulcore_pcout[33]));
AND2X1 mul_U4365(.A(n1843), .B(n3897), .Y(dpath_mulcore_pcout[32]));
AND2X1 mul_U4366(.A(n1844), .B(n3898), .Y(dpath_mulcore_pcout[31]));
AND2X1 mul_U4367(.A(n1845), .B(n3899), .Y(dpath_mulcore_pcout[30]));
INVX1 mul_U4368(.A(n9500), .Y(n9510));
INVX1 mul_U4369(.A(n9501), .Y(n9511));
INVX1 mul_U4370(.A(n9576), .Y(n9527));
INVX1 mul_U4371(.A(n9575), .Y(n9530));
INVX1 mul_U4372(.A(n9578), .Y(n9522));
INVX1 mul_U4373(.A(n9578), .Y(n9523));
INVX1 mul_U4374(.A(n9578), .Y(n9524));
INVX1 mul_U4375(.A(n9593), .Y(n9662));
INVX1 mul_U4376(.A(n9593), .Y(n9661));
INVX1 mul_U4377(.A(n9569), .Y(n9548));
INVX1 mul_U4378(.A(n9569), .Y(n9549));
AND2X1 mul_U4379(.A(n14968), .B(dpath_mulcore_array2_s1x2), .Y(dpath_mulcore_pcoutx2));
INVX1 mul_U4380(.A(n9493), .Y(n9568));
AND2X1 mul_U4381(.A(n1599), .B(n1), .Y(dpath_mulcore_ary1_a0_c_2[76]));
AND2X1 mul_U4382(.A(n2480), .B(n4406), .Y(dpath_mulcore_ary1_a0_co[71]));
AND2X1 mul_U4383(.A(n2072), .B(n4121), .Y(dpath_mulcore_ary1_a0_co[70]));
AND2X1 mul_U4384(.A(n2074), .B(n4122), .Y(dpath_mulcore_ary1_a0_co[69]));
AND2X1 mul_U4385(.A(n2076), .B(n4123), .Y(dpath_mulcore_ary1_a0_co[68]));
AND2X1 mul_U4386(.A(n2078), .B(n4124), .Y(dpath_mulcore_ary1_a0_co[67]));
AND2X1 mul_U4387(.A(n2080), .B(n4125), .Y(dpath_mulcore_ary1_a0_co[66]));
AND2X1 mul_U4388(.A(n2082), .B(n4126), .Y(dpath_mulcore_ary1_a0_co[65]));
AND2X1 mul_U4389(.A(n2084), .B(n4127), .Y(dpath_mulcore_ary1_a0_co[64]));
AND2X1 mul_U4390(.A(n2086), .B(n4128), .Y(dpath_mulcore_ary1_a0_co[63]));
AND2X1 mul_U4391(.A(n2088), .B(n4129), .Y(dpath_mulcore_ary1_a0_co[62]));
AND2X1 mul_U4392(.A(n2090), .B(n4130), .Y(dpath_mulcore_ary1_a0_co[61]));
AND2X1 mul_U4393(.A(n2092), .B(n4131), .Y(dpath_mulcore_ary1_a0_co[60]));
AND2X1 mul_U4394(.A(n2094), .B(n4132), .Y(dpath_mulcore_ary1_a0_co[59]));
AND2X1 mul_U4395(.A(n2096), .B(n4133), .Y(dpath_mulcore_ary1_a0_co[58]));
AND2X1 mul_U4396(.A(n2098), .B(n4134), .Y(dpath_mulcore_ary1_a0_co[57]));
AND2X1 mul_U4397(.A(n2100), .B(n4135), .Y(dpath_mulcore_ary1_a0_co[56]));
AND2X1 mul_U4398(.A(n2102), .B(n4136), .Y(dpath_mulcore_ary1_a0_co[55]));
AND2X1 mul_U4399(.A(n2104), .B(n4137), .Y(dpath_mulcore_ary1_a0_co[54]));
AND2X1 mul_U4400(.A(n2106), .B(n4138), .Y(dpath_mulcore_ary1_a0_co[53]));
AND2X1 mul_U4401(.A(n2108), .B(n4139), .Y(dpath_mulcore_ary1_a0_co[52]));
AND2X1 mul_U4402(.A(n2110), .B(n4140), .Y(dpath_mulcore_ary1_a0_co[51]));
INVX1 mul_U4403(.A(n9565), .Y(n9561));
AND2X1 mul_U4404(.A(n2112), .B(n4141), .Y(dpath_mulcore_ary1_a0_co[50]));
INVX1 mul_U4405(.A(n9583), .Y(n9502));
AND2X1 mul_U4406(.A(n2114), .B(n4142), .Y(dpath_mulcore_ary1_a0_co[49]));
INVX1 mul_U4407(.A(n9583), .Y(n9503));
AND2X1 mul_U4408(.A(n2116), .B(n4143), .Y(dpath_mulcore_ary1_a0_co[48]));
INVX1 mul_U4409(.A(n9582), .Y(n9504));
AND2X1 mul_U4410(.A(n2118), .B(n4144), .Y(dpath_mulcore_ary1_a0_co[47]));
INVX1 mul_U4411(.A(n9582), .Y(n9505));
AND2X1 mul_U4412(.A(n2120), .B(n4145), .Y(dpath_mulcore_ary1_a0_co[46]));
INVX1 mul_U4413(.A(n9582), .Y(n9506));
AND2X1 mul_U4414(.A(n2122), .B(n4146), .Y(dpath_mulcore_ary1_a0_co[45]));
INVX1 mul_U4415(.A(n9581), .Y(n9508));
AND2X1 mul_U4416(.A(n2124), .B(n4147), .Y(dpath_mulcore_ary1_a0_co[44]));
AND2X1 mul_U4417(.A(n2126), .B(n4148), .Y(dpath_mulcore_ary1_a0_co[43]));
AND2X1 mul_U4418(.A(n2128), .B(n4149), .Y(dpath_mulcore_ary1_a0_co[42]));
AND2X1 mul_U4419(.A(n2130), .B(n4150), .Y(dpath_mulcore_ary1_a0_co[41]));
AND2X1 mul_U4420(.A(n2132), .B(n4151), .Y(dpath_mulcore_ary1_a0_co[40]));
AND2X1 mul_U4421(.A(n2134), .B(n4152), .Y(dpath_mulcore_ary1_a0_co[39]));
AND2X1 mul_U4422(.A(n2136), .B(n4153), .Y(dpath_mulcore_ary1_a0_co[38]));
AND2X1 mul_U4423(.A(n2138), .B(n4154), .Y(dpath_mulcore_ary1_a0_co[37]));
AND2X1 mul_U4424(.A(n2140), .B(n4155), .Y(dpath_mulcore_ary1_a0_co[36]));
AND2X1 mul_U4425(.A(n2142), .B(n4156), .Y(dpath_mulcore_ary1_a0_co[35]));
AND2X1 mul_U4426(.A(n2144), .B(n4157), .Y(dpath_mulcore_ary1_a0_co[34]));
AND2X1 mul_U4427(.A(n2146), .B(n4158), .Y(dpath_mulcore_ary1_a0_co[33]));
AND2X1 mul_U4428(.A(n2148), .B(n4159), .Y(dpath_mulcore_ary1_a0_co[32]));
AND2X1 mul_U4429(.A(n2150), .B(n4160), .Y(dpath_mulcore_ary1_a0_co[31]));
AND2X1 mul_U4430(.A(n2152), .B(n4161), .Y(dpath_mulcore_ary1_a0_co[30]));
AND2X1 mul_U4431(.A(n2154), .B(n4162), .Y(dpath_mulcore_ary1_a0_co[29]));
AND2X1 mul_U4432(.A(n2156), .B(n4163), .Y(dpath_mulcore_ary1_a0_co[28]));
AND2X1 mul_U4433(.A(n2158), .B(n4164), .Y(dpath_mulcore_ary1_a0_co[27]));
AND2X1 mul_U4434(.A(n2160), .B(n4165), .Y(dpath_mulcore_ary1_a0_co[26]));
AND2X1 mul_U4435(.A(n2162), .B(n4166), .Y(dpath_mulcore_ary1_a0_co[25]));
AND2X1 mul_U4436(.A(n2164), .B(n4167), .Y(dpath_mulcore_ary1_a0_co[24]));
AND2X1 mul_U4437(.A(n2166), .B(n4168), .Y(dpath_mulcore_ary1_a0_co[23]));
AND2X1 mul_U4438(.A(n2168), .B(n4169), .Y(dpath_mulcore_ary1_a0_co[22]));
AND2X1 mul_U4439(.A(n2170), .B(n4170), .Y(dpath_mulcore_ary1_a0_co[21]));
AND2X1 mul_U4440(.A(n2172), .B(n4171), .Y(dpath_mulcore_ary1_a0_co[20]));
AND2X1 mul_U4441(.A(n2174), .B(n4172), .Y(dpath_mulcore_ary1_a0_co[19]));
AND2X1 mul_U4442(.A(n2176), .B(n4173), .Y(dpath_mulcore_ary1_a0_co[18]));
AND2X1 mul_U4443(.A(n2178), .B(n4174), .Y(dpath_mulcore_ary1_a0_co[17]));
AND2X1 mul_U4444(.A(n2180), .B(n4175), .Y(dpath_mulcore_ary1_a0_co[16]));
AND2X1 mul_U4445(.A(n2182), .B(n4176), .Y(dpath_mulcore_ary1_a0_co[15]));
AND2X1 mul_U4446(.A(n2184), .B(n4177), .Y(dpath_mulcore_ary1_a0_co[14]));
AND2X1 mul_U4447(.A(n2186), .B(n4178), .Y(dpath_mulcore_ary1_a0_co[13]));
AND2X1 mul_U4448(.A(n2188), .B(n4179), .Y(dpath_mulcore_ary1_a0_co[12]));
AND2X1 mul_U4449(.A(n2190), .B(n4180), .Y(dpath_mulcore_ary1_a0_co[11]));
AND2X1 mul_U4450(.A(n1125), .B(n3186), .Y(dpath_mulcore_ary1_a0_c1[2]));
INVX1 mul_U4451(.A(n9572), .Y(n9537));
AND2X1 mul_U4452(.A(n7397), .B(dpath_mulcore_ary1_a0_I1_I0_b0n), .Y(dpath_mulcore_ary1_a0_c1[1]));
INVX1 mul_U4453(.A(n9572), .Y(n9538));
INVX1 mul_U4454(.A(n9566), .Y(n9557));
INVX1 mul_U4455(.A(n9574), .Y(n9533));
AND2X1 mul_U4456(.A(dpath_mulcore_ary1_a0_s0[2]), .B(dpath_mulcore_ary1_a0_c0[1]), .Y(dpath_mulcore_ary1_a0_c_1[2]));
INVX1 mul_U4457(.A(n9573), .Y(n9534));
AND2X1 mul_U4458(.A(n7398), .B(dpath_mulcore_ary1_a0_I0_I0_b0n), .Y(dpath_mulcore_ary1_a0_c0[1]));
INVX1 mul_U4459(.A(n9581), .Y(n9507));
AND2X1 mul_U4460(.A(n604), .B(n12126), .Y(dpath_mulcore_ary1_a0_I0_I0_p0_1));
OR2X1 mul_U4461(.A(n6678), .B(dpath_mulcore_b0[0]), .Y(n12126));
OR2X1 mul_U4462(.A(n13701), .B(n5935), .Y(dpath_mulcore_ary1_a0_I0_I0_b0n));
AND2X1 mul_U4463(.A(n7403), .B(n9841), .Y(n13701));
INVX1 mul_U4464(.A(n9573), .Y(n9535));
INVX1 mul_U4465(.A(n12128), .Y(n9841));
OR2X1 mul_U4466(.A(n6679), .B(dpath_mulcore_b0[0]), .Y(n12128));
OR2X1 mul_U4467(.A(n9721), .B(n5934), .Y(dpath_mulcore_ary1_a0_I0_I0_b0n_0));
INVX1 mul_U4468(.A(n9572), .Y(n9536));
OR2X1 mul_U4469(.A(n9312), .B(dpath_mulcore_b7[0]), .Y(n13661));
INVX1 mul_U4470(.A(dpath_mulcore_ary1_a0_sc3_76__z), .Y(n10027));
INVX1 mul_U4471(.A(dpath_mulcore_ary1_a0_sc3_75__z), .Y(n10023));
INVX1 mul_U4472(.A(dpath_mulcore_ary1_a0_sc3_74__z), .Y(n10020));
INVX1 mul_U4473(.A(dpath_mulcore_ary1_a0_sc3_73__z), .Y(n10017));
INVX1 mul_U4474(.A(dpath_mulcore_ary1_a0_sc3_72__z), .Y(n10014));
INVX1 mul_U4475(.A(dpath_mulcore_ary1_a0_sc3_71__z), .Y(n10011));
INVX1 mul_U4476(.A(dpath_mulcore_ary1_a0_sc3_70__z), .Y(n10008));
INVX1 mul_U4477(.A(dpath_mulcore_ary1_a0_sc3_69__z), .Y(n9819));
INVX1 mul_U4478(.A(dpath_mulcore_ary1_a0_sc3_68__z), .Y(n9820));
INVX1 mul_U4479(.A(dpath_mulcore_ary1_a0_sc3_67__z), .Y(n9821));
INVX1 mul_U4480(.A(dpath_mulcore_ary1_a0_sc3_66__z), .Y(n9822));
INVX1 mul_U4481(.A(dpath_mulcore_ary1_a0_sc3_65__z), .Y(n9823));
INVX1 mul_U4482(.A(dpath_mulcore_ary1_a0_sc3_64__z), .Y(n9995));
INVX1 mul_U4483(.A(dpath_mulcore_ary1_a0_sc3_63__z), .Y(n9992));
INVX1 mul_U4484(.A(dpath_mulcore_ary1_a0_sc3_62__z), .Y(n9989));
INVX1 mul_U4485(.A(dpath_mulcore_ary1_a0_sc3_61__z), .Y(n9986));
INVX1 mul_U4486(.A(dpath_mulcore_ary1_a0_sc3_60__z), .Y(n9983));
INVX1 mul_U4487(.A(dpath_mulcore_ary1_a0_sc3_59__z), .Y(n9980));
INVX1 mul_U4488(.A(dpath_mulcore_ary1_a0_sc3_58__z), .Y(n9977));
INVX1 mul_U4489(.A(dpath_mulcore_ary1_a0_sc3_57__z), .Y(n9974));
INVX1 mul_U4490(.A(dpath_mulcore_ary1_a0_sc3_56__z), .Y(n9971));
INVX1 mul_U4491(.A(dpath_mulcore_ary1_a0_sc3_55__z), .Y(n9968));
INVX1 mul_U4492(.A(dpath_mulcore_ary1_a0_sc3_54__z), .Y(n9965));
INVX1 mul_U4493(.A(dpath_mulcore_ary1_a0_sc3_53__z), .Y(n9962));
INVX1 mul_U4494(.A(dpath_mulcore_ary1_a0_sc3_52__z), .Y(n9959));
INVX1 mul_U4495(.A(dpath_mulcore_ary1_a0_sc3_51__z), .Y(n9956));
INVX1 mul_U4496(.A(dpath_mulcore_ary1_a0_sc3_50__z), .Y(n9953));
INVX1 mul_U4497(.A(dpath_mulcore_ary1_a0_sc3_49__z), .Y(n9950));
INVX1 mul_U4498(.A(dpath_mulcore_ary1_a0_sc3_48__z), .Y(n9947));
INVX1 mul_U4499(.A(dpath_mulcore_ary1_a0_sc3_47__z), .Y(n9944));
INVX1 mul_U4500(.A(dpath_mulcore_ary1_a0_sc3_46__z), .Y(n9941));
INVX1 mul_U4501(.A(dpath_mulcore_ary1_a0_sc3_45__z), .Y(n9938));
INVX1 mul_U4502(.A(dpath_mulcore_ary1_a0_sc3_44__z), .Y(n9935));
INVX1 mul_U4503(.A(dpath_mulcore_ary1_a0_sc3_43__z), .Y(n9932));
INVX1 mul_U4504(.A(dpath_mulcore_ary1_a0_sc3_42__z), .Y(n9929));
INVX1 mul_U4505(.A(dpath_mulcore_ary1_a0_sc3_41__z), .Y(n9926));
INVX1 mul_U4506(.A(dpath_mulcore_ary1_a0_sc3_40__z), .Y(n9923));
INVX1 mul_U4507(.A(dpath_mulcore_ary1_a0_sc3_39__z), .Y(n9920));
INVX1 mul_U4508(.A(dpath_mulcore_ary1_a0_sc3_38__z), .Y(n9917));
INVX1 mul_U4509(.A(dpath_mulcore_ary1_a0_sc3_37__z), .Y(n9914));
INVX1 mul_U4510(.A(dpath_mulcore_ary1_a0_sc3_36__z), .Y(n9911));
INVX1 mul_U4511(.A(dpath_mulcore_ary1_a0_sc3_35__z), .Y(n9908));
INVX1 mul_U4512(.A(dpath_mulcore_ary1_a0_sc3_34__z), .Y(n9905));
INVX1 mul_U4513(.A(dpath_mulcore_ary1_a0_sc3_33__z), .Y(n9902));
INVX1 mul_U4514(.A(dpath_mulcore_ary1_a0_sc3_32__z), .Y(n9899));
INVX1 mul_U4515(.A(dpath_mulcore_ary1_a0_sc3_31__z), .Y(n9896));
INVX1 mul_U4516(.A(dpath_mulcore_ary1_a0_sc3_30__z), .Y(n9893));
INVX1 mul_U4517(.A(dpath_mulcore_ary1_a0_sc3_29__z), .Y(n9890));
INVX1 mul_U4518(.A(dpath_mulcore_ary1_a0_sc3_28__z), .Y(n9887));
INVX1 mul_U4519(.A(dpath_mulcore_ary1_a0_sc3_27__z), .Y(n9884));
INVX1 mul_U4520(.A(dpath_mulcore_ary1_a0_sc3_26__z), .Y(n9881));
INVX1 mul_U4521(.A(dpath_mulcore_ary1_a0_sc3_25__z), .Y(n9878));
INVX1 mul_U4522(.A(dpath_mulcore_ary1_a0_sc3_24__z), .Y(n9875));
INVX1 mul_U4523(.A(dpath_mulcore_ary1_a0_sc3_23__z), .Y(n9872));
INVX1 mul_U4524(.A(dpath_mulcore_ary1_a0_sc3_22__z), .Y(n9869));
INVX1 mul_U4525(.A(dpath_mulcore_ary1_a0_sc3_21__z), .Y(n9866));
INVX1 mul_U4526(.A(dpath_mulcore_ary1_a0_sc3_20__z), .Y(n9863));
INVX1 mul_U4527(.A(dpath_mulcore_ary1_a0_sc3_19__z), .Y(n9860));
INVX1 mul_U4528(.A(dpath_mulcore_ary1_a0_sc3_18__z), .Y(n9857));
INVX1 mul_U4529(.A(dpath_mulcore_ary1_a0_sc3_17__z), .Y(n9849));
INVX1 mul_U4530(.A(n9567), .Y(n9553));
INVX1 mul_U4531(.A(dpath_mulcore_ary1_a0_sc3_16__z), .Y(n9850));
INVX1 mul_U4532(.A(n9567), .Y(n9554));
INVX1 mul_U4533(.A(dpath_mulcore_ary1_a0_sc3_15__z), .Y(n9851));
INVX1 mul_U4534(.A(n9567), .Y(n9555));
INVX1 mul_U4535(.A(dpath_mulcore_ary1_a0_sc3_14__z), .Y(n9852));
INVX1 mul_U4536(.A(n9564), .Y(n9562));
INVX1 mul_U4537(.A(dpath_mulcore_ary1_a0_sc3_13__z), .Y(n9846));
INVX1 mul_U4538(.A(n9564), .Y(n9563));
INVX1 mul_U4539(.A(dpath_mulcore_ary1_a0_sc3_12__z), .Y(n9847));
INVX1 mul_U4540(.A(n9566), .Y(n9556));
AND2X1 mul_U4541(.A(n1598), .B(n3662), .Y(dpath_mulcore_ary1_a0_c_2[10]));
INVX1 mul_U4542(.A(n9566), .Y(n9558));
AND2X1 mul_U4543(.A(n1669), .B(n3728), .Y(dpath_mulcore_ary1_a0_c_1[6]));
AND2X1 mul_U4544(.A(n1670), .B(n3729), .Y(dpath_mulcore_ary1_a0_c_1[5]));
INVX1 mul_U4545(.A(n9570), .Y(n9546));
AND2X1 mul_U4546(.A(n1671), .B(n3730), .Y(dpath_mulcore_ary1_a0_c_1[4]));
INVX1 mul_U4547(.A(n9570), .Y(n9547));
AND2X1 mul_U4548(.A(n1603), .B(n3665), .Y(dpath_mulcore_ary1_a0_c_1[3]));
OR2X1 mul_U4549(.A(spu_mul_op1_data[63]), .B(n7198), .Y(dpath_n9));
OR2X1 mul_U4550(.A(spu_mul_op1_data[62]), .B(n9773), .Y(dpath_n11));
OR2X1 mul_U4551(.A(spu_mul_op1_data[61]), .B(n9773), .Y(dpath_n13));
OR2X1 mul_U4552(.A(spu_mul_op1_data[60]), .B(n7198), .Y(dpath_n15));
OR2X1 mul_U4553(.A(spu_mul_op1_data[59]), .B(n9773), .Y(dpath_n17));
OR2X1 mul_U4554(.A(spu_mul_op1_data[58]), .B(n7198), .Y(dpath_n19));
OR2X1 mul_U4555(.A(spu_mul_op1_data[57]), .B(n9772), .Y(dpath_n21));
OR2X1 mul_U4556(.A(spu_mul_op1_data[56]), .B(n9774), .Y(dpath_n23));
OR2X1 mul_U4557(.A(spu_mul_op1_data[55]), .B(n9772), .Y(dpath_n25));
OR2X1 mul_U4558(.A(spu_mul_op1_data[54]), .B(n9772), .Y(dpath_n27));
OR2X1 mul_U4559(.A(spu_mul_op1_data[53]), .B(n9774), .Y(dpath_n29));
OR2X1 mul_U4560(.A(spu_mul_op1_data[52]), .B(n9772), .Y(dpath_n31));
OR2X1 mul_U4561(.A(spu_mul_op1_data[51]), .B(n9773), .Y(dpath_n33));
OR2X1 mul_U4562(.A(spu_mul_op1_data[50]), .B(n7198), .Y(dpath_n35));
OR2X1 mul_U4563(.A(spu_mul_op1_data[49]), .B(n9774), .Y(dpath_n37));
OR2X1 mul_U4564(.A(spu_mul_op1_data[48]), .B(n9772), .Y(dpath_n39));
OR2X1 mul_U4565(.A(spu_mul_op1_data[47]), .B(n9773), .Y(dpath_n41));
OR2X1 mul_U4566(.A(spu_mul_op1_data[46]), .B(n7198), .Y(dpath_n43));
OR2X1 mul_U4567(.A(spu_mul_op1_data[45]), .B(n9774), .Y(dpath_n45));
OR2X1 mul_U4568(.A(spu_mul_op1_data[44]), .B(n9772), .Y(dpath_n47));
OR2X1 mul_U4569(.A(spu_mul_op1_data[43]), .B(n9773), .Y(dpath_n49));
OR2X1 mul_U4570(.A(spu_mul_op1_data[42]), .B(n7198), .Y(dpath_n51));
OR2X1 mul_U4571(.A(spu_mul_op1_data[41]), .B(n9774), .Y(dpath_n53));
INVX1 mul_U4572(.A(n9772), .Y(n9771));
OR2X1 mul_U4573(.A(spu_mul_op1_data[40]), .B(n9772), .Y(dpath_n55));
OR2X1 mul_U4574(.A(spu_mul_op1_data[39]), .B(n9773), .Y(dpath_n57));
OR2X1 mul_U4575(.A(spu_mul_op1_data[38]), .B(n7198), .Y(dpath_n59));
OR2X1 mul_U4576(.A(spu_mul_op1_data[37]), .B(n9772), .Y(dpath_n61));
OR2X1 mul_U4577(.A(spu_mul_op1_data[36]), .B(n9773), .Y(dpath_n63));
OR2X1 mul_U4578(.A(spu_mul_op1_data[35]), .B(n9772), .Y(dpath_n65));
OR2X1 mul_U4579(.A(spu_mul_op1_data[34]), .B(n9773), .Y(dpath_n67));
OR2X1 mul_U4580(.A(spu_mul_op1_data[33]), .B(n9772), .Y(dpath_n69));
OR2X1 mul_U4581(.A(spu_mul_op1_data[32]), .B(n9773), .Y(dpath_n71));
OR2X1 mul_U4582(.A(spu_mul_op1_data[31]), .B(n9772), .Y(dpath_n73));
OR2X1 mul_U4583(.A(spu_mul_op1_data[30]), .B(n9773), .Y(dpath_n75));
OR2X1 mul_U4584(.A(spu_mul_op1_data[29]), .B(n9772), .Y(dpath_n77));
OR2X1 mul_U4585(.A(spu_mul_op1_data[28]), .B(n9773), .Y(dpath_n79));
OR2X1 mul_U4586(.A(spu_mul_op1_data[27]), .B(n9774), .Y(dpath_n81));
OR2X1 mul_U4587(.A(spu_mul_op1_data[26]), .B(n9773), .Y(dpath_n83));
OR2X1 mul_U4588(.A(spu_mul_op1_data[25]), .B(n9772), .Y(dpath_n85));
OR2X1 mul_U4589(.A(spu_mul_op1_data[24]), .B(n9774), .Y(dpath_n87));
OR2X1 mul_U4590(.A(spu_mul_op1_data[23]), .B(n9772), .Y(dpath_n89));
OR2X1 mul_U4591(.A(spu_mul_op1_data[22]), .B(n9773), .Y(dpath_n91));
OR2X1 mul_U4592(.A(spu_mul_op1_data[21]), .B(n7198), .Y(dpath_n93));
OR2X1 mul_U4593(.A(spu_mul_op1_data[20]), .B(n9773), .Y(dpath_n95));
OR2X1 mul_U4594(.A(spu_mul_op1_data[19]), .B(n9774), .Y(dpath_n97));
OR2X1 mul_U4595(.A(spu_mul_op1_data[18]), .B(n9772), .Y(dpath_n99));
OR2X1 mul_U4596(.A(spu_mul_op1_data[17]), .B(n9773), .Y(dpath_n101));
INVX1 mul_U4597(.A(n9772), .Y(n9770));
OR2X1 mul_U4598(.A(spu_mul_op1_data[16]), .B(n7198), .Y(dpath_n103));
OR2X1 mul_U4599(.A(spu_mul_op1_data[15]), .B(n7198), .Y(dpath_n105));
OR2X1 mul_U4600(.A(spu_mul_op1_data[14]), .B(n9774), .Y(dpath_n107));
OR2X1 mul_U4601(.A(spu_mul_op1_data[13]), .B(n9772), .Y(dpath_n109));
INVX1 mul_U4602(.A(n9773), .Y(n9769));
OR2X1 mul_U4603(.A(spu_mul_op1_data[12]), .B(n9773), .Y(dpath_n111));
OR2X1 mul_U4604(.A(spu_mul_op1_data[11]), .B(n9774), .Y(dpath_n113));
OR2X1 mul_U4605(.A(spu_mul_op1_data[10]), .B(n9774), .Y(dpath_n115));
OR2X1 mul_U4606(.A(spu_mul_op1_data[9]), .B(n7198), .Y(dpath_n117));
OR2X1 mul_U4607(.A(spu_mul_op1_data[8]), .B(n9774), .Y(dpath_n119));
OR2X1 mul_U4608(.A(spu_mul_op1_data[7]), .B(n7198), .Y(dpath_n121));
OR2X1 mul_U4609(.A(spu_mul_op1_data[6]), .B(n9773), .Y(dpath_n123));
INVX1 mul_U4610(.A(n9571), .Y(n9543));
OR2X1 mul_U4611(.A(spu_mul_op1_data[5]), .B(n7198), .Y(dpath_n125));
OR2X1 mul_U4612(.A(spu_mul_op1_data[4]), .B(n9774), .Y(dpath_n127));
OR2X1 mul_U4613(.A(spu_mul_op1_data[3]), .B(n7198), .Y(dpath_n129));
OR2X1 mul_U4614(.A(spu_mul_op1_data[2]), .B(n9774), .Y(dpath_n131));
OR2X1 mul_U4615(.A(spu_mul_op1_data[1]), .B(n9772), .Y(dpath_n133));
OR2X1 mul_U4616(.A(spu_mul_op1_data[0]), .B(n9773), .Y(dpath_n135));
INVX1 mul_U4617(.A(n9571), .Y(n9542));
OR2X1 mul_U4618(.A(acc_reg_shf), .B(byp_imm), .Y(acc_reg_enb));
INVX1 mul_U4619(.A(n9574), .Y(n9532));
AND2X1 mul_U4620(.A(n3085), .B(n9816), .Y(control_n20));
INVX1 mul_U4621(.A(n9491), .Y(n9815));
AND2X1 mul_U4622(.A(n3084), .B(n4685), .Y(control_n13));
AND2X1 mul_U4623(.A(n3083), .B(spu_mul_areg_shf), .Y(control_n14));
INVX1 mul_U4624(.A(n9588), .Y(n9587));
INVX1 mul_U4625(.A(n9588), .Y(n9586));
INVX1 mul_U4626(.A(n9588), .Y(n9585));
INVX1 mul_U4627(.A(n9597), .Y(n9598));
INVX1 mul_U4628(.A(n9589), .Y(n9599));
INVX1 mul_U4629(.A(n9670), .Y(n9600));
INVX1 mul_U4630(.A(n9670), .Y(n9601));
INVX1 mul_U4631(.A(n9670), .Y(n9602));
INVX1 mul_U4632(.A(n9669), .Y(n9603));
AND2X1 mul_U4633(.A(dpath_mulcore_ary1_a1_s2[67]), .B(n7209), .Y(dpath_mulcore_a1cout[79]));
AND2X1 mul_U4634(.A(dpath_mulcore_ary1_a1_s2[66]), .B(n7208), .Y(dpath_mulcore_a1cout[78]));
INVX1 mul_U4635(.A(n9669), .Y(n9604));
INVX1 mul_U4636(.A(n9669), .Y(n9605));
INVX1 mul_U4637(.A(n9668), .Y(n9606));
INVX1 mul_U4638(.A(n9668), .Y(n9607));
INVX1 mul_U4639(.A(n9668), .Y(n9608));
INVX1 mul_U4640(.A(n9667), .Y(n9609));
AND2X1 mul_U4641(.A(n7413), .B(dpath_mulcore_ary1_a1_s_1[7]), .Y(dpath_mulcore_a1cout[7]));
AND2X1 mul_U4642(.A(n7414), .B(dpath_mulcore_ary1_a1_s_1[6]), .Y(dpath_mulcore_a1cout[6]));
AND2X1 mul_U4643(.A(n7415), .B(dpath_mulcore_ary1_a1_s_1[5]), .Y(dpath_mulcore_a1cout[5]));
AND2X1 mul_U4644(.A(n7412), .B(dpath_mulcore_ary1_a1_s_1[4]), .Y(dpath_mulcore_a1cout[4]));
AND2X1 mul_U4645(.A(spu_mul_mulres_lshft), .B(n9775), .Y(x2));
OR2X1 mul_U4646(.A(n5836), .B(n5964), .Y(dpath_mul_op2_d[63]));
OR2X1 mul_U4647(.A(n5837), .B(n5965), .Y(dpath_mul_op2_d[62]));
OR2X1 mul_U4648(.A(n5838), .B(n5966), .Y(dpath_mul_op2_d[61]));
OR2X1 mul_U4649(.A(n5839), .B(n5967), .Y(dpath_mul_op2_d[60]));
OR2X1 mul_U4650(.A(n5841), .B(n5969), .Y(dpath_mul_op2_d[59]));
OR2X1 mul_U4651(.A(n5842), .B(n5970), .Y(dpath_mul_op2_d[58]));
OR2X1 mul_U4652(.A(n5843), .B(n5971), .Y(dpath_mul_op2_d[57]));
OR2X1 mul_U4653(.A(n5844), .B(n5972), .Y(dpath_mul_op2_d[56]));
OR2X1 mul_U4654(.A(n5845), .B(n5973), .Y(dpath_mul_op2_d[55]));
OR2X1 mul_U4655(.A(n5846), .B(n5974), .Y(dpath_mul_op2_d[54]));
OR2X1 mul_U4656(.A(n5847), .B(n5975), .Y(dpath_mul_op2_d[53]));
OR2X1 mul_U4657(.A(n5848), .B(n5976), .Y(dpath_mul_op2_d[52]));
OR2X1 mul_U4658(.A(n5849), .B(n5977), .Y(dpath_mul_op2_d[51]));
OR2X1 mul_U4659(.A(n5850), .B(n5978), .Y(dpath_mul_op2_d[50]));
OR2X1 mul_U4660(.A(n5852), .B(n5980), .Y(dpath_mul_op2_d[49]));
OR2X1 mul_U4661(.A(n5853), .B(n5981), .Y(dpath_mul_op2_d[48]));
OR2X1 mul_U4662(.A(n5854), .B(n5982), .Y(dpath_mul_op2_d[47]));
OR2X1 mul_U4663(.A(n5855), .B(n5983), .Y(dpath_mul_op2_d[46]));
OR2X1 mul_U4664(.A(n5856), .B(n5984), .Y(dpath_mul_op2_d[45]));
OR2X1 mul_U4665(.A(n5857), .B(n5985), .Y(dpath_mul_op2_d[44]));
OR2X1 mul_U4666(.A(n5858), .B(n5986), .Y(dpath_mul_op2_d[43]));
OR2X1 mul_U4667(.A(n5859), .B(n5987), .Y(dpath_mul_op2_d[42]));
OR2X1 mul_U4668(.A(n5860), .B(n5988), .Y(dpath_mul_op2_d[41]));
OR2X1 mul_U4669(.A(n5861), .B(n5989), .Y(dpath_mul_op2_d[40]));
OR2X1 mul_U4670(.A(n5863), .B(n5991), .Y(dpath_mul_op2_d[39]));
OR2X1 mul_U4671(.A(n5864), .B(n5992), .Y(dpath_mul_op2_d[38]));
OR2X1 mul_U4672(.A(n5865), .B(n5993), .Y(dpath_mul_op2_d[37]));
OR2X1 mul_U4673(.A(n5866), .B(n5994), .Y(dpath_mul_op2_d[36]));
OR2X1 mul_U4674(.A(n5867), .B(n5995), .Y(dpath_mul_op2_d[35]));
OR2X1 mul_U4675(.A(n5868), .B(n5996), .Y(dpath_mul_op2_d[34]));
OR2X1 mul_U4676(.A(n5869), .B(n5997), .Y(dpath_mul_op2_d[33]));
OR2X1 mul_U4677(.A(n5870), .B(n5998), .Y(dpath_mul_op2_d[32]));
AND2X1 mul_U4678(.A(dpath_mulcore_psum[98]), .B(n9216), .Y(dpath_mulcore_add_cin));
INVX1 mul_U4679(.A(n9589), .Y(n9584));
INVX1 mul_U4680(.A(n9667), .Y(n9610));
INVX1 mul_U4681(.A(n9667), .Y(n9611));
INVX1 mul_U4682(.A(n9595), .Y(n9612));
AND2X1 mul_U4683(.A(n10602), .B(n3184), .Y(n10603));
INVX1 mul_U4684(.A(n9597), .Y(n9613));
INVX1 mul_U4685(.A(n9595), .Y(n9614));
INVX1 mul_U4686(.A(n9666), .Y(n9615));
INVX1 mul_U4687(.A(n9666), .Y(n9616));
INVX1 mul_U4688(.A(n9666), .Y(n9617));
INVX1 mul_U4689(.A(n9665), .Y(n9618));
INVX1 mul_U4690(.A(n9665), .Y(n9619));
INVX1 mul_U4691(.A(n9665), .Y(n9620));
AND2X1 mul_U4692(.A(n1886), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[97]));
AND2X1 mul_U4693(.A(n6072), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[96]));
AND2X1 mul_U4694(.A(n9188), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[95]));
AND2X1 mul_U4695(.A(n9189), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[94]));
AND2X1 mul_U4696(.A(n9190), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[93]));
AND2X1 mul_U4697(.A(n9191), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[92]));
AND2X1 mul_U4698(.A(n9192), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[91]));
AND2X1 mul_U4699(.A(n9193), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[90]));
INVX1 mul_U4700(.A(n9597), .Y(n9621));
AND2X1 mul_U4701(.A(n9194), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[89]));
AND2X1 mul_U4702(.A(n9195), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[88]));
AND2X1 mul_U4703(.A(n9196), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[87]));
AND2X1 mul_U4704(.A(n9197), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[86]));
AND2X1 mul_U4705(.A(n9198), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[85]));
AND2X1 mul_U4706(.A(n9199), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[84]));
AND2X1 mul_U4707(.A(n9213), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[83]));
AND2X1 mul_U4708(.A(n9148), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[82]));
AND2X1 mul_U4709(.A(n9200), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[81]));
AND2X1 mul_U4710(.A(n9201), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[80]));
AND2X1 mul_U4711(.A(n9202), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[79]));
AND2X1 mul_U4712(.A(n9203), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[78]));
AND2X1 mul_U4713(.A(n9204), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[77]));
INVX1 mul_U4714(.A(n9589), .Y(n9622));
AND2X1 mul_U4715(.A(n9205), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[76]));
AND2X1 mul_U4716(.A(n9206), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[75]));
AND2X1 mul_U4717(.A(n9207), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[74]));
AND2X1 mul_U4718(.A(n9208), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[73]));
AND2X1 mul_U4719(.A(n9209), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[72]));
AND2X1 mul_U4720(.A(n9210), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[71]));
AND2X1 mul_U4721(.A(n9211), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[70]));
AND2X1 mul_U4722(.A(n9212), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[69]));
AND2X1 mul_U4723(.A(n9149), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[68]));
AND2X1 mul_U4724(.A(n9150), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[67]));
AND2X1 mul_U4725(.A(n9151), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[66]));
AND2X1 mul_U4726(.A(n9152), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[65]));
AND2X1 mul_U4727(.A(n9153), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[64]));
INVX1 mul_U4728(.A(n9659), .Y(n9623));
AND2X1 mul_U4729(.A(n9154), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[63]));
AND2X1 mul_U4730(.A(n9155), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[62]));
AND2X1 mul_U4731(.A(n9156), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[61]));
AND2X1 mul_U4732(.A(n9157), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[60]));
AND2X1 mul_U4733(.A(n9158), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[59]));
AND2X1 mul_U4734(.A(n9159), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[58]));
AND2X1 mul_U4735(.A(n9160), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[57]));
AND2X1 mul_U4736(.A(n9161), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[56]));
AND2X1 mul_U4737(.A(n9162), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[55]));
AND2X1 mul_U4738(.A(n9163), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[54]));
AND2X1 mul_U4739(.A(n9164), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[53]));
AND2X1 mul_U4740(.A(n9165), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[52]));
AND2X1 mul_U4741(.A(n9166), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[51]));
INVX1 mul_U4742(.A(n9664), .Y(n9624));
AND2X1 mul_U4743(.A(n9167), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[50]));
AND2X1 mul_U4744(.A(n9168), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[49]));
AND2X1 mul_U4745(.A(n9169), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[48]));
AND2X1 mul_U4746(.A(n9170), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[47]));
AND2X1 mul_U4747(.A(n9171), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[46]));
AND2X1 mul_U4748(.A(n9172), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[45]));
AND2X1 mul_U4749(.A(n9173), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[44]));
AND2X1 mul_U4750(.A(n9174), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[43]));
AND2X1 mul_U4751(.A(n9175), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[42]));
AND2X1 mul_U4752(.A(n9176), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[41]));
AND2X1 mul_U4753(.A(n9177), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[40]));
AND2X1 mul_U4754(.A(n9178), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[39]));
AND2X1 mul_U4755(.A(n9179), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[38]));
INVX1 mul_U4756(.A(n9664), .Y(n9625));
AND2X1 mul_U4757(.A(n9180), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[37]));
AND2X1 mul_U4758(.A(n9181), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[36]));
AND2X1 mul_U4759(.A(n9182), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[35]));
AND2X1 mul_U4760(.A(n9183), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[34]));
AND2X1 mul_U4761(.A(n9184), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[33]));
AND2X1 mul_U4762(.A(n9185), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[32]));
AND2X1 mul_U4763(.A(n9186), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_pcout_in[31]));
AND2X1 mul_U4764(.A(n9187), .B(dpath_mulcore_x2_c2), .Y(dpath_mulcore_pcout_in[30]));
AND2X1 mul_U4765(.A(dpath_mulcore_psum[98]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[98]));
AND2X1 mul_U4766(.A(dpath_mulcore_psum[97]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[97]));
AND2X1 mul_U4767(.A(dpath_mulcore_psum[96]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[96]));
AND2X1 mul_U4768(.A(dpath_mulcore_psum[95]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[95]));
AND2X1 mul_U4769(.A(dpath_mulcore_psum[94]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[94]));
INVX1 mul_U4770(.A(n9664), .Y(n9626));
AND2X1 mul_U4771(.A(dpath_mulcore_psum[93]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[93]));
AND2X1 mul_U4772(.A(dpath_mulcore_psum[92]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[92]));
AND2X1 mul_U4773(.A(dpath_mulcore_psum[91]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[91]));
AND2X1 mul_U4774(.A(dpath_mulcore_psum[90]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[90]));
AND2X1 mul_U4775(.A(dpath_mulcore_psum[89]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[89]));
AND2X1 mul_U4776(.A(dpath_mulcore_psum[88]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[88]));
AND2X1 mul_U4777(.A(dpath_mulcore_psum[87]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[87]));
AND2X1 mul_U4778(.A(dpath_mulcore_psum[86]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[86]));
AND2X1 mul_U4779(.A(dpath_mulcore_psum[85]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[85]));
AND2X1 mul_U4780(.A(dpath_mulcore_psum[84]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[84]));
AND2X1 mul_U4781(.A(dpath_mulcore_psum[83]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[83]));
AND2X1 mul_U4782(.A(dpath_mulcore_psum[82]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[82]));
AND2X1 mul_U4783(.A(dpath_mulcore_psum[81]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[81]));
INVX1 mul_U4784(.A(n9663), .Y(n9627));
AND2X1 mul_U4785(.A(dpath_mulcore_psum[80]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[80]));
AND2X1 mul_U4786(.A(dpath_mulcore_psum[79]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[79]));
AND2X1 mul_U4787(.A(dpath_mulcore_psum[78]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[78]));
AND2X1 mul_U4788(.A(dpath_mulcore_psum[77]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[77]));
AND2X1 mul_U4789(.A(dpath_mulcore_psum[76]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[76]));
AND2X1 mul_U4790(.A(dpath_mulcore_psum[75]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[75]));
AND2X1 mul_U4791(.A(dpath_mulcore_psum[74]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[74]));
AND2X1 mul_U4792(.A(dpath_mulcore_psum[73]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[73]));
AND2X1 mul_U4793(.A(dpath_mulcore_psum[72]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[72]));
AND2X1 mul_U4794(.A(dpath_mulcore_psum[71]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[71]));
AND2X1 mul_U4795(.A(dpath_mulcore_psum[70]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[70]));
AND2X1 mul_U4796(.A(dpath_mulcore_psum[69]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[69]));
AND2X1 mul_U4797(.A(dpath_mulcore_psum[68]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[68]));
INVX1 mul_U4798(.A(n9663), .Y(n9628));
AND2X1 mul_U4799(.A(dpath_mulcore_psum[67]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[67]));
AND2X1 mul_U4800(.A(dpath_mulcore_psum[66]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[66]));
AND2X1 mul_U4801(.A(dpath_mulcore_psum[65]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[65]));
AND2X1 mul_U4802(.A(dpath_mulcore_psum[64]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[64]));
AND2X1 mul_U4803(.A(dpath_mulcore_psum[63]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[63]));
AND2X1 mul_U4804(.A(dpath_mulcore_psum[62]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[62]));
AND2X1 mul_U4805(.A(dpath_mulcore_psum[61]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[61]));
AND2X1 mul_U4806(.A(dpath_mulcore_psum[60]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[60]));
AND2X1 mul_U4807(.A(dpath_mulcore_psum[59]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[59]));
AND2X1 mul_U4808(.A(dpath_mulcore_psum[58]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[58]));
AND2X1 mul_U4809(.A(dpath_mulcore_psum[57]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[57]));
AND2X1 mul_U4810(.A(dpath_mulcore_psum[56]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[56]));
AND2X1 mul_U4811(.A(dpath_mulcore_psum[55]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[55]));
INVX1 mul_U4812(.A(n9663), .Y(n9629));
AND2X1 mul_U4813(.A(dpath_mulcore_psum[54]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[54]));
AND2X1 mul_U4814(.A(dpath_mulcore_psum[53]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[53]));
AND2X1 mul_U4815(.A(dpath_mulcore_psum[52]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[52]));
AND2X1 mul_U4816(.A(dpath_mulcore_psum[51]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[51]));
AND2X1 mul_U4817(.A(dpath_mulcore_psum[50]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[50]));
AND2X1 mul_U4818(.A(dpath_mulcore_psum[49]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[49]));
AND2X1 mul_U4819(.A(dpath_mulcore_psum[48]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[48]));
AND2X1 mul_U4820(.A(dpath_mulcore_psum[47]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[47]));
AND2X1 mul_U4821(.A(dpath_mulcore_psum[46]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[46]));
AND2X1 mul_U4822(.A(dpath_mulcore_psum[45]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[45]));
AND2X1 mul_U4823(.A(dpath_mulcore_psum[44]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[44]));
AND2X1 mul_U4824(.A(dpath_mulcore_psum[43]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[43]));
AND2X1 mul_U4825(.A(dpath_mulcore_psum[42]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[42]));
INVX1 mul_U4826(.A(n9596), .Y(n9630));
AND2X1 mul_U4827(.A(dpath_mulcore_psum[41]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[41]));
AND2X1 mul_U4828(.A(dpath_mulcore_psum[40]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[40]));
AND2X1 mul_U4829(.A(dpath_mulcore_psum[39]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[39]));
AND2X1 mul_U4830(.A(dpath_mulcore_psum[38]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[38]));
AND2X1 mul_U4831(.A(dpath_mulcore_psum[37]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[37]));
AND2X1 mul_U4832(.A(dpath_mulcore_psum[36]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[36]));
AND2X1 mul_U4833(.A(dpath_mulcore_psum[35]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[35]));
AND2X1 mul_U4834(.A(dpath_mulcore_psum[34]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[34]));
AND2X1 mul_U4835(.A(dpath_mulcore_psum[33]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[33]));
AND2X1 mul_U4836(.A(dpath_mulcore_psum[32]), .B(dpath_mulcore_cyc2), .Y(dpath_mulcore_psum_in[32]));
AND2X1 mul_U4837(.A(dpath_mulcore_x2_c2), .B(dpath_mulcore_psum[31]), .Y(dpath_mulcore_psum_in[31]));
INVX1 mul_U4838(.A(n9666), .Y(n9631));
INVX1 mul_U4839(.A(n9665), .Y(n9632));
INVX1 mul_U4840(.A(n9662), .Y(n9633));
INVX1 mul_U4841(.A(n9662), .Y(n9634));
INVX1 mul_U4842(.A(n9662), .Y(n9635));
INVX1 mul_U4843(.A(n9661), .Y(n9636));
INVX1 mul_U4844(.A(n9661), .Y(n9637));
INVX1 mul_U4845(.A(n9661), .Y(n9638));
INVX1 mul_U4846(.A(n9597), .Y(n9639));
INVX1 mul_U4847(.A(n9668), .Y(n9640));
INVX1 mul_U4848(.A(n9667), .Y(n9641));
INVX1 mul_U4849(.A(n9595), .Y(n9642));
INVX1 mul_U4850(.A(n9664), .Y(n9643));
INVX1 mul_U4851(.A(n9663), .Y(n9644));
INVX1 mul_U4852(.A(n9596), .Y(n9645));
INVX1 mul_U4853(.A(n9568), .Y(n9550));
INVX1 mul_U4854(.A(n9670), .Y(n9646));
INVX1 mul_U4855(.A(n9669), .Y(n9647));
INVX1 mul_U4856(.A(n9595), .Y(n9648));
INVX1 mul_U4857(.A(n9596), .Y(n9649));
INVX1 mul_U4858(.A(n9589), .Y(n9650));
INVX1 mul_U4859(.A(n9660), .Y(n9651));
INVX1 mul_U4860(.A(n9588), .Y(n9652));
AND2X1 mul_U4861(.A(n9312), .B(n9474), .Y(dpath_mulcore_a0cout[79]));
AND2X1 mul_U4862(.A(dpath_mulcore_ary1_a0_I2_I2_net38), .B(n16569), .Y(dpath_mulcore_a0cout[78]));
INVX1 mul_U4863(.A(n9659), .Y(n9653));
INVX1 mul_U4864(.A(n9660), .Y(n9654));
INVX1 mul_U4865(.A(n9660), .Y(n9655));
INVX1 mul_U4866(.A(n9660), .Y(n9656));
INVX1 mul_U4867(.A(n9659), .Y(n9657));
AND2X1 mul_U4868(.A(n7409), .B(dpath_mulcore_ary1_a0_s_1[7]), .Y(dpath_mulcore_a0cout[7]));
AND2X1 mul_U4869(.A(n7410), .B(dpath_mulcore_ary1_a0_s_1[6]), .Y(dpath_mulcore_a0cout[6]));
INVX1 mul_U4870(.A(n9659), .Y(n9658));
AND2X1 mul_U4871(.A(n7411), .B(dpath_mulcore_ary1_a0_s_1[5]), .Y(dpath_mulcore_a0cout[5]));
AND2X1 mul_U4872(.A(n7408), .B(dpath_mulcore_ary1_a0_s_1[4]), .Y(dpath_mulcore_a0cout[4]));
OR2X1 mul_U4873(.A(control_n7), .B(exu_mul_rs1_data[63]), .Y(dpath_n10));
OR2X1 mul_U4874(.A(control_n7), .B(exu_mul_rs1_data[62]), .Y(dpath_n12));
OR2X1 mul_U4875(.A(control_n7), .B(exu_mul_rs1_data[61]), .Y(dpath_n14));
OR2X1 mul_U4876(.A(control_n7), .B(exu_mul_rs1_data[60]), .Y(dpath_n16));
OR2X1 mul_U4877(.A(n9775), .B(exu_mul_rs1_data[59]), .Y(dpath_n18));
OR2X1 mul_U4878(.A(control_n7), .B(exu_mul_rs1_data[58]), .Y(dpath_n20));
OR2X1 mul_U4879(.A(n9775), .B(exu_mul_rs1_data[57]), .Y(dpath_n22));
OR2X1 mul_U4880(.A(control_n7), .B(exu_mul_rs1_data[56]), .Y(dpath_n24));
OR2X1 mul_U4881(.A(n9775), .B(exu_mul_rs1_data[55]), .Y(dpath_n26));
OR2X1 mul_U4882(.A(control_n7), .B(exu_mul_rs1_data[54]), .Y(dpath_n28));
OR2X1 mul_U4883(.A(n9771), .B(exu_mul_rs1_data[53]), .Y(dpath_n30));
OR2X1 mul_U4884(.A(n9771), .B(exu_mul_rs1_data[52]), .Y(dpath_n32));
OR2X1 mul_U4885(.A(n9771), .B(exu_mul_rs1_data[51]), .Y(dpath_n34));
OR2X1 mul_U4886(.A(n9771), .B(exu_mul_rs1_data[50]), .Y(dpath_n36));
OR2X1 mul_U4887(.A(n9771), .B(exu_mul_rs1_data[49]), .Y(dpath_n38));
OR2X1 mul_U4888(.A(n9771), .B(exu_mul_rs1_data[48]), .Y(dpath_n40));
OR2X1 mul_U4889(.A(n9771), .B(exu_mul_rs1_data[47]), .Y(dpath_n42));
OR2X1 mul_U4890(.A(n9771), .B(exu_mul_rs1_data[46]), .Y(dpath_n44));
OR2X1 mul_U4891(.A(n9771), .B(exu_mul_rs1_data[45]), .Y(dpath_n46));
OR2X1 mul_U4892(.A(n9771), .B(exu_mul_rs1_data[44]), .Y(dpath_n48));
OR2X1 mul_U4893(.A(n9771), .B(exu_mul_rs1_data[43]), .Y(dpath_n50));
OR2X1 mul_U4894(.A(n9771), .B(exu_mul_rs1_data[42]), .Y(dpath_n52));
OR2X1 mul_U4895(.A(n9771), .B(exu_mul_rs1_data[41]), .Y(dpath_n54));
OR2X1 mul_U4896(.A(n9771), .B(exu_mul_rs1_data[40]), .Y(dpath_n56));
OR2X1 mul_U4897(.A(n9770), .B(exu_mul_rs1_data[39]), .Y(dpath_n58));
OR2X1 mul_U4898(.A(n9770), .B(exu_mul_rs1_data[38]), .Y(dpath_n60));
OR2X1 mul_U4899(.A(n9770), .B(exu_mul_rs1_data[37]), .Y(dpath_n62));
OR2X1 mul_U4900(.A(n9770), .B(exu_mul_rs1_data[36]), .Y(dpath_n64));
OR2X1 mul_U4901(.A(n9770), .B(exu_mul_rs1_data[35]), .Y(dpath_n66));
OR2X1 mul_U4902(.A(n9770), .B(exu_mul_rs1_data[34]), .Y(dpath_n68));
OR2X1 mul_U4903(.A(n9770), .B(exu_mul_rs1_data[33]), .Y(dpath_n70));
OR2X1 mul_U4904(.A(n9770), .B(exu_mul_rs1_data[32]), .Y(dpath_n72));
OR2X1 mul_U4905(.A(n9770), .B(exu_mul_rs1_data[31]), .Y(dpath_n74));
OR2X1 mul_U4906(.A(n9770), .B(exu_mul_rs1_data[30]), .Y(dpath_n76));
OR2X1 mul_U4907(.A(n9770), .B(exu_mul_rs1_data[29]), .Y(dpath_n78));
OR2X1 mul_U4908(.A(n9770), .B(exu_mul_rs1_data[28]), .Y(dpath_n80));
OR2X1 mul_U4909(.A(n9770), .B(exu_mul_rs1_data[27]), .Y(dpath_n82));
OR2X1 mul_U4910(.A(n9769), .B(exu_mul_rs1_data[26]), .Y(dpath_n84));
OR2X1 mul_U4911(.A(n9769), .B(exu_mul_rs1_data[25]), .Y(dpath_n86));
OR2X1 mul_U4912(.A(n9769), .B(exu_mul_rs1_data[24]), .Y(dpath_n88));
OR2X1 mul_U4913(.A(n9769), .B(exu_mul_rs1_data[23]), .Y(dpath_n90));
OR2X1 mul_U4914(.A(n9769), .B(exu_mul_rs1_data[22]), .Y(dpath_n92));
OR2X1 mul_U4915(.A(n9769), .B(exu_mul_rs1_data[21]), .Y(dpath_n94));
OR2X1 mul_U4916(.A(n9769), .B(exu_mul_rs1_data[20]), .Y(dpath_n96));
OR2X1 mul_U4917(.A(n9769), .B(exu_mul_rs1_data[19]), .Y(dpath_n98));
OR2X1 mul_U4918(.A(n9769), .B(exu_mul_rs1_data[18]), .Y(dpath_n100));
OR2X1 mul_U4919(.A(n9769), .B(exu_mul_rs1_data[17]), .Y(dpath_n102));
OR2X1 mul_U4920(.A(n9770), .B(exu_mul_rs1_data[16]), .Y(dpath_n104));
OR2X1 mul_U4921(.A(n9769), .B(exu_mul_rs1_data[15]), .Y(dpath_n106));
OR2X1 mul_U4922(.A(n9769), .B(exu_mul_rs1_data[14]), .Y(dpath_n108));
OR2X1 mul_U4923(.A(n9769), .B(exu_mul_rs1_data[13]), .Y(dpath_n110));
OR2X1 mul_U4924(.A(n9769), .B(exu_mul_rs1_data[12]), .Y(dpath_n112));
OR2X1 mul_U4925(.A(n9775), .B(exu_mul_rs1_data[11]), .Y(dpath_n114));
OR2X1 mul_U4926(.A(control_n7), .B(exu_mul_rs1_data[10]), .Y(dpath_n116));
OR2X1 mul_U4927(.A(n9775), .B(exu_mul_rs1_data[9]), .Y(dpath_n118));
OR2X1 mul_U4928(.A(control_n7), .B(exu_mul_rs1_data[8]), .Y(dpath_n120));
OR2X1 mul_U4929(.A(n9775), .B(exu_mul_rs1_data[7]), .Y(dpath_n122));
OR2X1 mul_U4930(.A(control_n7), .B(exu_mul_rs1_data[6]), .Y(dpath_n124));
OR2X1 mul_U4931(.A(n9775), .B(exu_mul_rs1_data[5]), .Y(dpath_n126));
OR2X1 mul_U4932(.A(control_n7), .B(exu_mul_rs1_data[4]), .Y(dpath_n128));
OR2X1 mul_U4933(.A(n9775), .B(exu_mul_rs1_data[3]), .Y(dpath_n130));
OR2X1 mul_U4934(.A(n9775), .B(exu_mul_rs1_data[2]), .Y(dpath_n132));
OR2X1 mul_U4935(.A(n9775), .B(exu_mul_rs1_data[1]), .Y(dpath_n134));
OR2X1 mul_U4936(.A(n9775), .B(exu_mul_rs1_data[0]), .Y(dpath_n136));
INVX1 mul_U4937(.A(dpath_mulcore_clk_enb0), .Y(n9785));
AND2X1 mul_U4938(.A(dpath_mout[135]), .B(n9778), .Y(dpath_acc_reg_in[135]));
AND2X1 mul_U4939(.A(dpath_mout[134]), .B(n9783), .Y(dpath_acc_reg_in[134]));
AND2X1 mul_U4940(.A(dpath_mout[133]), .B(n9781), .Y(dpath_acc_reg_in[133]));
AND2X1 mul_U4941(.A(dpath_mout[132]), .B(n9779), .Y(dpath_acc_reg_in[132]));
AND2X1 mul_U4942(.A(dpath_mout[131]), .B(n9783), .Y(dpath_acc_reg_in[131]));
AND2X1 mul_U4943(.A(dpath_mout[130]), .B(n9781), .Y(dpath_acc_reg_in[130]));
AND2X1 mul_U4944(.A(dpath_mout[129]), .B(n9781), .Y(dpath_acc_reg_in[129]));
AND2X1 mul_U4945(.A(n9782), .B(dpath_mout[128]), .Y(dpath_acc_reg_in[128]));
AND2X1 mul_U4946(.A(n9782), .B(dpath_mout[127]), .Y(dpath_acc_reg_in[127]));
AND2X1 mul_U4947(.A(n9782), .B(dpath_mout[126]), .Y(dpath_acc_reg_in[126]));
AND2X1 mul_U4948(.A(n9782), .B(dpath_mout[125]), .Y(dpath_acc_reg_in[125]));
AND2X1 mul_U4949(.A(n9782), .B(dpath_mout[124]), .Y(dpath_acc_reg_in[124]));
AND2X1 mul_U4950(.A(n9782), .B(dpath_mout[123]), .Y(dpath_acc_reg_in[123]));
AND2X1 mul_U4951(.A(n9782), .B(dpath_mout[122]), .Y(dpath_acc_reg_in[122]));
AND2X1 mul_U4952(.A(n9782), .B(dpath_mout[121]), .Y(dpath_acc_reg_in[121]));
AND2X1 mul_U4953(.A(n9782), .B(dpath_mout[120]), .Y(dpath_acc_reg_in[120]));
AND2X1 mul_U4954(.A(n9782), .B(dpath_mout[119]), .Y(dpath_acc_reg_in[119]));
AND2X1 mul_U4955(.A(n9782), .B(dpath_mout[118]), .Y(dpath_acc_reg_in[118]));
AND2X1 mul_U4956(.A(n9782), .B(dpath_mout[117]), .Y(dpath_acc_reg_in[117]));
AND2X1 mul_U4957(.A(n9782), .B(dpath_mout[116]), .Y(dpath_acc_reg_in[116]));
AND2X1 mul_U4958(.A(n9783), .B(dpath_mout[115]), .Y(dpath_acc_reg_in[115]));
AND2X1 mul_U4959(.A(n9783), .B(dpath_mout[114]), .Y(dpath_acc_reg_in[114]));
AND2X1 mul_U4960(.A(n9783), .B(dpath_mout[113]), .Y(dpath_acc_reg_in[113]));
AND2X1 mul_U4961(.A(n9783), .B(dpath_mout[112]), .Y(dpath_acc_reg_in[112]));
AND2X1 mul_U4962(.A(n9783), .B(dpath_mout[111]), .Y(dpath_acc_reg_in[111]));
AND2X1 mul_U4963(.A(n9783), .B(dpath_mout[110]), .Y(dpath_acc_reg_in[110]));
AND2X1 mul_U4964(.A(n9783), .B(dpath_mout[109]), .Y(dpath_acc_reg_in[109]));
AND2X1 mul_U4965(.A(n9783), .B(dpath_mout[108]), .Y(dpath_acc_reg_in[108]));
AND2X1 mul_U4966(.A(n9783), .B(dpath_mout[107]), .Y(dpath_acc_reg_in[107]));
AND2X1 mul_U4967(.A(n9783), .B(dpath_mout[106]), .Y(dpath_acc_reg_in[106]));
AND2X1 mul_U4968(.A(n9783), .B(dpath_mout[105]), .Y(dpath_acc_reg_in[105]));
AND2X1 mul_U4969(.A(n9783), .B(dpath_mout[104]), .Y(dpath_acc_reg_in[104]));
AND2X1 mul_U4970(.A(n9783), .B(dpath_mout[103]), .Y(dpath_acc_reg_in[103]));
AND2X1 mul_U4971(.A(n9783), .B(dpath_mout[102]), .Y(dpath_acc_reg_in[102]));
AND2X1 mul_U4972(.A(n9783), .B(dpath_mout[101]), .Y(dpath_acc_reg_in[101]));
AND2X1 mul_U4973(.A(n9782), .B(dpath_mout[100]), .Y(dpath_acc_reg_in[100]));
AND2X1 mul_U4974(.A(n9781), .B(dpath_mout[99]), .Y(dpath_acc_reg_in[99]));
AND2X1 mul_U4975(.A(n9781), .B(dpath_mout[98]), .Y(dpath_acc_reg_in[98]));
AND2X1 mul_U4976(.A(n9781), .B(dpath_mout[97]), .Y(dpath_acc_reg_in[97]));
AND2X1 mul_U4977(.A(n9782), .B(dpath_mout[96]), .Y(dpath_acc_reg_in[96]));
AND2X1 mul_U4978(.A(n9781), .B(dpath_mout[95]), .Y(dpath_acc_reg_in[95]));
AND2X1 mul_U4979(.A(n9781), .B(dpath_mout[94]), .Y(dpath_acc_reg_in[94]));
AND2X1 mul_U4980(.A(n9781), .B(dpath_mout[93]), .Y(dpath_acc_reg_in[93]));
AND2X1 mul_U4981(.A(n9781), .B(dpath_mout[92]), .Y(dpath_acc_reg_in[92]));
AND2X1 mul_U4982(.A(n9782), .B(dpath_mout[91]), .Y(dpath_acc_reg_in[91]));
AND2X1 mul_U4983(.A(n9781), .B(dpath_mout[90]), .Y(dpath_acc_reg_in[90]));
AND2X1 mul_U4984(.A(n9781), .B(dpath_mout[89]), .Y(dpath_acc_reg_in[89]));
AND2X1 mul_U4985(.A(n9781), .B(dpath_mout[88]), .Y(dpath_acc_reg_in[88]));
AND2X1 mul_U4986(.A(n9781), .B(dpath_mout[87]), .Y(dpath_acc_reg_in[87]));
AND2X1 mul_U4987(.A(n9778), .B(dpath_mout[86]), .Y(dpath_acc_reg_in[86]));
AND2X1 mul_U4988(.A(n9781), .B(dpath_mout[85]), .Y(dpath_acc_reg_in[85]));
AND2X1 mul_U4989(.A(n9781), .B(dpath_mout[84]), .Y(dpath_acc_reg_in[84]));
AND2X1 mul_U4990(.A(n9781), .B(dpath_mout[83]), .Y(dpath_acc_reg_in[83]));
AND2X1 mul_U4991(.A(n9783), .B(dpath_mout[82]), .Y(dpath_acc_reg_in[82]));
AND2X1 mul_U4992(.A(n9778), .B(dpath_mout[81]), .Y(dpath_acc_reg_in[81]));
AND2X1 mul_U4993(.A(n9779), .B(dpath_mout[80]), .Y(dpath_acc_reg_in[80]));
AND2X1 mul_U4994(.A(n9782), .B(dpath_mout[79]), .Y(dpath_acc_reg_in[79]));
AND2X1 mul_U4995(.A(n9782), .B(dpath_mout[78]), .Y(dpath_acc_reg_in[78]));
AND2X1 mul_U4996(.A(n9780), .B(dpath_mout[77]), .Y(dpath_acc_reg_in[77]));
AND2X1 mul_U4997(.A(n9781), .B(dpath_mout[76]), .Y(dpath_acc_reg_in[76]));
AND2X1 mul_U4998(.A(n9781), .B(dpath_mout[75]), .Y(dpath_acc_reg_in[75]));
AND2X1 mul_U4999(.A(n9778), .B(dpath_mout[74]), .Y(dpath_acc_reg_in[74]));
AND2X1 mul_U5000(.A(n9783), .B(dpath_mout[73]), .Y(dpath_acc_reg_in[73]));
AND2X1 mul_U5001(.A(n9778), .B(dpath_mout[72]), .Y(dpath_acc_reg_in[72]));
AND2X1 mul_U5002(.A(control_acc_actc1), .B(n9491), .Y(control_N7));
AND2X1 mul_U5003(.A(acc_actc2), .B(n9491), .Y(control_N8));
AND2X1 mul_U5004(.A(acc_actc3), .B(n9491), .Y(control_N9));
AND2X1 mul_U5005(.A(n3082), .B(control_mul_spu_ack_d), .Y(control_N5));
AND2X1 mul_U5006(.A(n9784), .B(n9491), .Y(control_N2));
AND2X1 mul_U5007(.A(control_c1_act), .B(n9491), .Y(control_N3));
AND2X1 mul_U5008(.A(control_c2_act), .B(n9491), .Y(control_N4));
AND2X1 mul_U5009(.A(spu_mul_acc), .B(mul_spu_ack), .Y(control_N6));
AND2X1 mul_U5010(.A(control_acc_actc4), .B(n9491), .Y(control_N11));
INVX1 mul_U5011(.A(n9594), .Y(n9664));
INVX1 mul_U5012(.A(n9594), .Y(n9663));
INVX1 mul_U5013(.A(n9594), .Y(n9670));
INVX1 mul_U5014(.A(n9594), .Y(n9669));
INVX1 mul_U5015(.A(n9778), .Y(n9777));
INVX1 mul_U5016(.A(n9596), .Y(n9594));
INVX1 mul_U5017(.A(dpath_mulcore_clk_enb0), .Y(n9666));
INVX1 mul_U5018(.A(dpath_mulcore_clk_enb0), .Y(n9665));
INVX1 mul_U5019(.A(dpath_mulcore_b7[0]), .Y(n9736));
INVX1 mul_U5020(.A(dpath_mulcore_b6[0]), .Y(n9734));
INVX1 mul_U5021(.A(dpath_mulcore_b5[0]), .Y(n9732));
INVX1 mul_U5022(.A(dpath_mulcore_b4[0]), .Y(n9730));
INVX1 mul_U5023(.A(dpath_mulcore_b0[0]), .Y(n9722));
INVX1 mul_U5024(.A(dpath_mulcore_b15[0]), .Y(n9752));
INVX1 mul_U5025(.A(dpath_mulcore_b14[0]), .Y(n9750));
INVX1 mul_U5026(.A(dpath_mulcore_b13[0]), .Y(n9748));
INVX1 mul_U5027(.A(dpath_mulcore_b12[0]), .Y(n9746));
INVX1 mul_U5028(.A(dpath_mulcore_b11[0]), .Y(n9744));
INVX1 mul_U5029(.A(dpath_mulcore_b10[0]), .Y(n9742));
INVX1 mul_U5030(.A(dpath_mulcore_b9[0]), .Y(n9740));
INVX1 mul_U5031(.A(dpath_mulcore_b8[0]), .Y(n9738));
INVX1 mul_U5032(.A(dpath_mulcore_b3[0]), .Y(n9728));
INVX1 mul_U5033(.A(dpath_mulcore_b2[0]), .Y(n9726));
INVX1 mul_U5034(.A(dpath_mulcore_b1[0]), .Y(n9724));
INVX1 mul_U5035(.A(n9576), .Y(n9498));
INVX1 mul_U5036(.A(n9497), .Y(n9500));
INVX1 mul_U5037(.A(n9671), .Y(n9697));
INVX1 mul_U5038(.A(se), .Y(n9497));
INVX1 mul_U5039(.A(n9497), .Y(n9501));
INVX1 mul_U5040(.A(n9754), .Y(n9755));
INVX1 mul_U5041(.A(n9596), .Y(n9593));
INVX1 mul_U5042(.A(dpath_mulcore_clk_enb0), .Y(n9668));
INVX1 mul_U5043(.A(dpath_mulcore_clk_enb0), .Y(n9667));
INVX1 mul_U5044(.A(n9681), .Y(n9675));
INVX1 mul_U5045(.A(dpath_mulcore_x2_c2c3), .Y(n9681));
INVX1 mul_U5046(.A(n9576), .Y(n9528));
INVX1 mul_U5047(.A(n9680), .Y(n9678));
INVX1 mul_U5048(.A(dpath_mulcore_x2_c2c3), .Y(n9680));
INVX1 mul_U5049(.A(n9496), .Y(n9576));
INVX1 mul_U5050(.A(n9500), .Y(n9496));
INVX1 mul_U5051(.A(se), .Y(n9512));
INVX1 mul_U5052(.A(se), .Y(n9513));
INVX1 mul_U5053(.A(n9754), .Y(n9757));
INVX1 mul_U5054(.A(n9754), .Y(n9759));
INVX1 mul_U5055(.A(dpath_mulcore_clk_enb0), .Y(n9660));
INVX1 mul_U5056(.A(dpath_mulcore_clk_enb0), .Y(n9588));
INVX1 mul_U5057(.A(n9680), .Y(n9679));
INVX1 mul_U5058(.A(n9671), .Y(n9698));
INVX1 mul_U5059(.A(n9496), .Y(n9577));
INVX1 mul_U5060(.A(n9581), .Y(n9509));
INVX1 mul_U5061(.A(n9501), .Y(n9517));
INVX1 mul_U5062(.A(n9501), .Y(n9518));
INVX1 mul_U5063(.A(dpath_n145), .Y(n9763));
INVX1 mul_U5064(.A(n9754), .Y(n9756));
INVX1 mul_U5065(.A(n9754), .Y(n9758));
INVX1 mul_U5066(.A(c0_act), .Y(n9784));
INVX1 mul_U5067(.A(dpath_acc_reg_shf2), .Y(n9753));
INVX1 mul_U5068(.A(dpath_mulcore_clk_enb0), .Y(n9596));
INVX1 mul_U5069(.A(n9495), .Y(n9573));
INVX1 mul_U5070(.A(n9500), .Y(n9495));
INVX1 mul_U5071(.A(n9565), .Y(n9559));
INVX1 mul_U5072(.A(n9565), .Y(n9560));
INVX1 mul_U5073(.A(n9672), .Y(n9699));
INVX1 mul_U5074(.A(n9682), .Y(n9672));
INVX1 mul_U5075(.A(n9698), .Y(n9691));
INVX1 mul_U5076(.A(n9698), .Y(n9692));
INVX1 mul_U5077(.A(dpath_n665), .Y(n9766));
INVX1 mul_U5078(.A(dpath_mulcore_clk_enb0), .Y(n9595));
INVX1 mul_U5079(.A(n9495), .Y(n9574));
INVX1 mul_U5080(.A(n9568), .Y(n9551));
INVX1 mul_U5081(.A(n9568), .Y(n9552));
INVX1 mul_U5082(.A(n9672), .Y(n9700));
INVX1 mul_U5083(.A(n9681), .Y(n9676));
INVX1 mul_U5084(.A(n9680), .Y(n9677));
INVX1 mul_U5085(.A(acc_reg_shf), .Y(n9778));
INVX1 mul_U5086(.A(dpath_mulcore_b0[2]), .Y(n9721));
INVX1 mul_U5087(.A(dpath_mulcore_b14[2]), .Y(n9749));
INVX1 mul_U5088(.A(dpath_mulcore_b13[2]), .Y(n9747));
INVX1 mul_U5089(.A(dpath_mulcore_b6[2]), .Y(n9733));
INVX1 mul_U5090(.A(dpath_mulcore_b5[2]), .Y(n9731));
INVX1 mul_U5091(.A(dpath_mulcore_b11[2]), .Y(n9743));
INVX1 mul_U5092(.A(dpath_mulcore_b8[2]), .Y(n9737));
INVX1 mul_U5093(.A(dpath_mulcore_b3[2]), .Y(n9727));
AND2X1 mul_U5094(.A(n1120), .B(n13683), .Y(dpath_mulcore_ary1_a1_I1_I2_net38));
AND2X1 mul_U5095(.A(n1123), .B(n13689), .Y(dpath_mulcore_ary1_a1_I0_I2_net38));
AND2X1 mul_U5096(.A(n1112), .B(n13667), .Y(dpath_mulcore_ary1_a0_I1_I2_net38));
INVX1 mul_U5097(.A(n9775), .Y(n9772));
AND2X1 mul_U5098(.A(control_n18), .B(n4686), .Y(control_n7));
INVX1 mul_U5099(.A(dpath_mulcore_x2_c2c3), .Y(n9682));
INVX1 mul_U5100(.A(n9493), .Y(n9569));
INVX1 mul_U5101(.A(n9501), .Y(n9493));
INVX1 mul_U5102(.A(n9571), .Y(n9544));
INVX1 mul_U5103(.A(n9570), .Y(n9545));
INVX1 mul_U5104(.A(acc_reg_shf), .Y(n9779));
INVX1 mul_U5105(.A(mul_spu_shf_ack), .Y(n9780));
INVX1 mul_U5106(.A(n9720), .Y(n9718));
INVX1 mul_U5107(.A(n9720), .Y(n9719));
INVX1 mul_U5108(.A(n9591), .Y(n9590));
INVX1 mul_U5109(.A(n9768), .Y(n9767));
INVX1 mul_U5110(.A(dpath_n662), .Y(n9764));
AND2X1 mul_U5111(.A(n1117), .B(n13677), .Y(dpath_mulcore_ary1_a1_I2_I2_net38));
AND2X1 mul_U5112(.A(n1114), .B(n13671), .Y(dpath_mulcore_ary1_a0_I0_I2_net073));
AND2X1 mul_U5113(.A(n1122), .B(n13687), .Y(dpath_mulcore_ary1_a1_I0_I2_net073));
AND2X1 mul_U5114(.A(n3080), .B(control_n7), .Y(dpath_n522));
INVX1 mul_U5115(.A(dpath_mulcore_clk_enb0), .Y(n9597));
INVX1 mul_U5116(.A(dpath_mulcore_clk_enb0), .Y(n9589));
INVX1 mul_U5117(.A(n9775), .Y(n9773));
INVX1 mul_U5118(.A(dpath_accum_n3), .Y(n9592));
AND2X1 mul_U5119(.A(n2686), .B(n9784), .Y(dpath_mulcore_cyc1_dff_n2));
INVX1 mul_U5120(.A(n9499), .Y(n9583));
INVX1 mul_U5121(.A(n9576), .Y(n9499));
INVX1 mul_U5122(.A(n9501), .Y(n9492));
INVX1 mul_U5123(.A(n9682), .Y(n9673));
OR2X1 mul_U5124(.A(dpath_mulcore_x2_c2), .B(dpath_mulcore_x2_c3), .Y(dpath_mulcore_x2_c2c3));
INVX1 mul_U5125(.A(n9681), .Y(n9674));
AND2X1 mul_U5126(.A(n9774), .B(n6073), .Y(c0_act));
OR2X1 mul_U5127(.A(n7193), .B(acc_actc2), .Y(dpath_n657));
INVX1 mul_U5128(.A(dpath_mulcore_b12[2]), .Y(n9745));
INVX1 mul_U5129(.A(dpath_mulcore_b9[2]), .Y(n9739));
INVX1 mul_U5130(.A(dpath_mulcore_b10[2]), .Y(n9741));
INVX1 mul_U5131(.A(dpath_mulcore_b7[2]), .Y(n9735));
INVX1 mul_U5132(.A(dpath_mulcore_b15[2]), .Y(n9751));
INVX1 mul_U5133(.A(dpath_mulcore_b4[2]), .Y(n9729));
INVX1 mul_U5134(.A(dpath_mulcore_b1[2]), .Y(n9723));
INVX1 mul_U5135(.A(dpath_mulcore_b2[2]), .Y(n9725));
INVX1 mul_U5136(.A(dpath_mulcore_booth_clk_enb1), .Y(n9591));
AND2X1 mul_U5137(.A(dpath_mulcore_booth_ckbuf_1_clken), .B(dpath_mulcore_clk_enb0), .Y(dpath_mulcore_booth_clk_enb1));
AND2X1 mul_U5138(.A(dpath_ckbuf_1_clken), .B(dpath_mulcore_clk_enb0), .Y(dpath_clk_enb1));
XNOR2X1 mul_U5139(.A(n16570), .B(n16573), .Y(n1));
XNOR2X1 mul_U5140(.A(dpath_mulcore_ary1_a1_s2[64]), .B(n8821), .Y(n2));
AND2X1 mul_U5141(.A(dpath_mulcore_cyc1), .B(n9217), .Y(dpath_mulcore_ary1_a0_I0_I2_sc1_66__b));
AND2X1 mul_U5142(.A(byp_imm), .B(dpath_n522), .Y(dpath_n145));
INVX1 mul_U5143(.A(n9763), .Y(n9762));
INVX1 mul_U5144(.A(n9775), .Y(n9774));
AND2X1 mul_U5145(.A(n2414), .B(n9532), .Y(n17815));
AND2X1 mul_U5146(.A(n2417), .B(n9524), .Y(n17818));
AND2X1 mul_U5147(.A(n2420), .B(n9524), .Y(n17821));
AND2X1 mul_U5148(.A(n2423), .B(n9524), .Y(n17824));
AND2X1 mul_U5149(.A(n2426), .B(n9524), .Y(n17827));
AND2X1 mul_U5150(.A(n2429), .B(n9524), .Y(n17830));
AND2X1 mul_U5151(.A(n2432), .B(n9523), .Y(n17833));
AND2X1 mul_U5152(.A(n2435), .B(n9523), .Y(n17836));
AND2X1 mul_U5153(.A(n2438), .B(n9523), .Y(n17839));
AND2X1 mul_U5154(.A(n2441), .B(n9523), .Y(n17842));
AND2X1 mul_U5155(.A(n2444), .B(n9522), .Y(n17845));
AND2X1 mul_U5156(.A(n2447), .B(n9522), .Y(n17848));
AND2X1 mul_U5157(.A(n2450), .B(n9522), .Y(n17851));
AND2X1 mul_U5158(.A(n2453), .B(n9522), .Y(n17854));
AND2X1 mul_U5159(.A(n2456), .B(n9521), .Y(n17857));
AND2X1 mul_U5160(.A(n2484), .B(n9509), .Y(dpath_mulcore_booth_out_dff0_n7));
AND2X1 mul_U5161(.A(n2512), .B(n9539), .Y(dpath_mulcore_a2sum_dff_n39));
AND2X1 mul_U5162(.A(n2513), .B(n9540), .Y(dpath_mulcore_a2sum_dff_n41));
AND2X1 mul_U5163(.A(n2514), .B(n9541), .Y(dpath_mulcore_a2sum_dff_n43));
AND2X1 mul_U5164(.A(n2515), .B(n9543), .Y(dpath_mulcore_a2sum_dff_n47));
AND2X1 mul_U5165(.A(n2516), .B(n9527), .Y(dpath_mulcore_a2sum_dff_n49));
AND2X1 mul_U5166(.A(n2517), .B(n9530), .Y(dpath_mulcore_a2sum_dff_n51));
AND2X1 mul_U5167(.A(n2518), .B(n9522), .Y(dpath_mulcore_a2sum_dff_n53));
AND2X1 mul_U5168(.A(n2519), .B(n9523), .Y(dpath_mulcore_a2sum_dff_n55));
AND2X1 mul_U5169(.A(n2520), .B(n9524), .Y(dpath_mulcore_a2sum_dff_n57));
AND2X1 mul_U5170(.A(n2521), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n59));
AND2X1 mul_U5171(.A(n2523), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n61));
AND2X1 mul_U5172(.A(n2533), .B(n9542), .Y(dpath_mulcore_a2sum_dff_n45));
INVX1 mul_U5173(.A(mul_spu_shf_ack), .Y(n9781));
INVX1 mul_U5174(.A(n9672), .Y(n9701));
INVX1 mul_U5175(.A(n9682), .Y(n9671));
INVX1 mul_U5176(.A(n9682), .Y(n9683));
INVX1 mul_U5177(.A(n9701), .Y(n9684));
AND2X1 mul_U5178(.A(n3081), .B(n4684), .Y(acc_imm));
AND2X1 mul_U5179(.A(dpath_n979), .B(acc_actc2), .Y(dpath_n658));
INVX1 mul_U5180(.A(n9500), .Y(n9494));
AND2X1 mul_U5181(.A(dpath_n984), .B(n6140), .Y(dpath_n661));
OR2X1 mul_U5182(.A(n6140), .B(n7194), .Y(dpath_n662));
AND2X1 mul_U5183(.A(acc_actc3), .B(n9214), .Y(dpath_n666));
INVX1 mul_U5184(.A(dpath_n666), .Y(n9768));
AND2X1 mul_U5185(.A(dpath_mulcore_ckbuf_1_clken), .B(dpath_mulcore_clk_enb0), .Y(dpath_mulcore_clk_enb1));
INVX1 mul_U5186(.A(dpath_mulcore_clk_enb1), .Y(n9720));
AND2X1 mul_U5187(.A(n1111), .B(n13665), .Y(dpath_mulcore_ary1_a0_I1_I2_net073));
AND2X1 mul_U5188(.A(n1119), .B(n13681), .Y(dpath_mulcore_ary1_a1_I1_I2_net073));
AND2X1 mul_U5189(.A(n1109), .B(n13661), .Y(dpath_mulcore_ary1_a0_I2_I2_net38));
AND2X1 mul_U5190(.A(acc_actc3), .B(acc_imm), .Y(dpath_n665));
INVX1 mul_U5191(.A(n9766), .Y(n9765));
INVX1 mul_U5192(.A(dpath_n141), .Y(n9761));
AND2X1 mul_U5193(.A(control_n7), .B(n9215), .Y(dpath_n141));
INVX1 mul_U5194(.A(n9761), .Y(n9760));
AND2X1 mul_U5195(.A(n2412), .B(n9525), .Y(n17813));
AND2X1 mul_U5196(.A(n2413), .B(n9525), .Y(n17814));
AND2X1 mul_U5197(.A(n2415), .B(n9524), .Y(n17816));
AND2X1 mul_U5198(.A(n2416), .B(n9524), .Y(n17817));
AND2X1 mul_U5199(.A(n2418), .B(n9524), .Y(n17819));
AND2X1 mul_U5200(.A(n2419), .B(n9524), .Y(n17820));
AND2X1 mul_U5201(.A(n2421), .B(n9524), .Y(n17822));
AND2X1 mul_U5202(.A(n2422), .B(n9524), .Y(n17823));
AND2X1 mul_U5203(.A(n2424), .B(n9524), .Y(n17825));
AND2X1 mul_U5204(.A(n2425), .B(n9524), .Y(n17826));
AND2X1 mul_U5205(.A(n2427), .B(n9523), .Y(n17828));
AND2X1 mul_U5206(.A(n2428), .B(n9523), .Y(n17829));
AND2X1 mul_U5207(.A(n2430), .B(n9523), .Y(n17831));
AND2X1 mul_U5208(.A(n2431), .B(n9523), .Y(n17832));
AND2X1 mul_U5209(.A(n2433), .B(n9523), .Y(n17834));
AND2X1 mul_U5210(.A(n2434), .B(n9523), .Y(n17835));
AND2X1 mul_U5211(.A(n2436), .B(n9523), .Y(n17837));
AND2X1 mul_U5212(.A(n2437), .B(n9523), .Y(n17838));
AND2X1 mul_U5213(.A(n2439), .B(n9522), .Y(n17840));
AND2X1 mul_U5214(.A(n2440), .B(n9523), .Y(n17841));
AND2X1 mul_U5215(.A(n2442), .B(n9522), .Y(n17843));
AND2X1 mul_U5216(.A(n2443), .B(n9522), .Y(n17844));
AND2X1 mul_U5217(.A(n2445), .B(n9522), .Y(n17846));
AND2X1 mul_U5218(.A(n2446), .B(n9522), .Y(n17847));
AND2X1 mul_U5219(.A(n2448), .B(n9522), .Y(n17849));
AND2X1 mul_U5220(.A(n2449), .B(n9522), .Y(n17850));
AND2X1 mul_U5221(.A(n2451), .B(n9522), .Y(n17852));
AND2X1 mul_U5222(.A(n2452), .B(n9522), .Y(n17853));
AND2X1 mul_U5223(.A(n2454), .B(n9521), .Y(n17855));
AND2X1 mul_U5224(.A(n2455), .B(n9521), .Y(n17856));
AND2X1 mul_U5225(.A(n1734), .B(n9495), .Y(n18226));
AND2X1 mul_U5226(.A(n2197), .B(n9495), .Y(n18227));
AND2X1 mul_U5227(.A(n2193), .B(n9495), .Y(n18228));
AND2X1 mul_U5228(.A(n2194), .B(n9495), .Y(n18229));
AND2X1 mul_U5229(.A(n2195), .B(n9527), .Y(n18230));
AND2X1 mul_U5230(.A(n2196), .B(n9527), .Y(n18231));
AND2X1 mul_U5231(.A(n2192), .B(n9527), .Y(n18232));
AND2X1 mul_U5232(.A(n2199), .B(n9527), .Y(n18234));
AND2X1 mul_U5233(.A(n2201), .B(n9527), .Y(n18235));
AND2X1 mul_U5234(.A(n2203), .B(n9527), .Y(n18236));
AND2X1 mul_U5235(.A(n2205), .B(n9527), .Y(n18237));
AND2X1 mul_U5236(.A(n2207), .B(n9527), .Y(n18238));
AND2X1 mul_U5237(.A(n2209), .B(n9527), .Y(n18239));
AND2X1 mul_U5238(.A(n2211), .B(n9527), .Y(n18240));
AND2X1 mul_U5239(.A(n2213), .B(n9527), .Y(n18241));
AND2X1 mul_U5240(.A(n2215), .B(n9527), .Y(n18242));
AND2X1 mul_U5241(.A(n2217), .B(n9496), .Y(n18243));
AND2X1 mul_U5242(.A(n2219), .B(n9496), .Y(n18245));
AND2X1 mul_U5243(.A(n2221), .B(n9496), .Y(n18246));
AND2X1 mul_U5244(.A(n2223), .B(n9512), .Y(n18247));
AND2X1 mul_U5245(.A(n2225), .B(n9513), .Y(n18248));
AND2X1 mul_U5246(.A(n2227), .B(n9498), .Y(n18249));
AND2X1 mul_U5247(.A(n2229), .B(n9498), .Y(n18250));
AND2X1 mul_U5248(.A(n2231), .B(n9514), .Y(n18251));
AND2X1 mul_U5249(.A(n2233), .B(n9515), .Y(n18252));
AND2X1 mul_U5250(.A(n2235), .B(n9516), .Y(n18253));
AND2X1 mul_U5251(.A(n2237), .B(n9534), .Y(n18254));
AND2X1 mul_U5252(.A(n2239), .B(n9528), .Y(n18256));
AND2X1 mul_U5253(.A(n2241), .B(n9528), .Y(n18257));
AND2X1 mul_U5254(.A(n2243), .B(n9528), .Y(n18258));
AND2X1 mul_U5255(.A(n2245), .B(n9528), .Y(n18259));
AND2X1 mul_U5256(.A(n2247), .B(n9528), .Y(n18260));
AND2X1 mul_U5257(.A(n2249), .B(n9528), .Y(n18261));
AND2X1 mul_U5258(.A(n2251), .B(n9528), .Y(n18262));
AND2X1 mul_U5259(.A(n2253), .B(n9528), .Y(n18263));
AND2X1 mul_U5260(.A(n2255), .B(n9528), .Y(n18264));
AND2X1 mul_U5261(.A(n2257), .B(n9528), .Y(n18265));
AND2X1 mul_U5262(.A(n2259), .B(n9528), .Y(n18267));
AND2X1 mul_U5263(.A(n2261), .B(n9529), .Y(n18268));
AND2X1 mul_U5264(.A(n2263), .B(n9529), .Y(n18269));
AND2X1 mul_U5265(.A(n2265), .B(n9529), .Y(n18270));
AND2X1 mul_U5266(.A(n2267), .B(n9529), .Y(n18271));
AND2X1 mul_U5267(.A(n2269), .B(n9529), .Y(n18272));
AND2X1 mul_U5268(.A(n2271), .B(n9529), .Y(n18273));
AND2X1 mul_U5269(.A(n2273), .B(n9529), .Y(n18274));
AND2X1 mul_U5270(.A(n2275), .B(n9529), .Y(n18275));
AND2X1 mul_U5271(.A(n2277), .B(n9529), .Y(n18276));
AND2X1 mul_U5272(.A(n2279), .B(n9529), .Y(n18278));
AND2X1 mul_U5273(.A(n2281), .B(n9529), .Y(n18279));
AND2X1 mul_U5274(.A(n2283), .B(n9529), .Y(n18280));
AND2X1 mul_U5275(.A(n2285), .B(n9530), .Y(n18281));
AND2X1 mul_U5276(.A(n2287), .B(n9530), .Y(n18282));
AND2X1 mul_U5277(.A(n2289), .B(n9530), .Y(n18283));
AND2X1 mul_U5278(.A(n2291), .B(n9530), .Y(n18284));
AND2X1 mul_U5279(.A(n2293), .B(n9530), .Y(n18285));
AND2X1 mul_U5280(.A(n2295), .B(n9530), .Y(n18286));
AND2X1 mul_U5281(.A(n2297), .B(n9530), .Y(n18287));
AND2X1 mul_U5282(.A(n2299), .B(n9530), .Y(n18288));
AND2X1 mul_U5283(.A(n2301), .B(n9530), .Y(n18289));
AND2X1 mul_U5284(.A(n2303), .B(n9530), .Y(n18290));
AND2X1 mul_U5285(.A(n2305), .B(n9530), .Y(n18291));
AND2X1 mul_U5286(.A(n2307), .B(n9530), .Y(n18292));
AND2X1 mul_U5287(.A(n2309), .B(n9530), .Y(n18293));
AND2X1 mul_U5288(.A(n2311), .B(n9531), .Y(n18294));
AND2X1 mul_U5289(.A(n2313), .B(n9531), .Y(n18295));
AND2X1 mul_U5290(.A(n2315), .B(n9531), .Y(n18296));
AND2X1 mul_U5291(.A(n1738), .B(n9509), .Y(n18221));
AND2X1 mul_U5292(.A(n1739), .B(n9517), .Y(n18222));
AND2X1 mul_U5293(.A(n1740), .B(n9527), .Y(n18233));
AND2X1 mul_U5294(.A(n2686), .B(dpath_mulcore_cyc1), .Y(n18298));
AND2X1 mul_U5295(.A(n2686), .B(dpath_mulcore_cyc2), .Y(n18299));
AND2X1 mul_U5296(.A(n2686), .B(x2), .Y(n18300));
AND2X1 mul_U5297(.A(n2686), .B(dpath_mulcore_x2_c1), .Y(n18301));
AND2X1 mul_U5298(.A(n2686), .B(dpath_mulcore_x2_c2), .Y(n18302));
AND2X1 mul_U5299(.A(n2482), .B(n9509), .Y(dpath_mulcore_booth_out_dff0_n3));
AND2X1 mul_U5300(.A(n2483), .B(n9509), .Y(dpath_mulcore_booth_out_dff0_n5));
AND2X1 mul_U5301(.A(n2492), .B(n9552), .Y(dpath_mulcore_a2sum_dff_n195));
AND2X1 mul_U5302(.A(n2493), .B(n9562), .Y(dpath_mulcore_a2sum_dff_n3));
AND2X1 mul_U5303(.A(n2494), .B(n9562), .Y(dpath_mulcore_a2sum_dff_n5));
AND2X1 mul_U5304(.A(n2495), .B(n9562), .Y(dpath_mulcore_a2sum_dff_n7));
AND2X1 mul_U5305(.A(n2496), .B(n9562), .Y(dpath_mulcore_a2sum_dff_n9));
AND2X1 mul_U5306(.A(n2497), .B(n9562), .Y(dpath_mulcore_a2sum_dff_n11));
AND2X1 mul_U5307(.A(n2498), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n13));
AND2X1 mul_U5308(.A(n2499), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n15));
AND2X1 mul_U5309(.A(n2501), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n17));
AND2X1 mul_U5310(.A(n2502), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n19));
AND2X1 mul_U5311(.A(n2503), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n21));
AND2X1 mul_U5312(.A(n2504), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n25));
AND2X1 mul_U5313(.A(n2505), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n27));
AND2X1 mul_U5314(.A(n2506), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n29));
AND2X1 mul_U5315(.A(n2507), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n31));
AND2X1 mul_U5316(.A(n2508), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n33));
AND2X1 mul_U5317(.A(n2509), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n35));
AND2X1 mul_U5318(.A(n2510), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n37));
AND2X1 mul_U5319(.A(n2524), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n63));
AND2X1 mul_U5320(.A(n2525), .B(n9499), .Y(dpath_mulcore_a2sum_dff_n65));
AND2X1 mul_U5321(.A(n2526), .B(n9499), .Y(dpath_mulcore_a2sum_dff_n69));
AND2X1 mul_U5322(.A(n2527), .B(n9499), .Y(dpath_mulcore_a2sum_dff_n71));
AND2X1 mul_U5323(.A(n2528), .B(n9493), .Y(dpath_mulcore_a2sum_dff_n73));
AND2X1 mul_U5324(.A(n2529), .B(n9495), .Y(dpath_mulcore_a2sum_dff_n75));
AND2X1 mul_U5325(.A(n2530), .B(n9496), .Y(dpath_mulcore_a2sum_dff_n77));
AND2X1 mul_U5326(.A(n2531), .B(n9497), .Y(dpath_mulcore_a2sum_dff_n79));
AND2X1 mul_U5327(.A(n2532), .B(n9498), .Y(dpath_mulcore_a2sum_dff_n81));
AND2X1 mul_U5328(.A(n2534), .B(n9544), .Y(dpath_mulcore_a2sum_dff_n83));
AND2X1 mul_U5329(.A(n2535), .B(n9545), .Y(dpath_mulcore_a2sum_dff_n85));
AND2X1 mul_U5330(.A(n2536), .B(n9546), .Y(dpath_mulcore_a2sum_dff_n87));
AND2X1 mul_U5331(.A(n2537), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n91));
AND2X1 mul_U5332(.A(n2538), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n93));
AND2X1 mul_U5333(.A(n2539), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n95));
AND2X1 mul_U5334(.A(n2540), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n97));
AND2X1 mul_U5335(.A(n2541), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n99));
AND2X1 mul_U5336(.A(n2542), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n101));
AND2X1 mul_U5337(.A(n2543), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n103));
AND2X1 mul_U5338(.A(n2545), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n105));
AND2X1 mul_U5339(.A(n2546), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n107));
AND2X1 mul_U5340(.A(n2547), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n109));
AND2X1 mul_U5341(.A(n2548), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n113));
AND2X1 mul_U5342(.A(n2549), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n115));
AND2X1 mul_U5343(.A(n2550), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n117));
AND2X1 mul_U5344(.A(n2551), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n119));
AND2X1 mul_U5345(.A(n2552), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n121));
AND2X1 mul_U5346(.A(n2553), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n123));
AND2X1 mul_U5347(.A(n2554), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n125));
AND2X1 mul_U5348(.A(n2556), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n127));
AND2X1 mul_U5349(.A(n2557), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n129));
AND2X1 mul_U5350(.A(n2558), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n131));
AND2X1 mul_U5351(.A(n2559), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n135));
AND2X1 mul_U5352(.A(n2560), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n137));
AND2X1 mul_U5353(.A(n2561), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n139));
AND2X1 mul_U5354(.A(n2562), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n141));
AND2X1 mul_U5355(.A(n2563), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n143));
AND2X1 mul_U5356(.A(n2564), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n145));
AND2X1 mul_U5357(.A(n2565), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n147));
AND2X1 mul_U5358(.A(n2567), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n149));
AND2X1 mul_U5359(.A(n2568), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n151));
AND2X1 mul_U5360(.A(n2569), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n153));
AND2X1 mul_U5361(.A(n2570), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n157));
AND2X1 mul_U5362(.A(n2571), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n159));
AND2X1 mul_U5363(.A(n2572), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n161));
AND2X1 mul_U5364(.A(n2573), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n163));
AND2X1 mul_U5365(.A(n2574), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n165));
AND2X1 mul_U5366(.A(n2575), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n167));
AND2X1 mul_U5367(.A(n2576), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n169));
AND2X1 mul_U5368(.A(n2578), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n171));
AND2X1 mul_U5369(.A(n2579), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n173));
AND2X1 mul_U5370(.A(n2580), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n175));
AND2X1 mul_U5371(.A(n2581), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n177));
AND2X1 mul_U5372(.A(n2582), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n179));
AND2X1 mul_U5373(.A(n2583), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n181));
AND2X1 mul_U5374(.A(n2584), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n183));
AND2X1 mul_U5375(.A(n2585), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n185));
AND2X1 mul_U5376(.A(n2586), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n187));
AND2X1 mul_U5377(.A(n2587), .B(n9551), .Y(dpath_mulcore_a2sum_dff_n189));
AND2X1 mul_U5378(.A(n2491), .B(n9552), .Y(dpath_mulcore_a2sum_dff_n191));
AND2X1 mul_U5379(.A(n2500), .B(n9552), .Y(dpath_mulcore_a2sum_dff_n193));
AND2X1 mul_U5380(.A(n2511), .B(n9552), .Y(dpath_mulcore_a2sum_dff_n197));
AND2X1 mul_U5381(.A(n2522), .B(n9563), .Y(dpath_mulcore_a2sum_dff_n23));
AND2X1 mul_U5382(.A(n2544), .B(n9547), .Y(dpath_mulcore_a2sum_dff_n67));
AND2X1 mul_U5383(.A(n2555), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n89));
AND2X1 mul_U5384(.A(n2566), .B(n9548), .Y(dpath_mulcore_a2sum_dff_n111));
AND2X1 mul_U5385(.A(n2577), .B(n9549), .Y(dpath_mulcore_a2sum_dff_n133));
AND2X1 mul_U5386(.A(n2588), .B(n9550), .Y(dpath_mulcore_a2sum_dff_n155));
AND2X1 mul_U5387(.A(n2590), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n3));
AND2X1 mul_U5388(.A(n2591), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n5));
AND2X1 mul_U5389(.A(n2592), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n7));
AND2X1 mul_U5390(.A(n2593), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n9));
AND2X1 mul_U5391(.A(n2594), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n11));
AND2X1 mul_U5392(.A(n2595), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n13));
AND2X1 mul_U5393(.A(n2596), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n15));
AND2X1 mul_U5394(.A(n2598), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n17));
AND2X1 mul_U5395(.A(n2599), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n19));
AND2X1 mul_U5396(.A(n2600), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n21));
AND2X1 mul_U5397(.A(n2601), .B(n9539), .Y(dpath_mulcore_a2cot_dff_n25));
AND2X1 mul_U5398(.A(n2602), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n27));
AND2X1 mul_U5399(.A(n2603), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n29));
AND2X1 mul_U5400(.A(n2604), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n31));
AND2X1 mul_U5401(.A(n2605), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n33));
AND2X1 mul_U5402(.A(n2606), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n35));
AND2X1 mul_U5403(.A(n2607), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n37));
AND2X1 mul_U5404(.A(n2609), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n39));
AND2X1 mul_U5405(.A(n2610), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n41));
AND2X1 mul_U5406(.A(n2611), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n43));
AND2X1 mul_U5407(.A(n2612), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n47));
AND2X1 mul_U5408(.A(n2613), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n49));
AND2X1 mul_U5409(.A(n2614), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n51));
AND2X1 mul_U5410(.A(n2615), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n53));
AND2X1 mul_U5411(.A(n2616), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n55));
AND2X1 mul_U5412(.A(n2617), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n57));
AND2X1 mul_U5413(.A(n2618), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n59));
AND2X1 mul_U5414(.A(n2620), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n61));
AND2X1 mul_U5415(.A(n2621), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n63));
AND2X1 mul_U5416(.A(n2622), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n65));
AND2X1 mul_U5417(.A(n2623), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n69));
AND2X1 mul_U5418(.A(n2624), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n71));
AND2X1 mul_U5419(.A(n2625), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n73));
AND2X1 mul_U5420(.A(n2626), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n75));
AND2X1 mul_U5421(.A(n2627), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n77));
AND2X1 mul_U5422(.A(n2628), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n79));
AND2X1 mul_U5423(.A(n2629), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n81));
AND2X1 mul_U5424(.A(n2631), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n83));
AND2X1 mul_U5425(.A(n2632), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n85));
AND2X1 mul_U5426(.A(n2633), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n87));
AND2X1 mul_U5427(.A(n2634), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n91));
AND2X1 mul_U5428(.A(n2635), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n93));
AND2X1 mul_U5429(.A(n2636), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n95));
AND2X1 mul_U5430(.A(n2637), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n97));
AND2X1 mul_U5431(.A(n2638), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n99));
AND2X1 mul_U5432(.A(n2639), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n101));
AND2X1 mul_U5433(.A(n2640), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n103));
AND2X1 mul_U5434(.A(n2642), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n105));
AND2X1 mul_U5435(.A(n2643), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n107));
AND2X1 mul_U5436(.A(n2644), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n109));
AND2X1 mul_U5437(.A(n2645), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n113));
AND2X1 mul_U5438(.A(n2646), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n115));
AND2X1 mul_U5439(.A(n2647), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n117));
AND2X1 mul_U5440(.A(n2648), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n119));
AND2X1 mul_U5441(.A(n2649), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n121));
AND2X1 mul_U5442(.A(n2650), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n123));
AND2X1 mul_U5443(.A(n2651), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n125));
AND2X1 mul_U5444(.A(n2653), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n127));
AND2X1 mul_U5445(.A(n2654), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n129));
AND2X1 mul_U5446(.A(n2655), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n131));
AND2X1 mul_U5447(.A(n2656), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n135));
AND2X1 mul_U5448(.A(n2657), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n137));
AND2X1 mul_U5449(.A(n2658), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n139));
AND2X1 mul_U5450(.A(n2659), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n141));
AND2X1 mul_U5451(.A(n2660), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n143));
AND2X1 mul_U5452(.A(n2661), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n145));
AND2X1 mul_U5453(.A(n2662), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n147));
AND2X1 mul_U5454(.A(n2664), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n149));
AND2X1 mul_U5455(.A(n2665), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n151));
AND2X1 mul_U5456(.A(n2666), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n153));
AND2X1 mul_U5457(.A(n2667), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n157));
AND2X1 mul_U5458(.A(n2668), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n159));
AND2X1 mul_U5459(.A(n2669), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n161));
AND2X1 mul_U5460(.A(n2670), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n163));
AND2X1 mul_U5461(.A(n2671), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n165));
AND2X1 mul_U5462(.A(n2672), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n167));
AND2X1 mul_U5463(.A(n2673), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n169));
AND2X1 mul_U5464(.A(n2675), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n171));
AND2X1 mul_U5465(.A(n2676), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n173));
AND2X1 mul_U5466(.A(n2677), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n175));
AND2X1 mul_U5467(.A(n2678), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n177));
AND2X1 mul_U5468(.A(n2679), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n179));
AND2X1 mul_U5469(.A(n2680), .B(n9562), .Y(dpath_mulcore_a2cot_dff_n181));
AND2X1 mul_U5470(.A(n2681), .B(n9562), .Y(dpath_mulcore_a2cot_dff_n183));
AND2X1 mul_U5471(.A(n2682), .B(n9562), .Y(dpath_mulcore_a2cot_dff_n185));
AND2X1 mul_U5472(.A(n2683), .B(n9562), .Y(dpath_mulcore_a2cot_dff_n187));
AND2X1 mul_U5473(.A(n2684), .B(n9562), .Y(dpath_mulcore_a2cot_dff_n189));
AND2X1 mul_U5474(.A(n2589), .B(n9562), .Y(dpath_mulcore_a2cot_dff_n191));
AND2X1 mul_U5475(.A(n2597), .B(n9562), .Y(dpath_mulcore_a2cot_dff_n193));
AND2X1 mul_U5476(.A(n2608), .B(n9562), .Y(dpath_mulcore_a2cot_dff_n195));
AND2X1 mul_U5477(.A(n2619), .B(n9538), .Y(dpath_mulcore_a2cot_dff_n23));
AND2X1 mul_U5478(.A(n2630), .B(n9556), .Y(dpath_mulcore_a2cot_dff_n45));
AND2X1 mul_U5479(.A(n2641), .B(n9557), .Y(dpath_mulcore_a2cot_dff_n67));
AND2X1 mul_U5480(.A(n2652), .B(n9558), .Y(dpath_mulcore_a2cot_dff_n89));
AND2X1 mul_U5481(.A(n2663), .B(n9559), .Y(dpath_mulcore_a2cot_dff_n111));
AND2X1 mul_U5482(.A(n2674), .B(n9560), .Y(dpath_mulcore_a2cot_dff_n133));
AND2X1 mul_U5483(.A(n2685), .B(n9561), .Y(dpath_mulcore_a2cot_dff_n155));
AND2X1 mul_U5484(.A(n1600), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n15));
AND2X1 mul_U5485(.A(n2071), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n17));
AND2X1 mul_U5486(.A(n2067), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n19));
AND2X1 mul_U5487(.A(n2068), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n21));
AND2X1 mul_U5488(.A(n2069), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n23));
AND2X1 mul_U5489(.A(n2070), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n25));
AND2X1 mul_U5490(.A(n2481), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n27));
AND2X1 mul_U5491(.A(n2073), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n31));
AND2X1 mul_U5492(.A(n2075), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n33));
AND2X1 mul_U5493(.A(n2077), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n35));
AND2X1 mul_U5494(.A(n2079), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n37));
AND2X1 mul_U5495(.A(n2081), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n39));
AND2X1 mul_U5496(.A(n2083), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n41));
AND2X1 mul_U5497(.A(n2085), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n43));
AND2X1 mul_U5498(.A(n2087), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n45));
AND2X1 mul_U5499(.A(n2089), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n47));
AND2X1 mul_U5500(.A(n2091), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n49));
AND2X1 mul_U5501(.A(n2093), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n53));
AND2X1 mul_U5502(.A(n2095), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n55));
AND2X1 mul_U5503(.A(n2097), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n57));
AND2X1 mul_U5504(.A(n2099), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n59));
AND2X1 mul_U5505(.A(n2101), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n61));
AND2X1 mul_U5506(.A(n2103), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n63));
AND2X1 mul_U5507(.A(n2105), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n65));
AND2X1 mul_U5508(.A(n2107), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n67));
AND2X1 mul_U5509(.A(n2109), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n69));
AND2X1 mul_U5510(.A(n2111), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n71));
AND2X1 mul_U5511(.A(n2113), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n75));
AND2X1 mul_U5512(.A(n2115), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n77));
AND2X1 mul_U5513(.A(n2117), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n79));
AND2X1 mul_U5514(.A(n2119), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n81));
AND2X1 mul_U5515(.A(n2121), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n83));
AND2X1 mul_U5516(.A(n2123), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n85));
AND2X1 mul_U5517(.A(n2125), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n87));
AND2X1 mul_U5518(.A(n2127), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n89));
AND2X1 mul_U5519(.A(n2129), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n91));
AND2X1 mul_U5520(.A(n2131), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n93));
AND2X1 mul_U5521(.A(n2133), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n97));
AND2X1 mul_U5522(.A(n2135), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n99));
AND2X1 mul_U5523(.A(n2137), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n101));
AND2X1 mul_U5524(.A(n2139), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n103));
AND2X1 mul_U5525(.A(n2141), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n105));
AND2X1 mul_U5526(.A(n2143), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n107));
AND2X1 mul_U5527(.A(n2145), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n109));
AND2X1 mul_U5528(.A(n2147), .B(n9495), .Y(dpath_mulcore_a0cot_dff_n111));
AND2X1 mul_U5529(.A(n2149), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n113));
AND2X1 mul_U5530(.A(n2151), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n115));
AND2X1 mul_U5531(.A(n2153), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n119));
AND2X1 mul_U5532(.A(n2155), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n121));
AND2X1 mul_U5533(.A(n2157), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n123));
AND2X1 mul_U5534(.A(n2159), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n125));
AND2X1 mul_U5535(.A(n2161), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n127));
AND2X1 mul_U5536(.A(n2163), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n129));
AND2X1 mul_U5537(.A(n2165), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n131));
AND2X1 mul_U5538(.A(n2167), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n133));
AND2X1 mul_U5539(.A(n2169), .B(n9493), .Y(dpath_mulcore_a0cot_dff_n135));
AND2X1 mul_U5540(.A(n2171), .B(n9493), .Y(dpath_mulcore_a0cot_dff_n137));
AND2X1 mul_U5541(.A(n2173), .B(n9493), .Y(dpath_mulcore_a0cot_dff_n139));
AND2X1 mul_U5542(.A(n2175), .B(n9551), .Y(dpath_mulcore_a0cot_dff_n141));
AND2X1 mul_U5543(.A(n2177), .B(n9552), .Y(dpath_mulcore_a0cot_dff_n143));
AND2X1 mul_U5544(.A(n2179), .B(n9553), .Y(dpath_mulcore_a0cot_dff_n145));
AND2X1 mul_U5545(.A(n2181), .B(n9554), .Y(dpath_mulcore_a0cot_dff_n147));
AND2X1 mul_U5546(.A(n2183), .B(n9555), .Y(dpath_mulcore_a0cot_dff_n149));
AND2X1 mul_U5547(.A(n2185), .B(n9562), .Y(dpath_mulcore_a0cot_dff_n151));
AND2X1 mul_U5548(.A(n2187), .B(n9563), .Y(dpath_mulcore_a0cot_dff_n153));
AND2X1 mul_U5549(.A(n2189), .B(n9556), .Y(dpath_mulcore_a0cot_dff_n155));
AND2X1 mul_U5550(.A(n1604), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n3));
AND2X1 mul_U5551(.A(n1605), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n7));
AND2X1 mul_U5552(.A(n1606), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n29));
AND2X1 mul_U5553(.A(n2687), .B(n9539), .Y(dpath_mulcore_ffrs1_n9));
AND2X1 mul_U5554(.A(n2688), .B(n9539), .Y(dpath_mulcore_ffrs1_n11));
AND2X1 mul_U5555(.A(n2689), .B(n9539), .Y(dpath_mulcore_ffrs1_n13));
AND2X1 mul_U5556(.A(n2690), .B(n9539), .Y(dpath_mulcore_ffrs1_n15));
AND2X1 mul_U5557(.A(n2691), .B(n9539), .Y(dpath_mulcore_ffrs1_n17));
AND2X1 mul_U5558(.A(n2692), .B(n9539), .Y(dpath_mulcore_ffrs1_n19));
AND2X1 mul_U5559(.A(n2693), .B(n9539), .Y(dpath_mulcore_ffrs1_n21));
AND2X1 mul_U5560(.A(n2694), .B(n9539), .Y(dpath_mulcore_ffrs1_n25));
AND2X1 mul_U5561(.A(n2695), .B(n9539), .Y(dpath_mulcore_ffrs1_n27));
AND2X1 mul_U5562(.A(n2696), .B(n9540), .Y(dpath_mulcore_ffrs1_n29));
AND2X1 mul_U5563(.A(n2697), .B(n9540), .Y(dpath_mulcore_ffrs1_n31));
AND2X1 mul_U5564(.A(n2698), .B(n9540), .Y(dpath_mulcore_ffrs1_n33));
AND2X1 mul_U5565(.A(n2699), .B(n9540), .Y(dpath_mulcore_ffrs1_n35));
AND2X1 mul_U5566(.A(n2700), .B(n9540), .Y(dpath_mulcore_ffrs1_n37));
AND2X1 mul_U5567(.A(n2701), .B(n9540), .Y(dpath_mulcore_ffrs1_n39));
AND2X1 mul_U5568(.A(n2702), .B(n9540), .Y(dpath_mulcore_ffrs1_n41));
AND2X1 mul_U5569(.A(n2703), .B(n9540), .Y(dpath_mulcore_ffrs1_n43));
AND2X1 mul_U5570(.A(n2704), .B(n9540), .Y(dpath_mulcore_ffrs1_n47));
AND2X1 mul_U5571(.A(n2705), .B(n9540), .Y(dpath_mulcore_ffrs1_n49));
AND2X1 mul_U5572(.A(n2706), .B(n9540), .Y(dpath_mulcore_ffrs1_n51));
AND2X1 mul_U5573(.A(n2707), .B(n9540), .Y(dpath_mulcore_ffrs1_n53));
AND2X1 mul_U5574(.A(n2708), .B(n9541), .Y(dpath_mulcore_ffrs1_n55));
AND2X1 mul_U5575(.A(n2709), .B(n9541), .Y(dpath_mulcore_ffrs1_n57));
AND2X1 mul_U5576(.A(n2710), .B(n9541), .Y(dpath_mulcore_ffrs1_n59));
AND2X1 mul_U5577(.A(n2711), .B(n9541), .Y(dpath_mulcore_ffrs1_n61));
AND2X1 mul_U5578(.A(n2712), .B(n9541), .Y(dpath_mulcore_ffrs1_n63));
AND2X1 mul_U5579(.A(n2713), .B(n9541), .Y(dpath_mulcore_ffrs1_n65));
AND2X1 mul_U5580(.A(n2714), .B(n9541), .Y(dpath_mulcore_ffrs1_n69));
AND2X1 mul_U5581(.A(n2715), .B(n9541), .Y(dpath_mulcore_ffrs1_n71));
AND2X1 mul_U5582(.A(n2716), .B(n9541), .Y(dpath_mulcore_ffrs1_n73));
AND2X1 mul_U5583(.A(n2717), .B(n9541), .Y(dpath_mulcore_ffrs1_n75));
AND2X1 mul_U5584(.A(n2718), .B(n9541), .Y(dpath_mulcore_ffrs1_n77));
AND2X1 mul_U5585(.A(n2719), .B(n9541), .Y(dpath_mulcore_ffrs1_n79));
AND2X1 mul_U5586(.A(n2720), .B(n9542), .Y(dpath_mulcore_ffrs1_n81));
AND2X1 mul_U5587(.A(n2721), .B(n9542), .Y(dpath_mulcore_ffrs1_n83));
AND2X1 mul_U5588(.A(n2722), .B(n9542), .Y(dpath_mulcore_ffrs1_n85));
AND2X1 mul_U5589(.A(n2723), .B(n9542), .Y(dpath_mulcore_ffrs1_n87));
AND2X1 mul_U5590(.A(n2724), .B(n9542), .Y(dpath_mulcore_ffrs1_n91));
AND2X1 mul_U5591(.A(n2725), .B(n9542), .Y(dpath_mulcore_ffrs1_n93));
AND2X1 mul_U5592(.A(n2726), .B(n9542), .Y(dpath_mulcore_ffrs1_n95));
AND2X1 mul_U5593(.A(n2727), .B(n9542), .Y(dpath_mulcore_ffrs1_n97));
AND2X1 mul_U5594(.A(n2728), .B(n9542), .Y(dpath_mulcore_ffrs1_n99));
AND2X1 mul_U5595(.A(n2729), .B(n9542), .Y(dpath_mulcore_ffrs1_n101));
AND2X1 mul_U5596(.A(n2730), .B(n9542), .Y(dpath_mulcore_ffrs1_n103));
AND2X1 mul_U5597(.A(n2731), .B(n9542), .Y(dpath_mulcore_ffrs1_n105));
AND2X1 mul_U5598(.A(n2732), .B(n9543), .Y(dpath_mulcore_ffrs1_n107));
AND2X1 mul_U5599(.A(n2733), .B(n9543), .Y(dpath_mulcore_ffrs1_n109));
AND2X1 mul_U5600(.A(n2734), .B(n9543), .Y(dpath_mulcore_ffrs1_n111));
AND2X1 mul_U5601(.A(n2735), .B(n9543), .Y(dpath_mulcore_ffrs1_n113));
AND2X1 mul_U5602(.A(n2736), .B(n9543), .Y(dpath_mulcore_ffrs1_n115));
AND2X1 mul_U5603(.A(n2737), .B(n9543), .Y(dpath_mulcore_ffrs1_n117));
AND2X1 mul_U5604(.A(n2738), .B(n9543), .Y(dpath_mulcore_ffrs1_n119));
AND2X1 mul_U5605(.A(n2739), .B(n9543), .Y(dpath_mulcore_ffrs1_n121));
AND2X1 mul_U5606(.A(n2740), .B(n9543), .Y(dpath_mulcore_ffrs1_n123));
AND2X1 mul_U5607(.A(n2741), .B(n9543), .Y(dpath_mulcore_ffrs1_n125));
AND2X1 mul_U5608(.A(n2742), .B(n9543), .Y(dpath_mulcore_ffrs1_n127));
AND2X1 mul_U5609(.A(n2743), .B(n9543), .Y(dpath_mulcore_ffrs1_n129));
AND2X1 mul_U5610(.A(n2744), .B(n9543), .Y(dpath_mulcore_ffrs1_n3));
AND2X1 mul_U5611(.A(n2745), .B(n9539), .Y(dpath_mulcore_ffrs1_n5));
AND2X1 mul_U5612(.A(n2746), .B(n9539), .Y(dpath_mulcore_ffrs1_n7));
AND2X1 mul_U5613(.A(n2747), .B(n9539), .Y(dpath_mulcore_ffrs1_n23));
AND2X1 mul_U5614(.A(n2748), .B(n9540), .Y(dpath_mulcore_ffrs1_n45));
AND2X1 mul_U5615(.A(n2749), .B(n9541), .Y(dpath_mulcore_ffrs1_n67));
AND2X1 mul_U5616(.A(n2750), .B(n9542), .Y(dpath_mulcore_ffrs1_n89));
AND2X1 mul_U5617(.A(n3011), .B(n7195), .Y(dpath_accum_n131));
AND2X1 mul_U5618(.A(n3012), .B(n7195), .Y(dpath_accum_n133));
AND2X1 mul_U5619(.A(n3014), .B(n7195), .Y(dpath_accum_n135));
AND2X1 mul_U5620(.A(n3015), .B(n9592), .Y(dpath_accum_n137));
AND2X1 mul_U5621(.A(n3016), .B(n7195), .Y(dpath_accum_n139));
AND2X1 mul_U5622(.A(n3017), .B(n9592), .Y(dpath_accum_n141));
AND2X1 mul_U5623(.A(n3018), .B(n9592), .Y(dpath_accum_n143));
AND2X1 mul_U5624(.A(n3019), .B(n9592), .Y(dpath_accum_n145));
AND2X1 mul_U5625(.A(n3020), .B(n7195), .Y(dpath_accum_n147));
AND2X1 mul_U5626(.A(n3021), .B(n7195), .Y(dpath_accum_n149));
AND2X1 mul_U5627(.A(n3022), .B(n7195), .Y(dpath_accum_n151));
AND2X1 mul_U5628(.A(n3023), .B(n7195), .Y(dpath_accum_n153));
AND2X1 mul_U5629(.A(n3025), .B(n9592), .Y(dpath_accum_n155));
AND2X1 mul_U5630(.A(n3026), .B(n7195), .Y(dpath_accum_n157));
AND2X1 mul_U5631(.A(n3027), .B(n9592), .Y(dpath_accum_n159));
AND2X1 mul_U5632(.A(n3028), .B(n7195), .Y(dpath_accum_n161));
AND2X1 mul_U5633(.A(n3029), .B(n7195), .Y(dpath_accum_n163));
AND2X1 mul_U5634(.A(n3030), .B(n7195), .Y(dpath_accum_n165));
AND2X1 mul_U5635(.A(n3031), .B(n9592), .Y(dpath_accum_n167));
AND2X1 mul_U5636(.A(n3032), .B(n9592), .Y(dpath_accum_n169));
AND2X1 mul_U5637(.A(n3033), .B(n7195), .Y(dpath_accum_n171));
AND2X1 mul_U5638(.A(n3034), .B(n9592), .Y(dpath_accum_n173));
AND2X1 mul_U5639(.A(n3036), .B(n9592), .Y(dpath_accum_n175));
AND2X1 mul_U5640(.A(n3037), .B(n9592), .Y(dpath_accum_n177));
AND2X1 mul_U5641(.A(n3038), .B(n7195), .Y(dpath_accum_n179));
AND2X1 mul_U5642(.A(n3039), .B(n7195), .Y(dpath_accum_n181));
AND2X1 mul_U5643(.A(n3040), .B(n9592), .Y(dpath_accum_n183));
AND2X1 mul_U5644(.A(n3041), .B(n7195), .Y(dpath_accum_n185));
AND2X1 mul_U5645(.A(n3042), .B(n7195), .Y(dpath_accum_n187));
AND2X1 mul_U5646(.A(n3043), .B(n9592), .Y(dpath_accum_n189));
AND2X1 mul_U5647(.A(n3044), .B(n9592), .Y(dpath_accum_n191));
AND2X1 mul_U5648(.A(n3045), .B(n9592), .Y(dpath_accum_n193));
AND2X1 mul_U5649(.A(n3047), .B(n7195), .Y(dpath_accum_n195));
AND2X1 mul_U5650(.A(n3048), .B(n9592), .Y(dpath_accum_n197));
AND2X1 mul_U5651(.A(n3049), .B(n7195), .Y(dpath_accum_n199));
AND2X1 mul_U5652(.A(n3050), .B(n9592), .Y(dpath_accum_n201));
AND2X1 mul_U5653(.A(n3051), .B(n7195), .Y(dpath_accum_n203));
AND2X1 mul_U5654(.A(n3052), .B(n9592), .Y(dpath_accum_n205));
AND2X1 mul_U5655(.A(n3053), .B(n9592), .Y(dpath_accum_n207));
AND2X1 mul_U5656(.A(n3054), .B(n7195), .Y(dpath_accum_n209));
AND2X1 mul_U5657(.A(n3055), .B(n7195), .Y(dpath_accum_n211));
AND2X1 mul_U5658(.A(n3056), .B(n9592), .Y(dpath_accum_n213));
AND2X1 mul_U5659(.A(n3058), .B(n7195), .Y(dpath_accum_n215));
AND2X1 mul_U5660(.A(n3059), .B(n9592), .Y(dpath_accum_n217));
AND2X1 mul_U5661(.A(n3060), .B(n7195), .Y(dpath_accum_n219));
AND2X1 mul_U5662(.A(n3061), .B(n9592), .Y(dpath_accum_n221));
AND2X1 mul_U5663(.A(n3062), .B(n9592), .Y(dpath_accum_n223));
AND2X1 mul_U5664(.A(n3063), .B(n9592), .Y(dpath_accum_n225));
AND2X1 mul_U5665(.A(n3064), .B(n9592), .Y(dpath_accum_n227));
AND2X1 mul_U5666(.A(n3065), .B(n9592), .Y(dpath_accum_n229));
AND2X1 mul_U5667(.A(n3066), .B(n9592), .Y(dpath_accum_n231));
AND2X1 mul_U5668(.A(n3067), .B(n7195), .Y(dpath_accum_n233));
AND2X1 mul_U5669(.A(n3069), .B(n7195), .Y(dpath_accum_n235));
AND2X1 mul_U5670(.A(n3070), .B(n9592), .Y(dpath_accum_n237));
AND2X1 mul_U5671(.A(n3071), .B(n9592), .Y(dpath_accum_n239));
AND2X1 mul_U5672(.A(n3072), .B(n7195), .Y(dpath_accum_n241));
AND2X1 mul_U5673(.A(n3073), .B(n9592), .Y(dpath_accum_n243));
AND2X1 mul_U5674(.A(n3074), .B(n9592), .Y(dpath_accum_n245));
AND2X1 mul_U5675(.A(n3075), .B(n9592), .Y(dpath_accum_n247));
AND2X1 mul_U5676(.A(n3076), .B(n7195), .Y(dpath_accum_n249));
AND2X1 mul_U5677(.A(n3077), .B(n9592), .Y(dpath_accum_n251));
AND2X1 mul_U5678(.A(n3078), .B(n7195), .Y(dpath_accum_n253));
AND2X1 mul_U5679(.A(n3008), .B(n9592), .Y(dpath_accum_n255));
AND2X1 mul_U5680(.A(n3009), .B(n7195), .Y(dpath_accum_n257));
AND2X1 mul_U5681(.A(n3010), .B(n7195), .Y(dpath_accum_n259));
AND2X1 mul_U5682(.A(n3013), .B(n7195), .Y(dpath_accum_n261));
AND2X1 mul_U5683(.A(n3024), .B(n9592), .Y(dpath_accum_n263));
AND2X1 mul_U5684(.A(n3035), .B(n7195), .Y(dpath_accum_n265));
AND2X1 mul_U5685(.A(n3046), .B(n7195), .Y(dpath_accum_n267));
AND2X1 mul_U5686(.A(n3057), .B(n7195), .Y(dpath_accum_n269));
AND2X1 mul_U5687(.A(n3068), .B(n9592), .Y(dpath_accum_n271));
AND2X1 mul_U5688(.A(n3079), .B(n7195), .Y(dpath_accum_n273));
INVX1 mul_U5689(.A(n9492), .Y(n9564));
INVX1 mul_U5690(.A(se), .Y(n9539));
INVX1 mul_U5691(.A(se), .Y(n9540));
INVX1 mul_U5692(.A(se), .Y(n9541));
INVX1 mul_U5693(.A(n9779), .Y(mul_spu_shf_ack));
INVX1 mul_U5694(.A(acc_reg_shf), .Y(n9782));
INVX1 mul_U5695(.A(mul_spu_shf_ack), .Y(n9783));
INVX1 mul_U5696(.A(dpath_mulcore_clk_enb0), .Y(n9659));
INVX1 mul_U5697(.A(n9671), .Y(n9696));
INVX1 mul_U5698(.A(n9701), .Y(n9685));
INVX1 mul_U5699(.A(dpath_clk_enb1), .Y(n9754));
AND2X1 mul_U5700(.A(n9499), .B(c0_act), .Y(dpath_mulcore_booth_ckbuf_1_N1));
INVX1 mul_U5701(.A(dpath_mulcore_booth_ckbuf_1_N1), .Y(n3));
AND2X1 mul_U5702(.A(n9497), .B(n5071), .Y(dpath_ckbuf_1_N1));
INVX1 mul_U5703(.A(dpath_ckbuf_1_N1), .Y(n4));
AND2X1 mul_U5704(.A(n9037), .B(n9843), .Y(n17022));
INVX1 mul_U5705(.A(dpath_mulcore_ary1_a0_sc3_11__z), .Y(n9843));
AND2X1 mul_U5706(.A(n9098), .B(n9830), .Y(n17466));
INVX1 mul_U5707(.A(dpath_mulcore_ary1_a1_sc3_11__z), .Y(n9830));
AND2X1 mul_U5708(.A(dpath_mulcore_addin_sum[1]), .B(n10184), .Y(n10112));
INVX1 mul_U5709(.A(n10112), .Y(n5));
AND2X1 mul_U5710(.A(dpath_mulcore_addin_sum[2]), .B(n9218), .Y(n10115));
INVX1 mul_U5711(.A(n10115), .Y(n6));
AND2X1 mul_U5712(.A(dpath_mulcore_addin_sum[3]), .B(n9219), .Y(n10118));
INVX1 mul_U5713(.A(n10118), .Y(n7));
AND2X1 mul_U5714(.A(dpath_mulcore_addin_sum[4]), .B(n9220), .Y(n10121));
INVX1 mul_U5715(.A(n10121), .Y(n8));
AND2X1 mul_U5716(.A(dpath_mulcore_addin_sum[5]), .B(n9221), .Y(n10124));
INVX1 mul_U5717(.A(n10124), .Y(n9));
AND2X1 mul_U5718(.A(dpath_mulcore_addin_sum[6]), .B(n9222), .Y(n10127));
INVX1 mul_U5719(.A(n10127), .Y(n10));
AND2X1 mul_U5720(.A(dpath_mulcore_addin_sum[7]), .B(n9223), .Y(n10130));
INVX1 mul_U5721(.A(n10130), .Y(n11));
AND2X1 mul_U5722(.A(dpath_mulcore_addin_sum[8]), .B(n9224), .Y(n10133));
INVX1 mul_U5723(.A(n10133), .Y(n12));
AND2X1 mul_U5724(.A(dpath_mulcore_addin_sum[9]), .B(n9225), .Y(n10136));
INVX1 mul_U5725(.A(n10136), .Y(n13));
AND2X1 mul_U5726(.A(dpath_mulcore_addin_sum[10]), .B(n9235), .Y(n10141));
INVX1 mul_U5727(.A(n10141), .Y(n14));
AND2X1 mul_U5728(.A(dpath_mulcore_addin_sum[11]), .B(n9236), .Y(n10146));
INVX1 mul_U5729(.A(n10146), .Y(n15));
AND2X1 mul_U5730(.A(dpath_mulcore_addin_sum[12]), .B(n9237), .Y(n10151));
INVX1 mul_U5731(.A(n10151), .Y(n16));
AND2X1 mul_U5732(.A(dpath_mulcore_addin_sum[13]), .B(n9238), .Y(n10156));
INVX1 mul_U5733(.A(n10156), .Y(n17));
AND2X1 mul_U5734(.A(dpath_mulcore_addin_sum[14]), .B(n9239), .Y(n10161));
INVX1 mul_U5735(.A(n10161), .Y(n18));
AND2X1 mul_U5736(.A(dpath_mulcore_addin_sum[15]), .B(n9240), .Y(n10166));
INVX1 mul_U5737(.A(n10166), .Y(n19));
AND2X1 mul_U5738(.A(dpath_mulcore_addin_sum[16]), .B(n9241), .Y(n10171));
INVX1 mul_U5739(.A(n10171), .Y(n20));
AND2X1 mul_U5740(.A(dpath_mulcore_addin_sum[17]), .B(n9242), .Y(n10176));
INVX1 mul_U5741(.A(n10176), .Y(n21));
AND2X1 mul_U5742(.A(dpath_mulcore_addin_sum[18]), .B(n9243), .Y(n10181));
INVX1 mul_U5743(.A(n10181), .Y(n22));
AND2X1 mul_U5744(.A(dpath_mulcore_addin_sum[19]), .B(n9244), .Y(n10188));
INVX1 mul_U5745(.A(n10188), .Y(n23));
AND2X1 mul_U5746(.A(dpath_mulcore_addin_sum[20]), .B(n9245), .Y(n10193));
INVX1 mul_U5747(.A(n10193), .Y(n24));
AND2X1 mul_U5748(.A(dpath_mulcore_addin_sum[21]), .B(n9246), .Y(n10198));
INVX1 mul_U5749(.A(n10198), .Y(n25));
AND2X1 mul_U5750(.A(dpath_mulcore_addin_sum[22]), .B(n9247), .Y(n10203));
INVX1 mul_U5751(.A(n10203), .Y(n26));
AND2X1 mul_U5752(.A(dpath_mulcore_addin_sum[23]), .B(n9248), .Y(n10208));
INVX1 mul_U5753(.A(n10208), .Y(n27));
AND2X1 mul_U5754(.A(dpath_mulcore_addin_sum[24]), .B(n9249), .Y(n10213));
INVX1 mul_U5755(.A(n10213), .Y(n28));
AND2X1 mul_U5756(.A(dpath_mulcore_addin_sum[25]), .B(n9250), .Y(n10218));
INVX1 mul_U5757(.A(n10218), .Y(n29));
AND2X1 mul_U5758(.A(dpath_mulcore_addin_sum[26]), .B(n9251), .Y(n10223));
INVX1 mul_U5759(.A(n10223), .Y(n30));
AND2X1 mul_U5760(.A(dpath_mulcore_addin_sum[27]), .B(n9252), .Y(n10228));
INVX1 mul_U5761(.A(n10228), .Y(n31));
AND2X1 mul_U5762(.A(dpath_mulcore_addin_sum[28]), .B(n9253), .Y(n10233));
INVX1 mul_U5763(.A(n10233), .Y(n32));
AND2X1 mul_U5764(.A(dpath_mulcore_addin_sum[29]), .B(n9254), .Y(n10240));
INVX1 mul_U5765(.A(n10240), .Y(n33));
AND2X1 mul_U5766(.A(dpath_mulcore_addin_sum[30]), .B(n9255), .Y(n10245));
INVX1 mul_U5767(.A(n10245), .Y(n34));
AND2X1 mul_U5768(.A(dpath_mulcore_addin_sum[31]), .B(n9256), .Y(n10250));
INVX1 mul_U5769(.A(n10250), .Y(n35));
AND2X1 mul_U5770(.A(dpath_mulcore_addin_cout[31]), .B(dpath_mulcore_addin_sum[32]), .Y(n10268));
INVX1 mul_U5771(.A(n10268), .Y(n36));
AND2X1 mul_U5772(.A(dpath_mulcore_addin_sum[33]), .B(n9226), .Y(n10271));
INVX1 mul_U5773(.A(n10271), .Y(n37));
AND2X1 mul_U5774(.A(dpath_mulcore_addin_sum[34]), .B(n9227), .Y(n10274));
INVX1 mul_U5775(.A(n10274), .Y(n38));
AND2X1 mul_U5776(.A(dpath_mulcore_addin_sum[35]), .B(n9228), .Y(n10277));
INVX1 mul_U5777(.A(n10277), .Y(n39));
AND2X1 mul_U5778(.A(dpath_mulcore_addin_sum[36]), .B(n9229), .Y(n10280));
INVX1 mul_U5779(.A(n10280), .Y(n40));
AND2X1 mul_U5780(.A(dpath_mulcore_addin_sum[37]), .B(n9230), .Y(n10283));
INVX1 mul_U5781(.A(n10283), .Y(n41));
AND2X1 mul_U5782(.A(dpath_mulcore_addin_sum[38]), .B(n9231), .Y(n10286));
INVX1 mul_U5783(.A(n10286), .Y(n42));
AND2X1 mul_U5784(.A(dpath_mulcore_addin_sum[39]), .B(n9232), .Y(n10289));
INVX1 mul_U5785(.A(n10289), .Y(n43));
AND2X1 mul_U5786(.A(dpath_mulcore_addin_sum[40]), .B(n9233), .Y(n10292));
INVX1 mul_U5787(.A(n10292), .Y(n44));
AND2X1 mul_U5788(.A(dpath_mulcore_addin_sum[41]), .B(n9234), .Y(n10295));
INVX1 mul_U5789(.A(n10295), .Y(n45));
AND2X1 mul_U5790(.A(dpath_mulcore_addin_sum[42]), .B(n9257), .Y(n10300));
INVX1 mul_U5791(.A(n10300), .Y(n46));
AND2X1 mul_U5792(.A(dpath_mulcore_addin_sum[43]), .B(n9258), .Y(n10305));
INVX1 mul_U5793(.A(n10305), .Y(n47));
AND2X1 mul_U5794(.A(dpath_mulcore_addin_sum[44]), .B(n9259), .Y(n10310));
INVX1 mul_U5795(.A(n10310), .Y(n48));
AND2X1 mul_U5796(.A(dpath_mulcore_addin_sum[45]), .B(n9260), .Y(n10315));
INVX1 mul_U5797(.A(n10315), .Y(n49));
AND2X1 mul_U5798(.A(dpath_mulcore_addin_sum[46]), .B(n9261), .Y(n10320));
INVX1 mul_U5799(.A(n10320), .Y(n50));
AND2X1 mul_U5800(.A(dpath_mulcore_addin_sum[47]), .B(n9262), .Y(n10325));
INVX1 mul_U5801(.A(n10325), .Y(n51));
AND2X1 mul_U5802(.A(dpath_mulcore_addin_sum[48]), .B(n9263), .Y(n10330));
INVX1 mul_U5803(.A(n10330), .Y(n52));
AND2X1 mul_U5804(.A(dpath_mulcore_addin_sum[49]), .B(n9264), .Y(n10335));
INVX1 mul_U5805(.A(n10335), .Y(n53));
AND2X1 mul_U5806(.A(dpath_mulcore_addin_sum[50]), .B(n9265), .Y(n10340));
INVX1 mul_U5807(.A(n10340), .Y(n54));
AND2X1 mul_U5808(.A(dpath_mulcore_addin_sum[51]), .B(n9266), .Y(n10347));
INVX1 mul_U5809(.A(n10347), .Y(n55));
AND2X1 mul_U5810(.A(dpath_mulcore_addin_sum[52]), .B(n9267), .Y(n10352));
INVX1 mul_U5811(.A(n10352), .Y(n56));
AND2X1 mul_U5812(.A(dpath_mulcore_addin_sum[53]), .B(n9268), .Y(n10357));
INVX1 mul_U5813(.A(n10357), .Y(n57));
AND2X1 mul_U5814(.A(dpath_mulcore_addin_sum[54]), .B(n9269), .Y(n10362));
INVX1 mul_U5815(.A(n10362), .Y(n58));
AND2X1 mul_U5816(.A(dpath_mulcore_addin_sum[55]), .B(n9270), .Y(n10367));
INVX1 mul_U5817(.A(n10367), .Y(n59));
AND2X1 mul_U5818(.A(dpath_mulcore_addin_sum[56]), .B(n9271), .Y(n10372));
INVX1 mul_U5819(.A(n10372), .Y(n60));
AND2X1 mul_U5820(.A(dpath_mulcore_addin_sum[57]), .B(n9272), .Y(n10377));
INVX1 mul_U5821(.A(n10377), .Y(n61));
AND2X1 mul_U5822(.A(dpath_mulcore_addin_sum[58]), .B(n9273), .Y(n10382));
INVX1 mul_U5823(.A(n10382), .Y(n62));
AND2X1 mul_U5824(.A(dpath_mulcore_addin_sum[59]), .B(n9274), .Y(n10387));
INVX1 mul_U5825(.A(n10387), .Y(n63));
AND2X1 mul_U5826(.A(dpath_mulcore_addin_sum[60]), .B(n9275), .Y(n10392));
INVX1 mul_U5827(.A(n10392), .Y(n64));
AND2X1 mul_U5828(.A(dpath_mulcore_addin_sum[61]), .B(n9276), .Y(n10399));
INVX1 mul_U5829(.A(n10399), .Y(n65));
AND2X1 mul_U5830(.A(dpath_mulcore_addin_sum[62]), .B(n9277), .Y(n10404));
INVX1 mul_U5831(.A(n10404), .Y(n66));
AND2X1 mul_U5832(.A(dpath_mulcore_addin_sum[63]), .B(n9278), .Y(n10409));
INVX1 mul_U5833(.A(n10409), .Y(n67));
AND2X1 mul_U5834(.A(dpath_mulcore_addin_sum[64]), .B(n9279), .Y(n10414));
INVX1 mul_U5835(.A(n10414), .Y(n68));
AND2X1 mul_U5836(.A(dpath_mulcore_addin_sum[65]), .B(n9280), .Y(n10419));
INVX1 mul_U5837(.A(n10419), .Y(n69));
AND2X1 mul_U5838(.A(dpath_mulcore_addin_sum[66]), .B(n9281), .Y(n10424));
INVX1 mul_U5839(.A(n10424), .Y(n70));
AND2X1 mul_U5840(.A(dpath_mulcore_addin_sum[67]), .B(n9282), .Y(n10429));
INVX1 mul_U5841(.A(n10429), .Y(n71));
AND2X1 mul_U5842(.A(dpath_mulcore_addin_sum[68]), .B(n9283), .Y(n10434));
INVX1 mul_U5843(.A(n10434), .Y(n72));
AND2X1 mul_U5844(.A(dpath_mulcore_addin_sum[69]), .B(n9284), .Y(n10439));
INVX1 mul_U5845(.A(n10439), .Y(n73));
AND2X1 mul_U5846(.A(dpath_mulcore_addin_sum[70]), .B(n9285), .Y(n10444));
INVX1 mul_U5847(.A(n10444), .Y(n74));
AND2X1 mul_U5848(.A(dpath_mulcore_addin_sum[71]), .B(n9286), .Y(n10451));
INVX1 mul_U5849(.A(n10451), .Y(n75));
AND2X1 mul_U5850(.A(dpath_mulcore_addin_sum[72]), .B(n9287), .Y(n10456));
INVX1 mul_U5851(.A(n10456), .Y(n76));
AND2X1 mul_U5852(.A(dpath_mulcore_addin_sum[73]), .B(n9288), .Y(n10461));
INVX1 mul_U5853(.A(n10461), .Y(n77));
AND2X1 mul_U5854(.A(dpath_mulcore_addin_sum[74]), .B(n9289), .Y(n10466));
INVX1 mul_U5855(.A(n10466), .Y(n78));
AND2X1 mul_U5856(.A(dpath_mulcore_addin_sum[75]), .B(n9290), .Y(n10471));
INVX1 mul_U5857(.A(n10471), .Y(n79));
AND2X1 mul_U5858(.A(dpath_mulcore_addin_sum[76]), .B(n9291), .Y(n10476));
INVX1 mul_U5859(.A(n10476), .Y(n80));
AND2X1 mul_U5860(.A(dpath_mulcore_addin_sum[77]), .B(n9292), .Y(n10481));
INVX1 mul_U5861(.A(n10481), .Y(n81));
AND2X1 mul_U5862(.A(dpath_mulcore_addin_sum[78]), .B(n9293), .Y(n10486));
INVX1 mul_U5863(.A(n10486), .Y(n82));
AND2X1 mul_U5864(.A(dpath_mulcore_addin_sum[79]), .B(n9294), .Y(n10491));
INVX1 mul_U5865(.A(n10491), .Y(n83));
AND2X1 mul_U5866(.A(dpath_mulcore_addin_sum[80]), .B(n9295), .Y(n10496));
INVX1 mul_U5867(.A(n10496), .Y(n84));
AND2X1 mul_U5868(.A(dpath_mulcore_addin_sum[81]), .B(n9296), .Y(n10503));
INVX1 mul_U5869(.A(n10503), .Y(n85));
AND2X1 mul_U5870(.A(dpath_mulcore_addin_sum[82]), .B(n9297), .Y(n10508));
INVX1 mul_U5871(.A(n10508), .Y(n86));
AND2X1 mul_U5872(.A(dpath_mulcore_addin_sum[83]), .B(n9298), .Y(n10513));
INVX1 mul_U5873(.A(n10513), .Y(n87));
AND2X1 mul_U5874(.A(dpath_mulcore_addin_sum[84]), .B(n9299), .Y(n10518));
INVX1 mul_U5875(.A(n10518), .Y(n88));
AND2X1 mul_U5876(.A(dpath_mulcore_addin_sum[85]), .B(n9300), .Y(n10523));
INVX1 mul_U5877(.A(n10523), .Y(n89));
AND2X1 mul_U5878(.A(dpath_mulcore_addin_sum[86]), .B(n9301), .Y(n10528));
INVX1 mul_U5879(.A(n10528), .Y(n90));
AND2X1 mul_U5880(.A(dpath_mulcore_addin_sum[87]), .B(n9302), .Y(n10533));
INVX1 mul_U5881(.A(n10533), .Y(n91));
AND2X1 mul_U5882(.A(dpath_mulcore_addin_sum[88]), .B(n9303), .Y(n10538));
INVX1 mul_U5883(.A(n10538), .Y(n92));
AND2X1 mul_U5884(.A(dpath_mulcore_addin_sum[89]), .B(n9304), .Y(n10543));
INVX1 mul_U5885(.A(n10543), .Y(n93));
AND2X1 mul_U5886(.A(dpath_mulcore_addin_sum[90]), .B(n9305), .Y(n10548));
INVX1 mul_U5887(.A(n10548), .Y(n94));
AND2X1 mul_U5888(.A(dpath_mulcore_addin_sum[91]), .B(n9306), .Y(n10555));
INVX1 mul_U5889(.A(n10555), .Y(n95));
AND2X1 mul_U5890(.A(dpath_mulcore_addin_sum[92]), .B(n9307), .Y(n10560));
INVX1 mul_U5891(.A(n10560), .Y(n96));
AND2X1 mul_U5892(.A(dpath_mulcore_addin_sum[93]), .B(n9308), .Y(n10565));
INVX1 mul_U5893(.A(n10565), .Y(n97));
AND2X1 mul_U5894(.A(dpath_mulcore_addin_sum[94]), .B(n9309), .Y(n10570));
INVX1 mul_U5895(.A(n10570), .Y(n98));
AND2X1 mul_U5896(.A(dpath_mulcore_addin_sum[95]), .B(n9310), .Y(n10575));
INVX1 mul_U5897(.A(n10575), .Y(n99));
AND2X1 mul_U5898(.A(dpath_mulcore_addin_sum[96]), .B(n9311), .Y(n10580));
INVX1 mul_U5899(.A(n10580), .Y(n100));
AND2X1 mul_U5900(.A(dpath_mulcore_ary1_a0_I2_I2_p1_l_64), .B(dpath_mulcore_b7[0]), .Y(n10604));
INVX1 mul_U5901(.A(n10604), .Y(n101));
AND2X1 mul_U5902(.A(dpath_mulcore_ary1_a0_I2_p1_l[63]), .B(dpath_mulcore_b7[0]), .Y(n10607));
INVX1 mul_U5903(.A(n10607), .Y(n102));
AND2X1 mul_U5904(.A(dpath_mulcore_ary1_a0_I2_p1_l[62]), .B(dpath_mulcore_b7[0]), .Y(n10610));
INVX1 mul_U5905(.A(n10610), .Y(n103));
AND2X1 mul_U5906(.A(dpath_mulcore_ary1_a0_I2_p0_l[62]), .B(dpath_mulcore_b6[0]), .Y(n10613));
INVX1 mul_U5907(.A(n10613), .Y(n104));
AND2X1 mul_U5908(.A(dpath_mulcore_ary1_a0_I2_p1_l[61]), .B(dpath_mulcore_b7[0]), .Y(n10616));
INVX1 mul_U5909(.A(n10616), .Y(n105));
AND2X1 mul_U5910(.A(dpath_mulcore_ary1_a0_I2_p0_l[61]), .B(dpath_mulcore_b6[0]), .Y(n10619));
INVX1 mul_U5911(.A(n10619), .Y(n106));
AND2X1 mul_U5912(.A(dpath_mulcore_ary1_a0_I2_p1_l[60]), .B(dpath_mulcore_b7[0]), .Y(n10622));
INVX1 mul_U5913(.A(n10622), .Y(n107));
AND2X1 mul_U5914(.A(dpath_mulcore_ary1_a0_I2_p0_l[60]), .B(dpath_mulcore_b6[0]), .Y(n10625));
INVX1 mul_U5915(.A(n10625), .Y(n108));
AND2X1 mul_U5916(.A(dpath_mulcore_ary1_a0_I2_p1_l[59]), .B(dpath_mulcore_b7[0]), .Y(n10628));
INVX1 mul_U5917(.A(n10628), .Y(n109));
AND2X1 mul_U5918(.A(dpath_mulcore_ary1_a0_I2_p0_l[59]), .B(dpath_mulcore_b6[0]), .Y(n10631));
INVX1 mul_U5919(.A(n10631), .Y(n110));
AND2X1 mul_U5920(.A(dpath_mulcore_ary1_a0_I2_p1_l[58]), .B(dpath_mulcore_b7[0]), .Y(n10634));
INVX1 mul_U5921(.A(n10634), .Y(n111));
AND2X1 mul_U5922(.A(dpath_mulcore_ary1_a0_I2_p0_l[58]), .B(dpath_mulcore_b6[0]), .Y(n10637));
INVX1 mul_U5923(.A(n10637), .Y(n112));
AND2X1 mul_U5924(.A(dpath_mulcore_ary1_a0_I2_p1_l[57]), .B(dpath_mulcore_b7[0]), .Y(n10640));
INVX1 mul_U5925(.A(n10640), .Y(n113));
AND2X1 mul_U5926(.A(dpath_mulcore_ary1_a0_I2_p0_l[57]), .B(dpath_mulcore_b6[0]), .Y(n10643));
INVX1 mul_U5927(.A(n10643), .Y(n114));
AND2X1 mul_U5928(.A(dpath_mulcore_ary1_a0_I2_p1_l[56]), .B(dpath_mulcore_b7[0]), .Y(n10646));
INVX1 mul_U5929(.A(n10646), .Y(n115));
AND2X1 mul_U5930(.A(dpath_mulcore_ary1_a0_I2_p0_l[56]), .B(dpath_mulcore_b6[0]), .Y(n10649));
INVX1 mul_U5931(.A(n10649), .Y(n116));
AND2X1 mul_U5932(.A(dpath_mulcore_ary1_a0_I2_p1_l[55]), .B(dpath_mulcore_b7[0]), .Y(n10652));
INVX1 mul_U5933(.A(n10652), .Y(n117));
AND2X1 mul_U5934(.A(dpath_mulcore_ary1_a0_I2_p0_l[55]), .B(dpath_mulcore_b6[0]), .Y(n10655));
INVX1 mul_U5935(.A(n10655), .Y(n118));
AND2X1 mul_U5936(.A(dpath_mulcore_ary1_a0_I2_p1_l[54]), .B(dpath_mulcore_b7[0]), .Y(n10658));
INVX1 mul_U5937(.A(n10658), .Y(n119));
AND2X1 mul_U5938(.A(dpath_mulcore_ary1_a0_I2_p0_l[54]), .B(dpath_mulcore_b6[0]), .Y(n10661));
INVX1 mul_U5939(.A(n10661), .Y(n120));
AND2X1 mul_U5940(.A(dpath_mulcore_ary1_a0_I2_p1_l[53]), .B(dpath_mulcore_b7[0]), .Y(n10664));
INVX1 mul_U5941(.A(n10664), .Y(n121));
AND2X1 mul_U5942(.A(dpath_mulcore_ary1_a0_I2_p0_l[53]), .B(dpath_mulcore_b6[0]), .Y(n10667));
INVX1 mul_U5943(.A(n10667), .Y(n122));
AND2X1 mul_U5944(.A(dpath_mulcore_ary1_a0_I2_p1_l[52]), .B(dpath_mulcore_b7[0]), .Y(n10670));
INVX1 mul_U5945(.A(n10670), .Y(n123));
AND2X1 mul_U5946(.A(dpath_mulcore_ary1_a0_I2_p0_l[52]), .B(dpath_mulcore_b6[0]), .Y(n10673));
INVX1 mul_U5947(.A(n10673), .Y(n124));
AND2X1 mul_U5948(.A(dpath_mulcore_ary1_a0_I2_p1_l[51]), .B(dpath_mulcore_b7[0]), .Y(n10676));
INVX1 mul_U5949(.A(n10676), .Y(n125));
AND2X1 mul_U5950(.A(dpath_mulcore_ary1_a0_I2_p0_l[51]), .B(dpath_mulcore_b6[0]), .Y(n10679));
INVX1 mul_U5951(.A(n10679), .Y(n126));
AND2X1 mul_U5952(.A(dpath_mulcore_ary1_a0_I2_p1_l[50]), .B(dpath_mulcore_b7[0]), .Y(n10682));
INVX1 mul_U5953(.A(n10682), .Y(n127));
AND2X1 mul_U5954(.A(dpath_mulcore_ary1_a0_I2_p0_l[50]), .B(dpath_mulcore_b6[0]), .Y(n10685));
INVX1 mul_U5955(.A(n10685), .Y(n128));
AND2X1 mul_U5956(.A(dpath_mulcore_ary1_a0_I2_p1_l[49]), .B(dpath_mulcore_b7[0]), .Y(n10688));
INVX1 mul_U5957(.A(n10688), .Y(n129));
AND2X1 mul_U5958(.A(dpath_mulcore_ary1_a0_I2_p0_l[49]), .B(dpath_mulcore_b6[0]), .Y(n10691));
INVX1 mul_U5959(.A(n10691), .Y(n130));
AND2X1 mul_U5960(.A(dpath_mulcore_ary1_a0_I2_p1_l[48]), .B(dpath_mulcore_b7[0]), .Y(n10694));
INVX1 mul_U5961(.A(n10694), .Y(n131));
AND2X1 mul_U5962(.A(dpath_mulcore_ary1_a0_I2_p0_l[48]), .B(dpath_mulcore_b6[0]), .Y(n10697));
INVX1 mul_U5963(.A(n10697), .Y(n132));
AND2X1 mul_U5964(.A(dpath_mulcore_ary1_a0_I2_p1_l[47]), .B(dpath_mulcore_b7[0]), .Y(n10700));
INVX1 mul_U5965(.A(n10700), .Y(n133));
AND2X1 mul_U5966(.A(dpath_mulcore_ary1_a0_I2_p0_l[47]), .B(dpath_mulcore_b6[0]), .Y(n10703));
INVX1 mul_U5967(.A(n10703), .Y(n134));
AND2X1 mul_U5968(.A(dpath_mulcore_ary1_a0_I2_p1_l[46]), .B(dpath_mulcore_b7[0]), .Y(n10706));
INVX1 mul_U5969(.A(n10706), .Y(n135));
AND2X1 mul_U5970(.A(dpath_mulcore_ary1_a0_I2_p0_l[46]), .B(dpath_mulcore_b6[0]), .Y(n10709));
INVX1 mul_U5971(.A(n10709), .Y(n136));
AND2X1 mul_U5972(.A(dpath_mulcore_ary1_a0_I2_p1_l[45]), .B(dpath_mulcore_b7[0]), .Y(n10712));
INVX1 mul_U5973(.A(n10712), .Y(n137));
AND2X1 mul_U5974(.A(dpath_mulcore_ary1_a0_I2_p0_l[45]), .B(dpath_mulcore_b6[0]), .Y(n10715));
INVX1 mul_U5975(.A(n10715), .Y(n138));
AND2X1 mul_U5976(.A(dpath_mulcore_ary1_a0_I2_p1_l[44]), .B(dpath_mulcore_b7[0]), .Y(n10718));
INVX1 mul_U5977(.A(n10718), .Y(n139));
AND2X1 mul_U5978(.A(dpath_mulcore_ary1_a0_I2_p0_l[44]), .B(dpath_mulcore_b6[0]), .Y(n10721));
INVX1 mul_U5979(.A(n10721), .Y(n140));
AND2X1 mul_U5980(.A(dpath_mulcore_ary1_a0_I2_p1_l[43]), .B(dpath_mulcore_b7[0]), .Y(n10724));
INVX1 mul_U5981(.A(n10724), .Y(n141));
AND2X1 mul_U5982(.A(dpath_mulcore_ary1_a0_I2_p0_l[43]), .B(dpath_mulcore_b6[0]), .Y(n10727));
INVX1 mul_U5983(.A(n10727), .Y(n142));
AND2X1 mul_U5984(.A(dpath_mulcore_ary1_a0_I2_p1_l[42]), .B(dpath_mulcore_b7[0]), .Y(n10730));
INVX1 mul_U5985(.A(n10730), .Y(n143));
AND2X1 mul_U5986(.A(dpath_mulcore_ary1_a0_I2_p0_l[42]), .B(dpath_mulcore_b6[0]), .Y(n10733));
INVX1 mul_U5987(.A(n10733), .Y(n144));
AND2X1 mul_U5988(.A(dpath_mulcore_ary1_a0_I2_p1_l[41]), .B(dpath_mulcore_b7[0]), .Y(n10736));
INVX1 mul_U5989(.A(n10736), .Y(n145));
AND2X1 mul_U5990(.A(dpath_mulcore_ary1_a0_I2_p0_l[41]), .B(dpath_mulcore_b6[0]), .Y(n10739));
INVX1 mul_U5991(.A(n10739), .Y(n146));
AND2X1 mul_U5992(.A(dpath_mulcore_ary1_a0_I2_p1_l[40]), .B(dpath_mulcore_b7[0]), .Y(n10742));
INVX1 mul_U5993(.A(n10742), .Y(n147));
AND2X1 mul_U5994(.A(dpath_mulcore_ary1_a0_I2_p0_l[40]), .B(dpath_mulcore_b6[0]), .Y(n10745));
INVX1 mul_U5995(.A(n10745), .Y(n148));
AND2X1 mul_U5996(.A(dpath_mulcore_ary1_a0_I2_p1_l[39]), .B(dpath_mulcore_b7[0]), .Y(n10748));
INVX1 mul_U5997(.A(n10748), .Y(n149));
AND2X1 mul_U5998(.A(dpath_mulcore_ary1_a0_I2_p0_l[39]), .B(dpath_mulcore_b6[0]), .Y(n10751));
INVX1 mul_U5999(.A(n10751), .Y(n150));
AND2X1 mul_U6000(.A(dpath_mulcore_ary1_a0_I2_p1_l[38]), .B(dpath_mulcore_b7[0]), .Y(n10754));
INVX1 mul_U6001(.A(n10754), .Y(n151));
AND2X1 mul_U6002(.A(dpath_mulcore_ary1_a0_I2_p0_l[38]), .B(dpath_mulcore_b6[0]), .Y(n10757));
INVX1 mul_U6003(.A(n10757), .Y(n152));
AND2X1 mul_U6004(.A(dpath_mulcore_ary1_a0_I2_p1_l[37]), .B(dpath_mulcore_b7[0]), .Y(n10760));
INVX1 mul_U6005(.A(n10760), .Y(n153));
AND2X1 mul_U6006(.A(dpath_mulcore_ary1_a0_I2_p0_l[37]), .B(dpath_mulcore_b6[0]), .Y(n10763));
INVX1 mul_U6007(.A(n10763), .Y(n154));
AND2X1 mul_U6008(.A(dpath_mulcore_ary1_a0_I2_p1_l[36]), .B(dpath_mulcore_b7[0]), .Y(n10766));
INVX1 mul_U6009(.A(n10766), .Y(n155));
AND2X1 mul_U6010(.A(dpath_mulcore_ary1_a0_I2_p0_l[36]), .B(dpath_mulcore_b6[0]), .Y(n10769));
INVX1 mul_U6011(.A(n10769), .Y(n156));
AND2X1 mul_U6012(.A(dpath_mulcore_ary1_a0_I2_p1_l[35]), .B(dpath_mulcore_b7[0]), .Y(n10772));
INVX1 mul_U6013(.A(n10772), .Y(n157));
AND2X1 mul_U6014(.A(dpath_mulcore_ary1_a0_I2_p0_l[35]), .B(dpath_mulcore_b6[0]), .Y(n10775));
INVX1 mul_U6015(.A(n10775), .Y(n158));
AND2X1 mul_U6016(.A(dpath_mulcore_ary1_a0_I2_p1_l[34]), .B(dpath_mulcore_b7[0]), .Y(n10778));
INVX1 mul_U6017(.A(n10778), .Y(n159));
AND2X1 mul_U6018(.A(dpath_mulcore_ary1_a0_I2_p0_l[34]), .B(dpath_mulcore_b6[0]), .Y(n10781));
INVX1 mul_U6019(.A(n10781), .Y(n160));
AND2X1 mul_U6020(.A(dpath_mulcore_ary1_a0_I2_p1_l[33]), .B(dpath_mulcore_b7[0]), .Y(n10784));
INVX1 mul_U6021(.A(n10784), .Y(n161));
AND2X1 mul_U6022(.A(dpath_mulcore_ary1_a0_I2_p0_l[33]), .B(dpath_mulcore_b6[0]), .Y(n10787));
INVX1 mul_U6023(.A(n10787), .Y(n162));
AND2X1 mul_U6024(.A(dpath_mulcore_ary1_a0_I2_p1_l[32]), .B(dpath_mulcore_b7[0]), .Y(n10790));
INVX1 mul_U6025(.A(n10790), .Y(n163));
AND2X1 mul_U6026(.A(dpath_mulcore_ary1_a0_I2_p0_l[32]), .B(dpath_mulcore_b6[0]), .Y(n10793));
INVX1 mul_U6027(.A(n10793), .Y(n164));
AND2X1 mul_U6028(.A(dpath_mulcore_ary1_a0_I2_p1_l[31]), .B(dpath_mulcore_b7[0]), .Y(n10796));
INVX1 mul_U6029(.A(n10796), .Y(n165));
AND2X1 mul_U6030(.A(dpath_mulcore_ary1_a0_I2_p0_l[31]), .B(dpath_mulcore_b6[0]), .Y(n10799));
INVX1 mul_U6031(.A(n10799), .Y(n166));
AND2X1 mul_U6032(.A(dpath_mulcore_ary1_a0_I2_p1_l[30]), .B(dpath_mulcore_b7[0]), .Y(n10802));
INVX1 mul_U6033(.A(n10802), .Y(n167));
AND2X1 mul_U6034(.A(dpath_mulcore_ary1_a0_I2_p0_l[30]), .B(dpath_mulcore_b6[0]), .Y(n10805));
INVX1 mul_U6035(.A(n10805), .Y(n168));
AND2X1 mul_U6036(.A(dpath_mulcore_ary1_a0_I2_p1_l[29]), .B(dpath_mulcore_b7[0]), .Y(n10808));
INVX1 mul_U6037(.A(n10808), .Y(n169));
AND2X1 mul_U6038(.A(dpath_mulcore_ary1_a0_I2_p0_l[29]), .B(dpath_mulcore_b6[0]), .Y(n10811));
INVX1 mul_U6039(.A(n10811), .Y(n170));
AND2X1 mul_U6040(.A(dpath_mulcore_ary1_a0_I2_p1_l[28]), .B(dpath_mulcore_b7[0]), .Y(n10814));
INVX1 mul_U6041(.A(n10814), .Y(n171));
AND2X1 mul_U6042(.A(dpath_mulcore_ary1_a0_I2_p0_l[28]), .B(dpath_mulcore_b6[0]), .Y(n10817));
INVX1 mul_U6043(.A(n10817), .Y(n172));
AND2X1 mul_U6044(.A(dpath_mulcore_ary1_a0_I2_p1_l[27]), .B(dpath_mulcore_b7[0]), .Y(n10820));
INVX1 mul_U6045(.A(n10820), .Y(n173));
AND2X1 mul_U6046(.A(dpath_mulcore_ary1_a0_I2_p0_l[27]), .B(dpath_mulcore_b6[0]), .Y(n10823));
INVX1 mul_U6047(.A(n10823), .Y(n174));
AND2X1 mul_U6048(.A(dpath_mulcore_ary1_a0_I2_p1_l[26]), .B(dpath_mulcore_b7[0]), .Y(n10826));
INVX1 mul_U6049(.A(n10826), .Y(n175));
AND2X1 mul_U6050(.A(dpath_mulcore_ary1_a0_I2_p0_l[26]), .B(dpath_mulcore_b6[0]), .Y(n10829));
INVX1 mul_U6051(.A(n10829), .Y(n176));
AND2X1 mul_U6052(.A(dpath_mulcore_ary1_a0_I2_p1_l[25]), .B(dpath_mulcore_b7[0]), .Y(n10832));
INVX1 mul_U6053(.A(n10832), .Y(n177));
AND2X1 mul_U6054(.A(dpath_mulcore_ary1_a0_I2_p0_l[25]), .B(dpath_mulcore_b6[0]), .Y(n10835));
INVX1 mul_U6055(.A(n10835), .Y(n178));
AND2X1 mul_U6056(.A(dpath_mulcore_ary1_a0_I2_p1_l[24]), .B(dpath_mulcore_b7[0]), .Y(n10838));
INVX1 mul_U6057(.A(n10838), .Y(n179));
AND2X1 mul_U6058(.A(dpath_mulcore_ary1_a0_I2_p0_l[24]), .B(dpath_mulcore_b6[0]), .Y(n10841));
INVX1 mul_U6059(.A(n10841), .Y(n180));
AND2X1 mul_U6060(.A(dpath_mulcore_ary1_a0_I2_p1_l[23]), .B(dpath_mulcore_b7[0]), .Y(n10844));
INVX1 mul_U6061(.A(n10844), .Y(n181));
AND2X1 mul_U6062(.A(dpath_mulcore_ary1_a0_I2_p0_l[23]), .B(dpath_mulcore_b6[0]), .Y(n10847));
INVX1 mul_U6063(.A(n10847), .Y(n182));
AND2X1 mul_U6064(.A(dpath_mulcore_ary1_a0_I2_p1_l[22]), .B(dpath_mulcore_b7[0]), .Y(n10850));
INVX1 mul_U6065(.A(n10850), .Y(n183));
AND2X1 mul_U6066(.A(dpath_mulcore_ary1_a0_I2_p0_l[22]), .B(dpath_mulcore_b6[0]), .Y(n10853));
INVX1 mul_U6067(.A(n10853), .Y(n184));
AND2X1 mul_U6068(.A(dpath_mulcore_ary1_a0_I2_p1_l[21]), .B(dpath_mulcore_b7[0]), .Y(n10856));
INVX1 mul_U6069(.A(n10856), .Y(n185));
AND2X1 mul_U6070(.A(dpath_mulcore_ary1_a0_I2_p0_l[21]), .B(dpath_mulcore_b6[0]), .Y(n10859));
INVX1 mul_U6071(.A(n10859), .Y(n186));
AND2X1 mul_U6072(.A(dpath_mulcore_ary1_a0_I2_p1_l[20]), .B(dpath_mulcore_b7[0]), .Y(n10862));
INVX1 mul_U6073(.A(n10862), .Y(n187));
AND2X1 mul_U6074(.A(dpath_mulcore_ary1_a0_I2_p0_l[20]), .B(dpath_mulcore_b6[0]), .Y(n10865));
INVX1 mul_U6075(.A(n10865), .Y(n188));
AND2X1 mul_U6076(.A(dpath_mulcore_ary1_a0_I2_p1_l[19]), .B(dpath_mulcore_b7[0]), .Y(n10868));
INVX1 mul_U6077(.A(n10868), .Y(n189));
AND2X1 mul_U6078(.A(dpath_mulcore_ary1_a0_I2_p0_l[19]), .B(dpath_mulcore_b6[0]), .Y(n10871));
INVX1 mul_U6079(.A(n10871), .Y(n190));
AND2X1 mul_U6080(.A(dpath_mulcore_ary1_a0_I2_p1_l[18]), .B(dpath_mulcore_b7[0]), .Y(n10874));
INVX1 mul_U6081(.A(n10874), .Y(n191));
AND2X1 mul_U6082(.A(dpath_mulcore_ary1_a0_I2_p0_l[18]), .B(dpath_mulcore_b6[0]), .Y(n10877));
INVX1 mul_U6083(.A(n10877), .Y(n192));
AND2X1 mul_U6084(.A(dpath_mulcore_ary1_a0_I2_p1_l[17]), .B(dpath_mulcore_b7[0]), .Y(n10880));
INVX1 mul_U6085(.A(n10880), .Y(n193));
AND2X1 mul_U6086(.A(dpath_mulcore_ary1_a0_I2_p0_l[17]), .B(dpath_mulcore_b6[0]), .Y(n10883));
INVX1 mul_U6087(.A(n10883), .Y(n194));
AND2X1 mul_U6088(.A(dpath_mulcore_ary1_a0_I2_p1_l[16]), .B(dpath_mulcore_b7[0]), .Y(n10886));
INVX1 mul_U6089(.A(n10886), .Y(n195));
AND2X1 mul_U6090(.A(dpath_mulcore_ary1_a0_I2_p0_l[16]), .B(dpath_mulcore_b6[0]), .Y(n10889));
INVX1 mul_U6091(.A(n10889), .Y(n196));
AND2X1 mul_U6092(.A(dpath_mulcore_ary1_a0_I2_p1_l[15]), .B(dpath_mulcore_b7[0]), .Y(n10892));
INVX1 mul_U6093(.A(n10892), .Y(n197));
AND2X1 mul_U6094(.A(dpath_mulcore_ary1_a0_I2_p0_l[15]), .B(dpath_mulcore_b6[0]), .Y(n10895));
INVX1 mul_U6095(.A(n10895), .Y(n198));
AND2X1 mul_U6096(.A(dpath_mulcore_ary1_a0_I2_p1_l[14]), .B(dpath_mulcore_b7[0]), .Y(n10898));
INVX1 mul_U6097(.A(n10898), .Y(n199));
AND2X1 mul_U6098(.A(dpath_mulcore_ary1_a0_I2_p0_l[14]), .B(dpath_mulcore_b6[0]), .Y(n10901));
INVX1 mul_U6099(.A(n10901), .Y(n200));
AND2X1 mul_U6100(.A(dpath_mulcore_ary1_a0_I2_p1_l[13]), .B(dpath_mulcore_b7[0]), .Y(n10904));
INVX1 mul_U6101(.A(n10904), .Y(n201));
AND2X1 mul_U6102(.A(dpath_mulcore_ary1_a0_I2_p0_l[13]), .B(dpath_mulcore_b6[0]), .Y(n10907));
INVX1 mul_U6103(.A(n10907), .Y(n202));
AND2X1 mul_U6104(.A(dpath_mulcore_ary1_a0_I2_p1_l[12]), .B(dpath_mulcore_b7[0]), .Y(n10910));
INVX1 mul_U6105(.A(n10910), .Y(n203));
AND2X1 mul_U6106(.A(dpath_mulcore_ary1_a0_I2_p0_l[12]), .B(dpath_mulcore_b6[0]), .Y(n10913));
INVX1 mul_U6107(.A(n10913), .Y(n204));
AND2X1 mul_U6108(.A(dpath_mulcore_ary1_a0_I2_p1_l[11]), .B(dpath_mulcore_b7[0]), .Y(n10916));
INVX1 mul_U6109(.A(n10916), .Y(n205));
AND2X1 mul_U6110(.A(dpath_mulcore_ary1_a0_I2_p0_l[11]), .B(dpath_mulcore_b6[0]), .Y(n10919));
INVX1 mul_U6111(.A(n10919), .Y(n206));
AND2X1 mul_U6112(.A(dpath_mulcore_ary1_a0_I2_p1_l[10]), .B(dpath_mulcore_b7[0]), .Y(n10922));
INVX1 mul_U6113(.A(n10922), .Y(n207));
AND2X1 mul_U6114(.A(dpath_mulcore_ary1_a0_I2_p0_l[10]), .B(dpath_mulcore_b6[0]), .Y(n10925));
INVX1 mul_U6115(.A(n10925), .Y(n208));
AND2X1 mul_U6116(.A(dpath_mulcore_ary1_a0_I2_p1_l[9]), .B(dpath_mulcore_b7[0]), .Y(n10928));
INVX1 mul_U6117(.A(n10928), .Y(n209));
AND2X1 mul_U6118(.A(dpath_mulcore_ary1_a0_I2_p0_l[9]), .B(dpath_mulcore_b6[0]), .Y(n10931));
INVX1 mul_U6119(.A(n10931), .Y(n210));
AND2X1 mul_U6120(.A(dpath_mulcore_ary1_a0_I2_p1_l[8]), .B(dpath_mulcore_b7[0]), .Y(n10934));
INVX1 mul_U6121(.A(n10934), .Y(n211));
AND2X1 mul_U6122(.A(dpath_mulcore_ary1_a0_I2_p0_l[8]), .B(dpath_mulcore_b6[0]), .Y(n10937));
INVX1 mul_U6123(.A(n10937), .Y(n212));
AND2X1 mul_U6124(.A(dpath_mulcore_ary1_a0_I2_p1_l[7]), .B(dpath_mulcore_b7[0]), .Y(n10940));
INVX1 mul_U6125(.A(n10940), .Y(n213));
AND2X1 mul_U6126(.A(dpath_mulcore_ary1_a0_I2_p0_l[7]), .B(dpath_mulcore_b6[0]), .Y(n10943));
INVX1 mul_U6127(.A(n10943), .Y(n214));
AND2X1 mul_U6128(.A(dpath_mulcore_ary1_a0_I2_p1_l[6]), .B(dpath_mulcore_b7[0]), .Y(n10946));
INVX1 mul_U6129(.A(n10946), .Y(n215));
AND2X1 mul_U6130(.A(dpath_mulcore_ary1_a0_I2_p0_l[6]), .B(dpath_mulcore_b6[0]), .Y(n10949));
INVX1 mul_U6131(.A(n10949), .Y(n216));
AND2X1 mul_U6132(.A(dpath_mulcore_ary1_a0_I2_p1_l[5]), .B(dpath_mulcore_b7[0]), .Y(n10952));
INVX1 mul_U6133(.A(n10952), .Y(n217));
AND2X1 mul_U6134(.A(dpath_mulcore_ary1_a0_I2_p0_l[5]), .B(dpath_mulcore_b6[0]), .Y(n10955));
INVX1 mul_U6135(.A(n10955), .Y(n218));
AND2X1 mul_U6136(.A(dpath_mulcore_ary1_a0_I2_p1_l[4]), .B(dpath_mulcore_b7[0]), .Y(n10958));
INVX1 mul_U6137(.A(n10958), .Y(n219));
AND2X1 mul_U6138(.A(dpath_mulcore_ary1_a0_I2_p0_l[4]), .B(dpath_mulcore_b6[0]), .Y(n10961));
INVX1 mul_U6139(.A(n10961), .Y(n220));
AND2X1 mul_U6140(.A(dpath_mulcore_ary1_a0_I2_p1_l[3]), .B(dpath_mulcore_b7[0]), .Y(n10964));
INVX1 mul_U6141(.A(n10964), .Y(n221));
AND2X1 mul_U6142(.A(dpath_mulcore_ary1_a0_I2_p0_l[3]), .B(dpath_mulcore_b6[0]), .Y(n10967));
INVX1 mul_U6143(.A(n10967), .Y(n222));
AND2X1 mul_U6144(.A(dpath_mulcore_ary1_a0_I2_I0_p0_l_2), .B(dpath_mulcore_b6[0]), .Y(n10970));
INVX1 mul_U6145(.A(n10970), .Y(n223));
AND2X1 mul_U6146(.A(dpath_mulcore_ary1_a0_I2_I0_p1_l_2), .B(dpath_mulcore_b7[0]), .Y(n10973));
INVX1 mul_U6147(.A(n10973), .Y(n224));
AND2X1 mul_U6148(.A(dpath_mulcore_ary1_a0_I2_I0_p0_l_1), .B(dpath_mulcore_b6[0]), .Y(n10976));
INVX1 mul_U6149(.A(n10976), .Y(n225));
AND2X1 mul_U6150(.A(dpath_mulcore_ary1_a0_I2_I0_p0_l_0), .B(dpath_mulcore_b6[0]), .Y(n10979));
INVX1 mul_U6151(.A(n10979), .Y(n226));
AND2X1 mul_U6152(.A(dpath_mulcore_ary1_a0_I1_I2_p2_l_66), .B(dpath_mulcore_b5[0]), .Y(n10986));
INVX1 mul_U6153(.A(n10986), .Y(n227));
AND2X1 mul_U6154(.A(dpath_mulcore_ary1_a0_I1_I2_p2_l_65), .B(dpath_mulcore_b5[0]), .Y(n10989));
INVX1 mul_U6155(.A(n10989), .Y(n228));
AND2X1 mul_U6156(.A(dpath_mulcore_ary1_a0_I1_I2_p2_l_64), .B(dpath_mulcore_b5[0]), .Y(n10992));
INVX1 mul_U6157(.A(n10992), .Y(n229));
AND2X1 mul_U6158(.A(dpath_mulcore_ary1_a0_I1_I2_p1_l_64), .B(dpath_mulcore_b4[0]), .Y(n10995));
INVX1 mul_U6159(.A(n10995), .Y(n230));
AND2X1 mul_U6160(.A(dpath_mulcore_ary1_a0_I1_p1_l[63]), .B(dpath_mulcore_b4[0]), .Y(n10998));
INVX1 mul_U6161(.A(n10998), .Y(n231));
AND2X1 mul_U6162(.A(dpath_mulcore_ary1_a0_I1_p2_l[63]), .B(dpath_mulcore_b5[0]), .Y(n11001));
INVX1 mul_U6163(.A(n11001), .Y(n232));
AND2X1 mul_U6164(.A(dpath_mulcore_ary1_a0_I1_p2_l[62]), .B(dpath_mulcore_b5[0]), .Y(n11004));
INVX1 mul_U6165(.A(n11004), .Y(n233));
AND2X1 mul_U6166(.A(dpath_mulcore_ary1_a0_I1_p1_l[62]), .B(dpath_mulcore_b4[0]), .Y(n11007));
INVX1 mul_U6167(.A(n11007), .Y(n234));
AND2X1 mul_U6168(.A(dpath_mulcore_ary1_a0_I1_p0_l[62]), .B(dpath_mulcore_b3[0]), .Y(n11010));
INVX1 mul_U6169(.A(n11010), .Y(n235));
AND2X1 mul_U6170(.A(dpath_mulcore_ary1_a0_I1_p2_l[61]), .B(dpath_mulcore_b5[0]), .Y(n11013));
INVX1 mul_U6171(.A(n11013), .Y(n236));
AND2X1 mul_U6172(.A(dpath_mulcore_ary1_a0_I1_p1_l[61]), .B(dpath_mulcore_b4[0]), .Y(n11016));
INVX1 mul_U6173(.A(n11016), .Y(n237));
AND2X1 mul_U6174(.A(dpath_mulcore_ary1_a0_I1_p0_l[61]), .B(dpath_mulcore_b3[0]), .Y(n11019));
INVX1 mul_U6175(.A(n11019), .Y(n238));
AND2X1 mul_U6176(.A(dpath_mulcore_ary1_a0_I1_p2_l[60]), .B(dpath_mulcore_b5[0]), .Y(n11022));
INVX1 mul_U6177(.A(n11022), .Y(n239));
AND2X1 mul_U6178(.A(dpath_mulcore_ary1_a0_I1_p1_l[60]), .B(dpath_mulcore_b4[0]), .Y(n11025));
INVX1 mul_U6179(.A(n11025), .Y(n240));
AND2X1 mul_U6180(.A(dpath_mulcore_ary1_a0_I1_p0_l[60]), .B(dpath_mulcore_b3[0]), .Y(n11028));
INVX1 mul_U6181(.A(n11028), .Y(n241));
AND2X1 mul_U6182(.A(dpath_mulcore_ary1_a0_I1_p2_l[59]), .B(dpath_mulcore_b5[0]), .Y(n11031));
INVX1 mul_U6183(.A(n11031), .Y(n242));
AND2X1 mul_U6184(.A(dpath_mulcore_ary1_a0_I1_p1_l[59]), .B(dpath_mulcore_b4[0]), .Y(n11034));
INVX1 mul_U6185(.A(n11034), .Y(n243));
AND2X1 mul_U6186(.A(dpath_mulcore_ary1_a0_I1_p0_l[59]), .B(dpath_mulcore_b3[0]), .Y(n11037));
INVX1 mul_U6187(.A(n11037), .Y(n244));
AND2X1 mul_U6188(.A(dpath_mulcore_ary1_a0_I1_p2_l[58]), .B(dpath_mulcore_b5[0]), .Y(n11040));
INVX1 mul_U6189(.A(n11040), .Y(n245));
AND2X1 mul_U6190(.A(dpath_mulcore_ary1_a0_I1_p1_l[58]), .B(dpath_mulcore_b4[0]), .Y(n11043));
INVX1 mul_U6191(.A(n11043), .Y(n246));
AND2X1 mul_U6192(.A(dpath_mulcore_ary1_a0_I1_p0_l[58]), .B(dpath_mulcore_b3[0]), .Y(n11046));
INVX1 mul_U6193(.A(n11046), .Y(n247));
AND2X1 mul_U6194(.A(dpath_mulcore_ary1_a0_I1_p2_l[57]), .B(dpath_mulcore_b5[0]), .Y(n11049));
INVX1 mul_U6195(.A(n11049), .Y(n248));
AND2X1 mul_U6196(.A(dpath_mulcore_ary1_a0_I1_p1_l[57]), .B(dpath_mulcore_b4[0]), .Y(n11052));
INVX1 mul_U6197(.A(n11052), .Y(n249));
AND2X1 mul_U6198(.A(dpath_mulcore_ary1_a0_I1_p0_l[57]), .B(dpath_mulcore_b3[0]), .Y(n11055));
INVX1 mul_U6199(.A(n11055), .Y(n250));
AND2X1 mul_U6200(.A(dpath_mulcore_ary1_a0_I1_p2_l[56]), .B(dpath_mulcore_b5[0]), .Y(n11058));
INVX1 mul_U6201(.A(n11058), .Y(n251));
AND2X1 mul_U6202(.A(dpath_mulcore_ary1_a0_I1_p1_l[56]), .B(dpath_mulcore_b4[0]), .Y(n11061));
INVX1 mul_U6203(.A(n11061), .Y(n252));
AND2X1 mul_U6204(.A(dpath_mulcore_ary1_a0_I1_p0_l[56]), .B(dpath_mulcore_b3[0]), .Y(n11064));
INVX1 mul_U6205(.A(n11064), .Y(n253));
AND2X1 mul_U6206(.A(dpath_mulcore_ary1_a0_I1_p2_l[55]), .B(dpath_mulcore_b5[0]), .Y(n11067));
INVX1 mul_U6207(.A(n11067), .Y(n254));
AND2X1 mul_U6208(.A(dpath_mulcore_ary1_a0_I1_p1_l[55]), .B(dpath_mulcore_b4[0]), .Y(n11070));
INVX1 mul_U6209(.A(n11070), .Y(n255));
AND2X1 mul_U6210(.A(dpath_mulcore_ary1_a0_I1_p0_l[55]), .B(dpath_mulcore_b3[0]), .Y(n11073));
INVX1 mul_U6211(.A(n11073), .Y(n256));
AND2X1 mul_U6212(.A(dpath_mulcore_ary1_a0_I1_p2_l[54]), .B(dpath_mulcore_b5[0]), .Y(n11076));
INVX1 mul_U6213(.A(n11076), .Y(n257));
AND2X1 mul_U6214(.A(dpath_mulcore_ary1_a0_I1_p1_l[54]), .B(dpath_mulcore_b4[0]), .Y(n11079));
INVX1 mul_U6215(.A(n11079), .Y(n258));
AND2X1 mul_U6216(.A(dpath_mulcore_ary1_a0_I1_p0_l[54]), .B(dpath_mulcore_b3[0]), .Y(n11082));
INVX1 mul_U6217(.A(n11082), .Y(n259));
AND2X1 mul_U6218(.A(dpath_mulcore_ary1_a0_I1_p2_l[53]), .B(dpath_mulcore_b5[0]), .Y(n11085));
INVX1 mul_U6219(.A(n11085), .Y(n260));
AND2X1 mul_U6220(.A(dpath_mulcore_ary1_a0_I1_p1_l[53]), .B(dpath_mulcore_b4[0]), .Y(n11088));
INVX1 mul_U6221(.A(n11088), .Y(n261));
AND2X1 mul_U6222(.A(dpath_mulcore_ary1_a0_I1_p0_l[53]), .B(dpath_mulcore_b3[0]), .Y(n11091));
INVX1 mul_U6223(.A(n11091), .Y(n262));
AND2X1 mul_U6224(.A(dpath_mulcore_ary1_a0_I1_p2_l[52]), .B(dpath_mulcore_b5[0]), .Y(n11094));
INVX1 mul_U6225(.A(n11094), .Y(n263));
AND2X1 mul_U6226(.A(dpath_mulcore_ary1_a0_I1_p1_l[52]), .B(dpath_mulcore_b4[0]), .Y(n11097));
INVX1 mul_U6227(.A(n11097), .Y(n264));
AND2X1 mul_U6228(.A(dpath_mulcore_ary1_a0_I1_p0_l[52]), .B(dpath_mulcore_b3[0]), .Y(n11100));
INVX1 mul_U6229(.A(n11100), .Y(n265));
AND2X1 mul_U6230(.A(dpath_mulcore_ary1_a0_I1_p2_l[51]), .B(dpath_mulcore_b5[0]), .Y(n11103));
INVX1 mul_U6231(.A(n11103), .Y(n266));
AND2X1 mul_U6232(.A(dpath_mulcore_ary1_a0_I1_p1_l[51]), .B(dpath_mulcore_b4[0]), .Y(n11106));
INVX1 mul_U6233(.A(n11106), .Y(n267));
AND2X1 mul_U6234(.A(dpath_mulcore_ary1_a0_I1_p0_l[51]), .B(dpath_mulcore_b3[0]), .Y(n11109));
INVX1 mul_U6235(.A(n11109), .Y(n268));
AND2X1 mul_U6236(.A(dpath_mulcore_ary1_a0_I1_p2_l[50]), .B(dpath_mulcore_b5[0]), .Y(n11112));
INVX1 mul_U6237(.A(n11112), .Y(n269));
AND2X1 mul_U6238(.A(dpath_mulcore_ary1_a0_I1_p1_l[50]), .B(dpath_mulcore_b4[0]), .Y(n11115));
INVX1 mul_U6239(.A(n11115), .Y(n270));
AND2X1 mul_U6240(.A(dpath_mulcore_ary1_a0_I1_p0_l[50]), .B(dpath_mulcore_b3[0]), .Y(n11118));
INVX1 mul_U6241(.A(n11118), .Y(n271));
AND2X1 mul_U6242(.A(dpath_mulcore_ary1_a0_I1_p2_l[49]), .B(dpath_mulcore_b5[0]), .Y(n11121));
INVX1 mul_U6243(.A(n11121), .Y(n272));
AND2X1 mul_U6244(.A(dpath_mulcore_ary1_a0_I1_p1_l[49]), .B(dpath_mulcore_b4[0]), .Y(n11124));
INVX1 mul_U6245(.A(n11124), .Y(n273));
AND2X1 mul_U6246(.A(dpath_mulcore_ary1_a0_I1_p0_l[49]), .B(dpath_mulcore_b3[0]), .Y(n11127));
INVX1 mul_U6247(.A(n11127), .Y(n274));
AND2X1 mul_U6248(.A(dpath_mulcore_ary1_a0_I1_p2_l[48]), .B(dpath_mulcore_b5[0]), .Y(n11130));
INVX1 mul_U6249(.A(n11130), .Y(n275));
AND2X1 mul_U6250(.A(dpath_mulcore_ary1_a0_I1_p1_l[48]), .B(dpath_mulcore_b4[0]), .Y(n11133));
INVX1 mul_U6251(.A(n11133), .Y(n276));
AND2X1 mul_U6252(.A(dpath_mulcore_ary1_a0_I1_p0_l[48]), .B(dpath_mulcore_b3[0]), .Y(n11136));
INVX1 mul_U6253(.A(n11136), .Y(n277));
AND2X1 mul_U6254(.A(dpath_mulcore_ary1_a0_I1_p2_l[47]), .B(dpath_mulcore_b5[0]), .Y(n11139));
INVX1 mul_U6255(.A(n11139), .Y(n278));
AND2X1 mul_U6256(.A(dpath_mulcore_ary1_a0_I1_p1_l[47]), .B(dpath_mulcore_b4[0]), .Y(n11142));
INVX1 mul_U6257(.A(n11142), .Y(n279));
AND2X1 mul_U6258(.A(dpath_mulcore_ary1_a0_I1_p0_l[47]), .B(dpath_mulcore_b3[0]), .Y(n11145));
INVX1 mul_U6259(.A(n11145), .Y(n280));
AND2X1 mul_U6260(.A(dpath_mulcore_ary1_a0_I1_p2_l[46]), .B(dpath_mulcore_b5[0]), .Y(n11148));
INVX1 mul_U6261(.A(n11148), .Y(n281));
AND2X1 mul_U6262(.A(dpath_mulcore_ary1_a0_I1_p1_l[46]), .B(dpath_mulcore_b4[0]), .Y(n11151));
INVX1 mul_U6263(.A(n11151), .Y(n282));
AND2X1 mul_U6264(.A(dpath_mulcore_ary1_a0_I1_p0_l[46]), .B(dpath_mulcore_b3[0]), .Y(n11154));
INVX1 mul_U6265(.A(n11154), .Y(n283));
AND2X1 mul_U6266(.A(dpath_mulcore_ary1_a0_I1_p2_l[45]), .B(dpath_mulcore_b5[0]), .Y(n11157));
INVX1 mul_U6267(.A(n11157), .Y(n284));
AND2X1 mul_U6268(.A(dpath_mulcore_ary1_a0_I1_p1_l[45]), .B(dpath_mulcore_b4[0]), .Y(n11160));
INVX1 mul_U6269(.A(n11160), .Y(n285));
AND2X1 mul_U6270(.A(dpath_mulcore_ary1_a0_I1_p0_l[45]), .B(dpath_mulcore_b3[0]), .Y(n11163));
INVX1 mul_U6271(.A(n11163), .Y(n286));
AND2X1 mul_U6272(.A(dpath_mulcore_ary1_a0_I1_p2_l[44]), .B(dpath_mulcore_b5[0]), .Y(n11166));
INVX1 mul_U6273(.A(n11166), .Y(n287));
AND2X1 mul_U6274(.A(dpath_mulcore_ary1_a0_I1_p1_l[44]), .B(dpath_mulcore_b4[0]), .Y(n11169));
INVX1 mul_U6275(.A(n11169), .Y(n288));
AND2X1 mul_U6276(.A(dpath_mulcore_ary1_a0_I1_p0_l[44]), .B(dpath_mulcore_b3[0]), .Y(n11172));
INVX1 mul_U6277(.A(n11172), .Y(n289));
AND2X1 mul_U6278(.A(dpath_mulcore_ary1_a0_I1_p2_l[43]), .B(dpath_mulcore_b5[0]), .Y(n11175));
INVX1 mul_U6279(.A(n11175), .Y(n290));
AND2X1 mul_U6280(.A(dpath_mulcore_ary1_a0_I1_p1_l[43]), .B(dpath_mulcore_b4[0]), .Y(n11178));
INVX1 mul_U6281(.A(n11178), .Y(n291));
AND2X1 mul_U6282(.A(dpath_mulcore_ary1_a0_I1_p0_l[43]), .B(dpath_mulcore_b3[0]), .Y(n11181));
INVX1 mul_U6283(.A(n11181), .Y(n292));
AND2X1 mul_U6284(.A(dpath_mulcore_ary1_a0_I1_p2_l[42]), .B(dpath_mulcore_b5[0]), .Y(n11184));
INVX1 mul_U6285(.A(n11184), .Y(n293));
AND2X1 mul_U6286(.A(dpath_mulcore_ary1_a0_I1_p1_l[42]), .B(dpath_mulcore_b4[0]), .Y(n11187));
INVX1 mul_U6287(.A(n11187), .Y(n294));
AND2X1 mul_U6288(.A(dpath_mulcore_ary1_a0_I1_p0_l[42]), .B(dpath_mulcore_b3[0]), .Y(n11190));
INVX1 mul_U6289(.A(n11190), .Y(n295));
AND2X1 mul_U6290(.A(dpath_mulcore_ary1_a0_I1_p2_l[41]), .B(dpath_mulcore_b5[0]), .Y(n11193));
INVX1 mul_U6291(.A(n11193), .Y(n296));
AND2X1 mul_U6292(.A(dpath_mulcore_ary1_a0_I1_p1_l[41]), .B(dpath_mulcore_b4[0]), .Y(n11196));
INVX1 mul_U6293(.A(n11196), .Y(n297));
AND2X1 mul_U6294(.A(dpath_mulcore_ary1_a0_I1_p0_l[41]), .B(dpath_mulcore_b3[0]), .Y(n11199));
INVX1 mul_U6295(.A(n11199), .Y(n298));
AND2X1 mul_U6296(.A(dpath_mulcore_ary1_a0_I1_p2_l[40]), .B(dpath_mulcore_b5[0]), .Y(n11202));
INVX1 mul_U6297(.A(n11202), .Y(n299));
AND2X1 mul_U6298(.A(dpath_mulcore_ary1_a0_I1_p1_l[40]), .B(dpath_mulcore_b4[0]), .Y(n11205));
INVX1 mul_U6299(.A(n11205), .Y(n300));
AND2X1 mul_U6300(.A(dpath_mulcore_ary1_a0_I1_p0_l[40]), .B(dpath_mulcore_b3[0]), .Y(n11208));
INVX1 mul_U6301(.A(n11208), .Y(n301));
AND2X1 mul_U6302(.A(dpath_mulcore_ary1_a0_I1_p2_l[39]), .B(dpath_mulcore_b5[0]), .Y(n11211));
INVX1 mul_U6303(.A(n11211), .Y(n302));
AND2X1 mul_U6304(.A(dpath_mulcore_ary1_a0_I1_p1_l[39]), .B(dpath_mulcore_b4[0]), .Y(n11214));
INVX1 mul_U6305(.A(n11214), .Y(n303));
AND2X1 mul_U6306(.A(dpath_mulcore_ary1_a0_I1_p0_l[39]), .B(dpath_mulcore_b3[0]), .Y(n11217));
INVX1 mul_U6307(.A(n11217), .Y(n304));
AND2X1 mul_U6308(.A(dpath_mulcore_ary1_a0_I1_p2_l[38]), .B(dpath_mulcore_b5[0]), .Y(n11220));
INVX1 mul_U6309(.A(n11220), .Y(n305));
AND2X1 mul_U6310(.A(dpath_mulcore_ary1_a0_I1_p1_l[38]), .B(dpath_mulcore_b4[0]), .Y(n11223));
INVX1 mul_U6311(.A(n11223), .Y(n306));
AND2X1 mul_U6312(.A(dpath_mulcore_ary1_a0_I1_p0_l[38]), .B(dpath_mulcore_b3[0]), .Y(n11226));
INVX1 mul_U6313(.A(n11226), .Y(n307));
AND2X1 mul_U6314(.A(dpath_mulcore_ary1_a0_I1_p2_l[37]), .B(dpath_mulcore_b5[0]), .Y(n11229));
INVX1 mul_U6315(.A(n11229), .Y(n308));
AND2X1 mul_U6316(.A(dpath_mulcore_ary1_a0_I1_p1_l[37]), .B(dpath_mulcore_b4[0]), .Y(n11232));
INVX1 mul_U6317(.A(n11232), .Y(n309));
AND2X1 mul_U6318(.A(dpath_mulcore_ary1_a0_I1_p0_l[37]), .B(dpath_mulcore_b3[0]), .Y(n11235));
INVX1 mul_U6319(.A(n11235), .Y(n310));
AND2X1 mul_U6320(.A(dpath_mulcore_ary1_a0_I1_p2_l[36]), .B(dpath_mulcore_b5[0]), .Y(n11238));
INVX1 mul_U6321(.A(n11238), .Y(n311));
AND2X1 mul_U6322(.A(dpath_mulcore_ary1_a0_I1_p1_l[36]), .B(dpath_mulcore_b4[0]), .Y(n11241));
INVX1 mul_U6323(.A(n11241), .Y(n312));
AND2X1 mul_U6324(.A(dpath_mulcore_ary1_a0_I1_p0_l[36]), .B(dpath_mulcore_b3[0]), .Y(n11244));
INVX1 mul_U6325(.A(n11244), .Y(n313));
AND2X1 mul_U6326(.A(dpath_mulcore_ary1_a0_I1_p2_l[35]), .B(dpath_mulcore_b5[0]), .Y(n11247));
INVX1 mul_U6327(.A(n11247), .Y(n314));
AND2X1 mul_U6328(.A(dpath_mulcore_ary1_a0_I1_p1_l[35]), .B(dpath_mulcore_b4[0]), .Y(n11250));
INVX1 mul_U6329(.A(n11250), .Y(n315));
AND2X1 mul_U6330(.A(dpath_mulcore_ary1_a0_I1_p0_l[35]), .B(dpath_mulcore_b3[0]), .Y(n11253));
INVX1 mul_U6331(.A(n11253), .Y(n316));
AND2X1 mul_U6332(.A(dpath_mulcore_ary1_a0_I1_p2_l[34]), .B(dpath_mulcore_b5[0]), .Y(n11256));
INVX1 mul_U6333(.A(n11256), .Y(n317));
AND2X1 mul_U6334(.A(dpath_mulcore_ary1_a0_I1_p1_l[34]), .B(dpath_mulcore_b4[0]), .Y(n11259));
INVX1 mul_U6335(.A(n11259), .Y(n318));
AND2X1 mul_U6336(.A(dpath_mulcore_ary1_a0_I1_p0_l[34]), .B(dpath_mulcore_b3[0]), .Y(n11262));
INVX1 mul_U6337(.A(n11262), .Y(n319));
AND2X1 mul_U6338(.A(dpath_mulcore_ary1_a0_I1_p2_l[33]), .B(dpath_mulcore_b5[0]), .Y(n11265));
INVX1 mul_U6339(.A(n11265), .Y(n320));
AND2X1 mul_U6340(.A(dpath_mulcore_ary1_a0_I1_p1_l[33]), .B(dpath_mulcore_b4[0]), .Y(n11268));
INVX1 mul_U6341(.A(n11268), .Y(n321));
AND2X1 mul_U6342(.A(dpath_mulcore_ary1_a0_I1_p0_l[33]), .B(dpath_mulcore_b3[0]), .Y(n11271));
INVX1 mul_U6343(.A(n11271), .Y(n322));
AND2X1 mul_U6344(.A(dpath_mulcore_ary1_a0_I1_p2_l[32]), .B(dpath_mulcore_b5[0]), .Y(n11274));
INVX1 mul_U6345(.A(n11274), .Y(n323));
AND2X1 mul_U6346(.A(dpath_mulcore_ary1_a0_I1_p1_l[32]), .B(dpath_mulcore_b4[0]), .Y(n11277));
INVX1 mul_U6347(.A(n11277), .Y(n324));
AND2X1 mul_U6348(.A(dpath_mulcore_ary1_a0_I1_p0_l[32]), .B(dpath_mulcore_b3[0]), .Y(n11280));
INVX1 mul_U6349(.A(n11280), .Y(n325));
AND2X1 mul_U6350(.A(dpath_mulcore_ary1_a0_I1_p2_l[31]), .B(dpath_mulcore_b5[0]), .Y(n11283));
INVX1 mul_U6351(.A(n11283), .Y(n326));
AND2X1 mul_U6352(.A(dpath_mulcore_ary1_a0_I1_p1_l[31]), .B(dpath_mulcore_b4[0]), .Y(n11286));
INVX1 mul_U6353(.A(n11286), .Y(n327));
AND2X1 mul_U6354(.A(dpath_mulcore_ary1_a0_I1_p0_l[31]), .B(dpath_mulcore_b3[0]), .Y(n11289));
INVX1 mul_U6355(.A(n11289), .Y(n328));
AND2X1 mul_U6356(.A(dpath_mulcore_ary1_a0_I1_p2_l[30]), .B(dpath_mulcore_b5[0]), .Y(n11292));
INVX1 mul_U6357(.A(n11292), .Y(n329));
AND2X1 mul_U6358(.A(dpath_mulcore_ary1_a0_I1_p1_l[30]), .B(dpath_mulcore_b4[0]), .Y(n11295));
INVX1 mul_U6359(.A(n11295), .Y(n330));
AND2X1 mul_U6360(.A(dpath_mulcore_ary1_a0_I1_p0_l[30]), .B(dpath_mulcore_b3[0]), .Y(n11298));
INVX1 mul_U6361(.A(n11298), .Y(n331));
AND2X1 mul_U6362(.A(dpath_mulcore_ary1_a0_I1_p2_l[29]), .B(dpath_mulcore_b5[0]), .Y(n11301));
INVX1 mul_U6363(.A(n11301), .Y(n332));
AND2X1 mul_U6364(.A(dpath_mulcore_ary1_a0_I1_p1_l[29]), .B(dpath_mulcore_b4[0]), .Y(n11304));
INVX1 mul_U6365(.A(n11304), .Y(n333));
AND2X1 mul_U6366(.A(dpath_mulcore_ary1_a0_I1_p0_l[29]), .B(dpath_mulcore_b3[0]), .Y(n11307));
INVX1 mul_U6367(.A(n11307), .Y(n334));
AND2X1 mul_U6368(.A(dpath_mulcore_ary1_a0_I1_p2_l[28]), .B(dpath_mulcore_b5[0]), .Y(n11310));
INVX1 mul_U6369(.A(n11310), .Y(n335));
AND2X1 mul_U6370(.A(dpath_mulcore_ary1_a0_I1_p1_l[28]), .B(dpath_mulcore_b4[0]), .Y(n11313));
INVX1 mul_U6371(.A(n11313), .Y(n336));
AND2X1 mul_U6372(.A(dpath_mulcore_ary1_a0_I1_p0_l[28]), .B(dpath_mulcore_b3[0]), .Y(n11316));
INVX1 mul_U6373(.A(n11316), .Y(n337));
AND2X1 mul_U6374(.A(dpath_mulcore_ary1_a0_I1_p2_l[27]), .B(dpath_mulcore_b5[0]), .Y(n11319));
INVX1 mul_U6375(.A(n11319), .Y(n338));
AND2X1 mul_U6376(.A(dpath_mulcore_ary1_a0_I1_p1_l[27]), .B(dpath_mulcore_b4[0]), .Y(n11322));
INVX1 mul_U6377(.A(n11322), .Y(n339));
AND2X1 mul_U6378(.A(dpath_mulcore_ary1_a0_I1_p0_l[27]), .B(dpath_mulcore_b3[0]), .Y(n11325));
INVX1 mul_U6379(.A(n11325), .Y(n340));
AND2X1 mul_U6380(.A(dpath_mulcore_ary1_a0_I1_p2_l[26]), .B(dpath_mulcore_b5[0]), .Y(n11328));
INVX1 mul_U6381(.A(n11328), .Y(n341));
AND2X1 mul_U6382(.A(dpath_mulcore_ary1_a0_I1_p1_l[26]), .B(dpath_mulcore_b4[0]), .Y(n11331));
INVX1 mul_U6383(.A(n11331), .Y(n342));
AND2X1 mul_U6384(.A(dpath_mulcore_ary1_a0_I1_p0_l[26]), .B(dpath_mulcore_b3[0]), .Y(n11334));
INVX1 mul_U6385(.A(n11334), .Y(n343));
AND2X1 mul_U6386(.A(dpath_mulcore_ary1_a0_I1_p2_l[25]), .B(dpath_mulcore_b5[0]), .Y(n11337));
INVX1 mul_U6387(.A(n11337), .Y(n344));
AND2X1 mul_U6388(.A(dpath_mulcore_ary1_a0_I1_p1_l[25]), .B(dpath_mulcore_b4[0]), .Y(n11340));
INVX1 mul_U6389(.A(n11340), .Y(n345));
AND2X1 mul_U6390(.A(dpath_mulcore_ary1_a0_I1_p0_l[25]), .B(dpath_mulcore_b3[0]), .Y(n11343));
INVX1 mul_U6391(.A(n11343), .Y(n346));
AND2X1 mul_U6392(.A(dpath_mulcore_ary1_a0_I1_p2_l[24]), .B(dpath_mulcore_b5[0]), .Y(n11346));
INVX1 mul_U6393(.A(n11346), .Y(n347));
AND2X1 mul_U6394(.A(dpath_mulcore_ary1_a0_I1_p1_l[24]), .B(dpath_mulcore_b4[0]), .Y(n11349));
INVX1 mul_U6395(.A(n11349), .Y(n348));
AND2X1 mul_U6396(.A(dpath_mulcore_ary1_a0_I1_p0_l[24]), .B(dpath_mulcore_b3[0]), .Y(n11352));
INVX1 mul_U6397(.A(n11352), .Y(n349));
AND2X1 mul_U6398(.A(dpath_mulcore_ary1_a0_I1_p2_l[23]), .B(dpath_mulcore_b5[0]), .Y(n11355));
INVX1 mul_U6399(.A(n11355), .Y(n350));
AND2X1 mul_U6400(.A(dpath_mulcore_ary1_a0_I1_p1_l[23]), .B(dpath_mulcore_b4[0]), .Y(n11358));
INVX1 mul_U6401(.A(n11358), .Y(n351));
AND2X1 mul_U6402(.A(dpath_mulcore_ary1_a0_I1_p0_l[23]), .B(dpath_mulcore_b3[0]), .Y(n11361));
INVX1 mul_U6403(.A(n11361), .Y(n352));
AND2X1 mul_U6404(.A(dpath_mulcore_ary1_a0_I1_p2_l[22]), .B(dpath_mulcore_b5[0]), .Y(n11364));
INVX1 mul_U6405(.A(n11364), .Y(n353));
AND2X1 mul_U6406(.A(dpath_mulcore_ary1_a0_I1_p1_l[22]), .B(dpath_mulcore_b4[0]), .Y(n11367));
INVX1 mul_U6407(.A(n11367), .Y(n354));
AND2X1 mul_U6408(.A(dpath_mulcore_ary1_a0_I1_p0_l[22]), .B(dpath_mulcore_b3[0]), .Y(n11370));
INVX1 mul_U6409(.A(n11370), .Y(n355));
AND2X1 mul_U6410(.A(dpath_mulcore_ary1_a0_I1_p2_l[21]), .B(dpath_mulcore_b5[0]), .Y(n11373));
INVX1 mul_U6411(.A(n11373), .Y(n356));
AND2X1 mul_U6412(.A(dpath_mulcore_ary1_a0_I1_p1_l[21]), .B(dpath_mulcore_b4[0]), .Y(n11376));
INVX1 mul_U6413(.A(n11376), .Y(n357));
AND2X1 mul_U6414(.A(dpath_mulcore_ary1_a0_I1_p0_l[21]), .B(dpath_mulcore_b3[0]), .Y(n11379));
INVX1 mul_U6415(.A(n11379), .Y(n358));
AND2X1 mul_U6416(.A(dpath_mulcore_ary1_a0_I1_p2_l[20]), .B(dpath_mulcore_b5[0]), .Y(n11382));
INVX1 mul_U6417(.A(n11382), .Y(n359));
AND2X1 mul_U6418(.A(dpath_mulcore_ary1_a0_I1_p1_l[20]), .B(dpath_mulcore_b4[0]), .Y(n11385));
INVX1 mul_U6419(.A(n11385), .Y(n360));
AND2X1 mul_U6420(.A(dpath_mulcore_ary1_a0_I1_p0_l[20]), .B(dpath_mulcore_b3[0]), .Y(n11388));
INVX1 mul_U6421(.A(n11388), .Y(n361));
AND2X1 mul_U6422(.A(dpath_mulcore_ary1_a0_I1_p2_l[19]), .B(dpath_mulcore_b5[0]), .Y(n11391));
INVX1 mul_U6423(.A(n11391), .Y(n362));
AND2X1 mul_U6424(.A(dpath_mulcore_ary1_a0_I1_p1_l[19]), .B(dpath_mulcore_b4[0]), .Y(n11394));
INVX1 mul_U6425(.A(n11394), .Y(n363));
AND2X1 mul_U6426(.A(dpath_mulcore_ary1_a0_I1_p0_l[19]), .B(dpath_mulcore_b3[0]), .Y(n11397));
INVX1 mul_U6427(.A(n11397), .Y(n364));
AND2X1 mul_U6428(.A(dpath_mulcore_ary1_a0_I1_p2_l[18]), .B(dpath_mulcore_b5[0]), .Y(n11400));
INVX1 mul_U6429(.A(n11400), .Y(n365));
AND2X1 mul_U6430(.A(dpath_mulcore_ary1_a0_I1_p1_l[18]), .B(dpath_mulcore_b4[0]), .Y(n11403));
INVX1 mul_U6431(.A(n11403), .Y(n366));
AND2X1 mul_U6432(.A(dpath_mulcore_ary1_a0_I1_p0_l[18]), .B(dpath_mulcore_b3[0]), .Y(n11406));
INVX1 mul_U6433(.A(n11406), .Y(n367));
AND2X1 mul_U6434(.A(dpath_mulcore_ary1_a0_I1_p2_l[17]), .B(dpath_mulcore_b5[0]), .Y(n11409));
INVX1 mul_U6435(.A(n11409), .Y(n368));
AND2X1 mul_U6436(.A(dpath_mulcore_ary1_a0_I1_p1_l[17]), .B(dpath_mulcore_b4[0]), .Y(n11412));
INVX1 mul_U6437(.A(n11412), .Y(n369));
AND2X1 mul_U6438(.A(dpath_mulcore_ary1_a0_I1_p0_l[17]), .B(dpath_mulcore_b3[0]), .Y(n11415));
INVX1 mul_U6439(.A(n11415), .Y(n370));
AND2X1 mul_U6440(.A(dpath_mulcore_ary1_a0_I1_p2_l[16]), .B(dpath_mulcore_b5[0]), .Y(n11418));
INVX1 mul_U6441(.A(n11418), .Y(n371));
AND2X1 mul_U6442(.A(dpath_mulcore_ary1_a0_I1_p1_l[16]), .B(dpath_mulcore_b4[0]), .Y(n11421));
INVX1 mul_U6443(.A(n11421), .Y(n372));
AND2X1 mul_U6444(.A(dpath_mulcore_ary1_a0_I1_p0_l[16]), .B(dpath_mulcore_b3[0]), .Y(n11424));
INVX1 mul_U6445(.A(n11424), .Y(n373));
AND2X1 mul_U6446(.A(dpath_mulcore_ary1_a0_I1_p2_l[15]), .B(dpath_mulcore_b5[0]), .Y(n11427));
INVX1 mul_U6447(.A(n11427), .Y(n374));
AND2X1 mul_U6448(.A(dpath_mulcore_ary1_a0_I1_p1_l[15]), .B(dpath_mulcore_b4[0]), .Y(n11430));
INVX1 mul_U6449(.A(n11430), .Y(n375));
AND2X1 mul_U6450(.A(dpath_mulcore_ary1_a0_I1_p0_l[15]), .B(dpath_mulcore_b3[0]), .Y(n11433));
INVX1 mul_U6451(.A(n11433), .Y(n376));
AND2X1 mul_U6452(.A(dpath_mulcore_ary1_a0_I1_p2_l[14]), .B(dpath_mulcore_b5[0]), .Y(n11436));
INVX1 mul_U6453(.A(n11436), .Y(n377));
AND2X1 mul_U6454(.A(dpath_mulcore_ary1_a0_I1_p1_l[14]), .B(dpath_mulcore_b4[0]), .Y(n11439));
INVX1 mul_U6455(.A(n11439), .Y(n378));
AND2X1 mul_U6456(.A(dpath_mulcore_ary1_a0_I1_p0_l[14]), .B(dpath_mulcore_b3[0]), .Y(n11442));
INVX1 mul_U6457(.A(n11442), .Y(n379));
AND2X1 mul_U6458(.A(dpath_mulcore_ary1_a0_I1_p2_l[13]), .B(dpath_mulcore_b5[0]), .Y(n11445));
INVX1 mul_U6459(.A(n11445), .Y(n380));
AND2X1 mul_U6460(.A(dpath_mulcore_ary1_a0_I1_p1_l[13]), .B(dpath_mulcore_b4[0]), .Y(n11448));
INVX1 mul_U6461(.A(n11448), .Y(n381));
AND2X1 mul_U6462(.A(dpath_mulcore_ary1_a0_I1_p0_l[13]), .B(dpath_mulcore_b3[0]), .Y(n11451));
INVX1 mul_U6463(.A(n11451), .Y(n382));
AND2X1 mul_U6464(.A(dpath_mulcore_ary1_a0_I1_p2_l[12]), .B(dpath_mulcore_b5[0]), .Y(n11454));
INVX1 mul_U6465(.A(n11454), .Y(n383));
AND2X1 mul_U6466(.A(dpath_mulcore_ary1_a0_I1_p1_l[12]), .B(dpath_mulcore_b4[0]), .Y(n11457));
INVX1 mul_U6467(.A(n11457), .Y(n384));
AND2X1 mul_U6468(.A(dpath_mulcore_ary1_a0_I1_p0_l[12]), .B(dpath_mulcore_b3[0]), .Y(n11460));
INVX1 mul_U6469(.A(n11460), .Y(n385));
AND2X1 mul_U6470(.A(dpath_mulcore_ary1_a0_I1_p2_l[11]), .B(dpath_mulcore_b5[0]), .Y(n11463));
INVX1 mul_U6471(.A(n11463), .Y(n386));
AND2X1 mul_U6472(.A(dpath_mulcore_ary1_a0_I1_p1_l[11]), .B(dpath_mulcore_b4[0]), .Y(n11466));
INVX1 mul_U6473(.A(n11466), .Y(n387));
AND2X1 mul_U6474(.A(dpath_mulcore_ary1_a0_I1_p0_l[11]), .B(dpath_mulcore_b3[0]), .Y(n11469));
INVX1 mul_U6475(.A(n11469), .Y(n388));
AND2X1 mul_U6476(.A(dpath_mulcore_ary1_a0_I1_p2_l[10]), .B(dpath_mulcore_b5[0]), .Y(n11472));
INVX1 mul_U6477(.A(n11472), .Y(n389));
AND2X1 mul_U6478(.A(dpath_mulcore_ary1_a0_I1_p1_l[10]), .B(dpath_mulcore_b4[0]), .Y(n11475));
INVX1 mul_U6479(.A(n11475), .Y(n390));
AND2X1 mul_U6480(.A(dpath_mulcore_ary1_a0_I1_p0_l[10]), .B(dpath_mulcore_b3[0]), .Y(n11478));
INVX1 mul_U6481(.A(n11478), .Y(n391));
AND2X1 mul_U6482(.A(dpath_mulcore_ary1_a0_I1_p2_l[9]), .B(dpath_mulcore_b5[0]), .Y(n11481));
INVX1 mul_U6483(.A(n11481), .Y(n392));
AND2X1 mul_U6484(.A(dpath_mulcore_ary1_a0_I1_p1_l[9]), .B(dpath_mulcore_b4[0]), .Y(n11484));
INVX1 mul_U6485(.A(n11484), .Y(n393));
AND2X1 mul_U6486(.A(dpath_mulcore_ary1_a0_I1_p0_l[9]), .B(dpath_mulcore_b3[0]), .Y(n11487));
INVX1 mul_U6487(.A(n11487), .Y(n394));
AND2X1 mul_U6488(.A(dpath_mulcore_ary1_a0_I1_p2_l[8]), .B(dpath_mulcore_b5[0]), .Y(n11490));
INVX1 mul_U6489(.A(n11490), .Y(n395));
AND2X1 mul_U6490(.A(dpath_mulcore_ary1_a0_I1_p1_l[8]), .B(dpath_mulcore_b4[0]), .Y(n11493));
INVX1 mul_U6491(.A(n11493), .Y(n396));
AND2X1 mul_U6492(.A(dpath_mulcore_ary1_a0_I1_p0_l[8]), .B(dpath_mulcore_b3[0]), .Y(n11496));
INVX1 mul_U6493(.A(n11496), .Y(n397));
AND2X1 mul_U6494(.A(dpath_mulcore_ary1_a0_I1_p2_l[7]), .B(dpath_mulcore_b5[0]), .Y(n11499));
INVX1 mul_U6495(.A(n11499), .Y(n398));
AND2X1 mul_U6496(.A(dpath_mulcore_ary1_a0_I1_p1_l[7]), .B(dpath_mulcore_b4[0]), .Y(n11502));
INVX1 mul_U6497(.A(n11502), .Y(n399));
AND2X1 mul_U6498(.A(dpath_mulcore_ary1_a0_I1_p0_l[7]), .B(dpath_mulcore_b3[0]), .Y(n11505));
INVX1 mul_U6499(.A(n11505), .Y(n400));
AND2X1 mul_U6500(.A(dpath_mulcore_ary1_a0_I1_p2_l[6]), .B(dpath_mulcore_b5[0]), .Y(n11508));
INVX1 mul_U6501(.A(n11508), .Y(n401));
AND2X1 mul_U6502(.A(dpath_mulcore_ary1_a0_I1_p1_l[6]), .B(dpath_mulcore_b4[0]), .Y(n11511));
INVX1 mul_U6503(.A(n11511), .Y(n402));
AND2X1 mul_U6504(.A(dpath_mulcore_ary1_a0_I1_p0_l[6]), .B(dpath_mulcore_b3[0]), .Y(n11514));
INVX1 mul_U6505(.A(n11514), .Y(n403));
AND2X1 mul_U6506(.A(dpath_mulcore_ary1_a0_I1_p2_l[5]), .B(dpath_mulcore_b5[0]), .Y(n11517));
INVX1 mul_U6507(.A(n11517), .Y(n404));
AND2X1 mul_U6508(.A(dpath_mulcore_ary1_a0_I1_p1_l[5]), .B(dpath_mulcore_b4[0]), .Y(n11520));
INVX1 mul_U6509(.A(n11520), .Y(n405));
AND2X1 mul_U6510(.A(dpath_mulcore_ary1_a0_I1_p0_l[5]), .B(dpath_mulcore_b3[0]), .Y(n11523));
INVX1 mul_U6511(.A(n11523), .Y(n406));
AND2X1 mul_U6512(.A(dpath_mulcore_ary1_a0_I1_p2_l[4]), .B(dpath_mulcore_b5[0]), .Y(n11526));
INVX1 mul_U6513(.A(n11526), .Y(n407));
AND2X1 mul_U6514(.A(dpath_mulcore_ary1_a0_I1_p1_l[4]), .B(dpath_mulcore_b4[0]), .Y(n11529));
INVX1 mul_U6515(.A(n11529), .Y(n408));
AND2X1 mul_U6516(.A(dpath_mulcore_ary1_a0_I1_p0_l[4]), .B(dpath_mulcore_b3[0]), .Y(n11532));
INVX1 mul_U6517(.A(n11532), .Y(n409));
AND2X1 mul_U6518(.A(dpath_mulcore_ary1_a0_I1_p1_l[3]), .B(dpath_mulcore_b4[0]), .Y(n11537));
INVX1 mul_U6519(.A(n11537), .Y(n410));
AND2X1 mul_U6520(.A(dpath_mulcore_ary1_a0_I1_p0_l[3]), .B(dpath_mulcore_b3[0]), .Y(n11540));
INVX1 mul_U6521(.A(n11540), .Y(n411));
AND2X1 mul_U6522(.A(dpath_mulcore_ary1_a0_I1_I0_p0_l_2), .B(dpath_mulcore_b3[0]), .Y(n11543));
INVX1 mul_U6523(.A(n11543), .Y(n412));
AND2X1 mul_U6524(.A(dpath_mulcore_ary1_a0_I1_I0_p1_l_2), .B(dpath_mulcore_b4[0]), .Y(n11546));
INVX1 mul_U6525(.A(n11546), .Y(n413));
AND2X1 mul_U6526(.A(dpath_mulcore_ary1_a0_I1_I0_p0_l_1), .B(dpath_mulcore_b3[0]), .Y(n11549));
INVX1 mul_U6527(.A(n11549), .Y(n414));
AND2X1 mul_U6528(.A(dpath_mulcore_ary1_a0_I1_I0_p0_l_0), .B(dpath_mulcore_b3[0]), .Y(n11552));
INVX1 mul_U6529(.A(n11552), .Y(n415));
AND2X1 mul_U6530(.A(dpath_mulcore_ary1_a0_I0_I2_p2_l_66), .B(dpath_mulcore_b2[0]), .Y(n11559));
INVX1 mul_U6531(.A(n11559), .Y(n416));
AND2X1 mul_U6532(.A(dpath_mulcore_ary1_a0_I0_I2_p2_l_65), .B(dpath_mulcore_b2[0]), .Y(n11562));
INVX1 mul_U6533(.A(n11562), .Y(n417));
AND2X1 mul_U6534(.A(dpath_mulcore_ary1_a0_I0_I2_p2_l_64), .B(dpath_mulcore_b2[0]), .Y(n11565));
INVX1 mul_U6535(.A(n11565), .Y(n418));
AND2X1 mul_U6536(.A(dpath_mulcore_ary1_a0_I0_I2_p1_l_64), .B(dpath_mulcore_b1[0]), .Y(n11568));
INVX1 mul_U6537(.A(n11568), .Y(n419));
AND2X1 mul_U6538(.A(dpath_mulcore_ary1_a0_I0_p1_l[63]), .B(dpath_mulcore_b1[0]), .Y(n11571));
INVX1 mul_U6539(.A(n11571), .Y(n420));
AND2X1 mul_U6540(.A(dpath_mulcore_ary1_a0_I0_p2_l[63]), .B(dpath_mulcore_b2[0]), .Y(n11574));
INVX1 mul_U6541(.A(n11574), .Y(n421));
AND2X1 mul_U6542(.A(dpath_mulcore_ary1_a0_I0_p2_l[62]), .B(dpath_mulcore_b2[0]), .Y(n11577));
INVX1 mul_U6543(.A(n11577), .Y(n422));
AND2X1 mul_U6544(.A(dpath_mulcore_ary1_a0_I0_p1_l[62]), .B(dpath_mulcore_b1[0]), .Y(n11580));
INVX1 mul_U6545(.A(n11580), .Y(n423));
AND2X1 mul_U6546(.A(dpath_mulcore_ary1_a0_I0_p0_l[62]), .B(dpath_mulcore_b0[0]), .Y(n11583));
INVX1 mul_U6547(.A(n11583), .Y(n424));
AND2X1 mul_U6548(.A(dpath_mulcore_ary1_a0_I0_p2_l[61]), .B(dpath_mulcore_b2[0]), .Y(n11586));
INVX1 mul_U6549(.A(n11586), .Y(n425));
AND2X1 mul_U6550(.A(dpath_mulcore_ary1_a0_I0_p1_l[61]), .B(dpath_mulcore_b1[0]), .Y(n11589));
INVX1 mul_U6551(.A(n11589), .Y(n426));
AND2X1 mul_U6552(.A(dpath_mulcore_ary1_a0_I0_p0_l[61]), .B(dpath_mulcore_b0[0]), .Y(n11592));
INVX1 mul_U6553(.A(n11592), .Y(n427));
AND2X1 mul_U6554(.A(dpath_mulcore_ary1_a0_I0_p2_l[60]), .B(dpath_mulcore_b2[0]), .Y(n11595));
INVX1 mul_U6555(.A(n11595), .Y(n428));
AND2X1 mul_U6556(.A(dpath_mulcore_ary1_a0_I0_p1_l[60]), .B(dpath_mulcore_b1[0]), .Y(n11598));
INVX1 mul_U6557(.A(n11598), .Y(n429));
AND2X1 mul_U6558(.A(dpath_mulcore_ary1_a0_I0_p0_l[60]), .B(dpath_mulcore_b0[0]), .Y(n11601));
INVX1 mul_U6559(.A(n11601), .Y(n430));
AND2X1 mul_U6560(.A(dpath_mulcore_ary1_a0_I0_p2_l[59]), .B(dpath_mulcore_b2[0]), .Y(n11604));
INVX1 mul_U6561(.A(n11604), .Y(n431));
AND2X1 mul_U6562(.A(dpath_mulcore_ary1_a0_I0_p1_l[59]), .B(dpath_mulcore_b1[0]), .Y(n11607));
INVX1 mul_U6563(.A(n11607), .Y(n432));
AND2X1 mul_U6564(.A(dpath_mulcore_ary1_a0_I0_p0_l[59]), .B(dpath_mulcore_b0[0]), .Y(n11610));
INVX1 mul_U6565(.A(n11610), .Y(n433));
AND2X1 mul_U6566(.A(dpath_mulcore_ary1_a0_I0_p2_l[58]), .B(dpath_mulcore_b2[0]), .Y(n11613));
INVX1 mul_U6567(.A(n11613), .Y(n434));
AND2X1 mul_U6568(.A(dpath_mulcore_ary1_a0_I0_p1_l[58]), .B(dpath_mulcore_b1[0]), .Y(n11616));
INVX1 mul_U6569(.A(n11616), .Y(n435));
AND2X1 mul_U6570(.A(dpath_mulcore_ary1_a0_I0_p0_l[58]), .B(dpath_mulcore_b0[0]), .Y(n11619));
INVX1 mul_U6571(.A(n11619), .Y(n436));
AND2X1 mul_U6572(.A(dpath_mulcore_ary1_a0_I0_p2_l[57]), .B(dpath_mulcore_b2[0]), .Y(n11622));
INVX1 mul_U6573(.A(n11622), .Y(n437));
AND2X1 mul_U6574(.A(dpath_mulcore_ary1_a0_I0_p1_l[57]), .B(dpath_mulcore_b1[0]), .Y(n11625));
INVX1 mul_U6575(.A(n11625), .Y(n438));
AND2X1 mul_U6576(.A(dpath_mulcore_ary1_a0_I0_p0_l[57]), .B(dpath_mulcore_b0[0]), .Y(n11628));
INVX1 mul_U6577(.A(n11628), .Y(n439));
AND2X1 mul_U6578(.A(dpath_mulcore_ary1_a0_I0_p2_l[56]), .B(dpath_mulcore_b2[0]), .Y(n11631));
INVX1 mul_U6579(.A(n11631), .Y(n440));
AND2X1 mul_U6580(.A(dpath_mulcore_ary1_a0_I0_p1_l[56]), .B(dpath_mulcore_b1[0]), .Y(n11634));
INVX1 mul_U6581(.A(n11634), .Y(n441));
AND2X1 mul_U6582(.A(dpath_mulcore_ary1_a0_I0_p0_l[56]), .B(dpath_mulcore_b0[0]), .Y(n11637));
INVX1 mul_U6583(.A(n11637), .Y(n442));
AND2X1 mul_U6584(.A(dpath_mulcore_ary1_a0_I0_p2_l[55]), .B(dpath_mulcore_b2[0]), .Y(n11640));
INVX1 mul_U6585(.A(n11640), .Y(n443));
AND2X1 mul_U6586(.A(dpath_mulcore_ary1_a0_I0_p1_l[55]), .B(dpath_mulcore_b1[0]), .Y(n11643));
INVX1 mul_U6587(.A(n11643), .Y(n444));
AND2X1 mul_U6588(.A(dpath_mulcore_ary1_a0_I0_p0_l[55]), .B(dpath_mulcore_b0[0]), .Y(n11646));
INVX1 mul_U6589(.A(n11646), .Y(n445));
AND2X1 mul_U6590(.A(dpath_mulcore_ary1_a0_I0_p2_l[54]), .B(dpath_mulcore_b2[0]), .Y(n11649));
INVX1 mul_U6591(.A(n11649), .Y(n446));
AND2X1 mul_U6592(.A(dpath_mulcore_ary1_a0_I0_p1_l[54]), .B(dpath_mulcore_b1[0]), .Y(n11652));
INVX1 mul_U6593(.A(n11652), .Y(n447));
AND2X1 mul_U6594(.A(dpath_mulcore_ary1_a0_I0_p0_l[54]), .B(dpath_mulcore_b0[0]), .Y(n11655));
INVX1 mul_U6595(.A(n11655), .Y(n448));
AND2X1 mul_U6596(.A(dpath_mulcore_ary1_a0_I0_p2_l[53]), .B(dpath_mulcore_b2[0]), .Y(n11658));
INVX1 mul_U6597(.A(n11658), .Y(n449));
AND2X1 mul_U6598(.A(dpath_mulcore_ary1_a0_I0_p1_l[53]), .B(dpath_mulcore_b1[0]), .Y(n11661));
INVX1 mul_U6599(.A(n11661), .Y(n450));
AND2X1 mul_U6600(.A(dpath_mulcore_ary1_a0_I0_p0_l[53]), .B(dpath_mulcore_b0[0]), .Y(n11664));
INVX1 mul_U6601(.A(n11664), .Y(n451));
AND2X1 mul_U6602(.A(dpath_mulcore_ary1_a0_I0_p2_l[52]), .B(dpath_mulcore_b2[0]), .Y(n11667));
INVX1 mul_U6603(.A(n11667), .Y(n452));
AND2X1 mul_U6604(.A(dpath_mulcore_ary1_a0_I0_p1_l[52]), .B(dpath_mulcore_b1[0]), .Y(n11670));
INVX1 mul_U6605(.A(n11670), .Y(n453));
AND2X1 mul_U6606(.A(dpath_mulcore_ary1_a0_I0_p0_l[52]), .B(dpath_mulcore_b0[0]), .Y(n11673));
INVX1 mul_U6607(.A(n11673), .Y(n454));
AND2X1 mul_U6608(.A(dpath_mulcore_ary1_a0_I0_p2_l[51]), .B(dpath_mulcore_b2[0]), .Y(n11676));
INVX1 mul_U6609(.A(n11676), .Y(n455));
AND2X1 mul_U6610(.A(dpath_mulcore_ary1_a0_I0_p1_l[51]), .B(dpath_mulcore_b1[0]), .Y(n11679));
INVX1 mul_U6611(.A(n11679), .Y(n456));
AND2X1 mul_U6612(.A(dpath_mulcore_ary1_a0_I0_p0_l[51]), .B(dpath_mulcore_b0[0]), .Y(n11682));
INVX1 mul_U6613(.A(n11682), .Y(n457));
AND2X1 mul_U6614(.A(dpath_mulcore_ary1_a0_I0_p2_l[50]), .B(dpath_mulcore_b2[0]), .Y(n11685));
INVX1 mul_U6615(.A(n11685), .Y(n458));
AND2X1 mul_U6616(.A(dpath_mulcore_ary1_a0_I0_p1_l[50]), .B(dpath_mulcore_b1[0]), .Y(n11688));
INVX1 mul_U6617(.A(n11688), .Y(n459));
AND2X1 mul_U6618(.A(dpath_mulcore_ary1_a0_I0_p0_l[50]), .B(dpath_mulcore_b0[0]), .Y(n11691));
INVX1 mul_U6619(.A(n11691), .Y(n460));
AND2X1 mul_U6620(.A(dpath_mulcore_ary1_a0_I0_p2_l[49]), .B(dpath_mulcore_b2[0]), .Y(n11694));
INVX1 mul_U6621(.A(n11694), .Y(n461));
AND2X1 mul_U6622(.A(dpath_mulcore_ary1_a0_I0_p1_l[49]), .B(dpath_mulcore_b1[0]), .Y(n11697));
INVX1 mul_U6623(.A(n11697), .Y(n462));
AND2X1 mul_U6624(.A(dpath_mulcore_ary1_a0_I0_p0_l[49]), .B(dpath_mulcore_b0[0]), .Y(n11700));
INVX1 mul_U6625(.A(n11700), .Y(n463));
AND2X1 mul_U6626(.A(dpath_mulcore_ary1_a0_I0_p2_l[48]), .B(dpath_mulcore_b2[0]), .Y(n11703));
INVX1 mul_U6627(.A(n11703), .Y(n464));
AND2X1 mul_U6628(.A(dpath_mulcore_ary1_a0_I0_p1_l[48]), .B(dpath_mulcore_b1[0]), .Y(n11706));
INVX1 mul_U6629(.A(n11706), .Y(n465));
AND2X1 mul_U6630(.A(dpath_mulcore_ary1_a0_I0_p0_l[48]), .B(dpath_mulcore_b0[0]), .Y(n11709));
INVX1 mul_U6631(.A(n11709), .Y(n466));
AND2X1 mul_U6632(.A(dpath_mulcore_ary1_a0_I0_p2_l[47]), .B(dpath_mulcore_b2[0]), .Y(n11712));
INVX1 mul_U6633(.A(n11712), .Y(n467));
AND2X1 mul_U6634(.A(dpath_mulcore_ary1_a0_I0_p1_l[47]), .B(dpath_mulcore_b1[0]), .Y(n11715));
INVX1 mul_U6635(.A(n11715), .Y(n468));
AND2X1 mul_U6636(.A(dpath_mulcore_ary1_a0_I0_p0_l[47]), .B(dpath_mulcore_b0[0]), .Y(n11718));
INVX1 mul_U6637(.A(n11718), .Y(n469));
AND2X1 mul_U6638(.A(dpath_mulcore_ary1_a0_I0_p2_l[46]), .B(dpath_mulcore_b2[0]), .Y(n11721));
INVX1 mul_U6639(.A(n11721), .Y(n470));
AND2X1 mul_U6640(.A(dpath_mulcore_ary1_a0_I0_p1_l[46]), .B(dpath_mulcore_b1[0]), .Y(n11724));
INVX1 mul_U6641(.A(n11724), .Y(n471));
AND2X1 mul_U6642(.A(dpath_mulcore_ary1_a0_I0_p0_l[46]), .B(dpath_mulcore_b0[0]), .Y(n11727));
INVX1 mul_U6643(.A(n11727), .Y(n472));
AND2X1 mul_U6644(.A(dpath_mulcore_ary1_a0_I0_p2_l[45]), .B(dpath_mulcore_b2[0]), .Y(n11730));
INVX1 mul_U6645(.A(n11730), .Y(n473));
AND2X1 mul_U6646(.A(dpath_mulcore_ary1_a0_I0_p1_l[45]), .B(dpath_mulcore_b1[0]), .Y(n11733));
INVX1 mul_U6647(.A(n11733), .Y(n474));
AND2X1 mul_U6648(.A(dpath_mulcore_ary1_a0_I0_p0_l[45]), .B(dpath_mulcore_b0[0]), .Y(n11736));
INVX1 mul_U6649(.A(n11736), .Y(n475));
AND2X1 mul_U6650(.A(dpath_mulcore_ary1_a0_I0_p2_l[44]), .B(dpath_mulcore_b2[0]), .Y(n11739));
INVX1 mul_U6651(.A(n11739), .Y(n476));
AND2X1 mul_U6652(.A(dpath_mulcore_ary1_a0_I0_p1_l[44]), .B(dpath_mulcore_b1[0]), .Y(n11742));
INVX1 mul_U6653(.A(n11742), .Y(n477));
AND2X1 mul_U6654(.A(dpath_mulcore_ary1_a0_I0_p0_l[44]), .B(dpath_mulcore_b0[0]), .Y(n11745));
INVX1 mul_U6655(.A(n11745), .Y(n478));
AND2X1 mul_U6656(.A(dpath_mulcore_ary1_a0_I0_p2_l[43]), .B(dpath_mulcore_b2[0]), .Y(n11748));
INVX1 mul_U6657(.A(n11748), .Y(n479));
AND2X1 mul_U6658(.A(dpath_mulcore_ary1_a0_I0_p1_l[43]), .B(dpath_mulcore_b1[0]), .Y(n11751));
INVX1 mul_U6659(.A(n11751), .Y(n480));
AND2X1 mul_U6660(.A(dpath_mulcore_ary1_a0_I0_p0_l[43]), .B(dpath_mulcore_b0[0]), .Y(n11754));
INVX1 mul_U6661(.A(n11754), .Y(n481));
AND2X1 mul_U6662(.A(dpath_mulcore_ary1_a0_I0_p2_l[42]), .B(dpath_mulcore_b2[0]), .Y(n11757));
INVX1 mul_U6663(.A(n11757), .Y(n482));
AND2X1 mul_U6664(.A(dpath_mulcore_ary1_a0_I0_p1_l[42]), .B(dpath_mulcore_b1[0]), .Y(n11760));
INVX1 mul_U6665(.A(n11760), .Y(n483));
AND2X1 mul_U6666(.A(dpath_mulcore_ary1_a0_I0_p0_l[42]), .B(dpath_mulcore_b0[0]), .Y(n11763));
INVX1 mul_U6667(.A(n11763), .Y(n484));
AND2X1 mul_U6668(.A(dpath_mulcore_ary1_a0_I0_p2_l[41]), .B(dpath_mulcore_b2[0]), .Y(n11766));
INVX1 mul_U6669(.A(n11766), .Y(n485));
AND2X1 mul_U6670(.A(dpath_mulcore_ary1_a0_I0_p1_l[41]), .B(dpath_mulcore_b1[0]), .Y(n11769));
INVX1 mul_U6671(.A(n11769), .Y(n486));
AND2X1 mul_U6672(.A(dpath_mulcore_ary1_a0_I0_p0_l[41]), .B(dpath_mulcore_b0[0]), .Y(n11772));
INVX1 mul_U6673(.A(n11772), .Y(n487));
AND2X1 mul_U6674(.A(dpath_mulcore_ary1_a0_I0_p2_l[40]), .B(dpath_mulcore_b2[0]), .Y(n11775));
INVX1 mul_U6675(.A(n11775), .Y(n488));
AND2X1 mul_U6676(.A(dpath_mulcore_ary1_a0_I0_p1_l[40]), .B(dpath_mulcore_b1[0]), .Y(n11778));
INVX1 mul_U6677(.A(n11778), .Y(n489));
AND2X1 mul_U6678(.A(dpath_mulcore_ary1_a0_I0_p0_l[40]), .B(dpath_mulcore_b0[0]), .Y(n11781));
INVX1 mul_U6679(.A(n11781), .Y(n490));
AND2X1 mul_U6680(.A(dpath_mulcore_ary1_a0_I0_p2_l[39]), .B(dpath_mulcore_b2[0]), .Y(n11784));
INVX1 mul_U6681(.A(n11784), .Y(n491));
AND2X1 mul_U6682(.A(dpath_mulcore_ary1_a0_I0_p1_l[39]), .B(dpath_mulcore_b1[0]), .Y(n11787));
INVX1 mul_U6683(.A(n11787), .Y(n492));
AND2X1 mul_U6684(.A(dpath_mulcore_ary1_a0_I0_p0_l[39]), .B(dpath_mulcore_b0[0]), .Y(n11790));
INVX1 mul_U6685(.A(n11790), .Y(n493));
AND2X1 mul_U6686(.A(dpath_mulcore_ary1_a0_I0_p2_l[38]), .B(dpath_mulcore_b2[0]), .Y(n11793));
INVX1 mul_U6687(.A(n11793), .Y(n494));
AND2X1 mul_U6688(.A(dpath_mulcore_ary1_a0_I0_p1_l[38]), .B(dpath_mulcore_b1[0]), .Y(n11796));
INVX1 mul_U6689(.A(n11796), .Y(n495));
AND2X1 mul_U6690(.A(dpath_mulcore_ary1_a0_I0_p0_l[38]), .B(dpath_mulcore_b0[0]), .Y(n11799));
INVX1 mul_U6691(.A(n11799), .Y(n496));
AND2X1 mul_U6692(.A(dpath_mulcore_ary1_a0_I0_p2_l[37]), .B(dpath_mulcore_b2[0]), .Y(n11802));
INVX1 mul_U6693(.A(n11802), .Y(n497));
AND2X1 mul_U6694(.A(dpath_mulcore_ary1_a0_I0_p1_l[37]), .B(dpath_mulcore_b1[0]), .Y(n11805));
INVX1 mul_U6695(.A(n11805), .Y(n498));
AND2X1 mul_U6696(.A(dpath_mulcore_ary1_a0_I0_p0_l[37]), .B(dpath_mulcore_b0[0]), .Y(n11808));
INVX1 mul_U6697(.A(n11808), .Y(n499));
AND2X1 mul_U6698(.A(dpath_mulcore_ary1_a0_I0_p2_l[36]), .B(dpath_mulcore_b2[0]), .Y(n11811));
INVX1 mul_U6699(.A(n11811), .Y(n500));
AND2X1 mul_U6700(.A(dpath_mulcore_ary1_a0_I0_p1_l[36]), .B(dpath_mulcore_b1[0]), .Y(n11814));
INVX1 mul_U6701(.A(n11814), .Y(n501));
AND2X1 mul_U6702(.A(dpath_mulcore_ary1_a0_I0_p0_l[36]), .B(dpath_mulcore_b0[0]), .Y(n11817));
INVX1 mul_U6703(.A(n11817), .Y(n502));
AND2X1 mul_U6704(.A(dpath_mulcore_ary1_a0_I0_p2_l[35]), .B(dpath_mulcore_b2[0]), .Y(n11820));
INVX1 mul_U6705(.A(n11820), .Y(n503));
AND2X1 mul_U6706(.A(dpath_mulcore_ary1_a0_I0_p1_l[35]), .B(dpath_mulcore_b1[0]), .Y(n11823));
INVX1 mul_U6707(.A(n11823), .Y(n504));
AND2X1 mul_U6708(.A(dpath_mulcore_ary1_a0_I0_p0_l[35]), .B(dpath_mulcore_b0[0]), .Y(n11826));
INVX1 mul_U6709(.A(n11826), .Y(n505));
AND2X1 mul_U6710(.A(dpath_mulcore_ary1_a0_I0_p2_l[34]), .B(dpath_mulcore_b2[0]), .Y(n11829));
INVX1 mul_U6711(.A(n11829), .Y(n506));
AND2X1 mul_U6712(.A(dpath_mulcore_ary1_a0_I0_p1_l[34]), .B(dpath_mulcore_b1[0]), .Y(n11832));
INVX1 mul_U6713(.A(n11832), .Y(n507));
AND2X1 mul_U6714(.A(dpath_mulcore_ary1_a0_I0_p0_l[34]), .B(dpath_mulcore_b0[0]), .Y(n11835));
INVX1 mul_U6715(.A(n11835), .Y(n508));
AND2X1 mul_U6716(.A(dpath_mulcore_ary1_a0_I0_p2_l[33]), .B(dpath_mulcore_b2[0]), .Y(n11838));
INVX1 mul_U6717(.A(n11838), .Y(n509));
AND2X1 mul_U6718(.A(dpath_mulcore_ary1_a0_I0_p1_l[33]), .B(dpath_mulcore_b1[0]), .Y(n11841));
INVX1 mul_U6719(.A(n11841), .Y(n510));
AND2X1 mul_U6720(.A(dpath_mulcore_ary1_a0_I0_p0_l[33]), .B(dpath_mulcore_b0[0]), .Y(n11844));
INVX1 mul_U6721(.A(n11844), .Y(n511));
AND2X1 mul_U6722(.A(dpath_mulcore_ary1_a0_I0_p2_l[32]), .B(dpath_mulcore_b2[0]), .Y(n11847));
INVX1 mul_U6723(.A(n11847), .Y(n512));
AND2X1 mul_U6724(.A(dpath_mulcore_ary1_a0_I0_p1_l[32]), .B(dpath_mulcore_b1[0]), .Y(n11850));
INVX1 mul_U6725(.A(n11850), .Y(n513));
AND2X1 mul_U6726(.A(dpath_mulcore_ary1_a0_I0_p0_l[32]), .B(dpath_mulcore_b0[0]), .Y(n11853));
INVX1 mul_U6727(.A(n11853), .Y(n514));
AND2X1 mul_U6728(.A(dpath_mulcore_ary1_a0_I0_p2_l[31]), .B(dpath_mulcore_b2[0]), .Y(n11856));
INVX1 mul_U6729(.A(n11856), .Y(n515));
AND2X1 mul_U6730(.A(dpath_mulcore_ary1_a0_I0_p1_l[31]), .B(dpath_mulcore_b1[0]), .Y(n11859));
INVX1 mul_U6731(.A(n11859), .Y(n516));
AND2X1 mul_U6732(.A(dpath_mulcore_ary1_a0_I0_p0_l[31]), .B(dpath_mulcore_b0[0]), .Y(n11862));
INVX1 mul_U6733(.A(n11862), .Y(n517));
AND2X1 mul_U6734(.A(dpath_mulcore_ary1_a0_I0_p2_l[30]), .B(dpath_mulcore_b2[0]), .Y(n11865));
INVX1 mul_U6735(.A(n11865), .Y(n518));
AND2X1 mul_U6736(.A(dpath_mulcore_ary1_a0_I0_p1_l[30]), .B(dpath_mulcore_b1[0]), .Y(n11868));
INVX1 mul_U6737(.A(n11868), .Y(n519));
AND2X1 mul_U6738(.A(dpath_mulcore_ary1_a0_I0_p0_l[30]), .B(dpath_mulcore_b0[0]), .Y(n11871));
INVX1 mul_U6739(.A(n11871), .Y(n520));
AND2X1 mul_U6740(.A(dpath_mulcore_ary1_a0_I0_p2_l[29]), .B(dpath_mulcore_b2[0]), .Y(n11874));
INVX1 mul_U6741(.A(n11874), .Y(n521));
AND2X1 mul_U6742(.A(dpath_mulcore_ary1_a0_I0_p1_l[29]), .B(dpath_mulcore_b1[0]), .Y(n11877));
INVX1 mul_U6743(.A(n11877), .Y(n522));
AND2X1 mul_U6744(.A(dpath_mulcore_ary1_a0_I0_p0_l[29]), .B(dpath_mulcore_b0[0]), .Y(n11880));
INVX1 mul_U6745(.A(n11880), .Y(n523));
AND2X1 mul_U6746(.A(dpath_mulcore_ary1_a0_I0_p2_l[28]), .B(dpath_mulcore_b2[0]), .Y(n11883));
INVX1 mul_U6747(.A(n11883), .Y(n524));
AND2X1 mul_U6748(.A(dpath_mulcore_ary1_a0_I0_p1_l[28]), .B(dpath_mulcore_b1[0]), .Y(n11886));
INVX1 mul_U6749(.A(n11886), .Y(n525));
AND2X1 mul_U6750(.A(dpath_mulcore_ary1_a0_I0_p0_l[28]), .B(dpath_mulcore_b0[0]), .Y(n11889));
INVX1 mul_U6751(.A(n11889), .Y(n526));
AND2X1 mul_U6752(.A(dpath_mulcore_ary1_a0_I0_p2_l[27]), .B(dpath_mulcore_b2[0]), .Y(n11892));
INVX1 mul_U6753(.A(n11892), .Y(n527));
AND2X1 mul_U6754(.A(dpath_mulcore_ary1_a0_I0_p1_l[27]), .B(dpath_mulcore_b1[0]), .Y(n11895));
INVX1 mul_U6755(.A(n11895), .Y(n528));
AND2X1 mul_U6756(.A(dpath_mulcore_ary1_a0_I0_p0_l[27]), .B(dpath_mulcore_b0[0]), .Y(n11898));
INVX1 mul_U6757(.A(n11898), .Y(n529));
AND2X1 mul_U6758(.A(dpath_mulcore_ary1_a0_I0_p2_l[26]), .B(dpath_mulcore_b2[0]), .Y(n11901));
INVX1 mul_U6759(.A(n11901), .Y(n530));
AND2X1 mul_U6760(.A(dpath_mulcore_ary1_a0_I0_p1_l[26]), .B(dpath_mulcore_b1[0]), .Y(n11904));
INVX1 mul_U6761(.A(n11904), .Y(n531));
AND2X1 mul_U6762(.A(dpath_mulcore_ary1_a0_I0_p0_l[26]), .B(dpath_mulcore_b0[0]), .Y(n11907));
INVX1 mul_U6763(.A(n11907), .Y(n532));
AND2X1 mul_U6764(.A(dpath_mulcore_ary1_a0_I0_p2_l[25]), .B(dpath_mulcore_b2[0]), .Y(n11910));
INVX1 mul_U6765(.A(n11910), .Y(n533));
AND2X1 mul_U6766(.A(dpath_mulcore_ary1_a0_I0_p1_l[25]), .B(dpath_mulcore_b1[0]), .Y(n11913));
INVX1 mul_U6767(.A(n11913), .Y(n534));
AND2X1 mul_U6768(.A(dpath_mulcore_ary1_a0_I0_p0_l[25]), .B(dpath_mulcore_b0[0]), .Y(n11916));
INVX1 mul_U6769(.A(n11916), .Y(n535));
AND2X1 mul_U6770(.A(dpath_mulcore_ary1_a0_I0_p2_l[24]), .B(dpath_mulcore_b2[0]), .Y(n11919));
INVX1 mul_U6771(.A(n11919), .Y(n536));
AND2X1 mul_U6772(.A(dpath_mulcore_ary1_a0_I0_p1_l[24]), .B(dpath_mulcore_b1[0]), .Y(n11922));
INVX1 mul_U6773(.A(n11922), .Y(n537));
AND2X1 mul_U6774(.A(dpath_mulcore_ary1_a0_I0_p0_l[24]), .B(dpath_mulcore_b0[0]), .Y(n11925));
INVX1 mul_U6775(.A(n11925), .Y(n538));
AND2X1 mul_U6776(.A(dpath_mulcore_ary1_a0_I0_p2_l[23]), .B(dpath_mulcore_b2[0]), .Y(n11928));
INVX1 mul_U6777(.A(n11928), .Y(n539));
AND2X1 mul_U6778(.A(dpath_mulcore_ary1_a0_I0_p1_l[23]), .B(dpath_mulcore_b1[0]), .Y(n11931));
INVX1 mul_U6779(.A(n11931), .Y(n540));
AND2X1 mul_U6780(.A(dpath_mulcore_ary1_a0_I0_p0_l[23]), .B(dpath_mulcore_b0[0]), .Y(n11934));
INVX1 mul_U6781(.A(n11934), .Y(n541));
AND2X1 mul_U6782(.A(dpath_mulcore_ary1_a0_I0_p2_l[22]), .B(dpath_mulcore_b2[0]), .Y(n11937));
INVX1 mul_U6783(.A(n11937), .Y(n542));
AND2X1 mul_U6784(.A(dpath_mulcore_ary1_a0_I0_p1_l[22]), .B(dpath_mulcore_b1[0]), .Y(n11940));
INVX1 mul_U6785(.A(n11940), .Y(n543));
AND2X1 mul_U6786(.A(dpath_mulcore_ary1_a0_I0_p0_l[22]), .B(dpath_mulcore_b0[0]), .Y(n11943));
INVX1 mul_U6787(.A(n11943), .Y(n544));
AND2X1 mul_U6788(.A(dpath_mulcore_ary1_a0_I0_p2_l[21]), .B(dpath_mulcore_b2[0]), .Y(n11946));
INVX1 mul_U6789(.A(n11946), .Y(n545));
AND2X1 mul_U6790(.A(dpath_mulcore_ary1_a0_I0_p1_l[21]), .B(dpath_mulcore_b1[0]), .Y(n11949));
INVX1 mul_U6791(.A(n11949), .Y(n546));
AND2X1 mul_U6792(.A(dpath_mulcore_ary1_a0_I0_p0_l[21]), .B(dpath_mulcore_b0[0]), .Y(n11952));
INVX1 mul_U6793(.A(n11952), .Y(n547));
AND2X1 mul_U6794(.A(dpath_mulcore_ary1_a0_I0_p2_l[20]), .B(dpath_mulcore_b2[0]), .Y(n11955));
INVX1 mul_U6795(.A(n11955), .Y(n548));
AND2X1 mul_U6796(.A(dpath_mulcore_ary1_a0_I0_p1_l[20]), .B(dpath_mulcore_b1[0]), .Y(n11958));
INVX1 mul_U6797(.A(n11958), .Y(n549));
AND2X1 mul_U6798(.A(dpath_mulcore_ary1_a0_I0_p0_l[20]), .B(dpath_mulcore_b0[0]), .Y(n11961));
INVX1 mul_U6799(.A(n11961), .Y(n550));
AND2X1 mul_U6800(.A(dpath_mulcore_ary1_a0_I0_p2_l[19]), .B(dpath_mulcore_b2[0]), .Y(n11964));
INVX1 mul_U6801(.A(n11964), .Y(n551));
AND2X1 mul_U6802(.A(dpath_mulcore_ary1_a0_I0_p1_l[19]), .B(dpath_mulcore_b1[0]), .Y(n11967));
INVX1 mul_U6803(.A(n11967), .Y(n552));
AND2X1 mul_U6804(.A(dpath_mulcore_ary1_a0_I0_p0_l[19]), .B(dpath_mulcore_b0[0]), .Y(n11970));
INVX1 mul_U6805(.A(n11970), .Y(n553));
AND2X1 mul_U6806(.A(dpath_mulcore_ary1_a0_I0_p2_l[18]), .B(dpath_mulcore_b2[0]), .Y(n11973));
INVX1 mul_U6807(.A(n11973), .Y(n554));
AND2X1 mul_U6808(.A(dpath_mulcore_ary1_a0_I0_p1_l[18]), .B(dpath_mulcore_b1[0]), .Y(n11976));
INVX1 mul_U6809(.A(n11976), .Y(n555));
AND2X1 mul_U6810(.A(dpath_mulcore_ary1_a0_I0_p0_l[18]), .B(dpath_mulcore_b0[0]), .Y(n11979));
INVX1 mul_U6811(.A(n11979), .Y(n556));
AND2X1 mul_U6812(.A(dpath_mulcore_ary1_a0_I0_p2_l[17]), .B(dpath_mulcore_b2[0]), .Y(n11982));
INVX1 mul_U6813(.A(n11982), .Y(n557));
AND2X1 mul_U6814(.A(dpath_mulcore_ary1_a0_I0_p1_l[17]), .B(dpath_mulcore_b1[0]), .Y(n11985));
INVX1 mul_U6815(.A(n11985), .Y(n558));
AND2X1 mul_U6816(.A(dpath_mulcore_ary1_a0_I0_p0_l[17]), .B(dpath_mulcore_b0[0]), .Y(n11988));
INVX1 mul_U6817(.A(n11988), .Y(n559));
AND2X1 mul_U6818(.A(dpath_mulcore_ary1_a0_I0_p2_l[16]), .B(dpath_mulcore_b2[0]), .Y(n11991));
INVX1 mul_U6819(.A(n11991), .Y(n560));
AND2X1 mul_U6820(.A(dpath_mulcore_ary1_a0_I0_p1_l[16]), .B(dpath_mulcore_b1[0]), .Y(n11994));
INVX1 mul_U6821(.A(n11994), .Y(n561));
AND2X1 mul_U6822(.A(dpath_mulcore_ary1_a0_I0_p0_l[16]), .B(dpath_mulcore_b0[0]), .Y(n11997));
INVX1 mul_U6823(.A(n11997), .Y(n562));
AND2X1 mul_U6824(.A(dpath_mulcore_ary1_a0_I0_p2_l[15]), .B(dpath_mulcore_b2[0]), .Y(n12000));
INVX1 mul_U6825(.A(n12000), .Y(n563));
AND2X1 mul_U6826(.A(dpath_mulcore_ary1_a0_I0_p1_l[15]), .B(dpath_mulcore_b1[0]), .Y(n12003));
INVX1 mul_U6827(.A(n12003), .Y(n564));
AND2X1 mul_U6828(.A(dpath_mulcore_ary1_a0_I0_p0_l[15]), .B(dpath_mulcore_b0[0]), .Y(n12006));
INVX1 mul_U6829(.A(n12006), .Y(n565));
AND2X1 mul_U6830(.A(dpath_mulcore_ary1_a0_I0_p2_l[14]), .B(dpath_mulcore_b2[0]), .Y(n12009));
INVX1 mul_U6831(.A(n12009), .Y(n566));
AND2X1 mul_U6832(.A(dpath_mulcore_ary1_a0_I0_p1_l[14]), .B(dpath_mulcore_b1[0]), .Y(n12012));
INVX1 mul_U6833(.A(n12012), .Y(n567));
AND2X1 mul_U6834(.A(dpath_mulcore_ary1_a0_I0_p0_l[14]), .B(dpath_mulcore_b0[0]), .Y(n12015));
INVX1 mul_U6835(.A(n12015), .Y(n568));
AND2X1 mul_U6836(.A(dpath_mulcore_ary1_a0_I0_p2_l[13]), .B(dpath_mulcore_b2[0]), .Y(n12018));
INVX1 mul_U6837(.A(n12018), .Y(n569));
AND2X1 mul_U6838(.A(dpath_mulcore_ary1_a0_I0_p1_l[13]), .B(dpath_mulcore_b1[0]), .Y(n12021));
INVX1 mul_U6839(.A(n12021), .Y(n570));
AND2X1 mul_U6840(.A(dpath_mulcore_ary1_a0_I0_p0_l[13]), .B(dpath_mulcore_b0[0]), .Y(n12024));
INVX1 mul_U6841(.A(n12024), .Y(n571));
AND2X1 mul_U6842(.A(dpath_mulcore_ary1_a0_I0_p2_l[12]), .B(dpath_mulcore_b2[0]), .Y(n12027));
INVX1 mul_U6843(.A(n12027), .Y(n572));
AND2X1 mul_U6844(.A(dpath_mulcore_ary1_a0_I0_p1_l[12]), .B(dpath_mulcore_b1[0]), .Y(n12030));
INVX1 mul_U6845(.A(n12030), .Y(n573));
AND2X1 mul_U6846(.A(dpath_mulcore_ary1_a0_I0_p0_l[12]), .B(dpath_mulcore_b0[0]), .Y(n12033));
INVX1 mul_U6847(.A(n12033), .Y(n574));
AND2X1 mul_U6848(.A(dpath_mulcore_ary1_a0_I0_p2_l[11]), .B(dpath_mulcore_b2[0]), .Y(n12036));
INVX1 mul_U6849(.A(n12036), .Y(n575));
AND2X1 mul_U6850(.A(dpath_mulcore_ary1_a0_I0_p1_l[11]), .B(dpath_mulcore_b1[0]), .Y(n12039));
INVX1 mul_U6851(.A(n12039), .Y(n576));
AND2X1 mul_U6852(.A(dpath_mulcore_ary1_a0_I0_p0_l[11]), .B(dpath_mulcore_b0[0]), .Y(n12042));
INVX1 mul_U6853(.A(n12042), .Y(n577));
AND2X1 mul_U6854(.A(dpath_mulcore_ary1_a0_I0_p2_l[10]), .B(dpath_mulcore_b2[0]), .Y(n12045));
INVX1 mul_U6855(.A(n12045), .Y(n578));
AND2X1 mul_U6856(.A(dpath_mulcore_ary1_a0_I0_p1_l[10]), .B(dpath_mulcore_b1[0]), .Y(n12048));
INVX1 mul_U6857(.A(n12048), .Y(n579));
AND2X1 mul_U6858(.A(dpath_mulcore_ary1_a0_I0_p0_l[10]), .B(dpath_mulcore_b0[0]), .Y(n12051));
INVX1 mul_U6859(.A(n12051), .Y(n580));
AND2X1 mul_U6860(.A(dpath_mulcore_ary1_a0_I0_p2_l[9]), .B(dpath_mulcore_b2[0]), .Y(n12054));
INVX1 mul_U6861(.A(n12054), .Y(n581));
AND2X1 mul_U6862(.A(dpath_mulcore_ary1_a0_I0_p1_l[9]), .B(dpath_mulcore_b1[0]), .Y(n12057));
INVX1 mul_U6863(.A(n12057), .Y(n582));
AND2X1 mul_U6864(.A(dpath_mulcore_ary1_a0_I0_p0_l[9]), .B(dpath_mulcore_b0[0]), .Y(n12060));
INVX1 mul_U6865(.A(n12060), .Y(n583));
AND2X1 mul_U6866(.A(dpath_mulcore_ary1_a0_I0_p2_l[8]), .B(dpath_mulcore_b2[0]), .Y(n12063));
INVX1 mul_U6867(.A(n12063), .Y(n584));
AND2X1 mul_U6868(.A(dpath_mulcore_ary1_a0_I0_p1_l[8]), .B(dpath_mulcore_b1[0]), .Y(n12066));
INVX1 mul_U6869(.A(n12066), .Y(n585));
AND2X1 mul_U6870(.A(dpath_mulcore_ary1_a0_I0_p0_l[8]), .B(dpath_mulcore_b0[0]), .Y(n12069));
INVX1 mul_U6871(.A(n12069), .Y(n586));
AND2X1 mul_U6872(.A(dpath_mulcore_ary1_a0_I0_p2_l[7]), .B(dpath_mulcore_b2[0]), .Y(n12072));
INVX1 mul_U6873(.A(n12072), .Y(n587));
AND2X1 mul_U6874(.A(dpath_mulcore_ary1_a0_I0_p1_l[7]), .B(dpath_mulcore_b1[0]), .Y(n12075));
INVX1 mul_U6875(.A(n12075), .Y(n588));
AND2X1 mul_U6876(.A(dpath_mulcore_ary1_a0_I0_p0_l[7]), .B(dpath_mulcore_b0[0]), .Y(n12078));
INVX1 mul_U6877(.A(n12078), .Y(n589));
AND2X1 mul_U6878(.A(dpath_mulcore_ary1_a0_I0_p2_l[6]), .B(dpath_mulcore_b2[0]), .Y(n12081));
INVX1 mul_U6879(.A(n12081), .Y(n590));
AND2X1 mul_U6880(.A(dpath_mulcore_ary1_a0_I0_p1_l[6]), .B(dpath_mulcore_b1[0]), .Y(n12084));
INVX1 mul_U6881(.A(n12084), .Y(n591));
AND2X1 mul_U6882(.A(dpath_mulcore_ary1_a0_I0_p0_l[6]), .B(dpath_mulcore_b0[0]), .Y(n12087));
INVX1 mul_U6883(.A(n12087), .Y(n592));
AND2X1 mul_U6884(.A(dpath_mulcore_ary1_a0_I0_p2_l[5]), .B(dpath_mulcore_b2[0]), .Y(n12090));
INVX1 mul_U6885(.A(n12090), .Y(n593));
AND2X1 mul_U6886(.A(dpath_mulcore_ary1_a0_I0_p1_l[5]), .B(dpath_mulcore_b1[0]), .Y(n12093));
INVX1 mul_U6887(.A(n12093), .Y(n594));
AND2X1 mul_U6888(.A(dpath_mulcore_ary1_a0_I0_p0_l[5]), .B(dpath_mulcore_b0[0]), .Y(n12096));
INVX1 mul_U6889(.A(n12096), .Y(n595));
AND2X1 mul_U6890(.A(dpath_mulcore_ary1_a0_I0_p2_l[4]), .B(dpath_mulcore_b2[0]), .Y(n12099));
INVX1 mul_U6891(.A(n12099), .Y(n596));
AND2X1 mul_U6892(.A(dpath_mulcore_ary1_a0_I0_p1_l[4]), .B(dpath_mulcore_b1[0]), .Y(n12102));
INVX1 mul_U6893(.A(n12102), .Y(n597));
AND2X1 mul_U6894(.A(dpath_mulcore_ary1_a0_I0_p0_l[4]), .B(dpath_mulcore_b0[0]), .Y(n12105));
INVX1 mul_U6895(.A(n12105), .Y(n598));
AND2X1 mul_U6896(.A(dpath_mulcore_ary1_a0_I0_p1_l[3]), .B(dpath_mulcore_b1[0]), .Y(n12110));
INVX1 mul_U6897(.A(n12110), .Y(n599));
AND2X1 mul_U6898(.A(dpath_mulcore_ary1_a0_I0_p0_l[3]), .B(dpath_mulcore_b0[0]), .Y(n12113));
INVX1 mul_U6899(.A(n12113), .Y(n600));
AND2X1 mul_U6900(.A(dpath_mulcore_ary1_a0_I0_I0_p0_l_2), .B(dpath_mulcore_b0[0]), .Y(n12116));
INVX1 mul_U6901(.A(n12116), .Y(n601));
AND2X1 mul_U6902(.A(dpath_mulcore_ary1_a0_I0_I0_p1_l_2), .B(dpath_mulcore_b1[0]), .Y(n12119));
INVX1 mul_U6903(.A(n12119), .Y(n602));
AND2X1 mul_U6904(.A(dpath_mulcore_ary1_a0_I0_I0_p0_l_1), .B(dpath_mulcore_b0[0]), .Y(n12122));
INVX1 mul_U6905(.A(n12122), .Y(n603));
AND2X1 mul_U6906(.A(dpath_mulcore_ary1_a0_I0_I0_p0_l_0), .B(dpath_mulcore_b0[0]), .Y(n12125));
INVX1 mul_U6907(.A(n12125), .Y(n604));
AND2X1 mul_U6908(.A(dpath_mulcore_ary1_a1_I2_I2_p1_l_64), .B(dpath_mulcore_b15[0]), .Y(n12132));
INVX1 mul_U6909(.A(n12132), .Y(n605));
AND2X1 mul_U6910(.A(dpath_mulcore_ary1_a1_I2_p1_l[63]), .B(dpath_mulcore_b15[0]), .Y(n12135));
INVX1 mul_U6911(.A(n12135), .Y(n606));
AND2X1 mul_U6912(.A(dpath_mulcore_ary1_a1_I2_p1_l[62]), .B(dpath_mulcore_b15[0]), .Y(n12138));
INVX1 mul_U6913(.A(n12138), .Y(n607));
AND2X1 mul_U6914(.A(dpath_mulcore_ary1_a1_I2_p0_l[62]), .B(dpath_mulcore_b14[0]), .Y(n12141));
INVX1 mul_U6915(.A(n12141), .Y(n608));
AND2X1 mul_U6916(.A(dpath_mulcore_ary1_a1_I2_p1_l[61]), .B(dpath_mulcore_b15[0]), .Y(n12144));
INVX1 mul_U6917(.A(n12144), .Y(n609));
AND2X1 mul_U6918(.A(dpath_mulcore_ary1_a1_I2_p0_l[61]), .B(dpath_mulcore_b14[0]), .Y(n12147));
INVX1 mul_U6919(.A(n12147), .Y(n610));
AND2X1 mul_U6920(.A(dpath_mulcore_ary1_a1_I2_p1_l[60]), .B(dpath_mulcore_b15[0]), .Y(n12150));
INVX1 mul_U6921(.A(n12150), .Y(n611));
AND2X1 mul_U6922(.A(dpath_mulcore_ary1_a1_I2_p0_l[60]), .B(dpath_mulcore_b14[0]), .Y(n12153));
INVX1 mul_U6923(.A(n12153), .Y(n612));
AND2X1 mul_U6924(.A(dpath_mulcore_ary1_a1_I2_p1_l[59]), .B(dpath_mulcore_b15[0]), .Y(n12156));
INVX1 mul_U6925(.A(n12156), .Y(n613));
AND2X1 mul_U6926(.A(dpath_mulcore_ary1_a1_I2_p0_l[59]), .B(dpath_mulcore_b14[0]), .Y(n12159));
INVX1 mul_U6927(.A(n12159), .Y(n614));
AND2X1 mul_U6928(.A(dpath_mulcore_ary1_a1_I2_p1_l[58]), .B(dpath_mulcore_b15[0]), .Y(n12162));
INVX1 mul_U6929(.A(n12162), .Y(n615));
AND2X1 mul_U6930(.A(dpath_mulcore_ary1_a1_I2_p0_l[58]), .B(dpath_mulcore_b14[0]), .Y(n12165));
INVX1 mul_U6931(.A(n12165), .Y(n616));
AND2X1 mul_U6932(.A(dpath_mulcore_ary1_a1_I2_p1_l[57]), .B(dpath_mulcore_b15[0]), .Y(n12168));
INVX1 mul_U6933(.A(n12168), .Y(n617));
AND2X1 mul_U6934(.A(dpath_mulcore_ary1_a1_I2_p0_l[57]), .B(dpath_mulcore_b14[0]), .Y(n12171));
INVX1 mul_U6935(.A(n12171), .Y(n618));
AND2X1 mul_U6936(.A(dpath_mulcore_ary1_a1_I2_p1_l[56]), .B(dpath_mulcore_b15[0]), .Y(n12174));
INVX1 mul_U6937(.A(n12174), .Y(n619));
AND2X1 mul_U6938(.A(dpath_mulcore_ary1_a1_I2_p0_l[56]), .B(dpath_mulcore_b14[0]), .Y(n12177));
INVX1 mul_U6939(.A(n12177), .Y(n620));
AND2X1 mul_U6940(.A(dpath_mulcore_ary1_a1_I2_p1_l[55]), .B(dpath_mulcore_b15[0]), .Y(n12180));
INVX1 mul_U6941(.A(n12180), .Y(n621));
AND2X1 mul_U6942(.A(dpath_mulcore_ary1_a1_I2_p0_l[55]), .B(dpath_mulcore_b14[0]), .Y(n12183));
INVX1 mul_U6943(.A(n12183), .Y(n622));
AND2X1 mul_U6944(.A(dpath_mulcore_ary1_a1_I2_p1_l[54]), .B(dpath_mulcore_b15[0]), .Y(n12186));
INVX1 mul_U6945(.A(n12186), .Y(n623));
AND2X1 mul_U6946(.A(dpath_mulcore_ary1_a1_I2_p0_l[54]), .B(dpath_mulcore_b14[0]), .Y(n12189));
INVX1 mul_U6947(.A(n12189), .Y(n624));
AND2X1 mul_U6948(.A(dpath_mulcore_ary1_a1_I2_p1_l[53]), .B(dpath_mulcore_b15[0]), .Y(n12192));
INVX1 mul_U6949(.A(n12192), .Y(n625));
AND2X1 mul_U6950(.A(dpath_mulcore_ary1_a1_I2_p0_l[53]), .B(dpath_mulcore_b14[0]), .Y(n12195));
INVX1 mul_U6951(.A(n12195), .Y(n626));
AND2X1 mul_U6952(.A(dpath_mulcore_ary1_a1_I2_p1_l[52]), .B(dpath_mulcore_b15[0]), .Y(n12198));
INVX1 mul_U6953(.A(n12198), .Y(n627));
AND2X1 mul_U6954(.A(dpath_mulcore_ary1_a1_I2_p0_l[52]), .B(dpath_mulcore_b14[0]), .Y(n12201));
INVX1 mul_U6955(.A(n12201), .Y(n628));
AND2X1 mul_U6956(.A(dpath_mulcore_ary1_a1_I2_p1_l[51]), .B(dpath_mulcore_b15[0]), .Y(n12204));
INVX1 mul_U6957(.A(n12204), .Y(n629));
AND2X1 mul_U6958(.A(dpath_mulcore_ary1_a1_I2_p0_l[51]), .B(dpath_mulcore_b14[0]), .Y(n12207));
INVX1 mul_U6959(.A(n12207), .Y(n630));
AND2X1 mul_U6960(.A(dpath_mulcore_ary1_a1_I2_p1_l[50]), .B(dpath_mulcore_b15[0]), .Y(n12210));
INVX1 mul_U6961(.A(n12210), .Y(n631));
AND2X1 mul_U6962(.A(dpath_mulcore_ary1_a1_I2_p0_l[50]), .B(dpath_mulcore_b14[0]), .Y(n12213));
INVX1 mul_U6963(.A(n12213), .Y(n632));
AND2X1 mul_U6964(.A(dpath_mulcore_ary1_a1_I2_p1_l[49]), .B(dpath_mulcore_b15[0]), .Y(n12216));
INVX1 mul_U6965(.A(n12216), .Y(n633));
AND2X1 mul_U6966(.A(dpath_mulcore_ary1_a1_I2_p0_l[49]), .B(dpath_mulcore_b14[0]), .Y(n12219));
INVX1 mul_U6967(.A(n12219), .Y(n634));
AND2X1 mul_U6968(.A(dpath_mulcore_ary1_a1_I2_p1_l[48]), .B(dpath_mulcore_b15[0]), .Y(n12222));
INVX1 mul_U6969(.A(n12222), .Y(n635));
AND2X1 mul_U6970(.A(dpath_mulcore_ary1_a1_I2_p0_l[48]), .B(dpath_mulcore_b14[0]), .Y(n12225));
INVX1 mul_U6971(.A(n12225), .Y(n636));
AND2X1 mul_U6972(.A(dpath_mulcore_ary1_a1_I2_p1_l[47]), .B(dpath_mulcore_b15[0]), .Y(n12228));
INVX1 mul_U6973(.A(n12228), .Y(n637));
AND2X1 mul_U6974(.A(dpath_mulcore_ary1_a1_I2_p0_l[47]), .B(dpath_mulcore_b14[0]), .Y(n12231));
INVX1 mul_U6975(.A(n12231), .Y(n638));
AND2X1 mul_U6976(.A(dpath_mulcore_ary1_a1_I2_p1_l[46]), .B(dpath_mulcore_b15[0]), .Y(n12234));
INVX1 mul_U6977(.A(n12234), .Y(n639));
AND2X1 mul_U6978(.A(dpath_mulcore_ary1_a1_I2_p0_l[46]), .B(dpath_mulcore_b14[0]), .Y(n12237));
INVX1 mul_U6979(.A(n12237), .Y(n640));
AND2X1 mul_U6980(.A(dpath_mulcore_ary1_a1_I2_p1_l[45]), .B(dpath_mulcore_b15[0]), .Y(n12240));
INVX1 mul_U6981(.A(n12240), .Y(n641));
AND2X1 mul_U6982(.A(dpath_mulcore_ary1_a1_I2_p0_l[45]), .B(dpath_mulcore_b14[0]), .Y(n12243));
INVX1 mul_U6983(.A(n12243), .Y(n642));
AND2X1 mul_U6984(.A(dpath_mulcore_ary1_a1_I2_p1_l[44]), .B(dpath_mulcore_b15[0]), .Y(n12246));
INVX1 mul_U6985(.A(n12246), .Y(n643));
AND2X1 mul_U6986(.A(dpath_mulcore_ary1_a1_I2_p0_l[44]), .B(dpath_mulcore_b14[0]), .Y(n12249));
INVX1 mul_U6987(.A(n12249), .Y(n644));
AND2X1 mul_U6988(.A(dpath_mulcore_ary1_a1_I2_p1_l[43]), .B(dpath_mulcore_b15[0]), .Y(n12252));
INVX1 mul_U6989(.A(n12252), .Y(n645));
AND2X1 mul_U6990(.A(dpath_mulcore_ary1_a1_I2_p0_l[43]), .B(dpath_mulcore_b14[0]), .Y(n12255));
INVX1 mul_U6991(.A(n12255), .Y(n646));
AND2X1 mul_U6992(.A(dpath_mulcore_ary1_a1_I2_p1_l[42]), .B(dpath_mulcore_b15[0]), .Y(n12258));
INVX1 mul_U6993(.A(n12258), .Y(n647));
AND2X1 mul_U6994(.A(dpath_mulcore_ary1_a1_I2_p0_l[42]), .B(dpath_mulcore_b14[0]), .Y(n12261));
INVX1 mul_U6995(.A(n12261), .Y(n648));
AND2X1 mul_U6996(.A(dpath_mulcore_ary1_a1_I2_p1_l[41]), .B(dpath_mulcore_b15[0]), .Y(n12264));
INVX1 mul_U6997(.A(n12264), .Y(n649));
AND2X1 mul_U6998(.A(dpath_mulcore_ary1_a1_I2_p0_l[41]), .B(dpath_mulcore_b14[0]), .Y(n12267));
INVX1 mul_U6999(.A(n12267), .Y(n650));
AND2X1 mul_U7000(.A(dpath_mulcore_ary1_a1_I2_p1_l[40]), .B(dpath_mulcore_b15[0]), .Y(n12270));
INVX1 mul_U7001(.A(n12270), .Y(n651));
AND2X1 mul_U7002(.A(dpath_mulcore_ary1_a1_I2_p0_l[40]), .B(dpath_mulcore_b14[0]), .Y(n12273));
INVX1 mul_U7003(.A(n12273), .Y(n652));
AND2X1 mul_U7004(.A(dpath_mulcore_ary1_a1_I2_p1_l[39]), .B(dpath_mulcore_b15[0]), .Y(n12276));
INVX1 mul_U7005(.A(n12276), .Y(n653));
AND2X1 mul_U7006(.A(dpath_mulcore_ary1_a1_I2_p0_l[39]), .B(dpath_mulcore_b14[0]), .Y(n12279));
INVX1 mul_U7007(.A(n12279), .Y(n654));
AND2X1 mul_U7008(.A(dpath_mulcore_ary1_a1_I2_p1_l[38]), .B(dpath_mulcore_b15[0]), .Y(n12282));
INVX1 mul_U7009(.A(n12282), .Y(n655));
AND2X1 mul_U7010(.A(dpath_mulcore_ary1_a1_I2_p0_l[38]), .B(dpath_mulcore_b14[0]), .Y(n12285));
INVX1 mul_U7011(.A(n12285), .Y(n656));
AND2X1 mul_U7012(.A(dpath_mulcore_ary1_a1_I2_p1_l[37]), .B(dpath_mulcore_b15[0]), .Y(n12288));
INVX1 mul_U7013(.A(n12288), .Y(n657));
AND2X1 mul_U7014(.A(dpath_mulcore_ary1_a1_I2_p0_l[37]), .B(dpath_mulcore_b14[0]), .Y(n12291));
INVX1 mul_U7015(.A(n12291), .Y(n658));
AND2X1 mul_U7016(.A(dpath_mulcore_ary1_a1_I2_p1_l[36]), .B(dpath_mulcore_b15[0]), .Y(n12294));
INVX1 mul_U7017(.A(n12294), .Y(n659));
AND2X1 mul_U7018(.A(dpath_mulcore_ary1_a1_I2_p0_l[36]), .B(dpath_mulcore_b14[0]), .Y(n12297));
INVX1 mul_U7019(.A(n12297), .Y(n660));
AND2X1 mul_U7020(.A(dpath_mulcore_ary1_a1_I2_p1_l[35]), .B(dpath_mulcore_b15[0]), .Y(n12300));
INVX1 mul_U7021(.A(n12300), .Y(n661));
AND2X1 mul_U7022(.A(dpath_mulcore_ary1_a1_I2_p0_l[35]), .B(dpath_mulcore_b14[0]), .Y(n12303));
INVX1 mul_U7023(.A(n12303), .Y(n662));
AND2X1 mul_U7024(.A(dpath_mulcore_ary1_a1_I2_p1_l[34]), .B(dpath_mulcore_b15[0]), .Y(n12306));
INVX1 mul_U7025(.A(n12306), .Y(n663));
AND2X1 mul_U7026(.A(dpath_mulcore_ary1_a1_I2_p0_l[34]), .B(dpath_mulcore_b14[0]), .Y(n12309));
INVX1 mul_U7027(.A(n12309), .Y(n664));
AND2X1 mul_U7028(.A(dpath_mulcore_ary1_a1_I2_p1_l[33]), .B(dpath_mulcore_b15[0]), .Y(n12312));
INVX1 mul_U7029(.A(n12312), .Y(n665));
AND2X1 mul_U7030(.A(dpath_mulcore_ary1_a1_I2_p0_l[33]), .B(dpath_mulcore_b14[0]), .Y(n12315));
INVX1 mul_U7031(.A(n12315), .Y(n666));
AND2X1 mul_U7032(.A(dpath_mulcore_ary1_a1_I2_p1_l[32]), .B(dpath_mulcore_b15[0]), .Y(n12318));
INVX1 mul_U7033(.A(n12318), .Y(n667));
AND2X1 mul_U7034(.A(dpath_mulcore_ary1_a1_I2_p0_l[32]), .B(dpath_mulcore_b14[0]), .Y(n12321));
INVX1 mul_U7035(.A(n12321), .Y(n668));
AND2X1 mul_U7036(.A(dpath_mulcore_ary1_a1_I2_p1_l[31]), .B(dpath_mulcore_b15[0]), .Y(n12324));
INVX1 mul_U7037(.A(n12324), .Y(n669));
AND2X1 mul_U7038(.A(dpath_mulcore_ary1_a1_I2_p0_l[31]), .B(dpath_mulcore_b14[0]), .Y(n12327));
INVX1 mul_U7039(.A(n12327), .Y(n670));
AND2X1 mul_U7040(.A(dpath_mulcore_ary1_a1_I2_p1_l[30]), .B(dpath_mulcore_b15[0]), .Y(n12330));
INVX1 mul_U7041(.A(n12330), .Y(n671));
AND2X1 mul_U7042(.A(dpath_mulcore_ary1_a1_I2_p0_l[30]), .B(dpath_mulcore_b14[0]), .Y(n12333));
INVX1 mul_U7043(.A(n12333), .Y(n672));
AND2X1 mul_U7044(.A(dpath_mulcore_ary1_a1_I2_p1_l[29]), .B(dpath_mulcore_b15[0]), .Y(n12336));
INVX1 mul_U7045(.A(n12336), .Y(n673));
AND2X1 mul_U7046(.A(dpath_mulcore_ary1_a1_I2_p0_l[29]), .B(dpath_mulcore_b14[0]), .Y(n12339));
INVX1 mul_U7047(.A(n12339), .Y(n674));
AND2X1 mul_U7048(.A(dpath_mulcore_ary1_a1_I2_p1_l[28]), .B(dpath_mulcore_b15[0]), .Y(n12342));
INVX1 mul_U7049(.A(n12342), .Y(n675));
AND2X1 mul_U7050(.A(dpath_mulcore_ary1_a1_I2_p0_l[28]), .B(dpath_mulcore_b14[0]), .Y(n12345));
INVX1 mul_U7051(.A(n12345), .Y(n676));
AND2X1 mul_U7052(.A(dpath_mulcore_ary1_a1_I2_p1_l[27]), .B(dpath_mulcore_b15[0]), .Y(n12348));
INVX1 mul_U7053(.A(n12348), .Y(n677));
AND2X1 mul_U7054(.A(dpath_mulcore_ary1_a1_I2_p0_l[27]), .B(dpath_mulcore_b14[0]), .Y(n12351));
INVX1 mul_U7055(.A(n12351), .Y(n678));
AND2X1 mul_U7056(.A(dpath_mulcore_ary1_a1_I2_p1_l[26]), .B(dpath_mulcore_b15[0]), .Y(n12354));
INVX1 mul_U7057(.A(n12354), .Y(n679));
AND2X1 mul_U7058(.A(dpath_mulcore_ary1_a1_I2_p0_l[26]), .B(dpath_mulcore_b14[0]), .Y(n12357));
INVX1 mul_U7059(.A(n12357), .Y(n680));
AND2X1 mul_U7060(.A(dpath_mulcore_ary1_a1_I2_p1_l[25]), .B(dpath_mulcore_b15[0]), .Y(n12360));
INVX1 mul_U7061(.A(n12360), .Y(n681));
AND2X1 mul_U7062(.A(dpath_mulcore_ary1_a1_I2_p0_l[25]), .B(dpath_mulcore_b14[0]), .Y(n12363));
INVX1 mul_U7063(.A(n12363), .Y(n682));
AND2X1 mul_U7064(.A(dpath_mulcore_ary1_a1_I2_p1_l[24]), .B(dpath_mulcore_b15[0]), .Y(n12366));
INVX1 mul_U7065(.A(n12366), .Y(n683));
AND2X1 mul_U7066(.A(dpath_mulcore_ary1_a1_I2_p0_l[24]), .B(dpath_mulcore_b14[0]), .Y(n12369));
INVX1 mul_U7067(.A(n12369), .Y(n684));
AND2X1 mul_U7068(.A(dpath_mulcore_ary1_a1_I2_p1_l[23]), .B(dpath_mulcore_b15[0]), .Y(n12372));
INVX1 mul_U7069(.A(n12372), .Y(n685));
AND2X1 mul_U7070(.A(dpath_mulcore_ary1_a1_I2_p0_l[23]), .B(dpath_mulcore_b14[0]), .Y(n12375));
INVX1 mul_U7071(.A(n12375), .Y(n686));
AND2X1 mul_U7072(.A(dpath_mulcore_ary1_a1_I2_p1_l[22]), .B(dpath_mulcore_b15[0]), .Y(n12378));
INVX1 mul_U7073(.A(n12378), .Y(n687));
AND2X1 mul_U7074(.A(dpath_mulcore_ary1_a1_I2_p0_l[22]), .B(dpath_mulcore_b14[0]), .Y(n12381));
INVX1 mul_U7075(.A(n12381), .Y(n688));
AND2X1 mul_U7076(.A(dpath_mulcore_ary1_a1_I2_p1_l[21]), .B(dpath_mulcore_b15[0]), .Y(n12384));
INVX1 mul_U7077(.A(n12384), .Y(n689));
AND2X1 mul_U7078(.A(dpath_mulcore_ary1_a1_I2_p0_l[21]), .B(dpath_mulcore_b14[0]), .Y(n12387));
INVX1 mul_U7079(.A(n12387), .Y(n690));
AND2X1 mul_U7080(.A(dpath_mulcore_ary1_a1_I2_p1_l[20]), .B(dpath_mulcore_b15[0]), .Y(n12390));
INVX1 mul_U7081(.A(n12390), .Y(n691));
AND2X1 mul_U7082(.A(dpath_mulcore_ary1_a1_I2_p0_l[20]), .B(dpath_mulcore_b14[0]), .Y(n12393));
INVX1 mul_U7083(.A(n12393), .Y(n692));
AND2X1 mul_U7084(.A(dpath_mulcore_ary1_a1_I2_p1_l[19]), .B(dpath_mulcore_b15[0]), .Y(n12396));
INVX1 mul_U7085(.A(n12396), .Y(n693));
AND2X1 mul_U7086(.A(dpath_mulcore_ary1_a1_I2_p0_l[19]), .B(dpath_mulcore_b14[0]), .Y(n12399));
INVX1 mul_U7087(.A(n12399), .Y(n694));
AND2X1 mul_U7088(.A(dpath_mulcore_ary1_a1_I2_p1_l[18]), .B(dpath_mulcore_b15[0]), .Y(n12402));
INVX1 mul_U7089(.A(n12402), .Y(n695));
AND2X1 mul_U7090(.A(dpath_mulcore_ary1_a1_I2_p0_l[18]), .B(dpath_mulcore_b14[0]), .Y(n12405));
INVX1 mul_U7091(.A(n12405), .Y(n696));
AND2X1 mul_U7092(.A(dpath_mulcore_ary1_a1_I2_p1_l[17]), .B(dpath_mulcore_b15[0]), .Y(n12408));
INVX1 mul_U7093(.A(n12408), .Y(n697));
AND2X1 mul_U7094(.A(dpath_mulcore_ary1_a1_I2_p0_l[17]), .B(dpath_mulcore_b14[0]), .Y(n12411));
INVX1 mul_U7095(.A(n12411), .Y(n698));
AND2X1 mul_U7096(.A(dpath_mulcore_ary1_a1_I2_p1_l[16]), .B(dpath_mulcore_b15[0]), .Y(n12414));
INVX1 mul_U7097(.A(n12414), .Y(n699));
AND2X1 mul_U7098(.A(dpath_mulcore_ary1_a1_I2_p0_l[16]), .B(dpath_mulcore_b14[0]), .Y(n12417));
INVX1 mul_U7099(.A(n12417), .Y(n700));
AND2X1 mul_U7100(.A(dpath_mulcore_ary1_a1_I2_p1_l[15]), .B(dpath_mulcore_b15[0]), .Y(n12420));
INVX1 mul_U7101(.A(n12420), .Y(n701));
AND2X1 mul_U7102(.A(dpath_mulcore_ary1_a1_I2_p0_l[15]), .B(dpath_mulcore_b14[0]), .Y(n12423));
INVX1 mul_U7103(.A(n12423), .Y(n702));
AND2X1 mul_U7104(.A(dpath_mulcore_ary1_a1_I2_p1_l[14]), .B(dpath_mulcore_b15[0]), .Y(n12426));
INVX1 mul_U7105(.A(n12426), .Y(n703));
AND2X1 mul_U7106(.A(dpath_mulcore_ary1_a1_I2_p0_l[14]), .B(dpath_mulcore_b14[0]), .Y(n12429));
INVX1 mul_U7107(.A(n12429), .Y(n704));
AND2X1 mul_U7108(.A(dpath_mulcore_ary1_a1_I2_p1_l[13]), .B(dpath_mulcore_b15[0]), .Y(n12432));
INVX1 mul_U7109(.A(n12432), .Y(n705));
AND2X1 mul_U7110(.A(dpath_mulcore_ary1_a1_I2_p0_l[13]), .B(dpath_mulcore_b14[0]), .Y(n12435));
INVX1 mul_U7111(.A(n12435), .Y(n706));
AND2X1 mul_U7112(.A(dpath_mulcore_ary1_a1_I2_p1_l[12]), .B(dpath_mulcore_b15[0]), .Y(n12438));
INVX1 mul_U7113(.A(n12438), .Y(n707));
AND2X1 mul_U7114(.A(dpath_mulcore_ary1_a1_I2_p0_l[12]), .B(dpath_mulcore_b14[0]), .Y(n12441));
INVX1 mul_U7115(.A(n12441), .Y(n708));
AND2X1 mul_U7116(.A(dpath_mulcore_ary1_a1_I2_p1_l[11]), .B(dpath_mulcore_b15[0]), .Y(n12444));
INVX1 mul_U7117(.A(n12444), .Y(n709));
AND2X1 mul_U7118(.A(dpath_mulcore_ary1_a1_I2_p0_l[11]), .B(dpath_mulcore_b14[0]), .Y(n12447));
INVX1 mul_U7119(.A(n12447), .Y(n710));
AND2X1 mul_U7120(.A(dpath_mulcore_ary1_a1_I2_p1_l[10]), .B(dpath_mulcore_b15[0]), .Y(n12450));
INVX1 mul_U7121(.A(n12450), .Y(n711));
AND2X1 mul_U7122(.A(dpath_mulcore_ary1_a1_I2_p0_l[10]), .B(dpath_mulcore_b14[0]), .Y(n12453));
INVX1 mul_U7123(.A(n12453), .Y(n712));
AND2X1 mul_U7124(.A(dpath_mulcore_ary1_a1_I2_p1_l[9]), .B(dpath_mulcore_b15[0]), .Y(n12456));
INVX1 mul_U7125(.A(n12456), .Y(n713));
AND2X1 mul_U7126(.A(dpath_mulcore_ary1_a1_I2_p0_l[9]), .B(dpath_mulcore_b14[0]), .Y(n12459));
INVX1 mul_U7127(.A(n12459), .Y(n714));
AND2X1 mul_U7128(.A(dpath_mulcore_ary1_a1_I2_p1_l[8]), .B(dpath_mulcore_b15[0]), .Y(n12462));
INVX1 mul_U7129(.A(n12462), .Y(n715));
AND2X1 mul_U7130(.A(dpath_mulcore_ary1_a1_I2_p0_l[8]), .B(dpath_mulcore_b14[0]), .Y(n12465));
INVX1 mul_U7131(.A(n12465), .Y(n716));
AND2X1 mul_U7132(.A(dpath_mulcore_ary1_a1_I2_p1_l[7]), .B(dpath_mulcore_b15[0]), .Y(n12468));
INVX1 mul_U7133(.A(n12468), .Y(n717));
AND2X1 mul_U7134(.A(dpath_mulcore_ary1_a1_I2_p0_l[7]), .B(dpath_mulcore_b14[0]), .Y(n12471));
INVX1 mul_U7135(.A(n12471), .Y(n718));
AND2X1 mul_U7136(.A(dpath_mulcore_ary1_a1_I2_p1_l[6]), .B(dpath_mulcore_b15[0]), .Y(n12474));
INVX1 mul_U7137(.A(n12474), .Y(n719));
AND2X1 mul_U7138(.A(dpath_mulcore_ary1_a1_I2_p0_l[6]), .B(dpath_mulcore_b14[0]), .Y(n12477));
INVX1 mul_U7139(.A(n12477), .Y(n720));
AND2X1 mul_U7140(.A(dpath_mulcore_ary1_a1_I2_p1_l[5]), .B(dpath_mulcore_b15[0]), .Y(n12480));
INVX1 mul_U7141(.A(n12480), .Y(n721));
AND2X1 mul_U7142(.A(dpath_mulcore_ary1_a1_I2_p0_l[5]), .B(dpath_mulcore_b14[0]), .Y(n12483));
INVX1 mul_U7143(.A(n12483), .Y(n722));
AND2X1 mul_U7144(.A(dpath_mulcore_ary1_a1_I2_p1_l[4]), .B(dpath_mulcore_b15[0]), .Y(n12486));
INVX1 mul_U7145(.A(n12486), .Y(n723));
AND2X1 mul_U7146(.A(dpath_mulcore_ary1_a1_I2_p0_l[4]), .B(dpath_mulcore_b14[0]), .Y(n12489));
INVX1 mul_U7147(.A(n12489), .Y(n724));
AND2X1 mul_U7148(.A(dpath_mulcore_ary1_a1_I2_p1_l[3]), .B(dpath_mulcore_b15[0]), .Y(n12492));
INVX1 mul_U7149(.A(n12492), .Y(n725));
AND2X1 mul_U7150(.A(dpath_mulcore_ary1_a1_I2_p0_l[3]), .B(dpath_mulcore_b14[0]), .Y(n12495));
INVX1 mul_U7151(.A(n12495), .Y(n726));
AND2X1 mul_U7152(.A(dpath_mulcore_ary1_a1_I2_I0_p0_l_2), .B(dpath_mulcore_b14[0]), .Y(n12498));
INVX1 mul_U7153(.A(n12498), .Y(n727));
AND2X1 mul_U7154(.A(dpath_mulcore_ary1_a1_I2_I0_p1_l_2), .B(dpath_mulcore_b15[0]), .Y(n12501));
INVX1 mul_U7155(.A(n12501), .Y(n728));
AND2X1 mul_U7156(.A(dpath_mulcore_ary1_a1_I2_I0_p0_l_1), .B(dpath_mulcore_b14[0]), .Y(n12504));
INVX1 mul_U7157(.A(n12504), .Y(n729));
AND2X1 mul_U7158(.A(dpath_mulcore_ary1_a1_I2_I0_p0_l_0), .B(dpath_mulcore_b14[0]), .Y(n12507));
INVX1 mul_U7159(.A(n12507), .Y(n730));
AND2X1 mul_U7160(.A(dpath_mulcore_ary1_a1_I1_I2_p2_l_66), .B(dpath_mulcore_b13[0]), .Y(n12514));
INVX1 mul_U7161(.A(n12514), .Y(n731));
AND2X1 mul_U7162(.A(dpath_mulcore_ary1_a1_I1_I2_p2_l_65), .B(dpath_mulcore_b13[0]), .Y(n12517));
INVX1 mul_U7163(.A(n12517), .Y(n732));
AND2X1 mul_U7164(.A(dpath_mulcore_ary1_a1_I1_I2_p2_l_64), .B(dpath_mulcore_b13[0]), .Y(n12520));
INVX1 mul_U7165(.A(n12520), .Y(n733));
AND2X1 mul_U7166(.A(dpath_mulcore_ary1_a1_I1_I2_p1_l_64), .B(dpath_mulcore_b12[0]), .Y(n12523));
INVX1 mul_U7167(.A(n12523), .Y(n734));
AND2X1 mul_U7168(.A(dpath_mulcore_ary1_a1_I1_p1_l[63]), .B(dpath_mulcore_b12[0]), .Y(n12526));
INVX1 mul_U7169(.A(n12526), .Y(n735));
AND2X1 mul_U7170(.A(dpath_mulcore_ary1_a1_I1_p2_l[63]), .B(dpath_mulcore_b13[0]), .Y(n12529));
INVX1 mul_U7171(.A(n12529), .Y(n736));
AND2X1 mul_U7172(.A(dpath_mulcore_ary1_a1_I1_p2_l[62]), .B(dpath_mulcore_b13[0]), .Y(n12532));
INVX1 mul_U7173(.A(n12532), .Y(n737));
AND2X1 mul_U7174(.A(dpath_mulcore_ary1_a1_I1_p1_l[62]), .B(dpath_mulcore_b12[0]), .Y(n12535));
INVX1 mul_U7175(.A(n12535), .Y(n738));
AND2X1 mul_U7176(.A(dpath_mulcore_ary1_a1_I1_p0_l[62]), .B(dpath_mulcore_b11[0]), .Y(n12538));
INVX1 mul_U7177(.A(n12538), .Y(n739));
AND2X1 mul_U7178(.A(dpath_mulcore_ary1_a1_I1_p2_l[61]), .B(dpath_mulcore_b13[0]), .Y(n12541));
INVX1 mul_U7179(.A(n12541), .Y(n740));
AND2X1 mul_U7180(.A(dpath_mulcore_ary1_a1_I1_p1_l[61]), .B(dpath_mulcore_b12[0]), .Y(n12544));
INVX1 mul_U7181(.A(n12544), .Y(n741));
AND2X1 mul_U7182(.A(dpath_mulcore_ary1_a1_I1_p0_l[61]), .B(dpath_mulcore_b11[0]), .Y(n12547));
INVX1 mul_U7183(.A(n12547), .Y(n742));
AND2X1 mul_U7184(.A(dpath_mulcore_ary1_a1_I1_p2_l[60]), .B(dpath_mulcore_b13[0]), .Y(n12550));
INVX1 mul_U7185(.A(n12550), .Y(n743));
AND2X1 mul_U7186(.A(dpath_mulcore_ary1_a1_I1_p1_l[60]), .B(dpath_mulcore_b12[0]), .Y(n12553));
INVX1 mul_U7187(.A(n12553), .Y(n744));
AND2X1 mul_U7188(.A(dpath_mulcore_ary1_a1_I1_p0_l[60]), .B(dpath_mulcore_b11[0]), .Y(n12556));
INVX1 mul_U7189(.A(n12556), .Y(n745));
AND2X1 mul_U7190(.A(dpath_mulcore_ary1_a1_I1_p2_l[59]), .B(dpath_mulcore_b13[0]), .Y(n12559));
INVX1 mul_U7191(.A(n12559), .Y(n746));
AND2X1 mul_U7192(.A(dpath_mulcore_ary1_a1_I1_p1_l[59]), .B(dpath_mulcore_b12[0]), .Y(n12562));
INVX1 mul_U7193(.A(n12562), .Y(n747));
AND2X1 mul_U7194(.A(dpath_mulcore_ary1_a1_I1_p0_l[59]), .B(dpath_mulcore_b11[0]), .Y(n12565));
INVX1 mul_U7195(.A(n12565), .Y(n748));
AND2X1 mul_U7196(.A(dpath_mulcore_ary1_a1_I1_p2_l[58]), .B(dpath_mulcore_b13[0]), .Y(n12568));
INVX1 mul_U7197(.A(n12568), .Y(n749));
AND2X1 mul_U7198(.A(dpath_mulcore_ary1_a1_I1_p1_l[58]), .B(dpath_mulcore_b12[0]), .Y(n12571));
INVX1 mul_U7199(.A(n12571), .Y(n750));
AND2X1 mul_U7200(.A(dpath_mulcore_ary1_a1_I1_p0_l[58]), .B(dpath_mulcore_b11[0]), .Y(n12574));
INVX1 mul_U7201(.A(n12574), .Y(n751));
AND2X1 mul_U7202(.A(dpath_mulcore_ary1_a1_I1_p2_l[57]), .B(dpath_mulcore_b13[0]), .Y(n12577));
INVX1 mul_U7203(.A(n12577), .Y(n752));
AND2X1 mul_U7204(.A(dpath_mulcore_ary1_a1_I1_p1_l[57]), .B(dpath_mulcore_b12[0]), .Y(n12580));
INVX1 mul_U7205(.A(n12580), .Y(n753));
AND2X1 mul_U7206(.A(dpath_mulcore_ary1_a1_I1_p0_l[57]), .B(dpath_mulcore_b11[0]), .Y(n12583));
INVX1 mul_U7207(.A(n12583), .Y(n754));
AND2X1 mul_U7208(.A(dpath_mulcore_ary1_a1_I1_p2_l[56]), .B(dpath_mulcore_b13[0]), .Y(n12586));
INVX1 mul_U7209(.A(n12586), .Y(n755));
AND2X1 mul_U7210(.A(dpath_mulcore_ary1_a1_I1_p1_l[56]), .B(dpath_mulcore_b12[0]), .Y(n12589));
INVX1 mul_U7211(.A(n12589), .Y(n756));
AND2X1 mul_U7212(.A(dpath_mulcore_ary1_a1_I1_p0_l[56]), .B(dpath_mulcore_b11[0]), .Y(n12592));
INVX1 mul_U7213(.A(n12592), .Y(n757));
AND2X1 mul_U7214(.A(dpath_mulcore_ary1_a1_I1_p2_l[55]), .B(dpath_mulcore_b13[0]), .Y(n12595));
INVX1 mul_U7215(.A(n12595), .Y(n758));
AND2X1 mul_U7216(.A(dpath_mulcore_ary1_a1_I1_p1_l[55]), .B(dpath_mulcore_b12[0]), .Y(n12598));
INVX1 mul_U7217(.A(n12598), .Y(n759));
AND2X1 mul_U7218(.A(dpath_mulcore_ary1_a1_I1_p0_l[55]), .B(dpath_mulcore_b11[0]), .Y(n12601));
INVX1 mul_U7219(.A(n12601), .Y(n760));
AND2X1 mul_U7220(.A(dpath_mulcore_ary1_a1_I1_p2_l[54]), .B(dpath_mulcore_b13[0]), .Y(n12604));
INVX1 mul_U7221(.A(n12604), .Y(n761));
AND2X1 mul_U7222(.A(dpath_mulcore_ary1_a1_I1_p1_l[54]), .B(dpath_mulcore_b12[0]), .Y(n12607));
INVX1 mul_U7223(.A(n12607), .Y(n762));
AND2X1 mul_U7224(.A(dpath_mulcore_ary1_a1_I1_p0_l[54]), .B(dpath_mulcore_b11[0]), .Y(n12610));
INVX1 mul_U7225(.A(n12610), .Y(n763));
AND2X1 mul_U7226(.A(dpath_mulcore_ary1_a1_I1_p2_l[53]), .B(dpath_mulcore_b13[0]), .Y(n12613));
INVX1 mul_U7227(.A(n12613), .Y(n764));
AND2X1 mul_U7228(.A(dpath_mulcore_ary1_a1_I1_p1_l[53]), .B(dpath_mulcore_b12[0]), .Y(n12616));
INVX1 mul_U7229(.A(n12616), .Y(n765));
AND2X1 mul_U7230(.A(dpath_mulcore_ary1_a1_I1_p0_l[53]), .B(dpath_mulcore_b11[0]), .Y(n12619));
INVX1 mul_U7231(.A(n12619), .Y(n766));
AND2X1 mul_U7232(.A(dpath_mulcore_ary1_a1_I1_p2_l[52]), .B(dpath_mulcore_b13[0]), .Y(n12622));
INVX1 mul_U7233(.A(n12622), .Y(n767));
AND2X1 mul_U7234(.A(dpath_mulcore_ary1_a1_I1_p1_l[52]), .B(dpath_mulcore_b12[0]), .Y(n12625));
INVX1 mul_U7235(.A(n12625), .Y(n768));
AND2X1 mul_U7236(.A(dpath_mulcore_ary1_a1_I1_p0_l[52]), .B(dpath_mulcore_b11[0]), .Y(n12628));
INVX1 mul_U7237(.A(n12628), .Y(n769));
AND2X1 mul_U7238(.A(dpath_mulcore_ary1_a1_I1_p2_l[51]), .B(dpath_mulcore_b13[0]), .Y(n12631));
INVX1 mul_U7239(.A(n12631), .Y(n770));
AND2X1 mul_U7240(.A(dpath_mulcore_ary1_a1_I1_p1_l[51]), .B(dpath_mulcore_b12[0]), .Y(n12634));
INVX1 mul_U7241(.A(n12634), .Y(n771));
AND2X1 mul_U7242(.A(dpath_mulcore_ary1_a1_I1_p0_l[51]), .B(dpath_mulcore_b11[0]), .Y(n12637));
INVX1 mul_U7243(.A(n12637), .Y(n772));
AND2X1 mul_U7244(.A(dpath_mulcore_ary1_a1_I1_p2_l[50]), .B(dpath_mulcore_b13[0]), .Y(n12640));
INVX1 mul_U7245(.A(n12640), .Y(n773));
AND2X1 mul_U7246(.A(dpath_mulcore_ary1_a1_I1_p1_l[50]), .B(dpath_mulcore_b12[0]), .Y(n12643));
INVX1 mul_U7247(.A(n12643), .Y(n774));
AND2X1 mul_U7248(.A(dpath_mulcore_ary1_a1_I1_p0_l[50]), .B(dpath_mulcore_b11[0]), .Y(n12646));
INVX1 mul_U7249(.A(n12646), .Y(n775));
AND2X1 mul_U7250(.A(dpath_mulcore_ary1_a1_I1_p2_l[49]), .B(dpath_mulcore_b13[0]), .Y(n12649));
INVX1 mul_U7251(.A(n12649), .Y(n776));
AND2X1 mul_U7252(.A(dpath_mulcore_ary1_a1_I1_p1_l[49]), .B(dpath_mulcore_b12[0]), .Y(n12652));
INVX1 mul_U7253(.A(n12652), .Y(n777));
AND2X1 mul_U7254(.A(dpath_mulcore_ary1_a1_I1_p0_l[49]), .B(dpath_mulcore_b11[0]), .Y(n12655));
INVX1 mul_U7255(.A(n12655), .Y(n778));
AND2X1 mul_U7256(.A(dpath_mulcore_ary1_a1_I1_p2_l[48]), .B(dpath_mulcore_b13[0]), .Y(n12658));
INVX1 mul_U7257(.A(n12658), .Y(n779));
AND2X1 mul_U7258(.A(dpath_mulcore_ary1_a1_I1_p1_l[48]), .B(dpath_mulcore_b12[0]), .Y(n12661));
INVX1 mul_U7259(.A(n12661), .Y(n780));
AND2X1 mul_U7260(.A(dpath_mulcore_ary1_a1_I1_p0_l[48]), .B(dpath_mulcore_b11[0]), .Y(n12664));
INVX1 mul_U7261(.A(n12664), .Y(n781));
AND2X1 mul_U7262(.A(dpath_mulcore_ary1_a1_I1_p2_l[47]), .B(dpath_mulcore_b13[0]), .Y(n12667));
INVX1 mul_U7263(.A(n12667), .Y(n782));
AND2X1 mul_U7264(.A(dpath_mulcore_ary1_a1_I1_p1_l[47]), .B(dpath_mulcore_b12[0]), .Y(n12670));
INVX1 mul_U7265(.A(n12670), .Y(n783));
AND2X1 mul_U7266(.A(dpath_mulcore_ary1_a1_I1_p0_l[47]), .B(dpath_mulcore_b11[0]), .Y(n12673));
INVX1 mul_U7267(.A(n12673), .Y(n784));
AND2X1 mul_U7268(.A(dpath_mulcore_ary1_a1_I1_p2_l[46]), .B(dpath_mulcore_b13[0]), .Y(n12676));
INVX1 mul_U7269(.A(n12676), .Y(n785));
AND2X1 mul_U7270(.A(dpath_mulcore_ary1_a1_I1_p1_l[46]), .B(dpath_mulcore_b12[0]), .Y(n12679));
INVX1 mul_U7271(.A(n12679), .Y(n786));
AND2X1 mul_U7272(.A(dpath_mulcore_ary1_a1_I1_p0_l[46]), .B(dpath_mulcore_b11[0]), .Y(n12682));
INVX1 mul_U7273(.A(n12682), .Y(n787));
AND2X1 mul_U7274(.A(dpath_mulcore_ary1_a1_I1_p2_l[45]), .B(dpath_mulcore_b13[0]), .Y(n12685));
INVX1 mul_U7275(.A(n12685), .Y(n788));
AND2X1 mul_U7276(.A(dpath_mulcore_ary1_a1_I1_p1_l[45]), .B(dpath_mulcore_b12[0]), .Y(n12688));
INVX1 mul_U7277(.A(n12688), .Y(n789));
AND2X1 mul_U7278(.A(dpath_mulcore_ary1_a1_I1_p0_l[45]), .B(dpath_mulcore_b11[0]), .Y(n12691));
INVX1 mul_U7279(.A(n12691), .Y(n790));
AND2X1 mul_U7280(.A(dpath_mulcore_ary1_a1_I1_p2_l[44]), .B(dpath_mulcore_b13[0]), .Y(n12694));
INVX1 mul_U7281(.A(n12694), .Y(n791));
AND2X1 mul_U7282(.A(dpath_mulcore_ary1_a1_I1_p1_l[44]), .B(dpath_mulcore_b12[0]), .Y(n12697));
INVX1 mul_U7283(.A(n12697), .Y(n792));
AND2X1 mul_U7284(.A(dpath_mulcore_ary1_a1_I1_p0_l[44]), .B(dpath_mulcore_b11[0]), .Y(n12700));
INVX1 mul_U7285(.A(n12700), .Y(n793));
AND2X1 mul_U7286(.A(dpath_mulcore_ary1_a1_I1_p2_l[43]), .B(dpath_mulcore_b13[0]), .Y(n12703));
INVX1 mul_U7287(.A(n12703), .Y(n794));
AND2X1 mul_U7288(.A(dpath_mulcore_ary1_a1_I1_p1_l[43]), .B(dpath_mulcore_b12[0]), .Y(n12706));
INVX1 mul_U7289(.A(n12706), .Y(n795));
AND2X1 mul_U7290(.A(dpath_mulcore_ary1_a1_I1_p0_l[43]), .B(dpath_mulcore_b11[0]), .Y(n12709));
INVX1 mul_U7291(.A(n12709), .Y(n796));
AND2X1 mul_U7292(.A(dpath_mulcore_ary1_a1_I1_p2_l[42]), .B(dpath_mulcore_b13[0]), .Y(n12712));
INVX1 mul_U7293(.A(n12712), .Y(n797));
AND2X1 mul_U7294(.A(dpath_mulcore_ary1_a1_I1_p1_l[42]), .B(dpath_mulcore_b12[0]), .Y(n12715));
INVX1 mul_U7295(.A(n12715), .Y(n798));
AND2X1 mul_U7296(.A(dpath_mulcore_ary1_a1_I1_p0_l[42]), .B(dpath_mulcore_b11[0]), .Y(n12718));
INVX1 mul_U7297(.A(n12718), .Y(n799));
AND2X1 mul_U7298(.A(dpath_mulcore_ary1_a1_I1_p2_l[41]), .B(dpath_mulcore_b13[0]), .Y(n12721));
INVX1 mul_U7299(.A(n12721), .Y(n800));
AND2X1 mul_U7300(.A(dpath_mulcore_ary1_a1_I1_p1_l[41]), .B(dpath_mulcore_b12[0]), .Y(n12724));
INVX1 mul_U7301(.A(n12724), .Y(n801));
AND2X1 mul_U7302(.A(dpath_mulcore_ary1_a1_I1_p0_l[41]), .B(dpath_mulcore_b11[0]), .Y(n12727));
INVX1 mul_U7303(.A(n12727), .Y(n802));
AND2X1 mul_U7304(.A(dpath_mulcore_ary1_a1_I1_p2_l[40]), .B(dpath_mulcore_b13[0]), .Y(n12730));
INVX1 mul_U7305(.A(n12730), .Y(n803));
AND2X1 mul_U7306(.A(dpath_mulcore_ary1_a1_I1_p1_l[40]), .B(dpath_mulcore_b12[0]), .Y(n12733));
INVX1 mul_U7307(.A(n12733), .Y(n804));
AND2X1 mul_U7308(.A(dpath_mulcore_ary1_a1_I1_p0_l[40]), .B(dpath_mulcore_b11[0]), .Y(n12736));
INVX1 mul_U7309(.A(n12736), .Y(n805));
AND2X1 mul_U7310(.A(dpath_mulcore_ary1_a1_I1_p2_l[39]), .B(dpath_mulcore_b13[0]), .Y(n12739));
INVX1 mul_U7311(.A(n12739), .Y(n806));
AND2X1 mul_U7312(.A(dpath_mulcore_ary1_a1_I1_p1_l[39]), .B(dpath_mulcore_b12[0]), .Y(n12742));
INVX1 mul_U7313(.A(n12742), .Y(n807));
AND2X1 mul_U7314(.A(dpath_mulcore_ary1_a1_I1_p0_l[39]), .B(dpath_mulcore_b11[0]), .Y(n12745));
INVX1 mul_U7315(.A(n12745), .Y(n808));
AND2X1 mul_U7316(.A(dpath_mulcore_ary1_a1_I1_p2_l[38]), .B(dpath_mulcore_b13[0]), .Y(n12748));
INVX1 mul_U7317(.A(n12748), .Y(n809));
AND2X1 mul_U7318(.A(dpath_mulcore_ary1_a1_I1_p1_l[38]), .B(dpath_mulcore_b12[0]), .Y(n12751));
INVX1 mul_U7319(.A(n12751), .Y(n810));
AND2X1 mul_U7320(.A(dpath_mulcore_ary1_a1_I1_p0_l[38]), .B(dpath_mulcore_b11[0]), .Y(n12754));
INVX1 mul_U7321(.A(n12754), .Y(n811));
AND2X1 mul_U7322(.A(dpath_mulcore_ary1_a1_I1_p2_l[37]), .B(dpath_mulcore_b13[0]), .Y(n12757));
INVX1 mul_U7323(.A(n12757), .Y(n812));
AND2X1 mul_U7324(.A(dpath_mulcore_ary1_a1_I1_p1_l[37]), .B(dpath_mulcore_b12[0]), .Y(n12760));
INVX1 mul_U7325(.A(n12760), .Y(n813));
AND2X1 mul_U7326(.A(dpath_mulcore_ary1_a1_I1_p0_l[37]), .B(dpath_mulcore_b11[0]), .Y(n12763));
INVX1 mul_U7327(.A(n12763), .Y(n814));
AND2X1 mul_U7328(.A(dpath_mulcore_ary1_a1_I1_p2_l[36]), .B(dpath_mulcore_b13[0]), .Y(n12766));
INVX1 mul_U7329(.A(n12766), .Y(n815));
AND2X1 mul_U7330(.A(dpath_mulcore_ary1_a1_I1_p1_l[36]), .B(dpath_mulcore_b12[0]), .Y(n12769));
INVX1 mul_U7331(.A(n12769), .Y(n816));
AND2X1 mul_U7332(.A(dpath_mulcore_ary1_a1_I1_p0_l[36]), .B(dpath_mulcore_b11[0]), .Y(n12772));
INVX1 mul_U7333(.A(n12772), .Y(n817));
AND2X1 mul_U7334(.A(dpath_mulcore_ary1_a1_I1_p2_l[35]), .B(dpath_mulcore_b13[0]), .Y(n12775));
INVX1 mul_U7335(.A(n12775), .Y(n818));
AND2X1 mul_U7336(.A(dpath_mulcore_ary1_a1_I1_p1_l[35]), .B(dpath_mulcore_b12[0]), .Y(n12778));
INVX1 mul_U7337(.A(n12778), .Y(n819));
AND2X1 mul_U7338(.A(dpath_mulcore_ary1_a1_I1_p0_l[35]), .B(dpath_mulcore_b11[0]), .Y(n12781));
INVX1 mul_U7339(.A(n12781), .Y(n820));
AND2X1 mul_U7340(.A(dpath_mulcore_ary1_a1_I1_p2_l[34]), .B(dpath_mulcore_b13[0]), .Y(n12784));
INVX1 mul_U7341(.A(n12784), .Y(n821));
AND2X1 mul_U7342(.A(dpath_mulcore_ary1_a1_I1_p1_l[34]), .B(dpath_mulcore_b12[0]), .Y(n12787));
INVX1 mul_U7343(.A(n12787), .Y(n822));
AND2X1 mul_U7344(.A(dpath_mulcore_ary1_a1_I1_p0_l[34]), .B(dpath_mulcore_b11[0]), .Y(n12790));
INVX1 mul_U7345(.A(n12790), .Y(n823));
AND2X1 mul_U7346(.A(dpath_mulcore_ary1_a1_I1_p2_l[33]), .B(dpath_mulcore_b13[0]), .Y(n12793));
INVX1 mul_U7347(.A(n12793), .Y(n824));
AND2X1 mul_U7348(.A(dpath_mulcore_ary1_a1_I1_p1_l[33]), .B(dpath_mulcore_b12[0]), .Y(n12796));
INVX1 mul_U7349(.A(n12796), .Y(n825));
AND2X1 mul_U7350(.A(dpath_mulcore_ary1_a1_I1_p0_l[33]), .B(dpath_mulcore_b11[0]), .Y(n12799));
INVX1 mul_U7351(.A(n12799), .Y(n826));
AND2X1 mul_U7352(.A(dpath_mulcore_ary1_a1_I1_p2_l[32]), .B(dpath_mulcore_b13[0]), .Y(n12802));
INVX1 mul_U7353(.A(n12802), .Y(n827));
AND2X1 mul_U7354(.A(dpath_mulcore_ary1_a1_I1_p1_l[32]), .B(dpath_mulcore_b12[0]), .Y(n12805));
INVX1 mul_U7355(.A(n12805), .Y(n828));
AND2X1 mul_U7356(.A(dpath_mulcore_ary1_a1_I1_p0_l[32]), .B(dpath_mulcore_b11[0]), .Y(n12808));
INVX1 mul_U7357(.A(n12808), .Y(n829));
AND2X1 mul_U7358(.A(dpath_mulcore_ary1_a1_I1_p2_l[31]), .B(dpath_mulcore_b13[0]), .Y(n12811));
INVX1 mul_U7359(.A(n12811), .Y(n830));
AND2X1 mul_U7360(.A(dpath_mulcore_ary1_a1_I1_p1_l[31]), .B(dpath_mulcore_b12[0]), .Y(n12814));
INVX1 mul_U7361(.A(n12814), .Y(n831));
AND2X1 mul_U7362(.A(dpath_mulcore_ary1_a1_I1_p0_l[31]), .B(dpath_mulcore_b11[0]), .Y(n12817));
INVX1 mul_U7363(.A(n12817), .Y(n832));
AND2X1 mul_U7364(.A(dpath_mulcore_ary1_a1_I1_p2_l[30]), .B(dpath_mulcore_b13[0]), .Y(n12820));
INVX1 mul_U7365(.A(n12820), .Y(n833));
AND2X1 mul_U7366(.A(dpath_mulcore_ary1_a1_I1_p1_l[30]), .B(dpath_mulcore_b12[0]), .Y(n12823));
INVX1 mul_U7367(.A(n12823), .Y(n834));
AND2X1 mul_U7368(.A(dpath_mulcore_ary1_a1_I1_p0_l[30]), .B(dpath_mulcore_b11[0]), .Y(n12826));
INVX1 mul_U7369(.A(n12826), .Y(n835));
AND2X1 mul_U7370(.A(dpath_mulcore_ary1_a1_I1_p2_l[29]), .B(dpath_mulcore_b13[0]), .Y(n12829));
INVX1 mul_U7371(.A(n12829), .Y(n836));
AND2X1 mul_U7372(.A(dpath_mulcore_ary1_a1_I1_p1_l[29]), .B(dpath_mulcore_b12[0]), .Y(n12832));
INVX1 mul_U7373(.A(n12832), .Y(n837));
AND2X1 mul_U7374(.A(dpath_mulcore_ary1_a1_I1_p0_l[29]), .B(dpath_mulcore_b11[0]), .Y(n12835));
INVX1 mul_U7375(.A(n12835), .Y(n838));
AND2X1 mul_U7376(.A(dpath_mulcore_ary1_a1_I1_p2_l[28]), .B(dpath_mulcore_b13[0]), .Y(n12838));
INVX1 mul_U7377(.A(n12838), .Y(n839));
AND2X1 mul_U7378(.A(dpath_mulcore_ary1_a1_I1_p1_l[28]), .B(dpath_mulcore_b12[0]), .Y(n12841));
INVX1 mul_U7379(.A(n12841), .Y(n840));
AND2X1 mul_U7380(.A(dpath_mulcore_ary1_a1_I1_p0_l[28]), .B(dpath_mulcore_b11[0]), .Y(n12844));
INVX1 mul_U7381(.A(n12844), .Y(n841));
AND2X1 mul_U7382(.A(dpath_mulcore_ary1_a1_I1_p2_l[27]), .B(dpath_mulcore_b13[0]), .Y(n12847));
INVX1 mul_U7383(.A(n12847), .Y(n842));
AND2X1 mul_U7384(.A(dpath_mulcore_ary1_a1_I1_p1_l[27]), .B(dpath_mulcore_b12[0]), .Y(n12850));
INVX1 mul_U7385(.A(n12850), .Y(n843));
AND2X1 mul_U7386(.A(dpath_mulcore_ary1_a1_I1_p0_l[27]), .B(dpath_mulcore_b11[0]), .Y(n12853));
INVX1 mul_U7387(.A(n12853), .Y(n844));
AND2X1 mul_U7388(.A(dpath_mulcore_ary1_a1_I1_p2_l[26]), .B(dpath_mulcore_b13[0]), .Y(n12856));
INVX1 mul_U7389(.A(n12856), .Y(n845));
AND2X1 mul_U7390(.A(dpath_mulcore_ary1_a1_I1_p1_l[26]), .B(dpath_mulcore_b12[0]), .Y(n12859));
INVX1 mul_U7391(.A(n12859), .Y(n846));
AND2X1 mul_U7392(.A(dpath_mulcore_ary1_a1_I1_p0_l[26]), .B(dpath_mulcore_b11[0]), .Y(n12862));
INVX1 mul_U7393(.A(n12862), .Y(n847));
AND2X1 mul_U7394(.A(dpath_mulcore_ary1_a1_I1_p2_l[25]), .B(dpath_mulcore_b13[0]), .Y(n12865));
INVX1 mul_U7395(.A(n12865), .Y(n848));
AND2X1 mul_U7396(.A(dpath_mulcore_ary1_a1_I1_p1_l[25]), .B(dpath_mulcore_b12[0]), .Y(n12868));
INVX1 mul_U7397(.A(n12868), .Y(n849));
AND2X1 mul_U7398(.A(dpath_mulcore_ary1_a1_I1_p0_l[25]), .B(dpath_mulcore_b11[0]), .Y(n12871));
INVX1 mul_U7399(.A(n12871), .Y(n850));
AND2X1 mul_U7400(.A(dpath_mulcore_ary1_a1_I1_p2_l[24]), .B(dpath_mulcore_b13[0]), .Y(n12874));
INVX1 mul_U7401(.A(n12874), .Y(n851));
AND2X1 mul_U7402(.A(dpath_mulcore_ary1_a1_I1_p1_l[24]), .B(dpath_mulcore_b12[0]), .Y(n12877));
INVX1 mul_U7403(.A(n12877), .Y(n852));
AND2X1 mul_U7404(.A(dpath_mulcore_ary1_a1_I1_p0_l[24]), .B(dpath_mulcore_b11[0]), .Y(n12880));
INVX1 mul_U7405(.A(n12880), .Y(n853));
AND2X1 mul_U7406(.A(dpath_mulcore_ary1_a1_I1_p2_l[23]), .B(dpath_mulcore_b13[0]), .Y(n12883));
INVX1 mul_U7407(.A(n12883), .Y(n854));
AND2X1 mul_U7408(.A(dpath_mulcore_ary1_a1_I1_p1_l[23]), .B(dpath_mulcore_b12[0]), .Y(n12886));
INVX1 mul_U7409(.A(n12886), .Y(n855));
AND2X1 mul_U7410(.A(dpath_mulcore_ary1_a1_I1_p0_l[23]), .B(dpath_mulcore_b11[0]), .Y(n12889));
INVX1 mul_U7411(.A(n12889), .Y(n856));
AND2X1 mul_U7412(.A(dpath_mulcore_ary1_a1_I1_p2_l[22]), .B(dpath_mulcore_b13[0]), .Y(n12892));
INVX1 mul_U7413(.A(n12892), .Y(n857));
AND2X1 mul_U7414(.A(dpath_mulcore_ary1_a1_I1_p1_l[22]), .B(dpath_mulcore_b12[0]), .Y(n12895));
INVX1 mul_U7415(.A(n12895), .Y(n858));
AND2X1 mul_U7416(.A(dpath_mulcore_ary1_a1_I1_p0_l[22]), .B(dpath_mulcore_b11[0]), .Y(n12898));
INVX1 mul_U7417(.A(n12898), .Y(n859));
AND2X1 mul_U7418(.A(dpath_mulcore_ary1_a1_I1_p2_l[21]), .B(dpath_mulcore_b13[0]), .Y(n12901));
INVX1 mul_U7419(.A(n12901), .Y(n860));
AND2X1 mul_U7420(.A(dpath_mulcore_ary1_a1_I1_p1_l[21]), .B(dpath_mulcore_b12[0]), .Y(n12904));
INVX1 mul_U7421(.A(n12904), .Y(n861));
AND2X1 mul_U7422(.A(dpath_mulcore_ary1_a1_I1_p0_l[21]), .B(dpath_mulcore_b11[0]), .Y(n12907));
INVX1 mul_U7423(.A(n12907), .Y(n862));
AND2X1 mul_U7424(.A(dpath_mulcore_ary1_a1_I1_p2_l[20]), .B(dpath_mulcore_b13[0]), .Y(n12910));
INVX1 mul_U7425(.A(n12910), .Y(n863));
AND2X1 mul_U7426(.A(dpath_mulcore_ary1_a1_I1_p1_l[20]), .B(dpath_mulcore_b12[0]), .Y(n12913));
INVX1 mul_U7427(.A(n12913), .Y(n864));
AND2X1 mul_U7428(.A(dpath_mulcore_ary1_a1_I1_p0_l[20]), .B(dpath_mulcore_b11[0]), .Y(n12916));
INVX1 mul_U7429(.A(n12916), .Y(n865));
AND2X1 mul_U7430(.A(dpath_mulcore_ary1_a1_I1_p2_l[19]), .B(dpath_mulcore_b13[0]), .Y(n12919));
INVX1 mul_U7431(.A(n12919), .Y(n866));
AND2X1 mul_U7432(.A(dpath_mulcore_ary1_a1_I1_p1_l[19]), .B(dpath_mulcore_b12[0]), .Y(n12922));
INVX1 mul_U7433(.A(n12922), .Y(n867));
AND2X1 mul_U7434(.A(dpath_mulcore_ary1_a1_I1_p0_l[19]), .B(dpath_mulcore_b11[0]), .Y(n12925));
INVX1 mul_U7435(.A(n12925), .Y(n868));
AND2X1 mul_U7436(.A(dpath_mulcore_ary1_a1_I1_p2_l[18]), .B(dpath_mulcore_b13[0]), .Y(n12928));
INVX1 mul_U7437(.A(n12928), .Y(n869));
AND2X1 mul_U7438(.A(dpath_mulcore_ary1_a1_I1_p1_l[18]), .B(dpath_mulcore_b12[0]), .Y(n12931));
INVX1 mul_U7439(.A(n12931), .Y(n870));
AND2X1 mul_U7440(.A(dpath_mulcore_ary1_a1_I1_p0_l[18]), .B(dpath_mulcore_b11[0]), .Y(n12934));
INVX1 mul_U7441(.A(n12934), .Y(n871));
AND2X1 mul_U7442(.A(dpath_mulcore_ary1_a1_I1_p2_l[17]), .B(dpath_mulcore_b13[0]), .Y(n12937));
INVX1 mul_U7443(.A(n12937), .Y(n872));
AND2X1 mul_U7444(.A(dpath_mulcore_ary1_a1_I1_p1_l[17]), .B(dpath_mulcore_b12[0]), .Y(n12940));
INVX1 mul_U7445(.A(n12940), .Y(n873));
AND2X1 mul_U7446(.A(dpath_mulcore_ary1_a1_I1_p0_l[17]), .B(dpath_mulcore_b11[0]), .Y(n12943));
INVX1 mul_U7447(.A(n12943), .Y(n874));
AND2X1 mul_U7448(.A(dpath_mulcore_ary1_a1_I1_p2_l[16]), .B(dpath_mulcore_b13[0]), .Y(n12946));
INVX1 mul_U7449(.A(n12946), .Y(n875));
AND2X1 mul_U7450(.A(dpath_mulcore_ary1_a1_I1_p1_l[16]), .B(dpath_mulcore_b12[0]), .Y(n12949));
INVX1 mul_U7451(.A(n12949), .Y(n876));
AND2X1 mul_U7452(.A(dpath_mulcore_ary1_a1_I1_p0_l[16]), .B(dpath_mulcore_b11[0]), .Y(n12952));
INVX1 mul_U7453(.A(n12952), .Y(n877));
AND2X1 mul_U7454(.A(dpath_mulcore_ary1_a1_I1_p2_l[15]), .B(dpath_mulcore_b13[0]), .Y(n12955));
INVX1 mul_U7455(.A(n12955), .Y(n878));
AND2X1 mul_U7456(.A(dpath_mulcore_ary1_a1_I1_p1_l[15]), .B(dpath_mulcore_b12[0]), .Y(n12958));
INVX1 mul_U7457(.A(n12958), .Y(n879));
AND2X1 mul_U7458(.A(dpath_mulcore_ary1_a1_I1_p0_l[15]), .B(dpath_mulcore_b11[0]), .Y(n12961));
INVX1 mul_U7459(.A(n12961), .Y(n880));
AND2X1 mul_U7460(.A(dpath_mulcore_ary1_a1_I1_p2_l[14]), .B(dpath_mulcore_b13[0]), .Y(n12964));
INVX1 mul_U7461(.A(n12964), .Y(n881));
AND2X1 mul_U7462(.A(dpath_mulcore_ary1_a1_I1_p1_l[14]), .B(dpath_mulcore_b12[0]), .Y(n12967));
INVX1 mul_U7463(.A(n12967), .Y(n882));
AND2X1 mul_U7464(.A(dpath_mulcore_ary1_a1_I1_p0_l[14]), .B(dpath_mulcore_b11[0]), .Y(n12970));
INVX1 mul_U7465(.A(n12970), .Y(n883));
AND2X1 mul_U7466(.A(dpath_mulcore_ary1_a1_I1_p2_l[13]), .B(dpath_mulcore_b13[0]), .Y(n12973));
INVX1 mul_U7467(.A(n12973), .Y(n884));
AND2X1 mul_U7468(.A(dpath_mulcore_ary1_a1_I1_p1_l[13]), .B(dpath_mulcore_b12[0]), .Y(n12976));
INVX1 mul_U7469(.A(n12976), .Y(n885));
AND2X1 mul_U7470(.A(dpath_mulcore_ary1_a1_I1_p0_l[13]), .B(dpath_mulcore_b11[0]), .Y(n12979));
INVX1 mul_U7471(.A(n12979), .Y(n886));
AND2X1 mul_U7472(.A(dpath_mulcore_ary1_a1_I1_p2_l[12]), .B(dpath_mulcore_b13[0]), .Y(n12982));
INVX1 mul_U7473(.A(n12982), .Y(n887));
AND2X1 mul_U7474(.A(dpath_mulcore_ary1_a1_I1_p1_l[12]), .B(dpath_mulcore_b12[0]), .Y(n12985));
INVX1 mul_U7475(.A(n12985), .Y(n888));
AND2X1 mul_U7476(.A(dpath_mulcore_ary1_a1_I1_p0_l[12]), .B(dpath_mulcore_b11[0]), .Y(n12988));
INVX1 mul_U7477(.A(n12988), .Y(n889));
AND2X1 mul_U7478(.A(dpath_mulcore_ary1_a1_I1_p2_l[11]), .B(dpath_mulcore_b13[0]), .Y(n12991));
INVX1 mul_U7479(.A(n12991), .Y(n890));
AND2X1 mul_U7480(.A(dpath_mulcore_ary1_a1_I1_p1_l[11]), .B(dpath_mulcore_b12[0]), .Y(n12994));
INVX1 mul_U7481(.A(n12994), .Y(n891));
AND2X1 mul_U7482(.A(dpath_mulcore_ary1_a1_I1_p0_l[11]), .B(dpath_mulcore_b11[0]), .Y(n12997));
INVX1 mul_U7483(.A(n12997), .Y(n892));
AND2X1 mul_U7484(.A(dpath_mulcore_ary1_a1_I1_p2_l[10]), .B(dpath_mulcore_b13[0]), .Y(n13000));
INVX1 mul_U7485(.A(n13000), .Y(n893));
AND2X1 mul_U7486(.A(dpath_mulcore_ary1_a1_I1_p1_l[10]), .B(dpath_mulcore_b12[0]), .Y(n13003));
INVX1 mul_U7487(.A(n13003), .Y(n894));
AND2X1 mul_U7488(.A(dpath_mulcore_ary1_a1_I1_p0_l[10]), .B(dpath_mulcore_b11[0]), .Y(n13006));
INVX1 mul_U7489(.A(n13006), .Y(n895));
AND2X1 mul_U7490(.A(dpath_mulcore_ary1_a1_I1_p2_l[9]), .B(dpath_mulcore_b13[0]), .Y(n13009));
INVX1 mul_U7491(.A(n13009), .Y(n896));
AND2X1 mul_U7492(.A(dpath_mulcore_ary1_a1_I1_p1_l[9]), .B(dpath_mulcore_b12[0]), .Y(n13012));
INVX1 mul_U7493(.A(n13012), .Y(n897));
AND2X1 mul_U7494(.A(dpath_mulcore_ary1_a1_I1_p0_l[9]), .B(dpath_mulcore_b11[0]), .Y(n13015));
INVX1 mul_U7495(.A(n13015), .Y(n898));
AND2X1 mul_U7496(.A(dpath_mulcore_ary1_a1_I1_p2_l[8]), .B(dpath_mulcore_b13[0]), .Y(n13018));
INVX1 mul_U7497(.A(n13018), .Y(n899));
AND2X1 mul_U7498(.A(dpath_mulcore_ary1_a1_I1_p1_l[8]), .B(dpath_mulcore_b12[0]), .Y(n13021));
INVX1 mul_U7499(.A(n13021), .Y(n900));
AND2X1 mul_U7500(.A(dpath_mulcore_ary1_a1_I1_p0_l[8]), .B(dpath_mulcore_b11[0]), .Y(n13024));
INVX1 mul_U7501(.A(n13024), .Y(n901));
AND2X1 mul_U7502(.A(dpath_mulcore_ary1_a1_I1_p2_l[7]), .B(dpath_mulcore_b13[0]), .Y(n13027));
INVX1 mul_U7503(.A(n13027), .Y(n902));
AND2X1 mul_U7504(.A(dpath_mulcore_ary1_a1_I1_p1_l[7]), .B(dpath_mulcore_b12[0]), .Y(n13030));
INVX1 mul_U7505(.A(n13030), .Y(n903));
AND2X1 mul_U7506(.A(dpath_mulcore_ary1_a1_I1_p0_l[7]), .B(dpath_mulcore_b11[0]), .Y(n13033));
INVX1 mul_U7507(.A(n13033), .Y(n904));
AND2X1 mul_U7508(.A(dpath_mulcore_ary1_a1_I1_p2_l[6]), .B(dpath_mulcore_b13[0]), .Y(n13036));
INVX1 mul_U7509(.A(n13036), .Y(n905));
AND2X1 mul_U7510(.A(dpath_mulcore_ary1_a1_I1_p1_l[6]), .B(dpath_mulcore_b12[0]), .Y(n13039));
INVX1 mul_U7511(.A(n13039), .Y(n906));
AND2X1 mul_U7512(.A(dpath_mulcore_ary1_a1_I1_p0_l[6]), .B(dpath_mulcore_b11[0]), .Y(n13042));
INVX1 mul_U7513(.A(n13042), .Y(n907));
AND2X1 mul_U7514(.A(dpath_mulcore_ary1_a1_I1_p2_l[5]), .B(dpath_mulcore_b13[0]), .Y(n13045));
INVX1 mul_U7515(.A(n13045), .Y(n908));
AND2X1 mul_U7516(.A(dpath_mulcore_ary1_a1_I1_p1_l[5]), .B(dpath_mulcore_b12[0]), .Y(n13048));
INVX1 mul_U7517(.A(n13048), .Y(n909));
AND2X1 mul_U7518(.A(dpath_mulcore_ary1_a1_I1_p0_l[5]), .B(dpath_mulcore_b11[0]), .Y(n13051));
INVX1 mul_U7519(.A(n13051), .Y(n910));
AND2X1 mul_U7520(.A(dpath_mulcore_ary1_a1_I1_p2_l[4]), .B(dpath_mulcore_b13[0]), .Y(n13054));
INVX1 mul_U7521(.A(n13054), .Y(n911));
AND2X1 mul_U7522(.A(dpath_mulcore_ary1_a1_I1_p1_l[4]), .B(dpath_mulcore_b12[0]), .Y(n13057));
INVX1 mul_U7523(.A(n13057), .Y(n912));
AND2X1 mul_U7524(.A(dpath_mulcore_ary1_a1_I1_p0_l[4]), .B(dpath_mulcore_b11[0]), .Y(n13060));
INVX1 mul_U7525(.A(n13060), .Y(n913));
AND2X1 mul_U7526(.A(dpath_mulcore_ary1_a1_I1_p1_l[3]), .B(dpath_mulcore_b12[0]), .Y(n13065));
INVX1 mul_U7527(.A(n13065), .Y(n914));
AND2X1 mul_U7528(.A(dpath_mulcore_ary1_a1_I1_p0_l[3]), .B(dpath_mulcore_b11[0]), .Y(n13068));
INVX1 mul_U7529(.A(n13068), .Y(n915));
AND2X1 mul_U7530(.A(dpath_mulcore_ary1_a1_I1_I0_p0_l_2), .B(dpath_mulcore_b11[0]), .Y(n13071));
INVX1 mul_U7531(.A(n13071), .Y(n916));
AND2X1 mul_U7532(.A(dpath_mulcore_ary1_a1_I1_I0_p1_l_2), .B(dpath_mulcore_b12[0]), .Y(n13074));
INVX1 mul_U7533(.A(n13074), .Y(n917));
AND2X1 mul_U7534(.A(dpath_mulcore_ary1_a1_I1_I0_p0_l_1), .B(dpath_mulcore_b11[0]), .Y(n13077));
INVX1 mul_U7535(.A(n13077), .Y(n918));
AND2X1 mul_U7536(.A(dpath_mulcore_ary1_a1_I1_I0_p0_l_0), .B(dpath_mulcore_b11[0]), .Y(n13080));
INVX1 mul_U7537(.A(n13080), .Y(n919));
AND2X1 mul_U7538(.A(dpath_mulcore_ary1_a1_I0_I2_p2_l_66), .B(dpath_mulcore_b10[0]), .Y(n13087));
INVX1 mul_U7539(.A(n13087), .Y(n920));
AND2X1 mul_U7540(.A(dpath_mulcore_ary1_a1_I0_I2_p2_l_65), .B(dpath_mulcore_b10[0]), .Y(n13090));
INVX1 mul_U7541(.A(n13090), .Y(n921));
AND2X1 mul_U7542(.A(dpath_mulcore_ary1_a1_I0_I2_p2_l_64), .B(dpath_mulcore_b10[0]), .Y(n13093));
INVX1 mul_U7543(.A(n13093), .Y(n922));
AND2X1 mul_U7544(.A(dpath_mulcore_ary1_a1_I0_I2_p1_l_64), .B(dpath_mulcore_b9[0]), .Y(n13096));
INVX1 mul_U7545(.A(n13096), .Y(n923));
AND2X1 mul_U7546(.A(dpath_mulcore_ary1_a1_I0_p1_l[63]), .B(dpath_mulcore_b9[0]), .Y(n13099));
INVX1 mul_U7547(.A(n13099), .Y(n924));
AND2X1 mul_U7548(.A(dpath_mulcore_ary1_a1_I0_p2_l[63]), .B(dpath_mulcore_b10[0]), .Y(n13102));
INVX1 mul_U7549(.A(n13102), .Y(n925));
AND2X1 mul_U7550(.A(dpath_mulcore_ary1_a1_I0_p2_l[62]), .B(dpath_mulcore_b10[0]), .Y(n13105));
INVX1 mul_U7551(.A(n13105), .Y(n926));
AND2X1 mul_U7552(.A(dpath_mulcore_ary1_a1_I0_p1_l[62]), .B(dpath_mulcore_b9[0]), .Y(n13108));
INVX1 mul_U7553(.A(n13108), .Y(n927));
AND2X1 mul_U7554(.A(dpath_mulcore_ary1_a1_I0_p0_l[62]), .B(dpath_mulcore_b8[0]), .Y(n13111));
INVX1 mul_U7555(.A(n13111), .Y(n928));
AND2X1 mul_U7556(.A(dpath_mulcore_ary1_a1_I0_p2_l[61]), .B(dpath_mulcore_b10[0]), .Y(n13114));
INVX1 mul_U7557(.A(n13114), .Y(n929));
AND2X1 mul_U7558(.A(dpath_mulcore_ary1_a1_I0_p1_l[61]), .B(dpath_mulcore_b9[0]), .Y(n13117));
INVX1 mul_U7559(.A(n13117), .Y(n930));
AND2X1 mul_U7560(.A(dpath_mulcore_ary1_a1_I0_p0_l[61]), .B(dpath_mulcore_b8[0]), .Y(n13120));
INVX1 mul_U7561(.A(n13120), .Y(n931));
AND2X1 mul_U7562(.A(dpath_mulcore_ary1_a1_I0_p2_l[60]), .B(dpath_mulcore_b10[0]), .Y(n13123));
INVX1 mul_U7563(.A(n13123), .Y(n932));
AND2X1 mul_U7564(.A(dpath_mulcore_ary1_a1_I0_p1_l[60]), .B(dpath_mulcore_b9[0]), .Y(n13126));
INVX1 mul_U7565(.A(n13126), .Y(n933));
AND2X1 mul_U7566(.A(dpath_mulcore_ary1_a1_I0_p0_l[60]), .B(dpath_mulcore_b8[0]), .Y(n13129));
INVX1 mul_U7567(.A(n13129), .Y(n934));
AND2X1 mul_U7568(.A(dpath_mulcore_ary1_a1_I0_p2_l[59]), .B(dpath_mulcore_b10[0]), .Y(n13132));
INVX1 mul_U7569(.A(n13132), .Y(n935));
AND2X1 mul_U7570(.A(dpath_mulcore_ary1_a1_I0_p1_l[59]), .B(dpath_mulcore_b9[0]), .Y(n13135));
INVX1 mul_U7571(.A(n13135), .Y(n936));
AND2X1 mul_U7572(.A(dpath_mulcore_ary1_a1_I0_p0_l[59]), .B(dpath_mulcore_b8[0]), .Y(n13138));
INVX1 mul_U7573(.A(n13138), .Y(n937));
AND2X1 mul_U7574(.A(dpath_mulcore_ary1_a1_I0_p2_l[58]), .B(dpath_mulcore_b10[0]), .Y(n13141));
INVX1 mul_U7575(.A(n13141), .Y(n938));
AND2X1 mul_U7576(.A(dpath_mulcore_ary1_a1_I0_p1_l[58]), .B(dpath_mulcore_b9[0]), .Y(n13144));
INVX1 mul_U7577(.A(n13144), .Y(n939));
AND2X1 mul_U7578(.A(dpath_mulcore_ary1_a1_I0_p0_l[58]), .B(dpath_mulcore_b8[0]), .Y(n13147));
INVX1 mul_U7579(.A(n13147), .Y(n940));
AND2X1 mul_U7580(.A(dpath_mulcore_ary1_a1_I0_p2_l[57]), .B(dpath_mulcore_b10[0]), .Y(n13150));
INVX1 mul_U7581(.A(n13150), .Y(n941));
AND2X1 mul_U7582(.A(dpath_mulcore_ary1_a1_I0_p1_l[57]), .B(dpath_mulcore_b9[0]), .Y(n13153));
INVX1 mul_U7583(.A(n13153), .Y(n942));
AND2X1 mul_U7584(.A(dpath_mulcore_ary1_a1_I0_p0_l[57]), .B(dpath_mulcore_b8[0]), .Y(n13156));
INVX1 mul_U7585(.A(n13156), .Y(n943));
AND2X1 mul_U7586(.A(dpath_mulcore_ary1_a1_I0_p2_l[56]), .B(dpath_mulcore_b10[0]), .Y(n13159));
INVX1 mul_U7587(.A(n13159), .Y(n944));
AND2X1 mul_U7588(.A(dpath_mulcore_ary1_a1_I0_p1_l[56]), .B(dpath_mulcore_b9[0]), .Y(n13162));
INVX1 mul_U7589(.A(n13162), .Y(n945));
AND2X1 mul_U7590(.A(dpath_mulcore_ary1_a1_I0_p0_l[56]), .B(dpath_mulcore_b8[0]), .Y(n13165));
INVX1 mul_U7591(.A(n13165), .Y(n946));
AND2X1 mul_U7592(.A(dpath_mulcore_ary1_a1_I0_p2_l[55]), .B(dpath_mulcore_b10[0]), .Y(n13168));
INVX1 mul_U7593(.A(n13168), .Y(n947));
AND2X1 mul_U7594(.A(dpath_mulcore_ary1_a1_I0_p1_l[55]), .B(dpath_mulcore_b9[0]), .Y(n13171));
INVX1 mul_U7595(.A(n13171), .Y(n948));
AND2X1 mul_U7596(.A(dpath_mulcore_ary1_a1_I0_p0_l[55]), .B(dpath_mulcore_b8[0]), .Y(n13174));
INVX1 mul_U7597(.A(n13174), .Y(n949));
AND2X1 mul_U7598(.A(dpath_mulcore_ary1_a1_I0_p2_l[54]), .B(dpath_mulcore_b10[0]), .Y(n13177));
INVX1 mul_U7599(.A(n13177), .Y(n950));
AND2X1 mul_U7600(.A(dpath_mulcore_ary1_a1_I0_p1_l[54]), .B(dpath_mulcore_b9[0]), .Y(n13180));
INVX1 mul_U7601(.A(n13180), .Y(n951));
AND2X1 mul_U7602(.A(dpath_mulcore_ary1_a1_I0_p0_l[54]), .B(dpath_mulcore_b8[0]), .Y(n13183));
INVX1 mul_U7603(.A(n13183), .Y(n952));
AND2X1 mul_U7604(.A(dpath_mulcore_ary1_a1_I0_p2_l[53]), .B(dpath_mulcore_b10[0]), .Y(n13186));
INVX1 mul_U7605(.A(n13186), .Y(n953));
AND2X1 mul_U7606(.A(dpath_mulcore_ary1_a1_I0_p1_l[53]), .B(dpath_mulcore_b9[0]), .Y(n13189));
INVX1 mul_U7607(.A(n13189), .Y(n954));
AND2X1 mul_U7608(.A(dpath_mulcore_ary1_a1_I0_p0_l[53]), .B(dpath_mulcore_b8[0]), .Y(n13192));
INVX1 mul_U7609(.A(n13192), .Y(n955));
AND2X1 mul_U7610(.A(dpath_mulcore_ary1_a1_I0_p2_l[52]), .B(dpath_mulcore_b10[0]), .Y(n13195));
INVX1 mul_U7611(.A(n13195), .Y(n956));
AND2X1 mul_U7612(.A(dpath_mulcore_ary1_a1_I0_p1_l[52]), .B(dpath_mulcore_b9[0]), .Y(n13198));
INVX1 mul_U7613(.A(n13198), .Y(n957));
AND2X1 mul_U7614(.A(dpath_mulcore_ary1_a1_I0_p0_l[52]), .B(dpath_mulcore_b8[0]), .Y(n13201));
INVX1 mul_U7615(.A(n13201), .Y(n958));
AND2X1 mul_U7616(.A(dpath_mulcore_ary1_a1_I0_p2_l[51]), .B(dpath_mulcore_b10[0]), .Y(n13204));
INVX1 mul_U7617(.A(n13204), .Y(n959));
AND2X1 mul_U7618(.A(dpath_mulcore_ary1_a1_I0_p1_l[51]), .B(dpath_mulcore_b9[0]), .Y(n13207));
INVX1 mul_U7619(.A(n13207), .Y(n960));
AND2X1 mul_U7620(.A(dpath_mulcore_ary1_a1_I0_p0_l[51]), .B(dpath_mulcore_b8[0]), .Y(n13210));
INVX1 mul_U7621(.A(n13210), .Y(n961));
AND2X1 mul_U7622(.A(dpath_mulcore_ary1_a1_I0_p2_l[50]), .B(dpath_mulcore_b10[0]), .Y(n13213));
INVX1 mul_U7623(.A(n13213), .Y(n962));
AND2X1 mul_U7624(.A(dpath_mulcore_ary1_a1_I0_p1_l[50]), .B(dpath_mulcore_b9[0]), .Y(n13216));
INVX1 mul_U7625(.A(n13216), .Y(n963));
AND2X1 mul_U7626(.A(dpath_mulcore_ary1_a1_I0_p0_l[50]), .B(dpath_mulcore_b8[0]), .Y(n13219));
INVX1 mul_U7627(.A(n13219), .Y(n964));
AND2X1 mul_U7628(.A(dpath_mulcore_ary1_a1_I0_p2_l[49]), .B(dpath_mulcore_b10[0]), .Y(n13222));
INVX1 mul_U7629(.A(n13222), .Y(n965));
AND2X1 mul_U7630(.A(dpath_mulcore_ary1_a1_I0_p1_l[49]), .B(dpath_mulcore_b9[0]), .Y(n13225));
INVX1 mul_U7631(.A(n13225), .Y(n966));
AND2X1 mul_U7632(.A(dpath_mulcore_ary1_a1_I0_p0_l[49]), .B(dpath_mulcore_b8[0]), .Y(n13228));
INVX1 mul_U7633(.A(n13228), .Y(n967));
AND2X1 mul_U7634(.A(dpath_mulcore_ary1_a1_I0_p2_l[48]), .B(dpath_mulcore_b10[0]), .Y(n13231));
INVX1 mul_U7635(.A(n13231), .Y(n968));
AND2X1 mul_U7636(.A(dpath_mulcore_ary1_a1_I0_p1_l[48]), .B(dpath_mulcore_b9[0]), .Y(n13234));
INVX1 mul_U7637(.A(n13234), .Y(n969));
AND2X1 mul_U7638(.A(dpath_mulcore_ary1_a1_I0_p0_l[48]), .B(dpath_mulcore_b8[0]), .Y(n13237));
INVX1 mul_U7639(.A(n13237), .Y(n970));
AND2X1 mul_U7640(.A(dpath_mulcore_ary1_a1_I0_p2_l[47]), .B(dpath_mulcore_b10[0]), .Y(n13240));
INVX1 mul_U7641(.A(n13240), .Y(n971));
AND2X1 mul_U7642(.A(dpath_mulcore_ary1_a1_I0_p1_l[47]), .B(dpath_mulcore_b9[0]), .Y(n13243));
INVX1 mul_U7643(.A(n13243), .Y(n972));
AND2X1 mul_U7644(.A(dpath_mulcore_ary1_a1_I0_p0_l[47]), .B(dpath_mulcore_b8[0]), .Y(n13246));
INVX1 mul_U7645(.A(n13246), .Y(n973));
AND2X1 mul_U7646(.A(dpath_mulcore_ary1_a1_I0_p2_l[46]), .B(dpath_mulcore_b10[0]), .Y(n13249));
INVX1 mul_U7647(.A(n13249), .Y(n974));
AND2X1 mul_U7648(.A(dpath_mulcore_ary1_a1_I0_p1_l[46]), .B(dpath_mulcore_b9[0]), .Y(n13252));
INVX1 mul_U7649(.A(n13252), .Y(n975));
AND2X1 mul_U7650(.A(dpath_mulcore_ary1_a1_I0_p0_l[46]), .B(dpath_mulcore_b8[0]), .Y(n13255));
INVX1 mul_U7651(.A(n13255), .Y(n976));
AND2X1 mul_U7652(.A(dpath_mulcore_ary1_a1_I0_p2_l[45]), .B(dpath_mulcore_b10[0]), .Y(n13258));
INVX1 mul_U7653(.A(n13258), .Y(n977));
AND2X1 mul_U7654(.A(dpath_mulcore_ary1_a1_I0_p1_l[45]), .B(dpath_mulcore_b9[0]), .Y(n13261));
INVX1 mul_U7655(.A(n13261), .Y(n978));
AND2X1 mul_U7656(.A(dpath_mulcore_ary1_a1_I0_p0_l[45]), .B(dpath_mulcore_b8[0]), .Y(n13264));
INVX1 mul_U7657(.A(n13264), .Y(n979));
AND2X1 mul_U7658(.A(dpath_mulcore_ary1_a1_I0_p2_l[44]), .B(dpath_mulcore_b10[0]), .Y(n13267));
INVX1 mul_U7659(.A(n13267), .Y(n980));
AND2X1 mul_U7660(.A(dpath_mulcore_ary1_a1_I0_p1_l[44]), .B(dpath_mulcore_b9[0]), .Y(n13270));
INVX1 mul_U7661(.A(n13270), .Y(n981));
AND2X1 mul_U7662(.A(dpath_mulcore_ary1_a1_I0_p0_l[44]), .B(dpath_mulcore_b8[0]), .Y(n13273));
INVX1 mul_U7663(.A(n13273), .Y(n982));
AND2X1 mul_U7664(.A(dpath_mulcore_ary1_a1_I0_p2_l[43]), .B(dpath_mulcore_b10[0]), .Y(n13276));
INVX1 mul_U7665(.A(n13276), .Y(n983));
AND2X1 mul_U7666(.A(dpath_mulcore_ary1_a1_I0_p1_l[43]), .B(dpath_mulcore_b9[0]), .Y(n13279));
INVX1 mul_U7667(.A(n13279), .Y(n984));
AND2X1 mul_U7668(.A(dpath_mulcore_ary1_a1_I0_p0_l[43]), .B(dpath_mulcore_b8[0]), .Y(n13282));
INVX1 mul_U7669(.A(n13282), .Y(n985));
AND2X1 mul_U7670(.A(dpath_mulcore_ary1_a1_I0_p2_l[42]), .B(dpath_mulcore_b10[0]), .Y(n13285));
INVX1 mul_U7671(.A(n13285), .Y(n986));
AND2X1 mul_U7672(.A(dpath_mulcore_ary1_a1_I0_p1_l[42]), .B(dpath_mulcore_b9[0]), .Y(n13288));
INVX1 mul_U7673(.A(n13288), .Y(n987));
AND2X1 mul_U7674(.A(dpath_mulcore_ary1_a1_I0_p0_l[42]), .B(dpath_mulcore_b8[0]), .Y(n13291));
INVX1 mul_U7675(.A(n13291), .Y(n988));
AND2X1 mul_U7676(.A(dpath_mulcore_ary1_a1_I0_p2_l[41]), .B(dpath_mulcore_b10[0]), .Y(n13294));
INVX1 mul_U7677(.A(n13294), .Y(n989));
AND2X1 mul_U7678(.A(dpath_mulcore_ary1_a1_I0_p1_l[41]), .B(dpath_mulcore_b9[0]), .Y(n13297));
INVX1 mul_U7679(.A(n13297), .Y(n990));
AND2X1 mul_U7680(.A(dpath_mulcore_ary1_a1_I0_p0_l[41]), .B(dpath_mulcore_b8[0]), .Y(n13300));
INVX1 mul_U7681(.A(n13300), .Y(n991));
AND2X1 mul_U7682(.A(dpath_mulcore_ary1_a1_I0_p2_l[40]), .B(dpath_mulcore_b10[0]), .Y(n13303));
INVX1 mul_U7683(.A(n13303), .Y(n992));
AND2X1 mul_U7684(.A(dpath_mulcore_ary1_a1_I0_p1_l[40]), .B(dpath_mulcore_b9[0]), .Y(n13306));
INVX1 mul_U7685(.A(n13306), .Y(n993));
AND2X1 mul_U7686(.A(dpath_mulcore_ary1_a1_I0_p0_l[40]), .B(dpath_mulcore_b8[0]), .Y(n13309));
INVX1 mul_U7687(.A(n13309), .Y(n994));
AND2X1 mul_U7688(.A(dpath_mulcore_ary1_a1_I0_p2_l[39]), .B(dpath_mulcore_b10[0]), .Y(n13312));
INVX1 mul_U7689(.A(n13312), .Y(n995));
AND2X1 mul_U7690(.A(dpath_mulcore_ary1_a1_I0_p1_l[39]), .B(dpath_mulcore_b9[0]), .Y(n13315));
INVX1 mul_U7691(.A(n13315), .Y(n996));
AND2X1 mul_U7692(.A(dpath_mulcore_ary1_a1_I0_p0_l[39]), .B(dpath_mulcore_b8[0]), .Y(n13318));
INVX1 mul_U7693(.A(n13318), .Y(n997));
AND2X1 mul_U7694(.A(dpath_mulcore_ary1_a1_I0_p2_l[38]), .B(dpath_mulcore_b10[0]), .Y(n13321));
INVX1 mul_U7695(.A(n13321), .Y(n998));
AND2X1 mul_U7696(.A(dpath_mulcore_ary1_a1_I0_p1_l[38]), .B(dpath_mulcore_b9[0]), .Y(n13324));
INVX1 mul_U7697(.A(n13324), .Y(n999));
AND2X1 mul_U7698(.A(dpath_mulcore_ary1_a1_I0_p0_l[38]), .B(dpath_mulcore_b8[0]), .Y(n13327));
INVX1 mul_U7699(.A(n13327), .Y(n1000));
AND2X1 mul_U7700(.A(dpath_mulcore_ary1_a1_I0_p2_l[37]), .B(dpath_mulcore_b10[0]), .Y(n13330));
INVX1 mul_U7701(.A(n13330), .Y(n1001));
AND2X1 mul_U7702(.A(dpath_mulcore_ary1_a1_I0_p1_l[37]), .B(dpath_mulcore_b9[0]), .Y(n13333));
INVX1 mul_U7703(.A(n13333), .Y(n1002));
AND2X1 mul_U7704(.A(dpath_mulcore_ary1_a1_I0_p0_l[37]), .B(dpath_mulcore_b8[0]), .Y(n13336));
INVX1 mul_U7705(.A(n13336), .Y(n1003));
AND2X1 mul_U7706(.A(dpath_mulcore_ary1_a1_I0_p2_l[36]), .B(dpath_mulcore_b10[0]), .Y(n13339));
INVX1 mul_U7707(.A(n13339), .Y(n1004));
AND2X1 mul_U7708(.A(dpath_mulcore_ary1_a1_I0_p1_l[36]), .B(dpath_mulcore_b9[0]), .Y(n13342));
INVX1 mul_U7709(.A(n13342), .Y(n1005));
AND2X1 mul_U7710(.A(dpath_mulcore_ary1_a1_I0_p0_l[36]), .B(dpath_mulcore_b8[0]), .Y(n13345));
INVX1 mul_U7711(.A(n13345), .Y(n1006));
AND2X1 mul_U7712(.A(dpath_mulcore_ary1_a1_I0_p2_l[35]), .B(dpath_mulcore_b10[0]), .Y(n13348));
INVX1 mul_U7713(.A(n13348), .Y(n1007));
AND2X1 mul_U7714(.A(dpath_mulcore_ary1_a1_I0_p1_l[35]), .B(dpath_mulcore_b9[0]), .Y(n13351));
INVX1 mul_U7715(.A(n13351), .Y(n1008));
AND2X1 mul_U7716(.A(dpath_mulcore_ary1_a1_I0_p0_l[35]), .B(dpath_mulcore_b8[0]), .Y(n13354));
INVX1 mul_U7717(.A(n13354), .Y(n1009));
AND2X1 mul_U7718(.A(dpath_mulcore_ary1_a1_I0_p2_l[34]), .B(dpath_mulcore_b10[0]), .Y(n13357));
INVX1 mul_U7719(.A(n13357), .Y(n1010));
AND2X1 mul_U7720(.A(dpath_mulcore_ary1_a1_I0_p1_l[34]), .B(dpath_mulcore_b9[0]), .Y(n13360));
INVX1 mul_U7721(.A(n13360), .Y(n1011));
AND2X1 mul_U7722(.A(dpath_mulcore_ary1_a1_I0_p0_l[34]), .B(dpath_mulcore_b8[0]), .Y(n13363));
INVX1 mul_U7723(.A(n13363), .Y(n1012));
AND2X1 mul_U7724(.A(dpath_mulcore_ary1_a1_I0_p2_l[33]), .B(dpath_mulcore_b10[0]), .Y(n13366));
INVX1 mul_U7725(.A(n13366), .Y(n1013));
AND2X1 mul_U7726(.A(dpath_mulcore_ary1_a1_I0_p1_l[33]), .B(dpath_mulcore_b9[0]), .Y(n13369));
INVX1 mul_U7727(.A(n13369), .Y(n1014));
AND2X1 mul_U7728(.A(dpath_mulcore_ary1_a1_I0_p0_l[33]), .B(dpath_mulcore_b8[0]), .Y(n13372));
INVX1 mul_U7729(.A(n13372), .Y(n1015));
AND2X1 mul_U7730(.A(dpath_mulcore_ary1_a1_I0_p2_l[32]), .B(dpath_mulcore_b10[0]), .Y(n13375));
INVX1 mul_U7731(.A(n13375), .Y(n1016));
AND2X1 mul_U7732(.A(dpath_mulcore_ary1_a1_I0_p1_l[32]), .B(dpath_mulcore_b9[0]), .Y(n13378));
INVX1 mul_U7733(.A(n13378), .Y(n1017));
AND2X1 mul_U7734(.A(dpath_mulcore_ary1_a1_I0_p0_l[32]), .B(dpath_mulcore_b8[0]), .Y(n13381));
INVX1 mul_U7735(.A(n13381), .Y(n1018));
AND2X1 mul_U7736(.A(dpath_mulcore_ary1_a1_I0_p2_l[31]), .B(dpath_mulcore_b10[0]), .Y(n13384));
INVX1 mul_U7737(.A(n13384), .Y(n1019));
AND2X1 mul_U7738(.A(dpath_mulcore_ary1_a1_I0_p1_l[31]), .B(dpath_mulcore_b9[0]), .Y(n13387));
INVX1 mul_U7739(.A(n13387), .Y(n1020));
AND2X1 mul_U7740(.A(dpath_mulcore_ary1_a1_I0_p0_l[31]), .B(dpath_mulcore_b8[0]), .Y(n13390));
INVX1 mul_U7741(.A(n13390), .Y(n1021));
AND2X1 mul_U7742(.A(dpath_mulcore_ary1_a1_I0_p2_l[30]), .B(dpath_mulcore_b10[0]), .Y(n13393));
INVX1 mul_U7743(.A(n13393), .Y(n1022));
AND2X1 mul_U7744(.A(dpath_mulcore_ary1_a1_I0_p1_l[30]), .B(dpath_mulcore_b9[0]), .Y(n13396));
INVX1 mul_U7745(.A(n13396), .Y(n1023));
AND2X1 mul_U7746(.A(dpath_mulcore_ary1_a1_I0_p0_l[30]), .B(dpath_mulcore_b8[0]), .Y(n13399));
INVX1 mul_U7747(.A(n13399), .Y(n1024));
AND2X1 mul_U7748(.A(dpath_mulcore_ary1_a1_I0_p2_l[29]), .B(dpath_mulcore_b10[0]), .Y(n13402));
INVX1 mul_U7749(.A(n13402), .Y(n1025));
AND2X1 mul_U7750(.A(dpath_mulcore_ary1_a1_I0_p1_l[29]), .B(dpath_mulcore_b9[0]), .Y(n13405));
INVX1 mul_U7751(.A(n13405), .Y(n1026));
AND2X1 mul_U7752(.A(dpath_mulcore_ary1_a1_I0_p0_l[29]), .B(dpath_mulcore_b8[0]), .Y(n13408));
INVX1 mul_U7753(.A(n13408), .Y(n1027));
AND2X1 mul_U7754(.A(dpath_mulcore_ary1_a1_I0_p2_l[28]), .B(dpath_mulcore_b10[0]), .Y(n13411));
INVX1 mul_U7755(.A(n13411), .Y(n1028));
AND2X1 mul_U7756(.A(dpath_mulcore_ary1_a1_I0_p1_l[28]), .B(dpath_mulcore_b9[0]), .Y(n13414));
INVX1 mul_U7757(.A(n13414), .Y(n1029));
AND2X1 mul_U7758(.A(dpath_mulcore_ary1_a1_I0_p0_l[28]), .B(dpath_mulcore_b8[0]), .Y(n13417));
INVX1 mul_U7759(.A(n13417), .Y(n1030));
AND2X1 mul_U7760(.A(dpath_mulcore_ary1_a1_I0_p2_l[27]), .B(dpath_mulcore_b10[0]), .Y(n13420));
INVX1 mul_U7761(.A(n13420), .Y(n1031));
AND2X1 mul_U7762(.A(dpath_mulcore_ary1_a1_I0_p1_l[27]), .B(dpath_mulcore_b9[0]), .Y(n13423));
INVX1 mul_U7763(.A(n13423), .Y(n1032));
AND2X1 mul_U7764(.A(dpath_mulcore_ary1_a1_I0_p0_l[27]), .B(dpath_mulcore_b8[0]), .Y(n13426));
INVX1 mul_U7765(.A(n13426), .Y(n1033));
AND2X1 mul_U7766(.A(dpath_mulcore_ary1_a1_I0_p2_l[26]), .B(dpath_mulcore_b10[0]), .Y(n13429));
INVX1 mul_U7767(.A(n13429), .Y(n1034));
AND2X1 mul_U7768(.A(dpath_mulcore_ary1_a1_I0_p1_l[26]), .B(dpath_mulcore_b9[0]), .Y(n13432));
INVX1 mul_U7769(.A(n13432), .Y(n1035));
AND2X1 mul_U7770(.A(dpath_mulcore_ary1_a1_I0_p0_l[26]), .B(dpath_mulcore_b8[0]), .Y(n13435));
INVX1 mul_U7771(.A(n13435), .Y(n1036));
AND2X1 mul_U7772(.A(dpath_mulcore_ary1_a1_I0_p2_l[25]), .B(dpath_mulcore_b10[0]), .Y(n13438));
INVX1 mul_U7773(.A(n13438), .Y(n1037));
AND2X1 mul_U7774(.A(dpath_mulcore_ary1_a1_I0_p1_l[25]), .B(dpath_mulcore_b9[0]), .Y(n13441));
INVX1 mul_U7775(.A(n13441), .Y(n1038));
AND2X1 mul_U7776(.A(dpath_mulcore_ary1_a1_I0_p0_l[25]), .B(dpath_mulcore_b8[0]), .Y(n13444));
INVX1 mul_U7777(.A(n13444), .Y(n1039));
AND2X1 mul_U7778(.A(dpath_mulcore_ary1_a1_I0_p2_l[24]), .B(dpath_mulcore_b10[0]), .Y(n13447));
INVX1 mul_U7779(.A(n13447), .Y(n1040));
AND2X1 mul_U7780(.A(dpath_mulcore_ary1_a1_I0_p1_l[24]), .B(dpath_mulcore_b9[0]), .Y(n13450));
INVX1 mul_U7781(.A(n13450), .Y(n1041));
AND2X1 mul_U7782(.A(dpath_mulcore_ary1_a1_I0_p0_l[24]), .B(dpath_mulcore_b8[0]), .Y(n13453));
INVX1 mul_U7783(.A(n13453), .Y(n1042));
AND2X1 mul_U7784(.A(dpath_mulcore_ary1_a1_I0_p2_l[23]), .B(dpath_mulcore_b10[0]), .Y(n13456));
INVX1 mul_U7785(.A(n13456), .Y(n1043));
AND2X1 mul_U7786(.A(dpath_mulcore_ary1_a1_I0_p1_l[23]), .B(dpath_mulcore_b9[0]), .Y(n13459));
INVX1 mul_U7787(.A(n13459), .Y(n1044));
AND2X1 mul_U7788(.A(dpath_mulcore_ary1_a1_I0_p0_l[23]), .B(dpath_mulcore_b8[0]), .Y(n13462));
INVX1 mul_U7789(.A(n13462), .Y(n1045));
AND2X1 mul_U7790(.A(dpath_mulcore_ary1_a1_I0_p2_l[22]), .B(dpath_mulcore_b10[0]), .Y(n13465));
INVX1 mul_U7791(.A(n13465), .Y(n1046));
AND2X1 mul_U7792(.A(dpath_mulcore_ary1_a1_I0_p1_l[22]), .B(dpath_mulcore_b9[0]), .Y(n13468));
INVX1 mul_U7793(.A(n13468), .Y(n1047));
AND2X1 mul_U7794(.A(dpath_mulcore_ary1_a1_I0_p0_l[22]), .B(dpath_mulcore_b8[0]), .Y(n13471));
INVX1 mul_U7795(.A(n13471), .Y(n1048));
AND2X1 mul_U7796(.A(dpath_mulcore_ary1_a1_I0_p2_l[21]), .B(dpath_mulcore_b10[0]), .Y(n13474));
INVX1 mul_U7797(.A(n13474), .Y(n1049));
AND2X1 mul_U7798(.A(dpath_mulcore_ary1_a1_I0_p1_l[21]), .B(dpath_mulcore_b9[0]), .Y(n13477));
INVX1 mul_U7799(.A(n13477), .Y(n1050));
AND2X1 mul_U7800(.A(dpath_mulcore_ary1_a1_I0_p0_l[21]), .B(dpath_mulcore_b8[0]), .Y(n13480));
INVX1 mul_U7801(.A(n13480), .Y(n1051));
AND2X1 mul_U7802(.A(dpath_mulcore_ary1_a1_I0_p2_l[20]), .B(dpath_mulcore_b10[0]), .Y(n13483));
INVX1 mul_U7803(.A(n13483), .Y(n1052));
AND2X1 mul_U7804(.A(dpath_mulcore_ary1_a1_I0_p1_l[20]), .B(dpath_mulcore_b9[0]), .Y(n13486));
INVX1 mul_U7805(.A(n13486), .Y(n1053));
AND2X1 mul_U7806(.A(dpath_mulcore_ary1_a1_I0_p0_l[20]), .B(dpath_mulcore_b8[0]), .Y(n13489));
INVX1 mul_U7807(.A(n13489), .Y(n1054));
AND2X1 mul_U7808(.A(dpath_mulcore_ary1_a1_I0_p2_l[19]), .B(dpath_mulcore_b10[0]), .Y(n13492));
INVX1 mul_U7809(.A(n13492), .Y(n1055));
AND2X1 mul_U7810(.A(dpath_mulcore_ary1_a1_I0_p1_l[19]), .B(dpath_mulcore_b9[0]), .Y(n13495));
INVX1 mul_U7811(.A(n13495), .Y(n1056));
AND2X1 mul_U7812(.A(dpath_mulcore_ary1_a1_I0_p0_l[19]), .B(dpath_mulcore_b8[0]), .Y(n13498));
INVX1 mul_U7813(.A(n13498), .Y(n1057));
AND2X1 mul_U7814(.A(dpath_mulcore_ary1_a1_I0_p2_l[18]), .B(dpath_mulcore_b10[0]), .Y(n13501));
INVX1 mul_U7815(.A(n13501), .Y(n1058));
AND2X1 mul_U7816(.A(dpath_mulcore_ary1_a1_I0_p1_l[18]), .B(dpath_mulcore_b9[0]), .Y(n13504));
INVX1 mul_U7817(.A(n13504), .Y(n1059));
AND2X1 mul_U7818(.A(dpath_mulcore_ary1_a1_I0_p0_l[18]), .B(dpath_mulcore_b8[0]), .Y(n13507));
INVX1 mul_U7819(.A(n13507), .Y(n1060));
AND2X1 mul_U7820(.A(dpath_mulcore_ary1_a1_I0_p2_l[17]), .B(dpath_mulcore_b10[0]), .Y(n13510));
INVX1 mul_U7821(.A(n13510), .Y(n1061));
AND2X1 mul_U7822(.A(dpath_mulcore_ary1_a1_I0_p1_l[17]), .B(dpath_mulcore_b9[0]), .Y(n13513));
INVX1 mul_U7823(.A(n13513), .Y(n1062));
AND2X1 mul_U7824(.A(dpath_mulcore_ary1_a1_I0_p0_l[17]), .B(dpath_mulcore_b8[0]), .Y(n13516));
INVX1 mul_U7825(.A(n13516), .Y(n1063));
AND2X1 mul_U7826(.A(dpath_mulcore_ary1_a1_I0_p2_l[16]), .B(dpath_mulcore_b10[0]), .Y(n13519));
INVX1 mul_U7827(.A(n13519), .Y(n1064));
AND2X1 mul_U7828(.A(dpath_mulcore_ary1_a1_I0_p1_l[16]), .B(dpath_mulcore_b9[0]), .Y(n13522));
INVX1 mul_U7829(.A(n13522), .Y(n1065));
AND2X1 mul_U7830(.A(dpath_mulcore_ary1_a1_I0_p0_l[16]), .B(dpath_mulcore_b8[0]), .Y(n13525));
INVX1 mul_U7831(.A(n13525), .Y(n1066));
AND2X1 mul_U7832(.A(dpath_mulcore_ary1_a1_I0_p2_l[15]), .B(dpath_mulcore_b10[0]), .Y(n13528));
INVX1 mul_U7833(.A(n13528), .Y(n1067));
AND2X1 mul_U7834(.A(dpath_mulcore_ary1_a1_I0_p1_l[15]), .B(dpath_mulcore_b9[0]), .Y(n13531));
INVX1 mul_U7835(.A(n13531), .Y(n1068));
AND2X1 mul_U7836(.A(dpath_mulcore_ary1_a1_I0_p0_l[15]), .B(dpath_mulcore_b8[0]), .Y(n13534));
INVX1 mul_U7837(.A(n13534), .Y(n1069));
AND2X1 mul_U7838(.A(dpath_mulcore_ary1_a1_I0_p2_l[14]), .B(dpath_mulcore_b10[0]), .Y(n13537));
INVX1 mul_U7839(.A(n13537), .Y(n1070));
AND2X1 mul_U7840(.A(dpath_mulcore_ary1_a1_I0_p1_l[14]), .B(dpath_mulcore_b9[0]), .Y(n13540));
INVX1 mul_U7841(.A(n13540), .Y(n1071));
AND2X1 mul_U7842(.A(dpath_mulcore_ary1_a1_I0_p0_l[14]), .B(dpath_mulcore_b8[0]), .Y(n13543));
INVX1 mul_U7843(.A(n13543), .Y(n1072));
AND2X1 mul_U7844(.A(dpath_mulcore_ary1_a1_I0_p2_l[13]), .B(dpath_mulcore_b10[0]), .Y(n13546));
INVX1 mul_U7845(.A(n13546), .Y(n1073));
AND2X1 mul_U7846(.A(dpath_mulcore_ary1_a1_I0_p1_l[13]), .B(dpath_mulcore_b9[0]), .Y(n13549));
INVX1 mul_U7847(.A(n13549), .Y(n1074));
AND2X1 mul_U7848(.A(dpath_mulcore_ary1_a1_I0_p0_l[13]), .B(dpath_mulcore_b8[0]), .Y(n13552));
INVX1 mul_U7849(.A(n13552), .Y(n1075));
AND2X1 mul_U7850(.A(dpath_mulcore_ary1_a1_I0_p2_l[12]), .B(dpath_mulcore_b10[0]), .Y(n13555));
INVX1 mul_U7851(.A(n13555), .Y(n1076));
AND2X1 mul_U7852(.A(dpath_mulcore_ary1_a1_I0_p1_l[12]), .B(dpath_mulcore_b9[0]), .Y(n13558));
INVX1 mul_U7853(.A(n13558), .Y(n1077));
AND2X1 mul_U7854(.A(dpath_mulcore_ary1_a1_I0_p0_l[12]), .B(dpath_mulcore_b8[0]), .Y(n13561));
INVX1 mul_U7855(.A(n13561), .Y(n1078));
AND2X1 mul_U7856(.A(dpath_mulcore_ary1_a1_I0_p2_l[11]), .B(dpath_mulcore_b10[0]), .Y(n13564));
INVX1 mul_U7857(.A(n13564), .Y(n1079));
AND2X1 mul_U7858(.A(dpath_mulcore_ary1_a1_I0_p1_l[11]), .B(dpath_mulcore_b9[0]), .Y(n13567));
INVX1 mul_U7859(.A(n13567), .Y(n1080));
AND2X1 mul_U7860(.A(dpath_mulcore_ary1_a1_I0_p0_l[11]), .B(dpath_mulcore_b8[0]), .Y(n13570));
INVX1 mul_U7861(.A(n13570), .Y(n1081));
AND2X1 mul_U7862(.A(dpath_mulcore_ary1_a1_I0_p2_l[10]), .B(dpath_mulcore_b10[0]), .Y(n13573));
INVX1 mul_U7863(.A(n13573), .Y(n1082));
AND2X1 mul_U7864(.A(dpath_mulcore_ary1_a1_I0_p1_l[10]), .B(dpath_mulcore_b9[0]), .Y(n13576));
INVX1 mul_U7865(.A(n13576), .Y(n1083));
AND2X1 mul_U7866(.A(dpath_mulcore_ary1_a1_I0_p0_l[10]), .B(dpath_mulcore_b8[0]), .Y(n13579));
INVX1 mul_U7867(.A(n13579), .Y(n1084));
AND2X1 mul_U7868(.A(dpath_mulcore_ary1_a1_I0_p2_l[9]), .B(dpath_mulcore_b10[0]), .Y(n13582));
INVX1 mul_U7869(.A(n13582), .Y(n1085));
AND2X1 mul_U7870(.A(dpath_mulcore_ary1_a1_I0_p1_l[9]), .B(dpath_mulcore_b9[0]), .Y(n13585));
INVX1 mul_U7871(.A(n13585), .Y(n1086));
AND2X1 mul_U7872(.A(dpath_mulcore_ary1_a1_I0_p0_l[9]), .B(dpath_mulcore_b8[0]), .Y(n13588));
INVX1 mul_U7873(.A(n13588), .Y(n1087));
AND2X1 mul_U7874(.A(dpath_mulcore_ary1_a1_I0_p2_l[8]), .B(dpath_mulcore_b10[0]), .Y(n13591));
INVX1 mul_U7875(.A(n13591), .Y(n1088));
AND2X1 mul_U7876(.A(dpath_mulcore_ary1_a1_I0_p1_l[8]), .B(dpath_mulcore_b9[0]), .Y(n13594));
INVX1 mul_U7877(.A(n13594), .Y(n1089));
AND2X1 mul_U7878(.A(dpath_mulcore_ary1_a1_I0_p0_l[8]), .B(dpath_mulcore_b8[0]), .Y(n13597));
INVX1 mul_U7879(.A(n13597), .Y(n1090));
AND2X1 mul_U7880(.A(dpath_mulcore_ary1_a1_I0_p2_l[7]), .B(dpath_mulcore_b10[0]), .Y(n13600));
INVX1 mul_U7881(.A(n13600), .Y(n1091));
AND2X1 mul_U7882(.A(dpath_mulcore_ary1_a1_I0_p1_l[7]), .B(dpath_mulcore_b9[0]), .Y(n13603));
INVX1 mul_U7883(.A(n13603), .Y(n1092));
AND2X1 mul_U7884(.A(dpath_mulcore_ary1_a1_I0_p0_l[7]), .B(dpath_mulcore_b8[0]), .Y(n13606));
INVX1 mul_U7885(.A(n13606), .Y(n1093));
AND2X1 mul_U7886(.A(dpath_mulcore_ary1_a1_I0_p2_l[6]), .B(dpath_mulcore_b10[0]), .Y(n13609));
INVX1 mul_U7887(.A(n13609), .Y(n1094));
AND2X1 mul_U7888(.A(dpath_mulcore_ary1_a1_I0_p1_l[6]), .B(dpath_mulcore_b9[0]), .Y(n13612));
INVX1 mul_U7889(.A(n13612), .Y(n1095));
AND2X1 mul_U7890(.A(dpath_mulcore_ary1_a1_I0_p0_l[6]), .B(dpath_mulcore_b8[0]), .Y(n13615));
INVX1 mul_U7891(.A(n13615), .Y(n1096));
AND2X1 mul_U7892(.A(dpath_mulcore_ary1_a1_I0_p2_l[5]), .B(dpath_mulcore_b10[0]), .Y(n13618));
INVX1 mul_U7893(.A(n13618), .Y(n1097));
AND2X1 mul_U7894(.A(dpath_mulcore_ary1_a1_I0_p1_l[5]), .B(dpath_mulcore_b9[0]), .Y(n13621));
INVX1 mul_U7895(.A(n13621), .Y(n1098));
AND2X1 mul_U7896(.A(dpath_mulcore_ary1_a1_I0_p0_l[5]), .B(dpath_mulcore_b8[0]), .Y(n13624));
INVX1 mul_U7897(.A(n13624), .Y(n1099));
AND2X1 mul_U7898(.A(dpath_mulcore_ary1_a1_I0_p2_l[4]), .B(dpath_mulcore_b10[0]), .Y(n13627));
INVX1 mul_U7899(.A(n13627), .Y(n1100));
AND2X1 mul_U7900(.A(dpath_mulcore_ary1_a1_I0_p1_l[4]), .B(dpath_mulcore_b9[0]), .Y(n13630));
INVX1 mul_U7901(.A(n13630), .Y(n1101));
AND2X1 mul_U7902(.A(dpath_mulcore_ary1_a1_I0_p0_l[4]), .B(dpath_mulcore_b8[0]), .Y(n13633));
INVX1 mul_U7903(.A(n13633), .Y(n1102));
AND2X1 mul_U7904(.A(dpath_mulcore_ary1_a1_I0_p1_l[3]), .B(dpath_mulcore_b9[0]), .Y(n13638));
INVX1 mul_U7905(.A(n13638), .Y(n1103));
AND2X1 mul_U7906(.A(dpath_mulcore_ary1_a1_I0_p0_l[3]), .B(dpath_mulcore_b8[0]), .Y(n13641));
INVX1 mul_U7907(.A(n13641), .Y(n1104));
AND2X1 mul_U7908(.A(dpath_mulcore_ary1_a1_I0_I0_p0_l_2), .B(dpath_mulcore_b8[0]), .Y(n13644));
INVX1 mul_U7909(.A(n13644), .Y(n1105));
AND2X1 mul_U7910(.A(dpath_mulcore_ary1_a1_I0_I0_p1_l_2), .B(dpath_mulcore_b9[0]), .Y(n13647));
INVX1 mul_U7911(.A(n13647), .Y(n1106));
AND2X1 mul_U7912(.A(dpath_mulcore_ary1_a1_I0_I0_p0_l_1), .B(dpath_mulcore_b8[0]), .Y(n13650));
INVX1 mul_U7913(.A(n13650), .Y(n1107));
AND2X1 mul_U7914(.A(dpath_mulcore_ary1_a1_I0_I0_p0_l_0), .B(dpath_mulcore_b8[0]), .Y(n13653));
INVX1 mul_U7915(.A(n13653), .Y(n1108));
AND2X1 mul_U7916(.A(dpath_mulcore_ary1_a0_I2_I2_p1_l_65), .B(dpath_mulcore_b7[0]), .Y(n13660));
INVX1 mul_U7917(.A(n13660), .Y(n1109));
AND2X1 mul_U7918(.A(dpath_mulcore_ary1_a0_I1_p0_l[63]), .B(dpath_mulcore_b3[0]), .Y(n13662));
INVX1 mul_U7919(.A(n13662), .Y(n1110));
AND2X1 mul_U7920(.A(dpath_mulcore_ary1_a0_I1_I2_p2_l_67), .B(dpath_mulcore_b5[0]), .Y(n13664));
INVX1 mul_U7921(.A(n13664), .Y(n1111));
AND2X1 mul_U7922(.A(dpath_mulcore_ary1_a0_I1_I2_p1_l_65), .B(dpath_mulcore_b4[0]), .Y(n13666));
INVX1 mul_U7923(.A(n13666), .Y(n1112));
AND2X1 mul_U7924(.A(dpath_mulcore_ary1_a0_I0_p0_l[63]), .B(dpath_mulcore_b0[0]), .Y(n13668));
INVX1 mul_U7925(.A(n13668), .Y(n1113));
AND2X1 mul_U7926(.A(dpath_mulcore_ary1_a0_I0_I2_p2_l_67), .B(dpath_mulcore_b2[0]), .Y(n13670));
INVX1 mul_U7927(.A(n13670), .Y(n1114));
AND2X1 mul_U7928(.A(dpath_mulcore_ary1_a0_I0_I2_p1_l_65), .B(dpath_mulcore_b1[0]), .Y(n13672));
INVX1 mul_U7929(.A(n13672), .Y(n1115));
AND2X1 mul_U7930(.A(dpath_mulcore_ary1_a1_I2_p0_l[63]), .B(dpath_mulcore_b14[0]), .Y(n13674));
INVX1 mul_U7931(.A(n13674), .Y(n1116));
AND2X1 mul_U7932(.A(dpath_mulcore_ary1_a1_I2_I2_p1_l_65), .B(dpath_mulcore_b15[0]), .Y(n13676));
INVX1 mul_U7933(.A(n13676), .Y(n1117));
AND2X1 mul_U7934(.A(dpath_mulcore_ary1_a1_I1_p0_l[63]), .B(dpath_mulcore_b11[0]), .Y(n13678));
INVX1 mul_U7935(.A(n13678), .Y(n1118));
AND2X1 mul_U7936(.A(dpath_mulcore_ary1_a1_I1_I2_p2_l_67), .B(dpath_mulcore_b13[0]), .Y(n13680));
INVX1 mul_U7937(.A(n13680), .Y(n1119));
AND2X1 mul_U7938(.A(dpath_mulcore_ary1_a1_I1_I2_p1_l_65), .B(dpath_mulcore_b12[0]), .Y(n13682));
INVX1 mul_U7939(.A(n13682), .Y(n1120));
AND2X1 mul_U7940(.A(dpath_mulcore_ary1_a1_I0_p0_l[63]), .B(dpath_mulcore_b8[0]), .Y(n13684));
INVX1 mul_U7941(.A(n13684), .Y(n1121));
AND2X1 mul_U7942(.A(dpath_mulcore_ary1_a1_I0_I2_p2_l_67), .B(dpath_mulcore_b10[0]), .Y(n13686));
INVX1 mul_U7943(.A(n13686), .Y(n1122));
AND2X1 mul_U7944(.A(dpath_mulcore_ary1_a1_I0_I2_p1_l_65), .B(dpath_mulcore_b9[0]), .Y(n13688));
INVX1 mul_U7945(.A(n13688), .Y(n1123));
AND2X1 mul_U7946(.A(n7606), .B(n8509), .Y(n13696));
INVX1 mul_U7947(.A(n13696), .Y(n1124));
AND2X1 mul_U7948(.A(n7607), .B(n9844), .Y(n13699));
INVX1 mul_U7949(.A(n13699), .Y(n1125));
AND2X1 mul_U7950(.A(n7733), .B(n8570), .Y(n13707));
INVX1 mul_U7951(.A(n13707), .Y(n1126));
AND2X1 mul_U7952(.A(n7734), .B(n9840), .Y(n13710));
INVX1 mul_U7953(.A(n13710), .Y(n1127));
AND2X1 mul_U7954(.A(n7797), .B(n8631), .Y(n13718));
INVX1 mul_U7955(.A(n13718), .Y(n1128));
AND2X1 mul_U7956(.A(n7798), .B(n9838), .Y(n13721));
INVX1 mul_U7957(.A(n13721), .Y(n1129));
AND2X1 mul_U7958(.A(n7924), .B(n8692), .Y(n13729));
INVX1 mul_U7959(.A(n13729), .Y(n1130));
AND2X1 mul_U7960(.A(n7925), .B(n9831), .Y(n13732));
INVX1 mul_U7961(.A(n13732), .Y(n1131));
AND2X1 mul_U7962(.A(n8051), .B(n8753), .Y(n13740));
INVX1 mul_U7963(.A(n13740), .Y(n1132));
AND2X1 mul_U7964(.A(n8052), .B(n9827), .Y(n13743));
INVX1 mul_U7965(.A(n13743), .Y(n1133));
AND2X1 mul_U7966(.A(n7488), .B(n8449), .Y(n13864));
INVX1 mul_U7967(.A(n13864), .Y(n1134));
AND2X1 mul_U7968(.A(n7490), .B(n8450), .Y(n13867));
INVX1 mul_U7969(.A(n13867), .Y(n1135));
AND2X1 mul_U7970(.A(n7492), .B(n8451), .Y(n13870));
INVX1 mul_U7971(.A(n13870), .Y(n1136));
AND2X1 mul_U7972(.A(n7494), .B(n8452), .Y(n13873));
INVX1 mul_U7973(.A(n13873), .Y(n1137));
AND2X1 mul_U7974(.A(n7496), .B(n8453), .Y(n13876));
INVX1 mul_U7975(.A(n13876), .Y(n1138));
AND2X1 mul_U7976(.A(n7498), .B(n8454), .Y(n13879));
INVX1 mul_U7977(.A(n13879), .Y(n1139));
AND2X1 mul_U7978(.A(n7500), .B(n8455), .Y(n13882));
INVX1 mul_U7979(.A(n13882), .Y(n1140));
AND2X1 mul_U7980(.A(n7502), .B(n8456), .Y(n13885));
INVX1 mul_U7981(.A(n13885), .Y(n1141));
AND2X1 mul_U7982(.A(n7504), .B(n8457), .Y(n13888));
INVX1 mul_U7983(.A(n13888), .Y(n1142));
AND2X1 mul_U7984(.A(n7506), .B(n8458), .Y(n13891));
INVX1 mul_U7985(.A(n13891), .Y(n1143));
AND2X1 mul_U7986(.A(n7508), .B(n8459), .Y(n13894));
INVX1 mul_U7987(.A(n13894), .Y(n1144));
AND2X1 mul_U7988(.A(n7510), .B(n8460), .Y(n13897));
INVX1 mul_U7989(.A(n13897), .Y(n1145));
AND2X1 mul_U7990(.A(n7512), .B(n8461), .Y(n13900));
INVX1 mul_U7991(.A(n13900), .Y(n1146));
AND2X1 mul_U7992(.A(n7514), .B(n8462), .Y(n13903));
INVX1 mul_U7993(.A(n13903), .Y(n1147));
AND2X1 mul_U7994(.A(n7516), .B(n8463), .Y(n13906));
INVX1 mul_U7995(.A(n13906), .Y(n1148));
AND2X1 mul_U7996(.A(n7518), .B(n8464), .Y(n13909));
INVX1 mul_U7997(.A(n13909), .Y(n1149));
AND2X1 mul_U7998(.A(n7520), .B(n8465), .Y(n13912));
INVX1 mul_U7999(.A(n13912), .Y(n1150));
AND2X1 mul_U8000(.A(n7522), .B(n8466), .Y(n13915));
INVX1 mul_U8001(.A(n13915), .Y(n1151));
AND2X1 mul_U8002(.A(n7524), .B(n8467), .Y(n13918));
INVX1 mul_U8003(.A(n13918), .Y(n1152));
AND2X1 mul_U8004(.A(n7526), .B(n8468), .Y(n13921));
INVX1 mul_U8005(.A(n13921), .Y(n1153));
AND2X1 mul_U8006(.A(n7528), .B(n8469), .Y(n13924));
INVX1 mul_U8007(.A(n13924), .Y(n1154));
AND2X1 mul_U8008(.A(n7530), .B(n8470), .Y(n13927));
INVX1 mul_U8009(.A(n13927), .Y(n1155));
AND2X1 mul_U8010(.A(n7532), .B(n8471), .Y(n13930));
INVX1 mul_U8011(.A(n13930), .Y(n1156));
AND2X1 mul_U8012(.A(n7534), .B(n8472), .Y(n13933));
INVX1 mul_U8013(.A(n13933), .Y(n1157));
AND2X1 mul_U8014(.A(n7536), .B(n8473), .Y(n13936));
INVX1 mul_U8015(.A(n13936), .Y(n1158));
AND2X1 mul_U8016(.A(n7538), .B(n8474), .Y(n13939));
INVX1 mul_U8017(.A(n13939), .Y(n1159));
AND2X1 mul_U8018(.A(n7540), .B(n8475), .Y(n13942));
INVX1 mul_U8019(.A(n13942), .Y(n1160));
AND2X1 mul_U8020(.A(n7542), .B(n8476), .Y(n13945));
INVX1 mul_U8021(.A(n13945), .Y(n1161));
AND2X1 mul_U8022(.A(n7544), .B(n8477), .Y(n13948));
INVX1 mul_U8023(.A(n13948), .Y(n1162));
AND2X1 mul_U8024(.A(n7546), .B(n8478), .Y(n13951));
INVX1 mul_U8025(.A(n13951), .Y(n1163));
AND2X1 mul_U8026(.A(n7548), .B(n8479), .Y(n13954));
INVX1 mul_U8027(.A(n13954), .Y(n1164));
AND2X1 mul_U8028(.A(n7550), .B(n8480), .Y(n13957));
INVX1 mul_U8029(.A(n13957), .Y(n1165));
AND2X1 mul_U8030(.A(n7552), .B(n8481), .Y(n13960));
INVX1 mul_U8031(.A(n13960), .Y(n1166));
AND2X1 mul_U8032(.A(n7554), .B(n8482), .Y(n13963));
INVX1 mul_U8033(.A(n13963), .Y(n1167));
AND2X1 mul_U8034(.A(n7556), .B(n8483), .Y(n13966));
INVX1 mul_U8035(.A(n13966), .Y(n1168));
AND2X1 mul_U8036(.A(n7558), .B(n8484), .Y(n13969));
INVX1 mul_U8037(.A(n13969), .Y(n1169));
AND2X1 mul_U8038(.A(n7560), .B(n8485), .Y(n13972));
INVX1 mul_U8039(.A(n13972), .Y(n1170));
AND2X1 mul_U8040(.A(n7562), .B(n8486), .Y(n13975));
INVX1 mul_U8041(.A(n13975), .Y(n1171));
AND2X1 mul_U8042(.A(n7564), .B(n8487), .Y(n13978));
INVX1 mul_U8043(.A(n13978), .Y(n1172));
AND2X1 mul_U8044(.A(n7566), .B(n8488), .Y(n13981));
INVX1 mul_U8045(.A(n13981), .Y(n1173));
AND2X1 mul_U8046(.A(n7568), .B(n8489), .Y(n13984));
INVX1 mul_U8047(.A(n13984), .Y(n1174));
AND2X1 mul_U8048(.A(n7570), .B(n8490), .Y(n13987));
INVX1 mul_U8049(.A(n13987), .Y(n1175));
AND2X1 mul_U8050(.A(n7572), .B(n8491), .Y(n13990));
INVX1 mul_U8051(.A(n13990), .Y(n1176));
AND2X1 mul_U8052(.A(n7574), .B(n8492), .Y(n13993));
INVX1 mul_U8053(.A(n13993), .Y(n1177));
AND2X1 mul_U8054(.A(n7576), .B(n8493), .Y(n13996));
INVX1 mul_U8055(.A(n13996), .Y(n1178));
AND2X1 mul_U8056(.A(n7578), .B(n8494), .Y(n13999));
INVX1 mul_U8057(.A(n13999), .Y(n1179));
AND2X1 mul_U8058(.A(n7580), .B(n8495), .Y(n14002));
INVX1 mul_U8059(.A(n14002), .Y(n1180));
AND2X1 mul_U8060(.A(n7582), .B(n8496), .Y(n14005));
INVX1 mul_U8061(.A(n14005), .Y(n1181));
AND2X1 mul_U8062(.A(n7584), .B(n8497), .Y(n14008));
INVX1 mul_U8063(.A(n14008), .Y(n1182));
AND2X1 mul_U8064(.A(n7586), .B(n8498), .Y(n14011));
INVX1 mul_U8065(.A(n14011), .Y(n1183));
AND2X1 mul_U8066(.A(n7588), .B(n8499), .Y(n14014));
INVX1 mul_U8067(.A(n14014), .Y(n1184));
AND2X1 mul_U8068(.A(n7590), .B(n8500), .Y(n14017));
INVX1 mul_U8069(.A(n14017), .Y(n1185));
AND2X1 mul_U8070(.A(n7592), .B(n8501), .Y(n14020));
INVX1 mul_U8071(.A(n14020), .Y(n1186));
AND2X1 mul_U8072(.A(n7594), .B(n8502), .Y(n14023));
INVX1 mul_U8073(.A(n14023), .Y(n1187));
AND2X1 mul_U8074(.A(n7596), .B(n8503), .Y(n14026));
INVX1 mul_U8075(.A(n14026), .Y(n1188));
AND2X1 mul_U8076(.A(n7598), .B(n8504), .Y(n14029));
INVX1 mul_U8077(.A(n14029), .Y(n1189));
AND2X1 mul_U8078(.A(n7600), .B(n8505), .Y(n14032));
INVX1 mul_U8079(.A(n14032), .Y(n1190));
AND2X1 mul_U8080(.A(n7602), .B(n8506), .Y(n14035));
INVX1 mul_U8081(.A(n14035), .Y(n1191));
AND2X1 mul_U8082(.A(n7604), .B(n8507), .Y(n14038));
INVX1 mul_U8083(.A(n14038), .Y(n1192));
AND2X1 mul_U8084(.A(n7605), .B(n8508), .Y(n14041));
INVX1 mul_U8085(.A(n14041), .Y(n1193));
AND2X1 mul_U8086(.A(n7615), .B(n8510), .Y(n14044));
INVX1 mul_U8087(.A(n14044), .Y(n1194));
AND2X1 mul_U8088(.A(n7617), .B(n8511), .Y(n14047));
INVX1 mul_U8089(.A(n14047), .Y(n1195));
AND2X1 mul_U8090(.A(n7619), .B(n8512), .Y(n14050));
INVX1 mul_U8091(.A(n14050), .Y(n1196));
AND2X1 mul_U8092(.A(n7621), .B(n8513), .Y(n14053));
INVX1 mul_U8093(.A(n14053), .Y(n1197));
AND2X1 mul_U8094(.A(n7623), .B(n8514), .Y(n14056));
INVX1 mul_U8095(.A(n14056), .Y(n1198));
AND2X1 mul_U8096(.A(n7625), .B(n8515), .Y(n14059));
INVX1 mul_U8097(.A(n14059), .Y(n1199));
AND2X1 mul_U8098(.A(n7627), .B(n8516), .Y(n14062));
INVX1 mul_U8099(.A(n14062), .Y(n1200));
AND2X1 mul_U8100(.A(n7629), .B(n8517), .Y(n14065));
INVX1 mul_U8101(.A(n14065), .Y(n1201));
AND2X1 mul_U8102(.A(n7631), .B(n8518), .Y(n14068));
INVX1 mul_U8103(.A(n14068), .Y(n1202));
AND2X1 mul_U8104(.A(n7633), .B(n8519), .Y(n14071));
INVX1 mul_U8105(.A(n14071), .Y(n1203));
AND2X1 mul_U8106(.A(n7635), .B(n8520), .Y(n14074));
INVX1 mul_U8107(.A(n14074), .Y(n1204));
AND2X1 mul_U8108(.A(n7637), .B(n8521), .Y(n14077));
INVX1 mul_U8109(.A(n14077), .Y(n1205));
AND2X1 mul_U8110(.A(n7639), .B(n8522), .Y(n14080));
INVX1 mul_U8111(.A(n14080), .Y(n1206));
AND2X1 mul_U8112(.A(n7641), .B(n8523), .Y(n14083));
INVX1 mul_U8113(.A(n14083), .Y(n1207));
AND2X1 mul_U8114(.A(n7643), .B(n8524), .Y(n14086));
INVX1 mul_U8115(.A(n14086), .Y(n1208));
AND2X1 mul_U8116(.A(n7645), .B(n8525), .Y(n14089));
INVX1 mul_U8117(.A(n14089), .Y(n1209));
AND2X1 mul_U8118(.A(n7647), .B(n8526), .Y(n14092));
INVX1 mul_U8119(.A(n14092), .Y(n1210));
AND2X1 mul_U8120(.A(n7649), .B(n8527), .Y(n14095));
INVX1 mul_U8121(.A(n14095), .Y(n1211));
AND2X1 mul_U8122(.A(n7651), .B(n8528), .Y(n14098));
INVX1 mul_U8123(.A(n14098), .Y(n1212));
AND2X1 mul_U8124(.A(n7653), .B(n8529), .Y(n14101));
INVX1 mul_U8125(.A(n14101), .Y(n1213));
AND2X1 mul_U8126(.A(n7655), .B(n8530), .Y(n14104));
INVX1 mul_U8127(.A(n14104), .Y(n1214));
AND2X1 mul_U8128(.A(n7657), .B(n8531), .Y(n14107));
INVX1 mul_U8129(.A(n14107), .Y(n1215));
AND2X1 mul_U8130(.A(n7659), .B(n8532), .Y(n14110));
INVX1 mul_U8131(.A(n14110), .Y(n1216));
AND2X1 mul_U8132(.A(n7661), .B(n8533), .Y(n14113));
INVX1 mul_U8133(.A(n14113), .Y(n1217));
AND2X1 mul_U8134(.A(n7663), .B(n8534), .Y(n14116));
INVX1 mul_U8135(.A(n14116), .Y(n1218));
AND2X1 mul_U8136(.A(n7665), .B(n8535), .Y(n14119));
INVX1 mul_U8137(.A(n14119), .Y(n1219));
AND2X1 mul_U8138(.A(n7667), .B(n8536), .Y(n14122));
INVX1 mul_U8139(.A(n14122), .Y(n1220));
AND2X1 mul_U8140(.A(n7669), .B(n8537), .Y(n14125));
INVX1 mul_U8141(.A(n14125), .Y(n1221));
AND2X1 mul_U8142(.A(n7671), .B(n8538), .Y(n14128));
INVX1 mul_U8143(.A(n14128), .Y(n1222));
AND2X1 mul_U8144(.A(n7673), .B(n8539), .Y(n14131));
INVX1 mul_U8145(.A(n14131), .Y(n1223));
AND2X1 mul_U8146(.A(n7675), .B(n8540), .Y(n14134));
INVX1 mul_U8147(.A(n14134), .Y(n1224));
AND2X1 mul_U8148(.A(n7677), .B(n8541), .Y(n14137));
INVX1 mul_U8149(.A(n14137), .Y(n1225));
AND2X1 mul_U8150(.A(n7679), .B(n8542), .Y(n14140));
INVX1 mul_U8151(.A(n14140), .Y(n1226));
AND2X1 mul_U8152(.A(n7681), .B(n8543), .Y(n14143));
INVX1 mul_U8153(.A(n14143), .Y(n1227));
AND2X1 mul_U8154(.A(n7683), .B(n8544), .Y(n14146));
INVX1 mul_U8155(.A(n14146), .Y(n1228));
AND2X1 mul_U8156(.A(n7685), .B(n8545), .Y(n14149));
INVX1 mul_U8157(.A(n14149), .Y(n1229));
AND2X1 mul_U8158(.A(n7687), .B(n8546), .Y(n14152));
INVX1 mul_U8159(.A(n14152), .Y(n1230));
AND2X1 mul_U8160(.A(n7689), .B(n8547), .Y(n14155));
INVX1 mul_U8161(.A(n14155), .Y(n1231));
AND2X1 mul_U8162(.A(n7691), .B(n8548), .Y(n14158));
INVX1 mul_U8163(.A(n14158), .Y(n1232));
AND2X1 mul_U8164(.A(n7693), .B(n8549), .Y(n14161));
INVX1 mul_U8165(.A(n14161), .Y(n1233));
AND2X1 mul_U8166(.A(n7695), .B(n8550), .Y(n14164));
INVX1 mul_U8167(.A(n14164), .Y(n1234));
AND2X1 mul_U8168(.A(n7697), .B(n8551), .Y(n14167));
INVX1 mul_U8169(.A(n14167), .Y(n1235));
AND2X1 mul_U8170(.A(n7699), .B(n8552), .Y(n14170));
INVX1 mul_U8171(.A(n14170), .Y(n1236));
AND2X1 mul_U8172(.A(n7701), .B(n8553), .Y(n14173));
INVX1 mul_U8173(.A(n14173), .Y(n1237));
AND2X1 mul_U8174(.A(n7703), .B(n8554), .Y(n14176));
INVX1 mul_U8175(.A(n14176), .Y(n1238));
AND2X1 mul_U8176(.A(n7705), .B(n8555), .Y(n14179));
INVX1 mul_U8177(.A(n14179), .Y(n1239));
AND2X1 mul_U8178(.A(n7707), .B(n8556), .Y(n14182));
INVX1 mul_U8179(.A(n14182), .Y(n1240));
AND2X1 mul_U8180(.A(n7709), .B(n8557), .Y(n14185));
INVX1 mul_U8181(.A(n14185), .Y(n1241));
AND2X1 mul_U8182(.A(n7711), .B(n8558), .Y(n14188));
INVX1 mul_U8183(.A(n14188), .Y(n1242));
AND2X1 mul_U8184(.A(n7713), .B(n8559), .Y(n14191));
INVX1 mul_U8185(.A(n14191), .Y(n1243));
AND2X1 mul_U8186(.A(n7715), .B(n8560), .Y(n14194));
INVX1 mul_U8187(.A(n14194), .Y(n1244));
AND2X1 mul_U8188(.A(n7717), .B(n8561), .Y(n14197));
INVX1 mul_U8189(.A(n14197), .Y(n1245));
AND2X1 mul_U8190(.A(n7719), .B(n8562), .Y(n14200));
INVX1 mul_U8191(.A(n14200), .Y(n1246));
AND2X1 mul_U8192(.A(n7721), .B(n8563), .Y(n14203));
INVX1 mul_U8193(.A(n14203), .Y(n1247));
AND2X1 mul_U8194(.A(n7723), .B(n8564), .Y(n14206));
INVX1 mul_U8195(.A(n14206), .Y(n1248));
AND2X1 mul_U8196(.A(n7725), .B(n8565), .Y(n14209));
INVX1 mul_U8197(.A(n14209), .Y(n1249));
AND2X1 mul_U8198(.A(n7727), .B(n8566), .Y(n14212));
INVX1 mul_U8199(.A(n14212), .Y(n1250));
AND2X1 mul_U8200(.A(n7729), .B(n8567), .Y(n14215));
INVX1 mul_U8201(.A(n14215), .Y(n1251));
AND2X1 mul_U8202(.A(n7731), .B(n8568), .Y(n14218));
INVX1 mul_U8203(.A(n14218), .Y(n1252));
AND2X1 mul_U8204(.A(n7732), .B(n8569), .Y(n14221));
INVX1 mul_U8205(.A(n14221), .Y(n1253));
AND2X1 mul_U8206(.A(n7737), .B(n8571), .Y(n14224));
INVX1 mul_U8207(.A(n14224), .Y(n1254));
AND2X1 mul_U8208(.A(n7738), .B(n8572), .Y(n14227));
INVX1 mul_U8209(.A(n14227), .Y(n1255));
AND2X1 mul_U8210(.A(n7739), .B(n8573), .Y(n14230));
INVX1 mul_U8211(.A(n14230), .Y(n1256));
AND2X1 mul_U8212(.A(n7740), .B(n8574), .Y(n14233));
INVX1 mul_U8213(.A(n14233), .Y(n1257));
AND2X1 mul_U8214(.A(n7741), .B(n8575), .Y(n14236));
INVX1 mul_U8215(.A(n14236), .Y(n1258));
AND2X1 mul_U8216(.A(n7742), .B(n8576), .Y(n14239));
INVX1 mul_U8217(.A(n14239), .Y(n1259));
AND2X1 mul_U8218(.A(n7743), .B(n8577), .Y(n14242));
INVX1 mul_U8219(.A(n14242), .Y(n1260));
AND2X1 mul_U8220(.A(n7744), .B(n8578), .Y(n14245));
INVX1 mul_U8221(.A(n14245), .Y(n1261));
AND2X1 mul_U8222(.A(n7745), .B(n8579), .Y(n14248));
INVX1 mul_U8223(.A(n14248), .Y(n1262));
AND2X1 mul_U8224(.A(n7746), .B(n8580), .Y(n14251));
INVX1 mul_U8225(.A(n14251), .Y(n1263));
AND2X1 mul_U8226(.A(n7747), .B(n8581), .Y(n14254));
INVX1 mul_U8227(.A(n14254), .Y(n1264));
AND2X1 mul_U8228(.A(n7748), .B(n8582), .Y(n14257));
INVX1 mul_U8229(.A(n14257), .Y(n1265));
AND2X1 mul_U8230(.A(n7749), .B(n8583), .Y(n14260));
INVX1 mul_U8231(.A(n14260), .Y(n1266));
AND2X1 mul_U8232(.A(n7750), .B(n8584), .Y(n14263));
INVX1 mul_U8233(.A(n14263), .Y(n1267));
AND2X1 mul_U8234(.A(n7751), .B(n8585), .Y(n14266));
INVX1 mul_U8235(.A(n14266), .Y(n1268));
AND2X1 mul_U8236(.A(n7752), .B(n8586), .Y(n14269));
INVX1 mul_U8237(.A(n14269), .Y(n1269));
AND2X1 mul_U8238(.A(n7753), .B(n8587), .Y(n14272));
INVX1 mul_U8239(.A(n14272), .Y(n1270));
AND2X1 mul_U8240(.A(n7754), .B(n8588), .Y(n14275));
INVX1 mul_U8241(.A(n14275), .Y(n1271));
AND2X1 mul_U8242(.A(n7755), .B(n8589), .Y(n14278));
INVX1 mul_U8243(.A(n14278), .Y(n1272));
AND2X1 mul_U8244(.A(n7756), .B(n8590), .Y(n14281));
INVX1 mul_U8245(.A(n14281), .Y(n1273));
AND2X1 mul_U8246(.A(n7757), .B(n8591), .Y(n14284));
INVX1 mul_U8247(.A(n14284), .Y(n1274));
AND2X1 mul_U8248(.A(n7758), .B(n8592), .Y(n14287));
INVX1 mul_U8249(.A(n14287), .Y(n1275));
AND2X1 mul_U8250(.A(n7759), .B(n8593), .Y(n14290));
INVX1 mul_U8251(.A(n14290), .Y(n1276));
AND2X1 mul_U8252(.A(n7760), .B(n8594), .Y(n14293));
INVX1 mul_U8253(.A(n14293), .Y(n1277));
AND2X1 mul_U8254(.A(n7761), .B(n8595), .Y(n14296));
INVX1 mul_U8255(.A(n14296), .Y(n1278));
AND2X1 mul_U8256(.A(n7762), .B(n8596), .Y(n14299));
INVX1 mul_U8257(.A(n14299), .Y(n1279));
AND2X1 mul_U8258(.A(n7763), .B(n8597), .Y(n14302));
INVX1 mul_U8259(.A(n14302), .Y(n1280));
AND2X1 mul_U8260(.A(n7764), .B(n8598), .Y(n14305));
INVX1 mul_U8261(.A(n14305), .Y(n1281));
AND2X1 mul_U8262(.A(n7765), .B(n8599), .Y(n14308));
INVX1 mul_U8263(.A(n14308), .Y(n1282));
AND2X1 mul_U8264(.A(n7766), .B(n8600), .Y(n14311));
INVX1 mul_U8265(.A(n14311), .Y(n1283));
AND2X1 mul_U8266(.A(n7767), .B(n8601), .Y(n14314));
INVX1 mul_U8267(.A(n14314), .Y(n1284));
AND2X1 mul_U8268(.A(n7768), .B(n8602), .Y(n14317));
INVX1 mul_U8269(.A(n14317), .Y(n1285));
AND2X1 mul_U8270(.A(n7769), .B(n8603), .Y(n14320));
INVX1 mul_U8271(.A(n14320), .Y(n1286));
AND2X1 mul_U8272(.A(n7770), .B(n8604), .Y(n14323));
INVX1 mul_U8273(.A(n14323), .Y(n1287));
AND2X1 mul_U8274(.A(n7771), .B(n8605), .Y(n14326));
INVX1 mul_U8275(.A(n14326), .Y(n1288));
AND2X1 mul_U8276(.A(n7772), .B(n8606), .Y(n14329));
INVX1 mul_U8277(.A(n14329), .Y(n1289));
AND2X1 mul_U8278(.A(n7773), .B(n8607), .Y(n14332));
INVX1 mul_U8279(.A(n14332), .Y(n1290));
AND2X1 mul_U8280(.A(n7774), .B(n8608), .Y(n14335));
INVX1 mul_U8281(.A(n14335), .Y(n1291));
AND2X1 mul_U8282(.A(n7775), .B(n8609), .Y(n14338));
INVX1 mul_U8283(.A(n14338), .Y(n1292));
AND2X1 mul_U8284(.A(n7776), .B(n8610), .Y(n14341));
INVX1 mul_U8285(.A(n14341), .Y(n1293));
AND2X1 mul_U8286(.A(n7777), .B(n8611), .Y(n14344));
INVX1 mul_U8287(.A(n14344), .Y(n1294));
AND2X1 mul_U8288(.A(n7778), .B(n8612), .Y(n14347));
INVX1 mul_U8289(.A(n14347), .Y(n1295));
AND2X1 mul_U8290(.A(n7779), .B(n8613), .Y(n14350));
INVX1 mul_U8291(.A(n14350), .Y(n1296));
AND2X1 mul_U8292(.A(n7780), .B(n8614), .Y(n14353));
INVX1 mul_U8293(.A(n14353), .Y(n1297));
AND2X1 mul_U8294(.A(n7781), .B(n8615), .Y(n14356));
INVX1 mul_U8295(.A(n14356), .Y(n1298));
AND2X1 mul_U8296(.A(n7782), .B(n8616), .Y(n14359));
INVX1 mul_U8297(.A(n14359), .Y(n1299));
AND2X1 mul_U8298(.A(n7783), .B(n8617), .Y(n14362));
INVX1 mul_U8299(.A(n14362), .Y(n1300));
AND2X1 mul_U8300(.A(n7784), .B(n8618), .Y(n14365));
INVX1 mul_U8301(.A(n14365), .Y(n1301));
AND2X1 mul_U8302(.A(n7785), .B(n8619), .Y(n14368));
INVX1 mul_U8303(.A(n14368), .Y(n1302));
AND2X1 mul_U8304(.A(n7786), .B(n8620), .Y(n14371));
INVX1 mul_U8305(.A(n14371), .Y(n1303));
AND2X1 mul_U8306(.A(n7787), .B(n8621), .Y(n14374));
INVX1 mul_U8307(.A(n14374), .Y(n1304));
AND2X1 mul_U8308(.A(n7788), .B(n8622), .Y(n14377));
INVX1 mul_U8309(.A(n14377), .Y(n1305));
AND2X1 mul_U8310(.A(n7789), .B(n8623), .Y(n14380));
INVX1 mul_U8311(.A(n14380), .Y(n1306));
AND2X1 mul_U8312(.A(n7790), .B(n8624), .Y(n14383));
INVX1 mul_U8313(.A(n14383), .Y(n1307));
AND2X1 mul_U8314(.A(n7791), .B(n8625), .Y(n14386));
INVX1 mul_U8315(.A(n14386), .Y(n1308));
AND2X1 mul_U8316(.A(n7792), .B(n8626), .Y(n14389));
INVX1 mul_U8317(.A(n14389), .Y(n1309));
AND2X1 mul_U8318(.A(n7793), .B(n8627), .Y(n14392));
INVX1 mul_U8319(.A(n14392), .Y(n1310));
AND2X1 mul_U8320(.A(n7794), .B(n8628), .Y(n14395));
INVX1 mul_U8321(.A(n14395), .Y(n1311));
AND2X1 mul_U8322(.A(n7795), .B(n8629), .Y(n14398));
INVX1 mul_U8323(.A(n14398), .Y(n1312));
AND2X1 mul_U8324(.A(n7796), .B(n8630), .Y(n14401));
INVX1 mul_U8325(.A(n14401), .Y(n1313));
AND2X1 mul_U8326(.A(n7806), .B(n8632), .Y(n14404));
INVX1 mul_U8327(.A(n14404), .Y(n1314));
AND2X1 mul_U8328(.A(n7808), .B(n8633), .Y(n14407));
INVX1 mul_U8329(.A(n14407), .Y(n1315));
AND2X1 mul_U8330(.A(n7810), .B(n8634), .Y(n14410));
INVX1 mul_U8331(.A(n14410), .Y(n1316));
AND2X1 mul_U8332(.A(n7812), .B(n8635), .Y(n14413));
INVX1 mul_U8333(.A(n14413), .Y(n1317));
AND2X1 mul_U8334(.A(n7814), .B(n8636), .Y(n14416));
INVX1 mul_U8335(.A(n14416), .Y(n1318));
AND2X1 mul_U8336(.A(n7816), .B(n8637), .Y(n14419));
INVX1 mul_U8337(.A(n14419), .Y(n1319));
AND2X1 mul_U8338(.A(n7818), .B(n8638), .Y(n14422));
INVX1 mul_U8339(.A(n14422), .Y(n1320));
AND2X1 mul_U8340(.A(n7820), .B(n8639), .Y(n14425));
INVX1 mul_U8341(.A(n14425), .Y(n1321));
AND2X1 mul_U8342(.A(n7822), .B(n8640), .Y(n14428));
INVX1 mul_U8343(.A(n14428), .Y(n1322));
AND2X1 mul_U8344(.A(n7824), .B(n8641), .Y(n14431));
INVX1 mul_U8345(.A(n14431), .Y(n1323));
AND2X1 mul_U8346(.A(n7826), .B(n8642), .Y(n14434));
INVX1 mul_U8347(.A(n14434), .Y(n1324));
AND2X1 mul_U8348(.A(n7828), .B(n8643), .Y(n14437));
INVX1 mul_U8349(.A(n14437), .Y(n1325));
AND2X1 mul_U8350(.A(n7830), .B(n8644), .Y(n14440));
INVX1 mul_U8351(.A(n14440), .Y(n1326));
AND2X1 mul_U8352(.A(n7832), .B(n8645), .Y(n14443));
INVX1 mul_U8353(.A(n14443), .Y(n1327));
AND2X1 mul_U8354(.A(n7834), .B(n8646), .Y(n14446));
INVX1 mul_U8355(.A(n14446), .Y(n1328));
AND2X1 mul_U8356(.A(n7836), .B(n8647), .Y(n14449));
INVX1 mul_U8357(.A(n14449), .Y(n1329));
AND2X1 mul_U8358(.A(n7838), .B(n8648), .Y(n14452));
INVX1 mul_U8359(.A(n14452), .Y(n1330));
AND2X1 mul_U8360(.A(n7840), .B(n8649), .Y(n14455));
INVX1 mul_U8361(.A(n14455), .Y(n1331));
AND2X1 mul_U8362(.A(n7842), .B(n8650), .Y(n14458));
INVX1 mul_U8363(.A(n14458), .Y(n1332));
AND2X1 mul_U8364(.A(n7844), .B(n8651), .Y(n14461));
INVX1 mul_U8365(.A(n14461), .Y(n1333));
AND2X1 mul_U8366(.A(n7846), .B(n8652), .Y(n14464));
INVX1 mul_U8367(.A(n14464), .Y(n1334));
AND2X1 mul_U8368(.A(n7848), .B(n8653), .Y(n14467));
INVX1 mul_U8369(.A(n14467), .Y(n1335));
AND2X1 mul_U8370(.A(n7850), .B(n8654), .Y(n14470));
INVX1 mul_U8371(.A(n14470), .Y(n1336));
AND2X1 mul_U8372(.A(n7852), .B(n8655), .Y(n14473));
INVX1 mul_U8373(.A(n14473), .Y(n1337));
AND2X1 mul_U8374(.A(n7854), .B(n8656), .Y(n14476));
INVX1 mul_U8375(.A(n14476), .Y(n1338));
AND2X1 mul_U8376(.A(n7856), .B(n8657), .Y(n14479));
INVX1 mul_U8377(.A(n14479), .Y(n1339));
AND2X1 mul_U8378(.A(n7858), .B(n8658), .Y(n14482));
INVX1 mul_U8379(.A(n14482), .Y(n1340));
AND2X1 mul_U8380(.A(n7860), .B(n8659), .Y(n14485));
INVX1 mul_U8381(.A(n14485), .Y(n1341));
AND2X1 mul_U8382(.A(n7862), .B(n8660), .Y(n14488));
INVX1 mul_U8383(.A(n14488), .Y(n1342));
AND2X1 mul_U8384(.A(n7864), .B(n8661), .Y(n14491));
INVX1 mul_U8385(.A(n14491), .Y(n1343));
AND2X1 mul_U8386(.A(n7866), .B(n8662), .Y(n14494));
INVX1 mul_U8387(.A(n14494), .Y(n1344));
AND2X1 mul_U8388(.A(n7868), .B(n8663), .Y(n14497));
INVX1 mul_U8389(.A(n14497), .Y(n1345));
AND2X1 mul_U8390(.A(n7870), .B(n8664), .Y(n14500));
INVX1 mul_U8391(.A(n14500), .Y(n1346));
AND2X1 mul_U8392(.A(n7872), .B(n8665), .Y(n14503));
INVX1 mul_U8393(.A(n14503), .Y(n1347));
AND2X1 mul_U8394(.A(n7874), .B(n8666), .Y(n14506));
INVX1 mul_U8395(.A(n14506), .Y(n1348));
AND2X1 mul_U8396(.A(n7876), .B(n8667), .Y(n14509));
INVX1 mul_U8397(.A(n14509), .Y(n1349));
AND2X1 mul_U8398(.A(n7878), .B(n8668), .Y(n14512));
INVX1 mul_U8399(.A(n14512), .Y(n1350));
AND2X1 mul_U8400(.A(n7880), .B(n8669), .Y(n14515));
INVX1 mul_U8401(.A(n14515), .Y(n1351));
AND2X1 mul_U8402(.A(n7882), .B(n8670), .Y(n14518));
INVX1 mul_U8403(.A(n14518), .Y(n1352));
AND2X1 mul_U8404(.A(n7884), .B(n8671), .Y(n14521));
INVX1 mul_U8405(.A(n14521), .Y(n1353));
AND2X1 mul_U8406(.A(n7886), .B(n8672), .Y(n14524));
INVX1 mul_U8407(.A(n14524), .Y(n1354));
AND2X1 mul_U8408(.A(n7888), .B(n8673), .Y(n14527));
INVX1 mul_U8409(.A(n14527), .Y(n1355));
AND2X1 mul_U8410(.A(n7890), .B(n8674), .Y(n14530));
INVX1 mul_U8411(.A(n14530), .Y(n1356));
AND2X1 mul_U8412(.A(n7892), .B(n8675), .Y(n14533));
INVX1 mul_U8413(.A(n14533), .Y(n1357));
AND2X1 mul_U8414(.A(n7894), .B(n8676), .Y(n14536));
INVX1 mul_U8415(.A(n14536), .Y(n1358));
AND2X1 mul_U8416(.A(n7896), .B(n8677), .Y(n14539));
INVX1 mul_U8417(.A(n14539), .Y(n1359));
AND2X1 mul_U8418(.A(n7898), .B(n8678), .Y(n14542));
INVX1 mul_U8419(.A(n14542), .Y(n1360));
AND2X1 mul_U8420(.A(n7900), .B(n8679), .Y(n14545));
INVX1 mul_U8421(.A(n14545), .Y(n1361));
AND2X1 mul_U8422(.A(n7902), .B(n8680), .Y(n14548));
INVX1 mul_U8423(.A(n14548), .Y(n1362));
AND2X1 mul_U8424(.A(n7904), .B(n8681), .Y(n14551));
INVX1 mul_U8425(.A(n14551), .Y(n1363));
AND2X1 mul_U8426(.A(n7906), .B(n8682), .Y(n14554));
INVX1 mul_U8427(.A(n14554), .Y(n1364));
AND2X1 mul_U8428(.A(n7908), .B(n8683), .Y(n14557));
INVX1 mul_U8429(.A(n14557), .Y(n1365));
AND2X1 mul_U8430(.A(n7910), .B(n8684), .Y(n14560));
INVX1 mul_U8431(.A(n14560), .Y(n1366));
AND2X1 mul_U8432(.A(n7912), .B(n8685), .Y(n14563));
INVX1 mul_U8433(.A(n14563), .Y(n1367));
AND2X1 mul_U8434(.A(n7914), .B(n8686), .Y(n14566));
INVX1 mul_U8435(.A(n14566), .Y(n1368));
AND2X1 mul_U8436(.A(n7916), .B(n8687), .Y(n14569));
INVX1 mul_U8437(.A(n14569), .Y(n1369));
AND2X1 mul_U8438(.A(n7918), .B(n8688), .Y(n14572));
INVX1 mul_U8439(.A(n14572), .Y(n1370));
AND2X1 mul_U8440(.A(n7920), .B(n8689), .Y(n14575));
INVX1 mul_U8441(.A(n14575), .Y(n1371));
AND2X1 mul_U8442(.A(n7922), .B(n8690), .Y(n14578));
INVX1 mul_U8443(.A(n14578), .Y(n1372));
AND2X1 mul_U8444(.A(n7923), .B(n8691), .Y(n14581));
INVX1 mul_U8445(.A(n14581), .Y(n1373));
AND2X1 mul_U8446(.A(n7933), .B(n8693), .Y(n14584));
INVX1 mul_U8447(.A(n14584), .Y(n1374));
AND2X1 mul_U8448(.A(n7935), .B(n8694), .Y(n14587));
INVX1 mul_U8449(.A(n14587), .Y(n1375));
AND2X1 mul_U8450(.A(n7937), .B(n8695), .Y(n14590));
INVX1 mul_U8451(.A(n14590), .Y(n1376));
AND2X1 mul_U8452(.A(n7939), .B(n8696), .Y(n14593));
INVX1 mul_U8453(.A(n14593), .Y(n1377));
AND2X1 mul_U8454(.A(n7941), .B(n8697), .Y(n14596));
INVX1 mul_U8455(.A(n14596), .Y(n1378));
AND2X1 mul_U8456(.A(n7943), .B(n8698), .Y(n14599));
INVX1 mul_U8457(.A(n14599), .Y(n1379));
AND2X1 mul_U8458(.A(n7945), .B(n8699), .Y(n14602));
INVX1 mul_U8459(.A(n14602), .Y(n1380));
AND2X1 mul_U8460(.A(n7947), .B(n8700), .Y(n14605));
INVX1 mul_U8461(.A(n14605), .Y(n1381));
AND2X1 mul_U8462(.A(n7949), .B(n8701), .Y(n14608));
INVX1 mul_U8463(.A(n14608), .Y(n1382));
AND2X1 mul_U8464(.A(n7951), .B(n8702), .Y(n14611));
INVX1 mul_U8465(.A(n14611), .Y(n1383));
AND2X1 mul_U8466(.A(n7953), .B(n8703), .Y(n14614));
INVX1 mul_U8467(.A(n14614), .Y(n1384));
AND2X1 mul_U8468(.A(n7955), .B(n8704), .Y(n14617));
INVX1 mul_U8469(.A(n14617), .Y(n1385));
AND2X1 mul_U8470(.A(n7957), .B(n8705), .Y(n14620));
INVX1 mul_U8471(.A(n14620), .Y(n1386));
AND2X1 mul_U8472(.A(n7959), .B(n8706), .Y(n14623));
INVX1 mul_U8473(.A(n14623), .Y(n1387));
AND2X1 mul_U8474(.A(n7961), .B(n8707), .Y(n14626));
INVX1 mul_U8475(.A(n14626), .Y(n1388));
AND2X1 mul_U8476(.A(n7963), .B(n8708), .Y(n14629));
INVX1 mul_U8477(.A(n14629), .Y(n1389));
AND2X1 mul_U8478(.A(n7965), .B(n8709), .Y(n14632));
INVX1 mul_U8479(.A(n14632), .Y(n1390));
AND2X1 mul_U8480(.A(n7967), .B(n8710), .Y(n14635));
INVX1 mul_U8481(.A(n14635), .Y(n1391));
AND2X1 mul_U8482(.A(n7969), .B(n8711), .Y(n14638));
INVX1 mul_U8483(.A(n14638), .Y(n1392));
AND2X1 mul_U8484(.A(n7971), .B(n8712), .Y(n14641));
INVX1 mul_U8485(.A(n14641), .Y(n1393));
AND2X1 mul_U8486(.A(n7973), .B(n8713), .Y(n14644));
INVX1 mul_U8487(.A(n14644), .Y(n1394));
AND2X1 mul_U8488(.A(n7975), .B(n8714), .Y(n14647));
INVX1 mul_U8489(.A(n14647), .Y(n1395));
AND2X1 mul_U8490(.A(n7977), .B(n8715), .Y(n14650));
INVX1 mul_U8491(.A(n14650), .Y(n1396));
AND2X1 mul_U8492(.A(n7979), .B(n8716), .Y(n14653));
INVX1 mul_U8493(.A(n14653), .Y(n1397));
AND2X1 mul_U8494(.A(n7981), .B(n8717), .Y(n14656));
INVX1 mul_U8495(.A(n14656), .Y(n1398));
AND2X1 mul_U8496(.A(n7983), .B(n8718), .Y(n14659));
INVX1 mul_U8497(.A(n14659), .Y(n1399));
AND2X1 mul_U8498(.A(n7985), .B(n8719), .Y(n14662));
INVX1 mul_U8499(.A(n14662), .Y(n1400));
AND2X1 mul_U8500(.A(n7987), .B(n8720), .Y(n14665));
INVX1 mul_U8501(.A(n14665), .Y(n1401));
AND2X1 mul_U8502(.A(n7989), .B(n8721), .Y(n14668));
INVX1 mul_U8503(.A(n14668), .Y(n1402));
AND2X1 mul_U8504(.A(n7991), .B(n8722), .Y(n14671));
INVX1 mul_U8505(.A(n14671), .Y(n1403));
AND2X1 mul_U8506(.A(n7993), .B(n8723), .Y(n14674));
INVX1 mul_U8507(.A(n14674), .Y(n1404));
AND2X1 mul_U8508(.A(n7995), .B(n8724), .Y(n14677));
INVX1 mul_U8509(.A(n14677), .Y(n1405));
AND2X1 mul_U8510(.A(n7997), .B(n8725), .Y(n14680));
INVX1 mul_U8511(.A(n14680), .Y(n1406));
AND2X1 mul_U8512(.A(n7999), .B(n8726), .Y(n14683));
INVX1 mul_U8513(.A(n14683), .Y(n1407));
AND2X1 mul_U8514(.A(n8001), .B(n8727), .Y(n14686));
INVX1 mul_U8515(.A(n14686), .Y(n1408));
AND2X1 mul_U8516(.A(n8003), .B(n8728), .Y(n14689));
INVX1 mul_U8517(.A(n14689), .Y(n1409));
AND2X1 mul_U8518(.A(n8005), .B(n8729), .Y(n14692));
INVX1 mul_U8519(.A(n14692), .Y(n1410));
AND2X1 mul_U8520(.A(n8007), .B(n8730), .Y(n14695));
INVX1 mul_U8521(.A(n14695), .Y(n1411));
AND2X1 mul_U8522(.A(n8009), .B(n8731), .Y(n14698));
INVX1 mul_U8523(.A(n14698), .Y(n1412));
AND2X1 mul_U8524(.A(n8011), .B(n8732), .Y(n14701));
INVX1 mul_U8525(.A(n14701), .Y(n1413));
AND2X1 mul_U8526(.A(n8013), .B(n8733), .Y(n14704));
INVX1 mul_U8527(.A(n14704), .Y(n1414));
AND2X1 mul_U8528(.A(n8015), .B(n8734), .Y(n14707));
INVX1 mul_U8529(.A(n14707), .Y(n1415));
AND2X1 mul_U8530(.A(n8017), .B(n8735), .Y(n14710));
INVX1 mul_U8531(.A(n14710), .Y(n1416));
AND2X1 mul_U8532(.A(n8019), .B(n8736), .Y(n14713));
INVX1 mul_U8533(.A(n14713), .Y(n1417));
AND2X1 mul_U8534(.A(n8021), .B(n8737), .Y(n14716));
INVX1 mul_U8535(.A(n14716), .Y(n1418));
AND2X1 mul_U8536(.A(n8023), .B(n8738), .Y(n14719));
INVX1 mul_U8537(.A(n14719), .Y(n1419));
AND2X1 mul_U8538(.A(n8025), .B(n8739), .Y(n14722));
INVX1 mul_U8539(.A(n14722), .Y(n1420));
AND2X1 mul_U8540(.A(n8027), .B(n8740), .Y(n14725));
INVX1 mul_U8541(.A(n14725), .Y(n1421));
AND2X1 mul_U8542(.A(n8029), .B(n8741), .Y(n14728));
INVX1 mul_U8543(.A(n14728), .Y(n1422));
AND2X1 mul_U8544(.A(n8031), .B(n8742), .Y(n14731));
INVX1 mul_U8545(.A(n14731), .Y(n1423));
AND2X1 mul_U8546(.A(n8033), .B(n8743), .Y(n14734));
INVX1 mul_U8547(.A(n14734), .Y(n1424));
AND2X1 mul_U8548(.A(n8035), .B(n8744), .Y(n14737));
INVX1 mul_U8549(.A(n14737), .Y(n1425));
AND2X1 mul_U8550(.A(n8037), .B(n8745), .Y(n14740));
INVX1 mul_U8551(.A(n14740), .Y(n1426));
AND2X1 mul_U8552(.A(n8039), .B(n8746), .Y(n14743));
INVX1 mul_U8553(.A(n14743), .Y(n1427));
AND2X1 mul_U8554(.A(n8041), .B(n8747), .Y(n14746));
INVX1 mul_U8555(.A(n14746), .Y(n1428));
AND2X1 mul_U8556(.A(n8043), .B(n8748), .Y(n14749));
INVX1 mul_U8557(.A(n14749), .Y(n1429));
AND2X1 mul_U8558(.A(n8045), .B(n8749), .Y(n14752));
INVX1 mul_U8559(.A(n14752), .Y(n1430));
AND2X1 mul_U8560(.A(n8047), .B(n8750), .Y(n14755));
INVX1 mul_U8561(.A(n14755), .Y(n1431));
AND2X1 mul_U8562(.A(n8049), .B(n8751), .Y(n14758));
INVX1 mul_U8563(.A(n14758), .Y(n1432));
AND2X1 mul_U8564(.A(n8050), .B(n8752), .Y(n14761));
INVX1 mul_U8565(.A(n14761), .Y(n1433));
AND2X1 mul_U8566(.A(n7612), .B(n8755), .Y(n14764));
INVX1 mul_U8567(.A(n14764), .Y(n1434));
AND2X1 mul_U8568(.A(n7611), .B(dpath_mulcore_ary1_a0_I0_I2_net42), .Y(n14767));
INVX1 mul_U8569(.A(n14767), .Y(n1435));
AND2X1 mul_U8570(.A(n8053), .B(n9490), .Y(n14770));
INVX1 mul_U8571(.A(n14770), .Y(n1436));
AND2X1 mul_U8572(.A(n9426), .B(dpath_mulcore_ary1_a0_I0_I2_sc1_66__b), .Y(n14773));
INVX1 mul_U8573(.A(n14773), .Y(n1437));
AND2X1 mul_U8574(.A(n7736), .B(n8756), .Y(n14776));
INVX1 mul_U8575(.A(n14776), .Y(n1438));
AND2X1 mul_U8576(.A(n7735), .B(n9477), .Y(n14779));
INVX1 mul_U8577(.A(n14779), .Y(n1439));
AND2X1 mul_U8578(.A(n7803), .B(n8757), .Y(n14784));
INVX1 mul_U8579(.A(n14784), .Y(n1440));
AND2X1 mul_U8580(.A(n7802), .B(n9479), .Y(n14787));
INVX1 mul_U8581(.A(n14787), .Y(n1441));
AND2X1 mul_U8582(.A(n7930), .B(n8758), .Y(n14792));
INVX1 mul_U8583(.A(n14792), .Y(n1442));
AND2X1 mul_U8584(.A(n7929), .B(n9481), .Y(n14795));
INVX1 mul_U8585(.A(n14795), .Y(n1443));
AND2X1 mul_U8586(.A(n9673), .B(n6102), .Y(n14799));
INVX1 mul_U8587(.A(n14799), .Y(n1444));
AND2X1 mul_U8588(.A(n9686), .B(n6103), .Y(n14801));
INVX1 mul_U8589(.A(n14801), .Y(n1445));
AND2X1 mul_U8590(.A(n9686), .B(n6104), .Y(n14803));
INVX1 mul_U8591(.A(n14803), .Y(n1446));
AND2X1 mul_U8592(.A(n9686), .B(n6105), .Y(n14805));
INVX1 mul_U8593(.A(n14805), .Y(n1447));
AND2X1 mul_U8594(.A(n9671), .B(n6106), .Y(n14807));
INVX1 mul_U8595(.A(n14807), .Y(n1448));
AND2X1 mul_U8596(.A(n9671), .B(n6107), .Y(n14809));
INVX1 mul_U8597(.A(n14809), .Y(n1449));
AND2X1 mul_U8598(.A(n9671), .B(n6108), .Y(n14811));
INVX1 mul_U8599(.A(n14811), .Y(n1450));
AND2X1 mul_U8600(.A(n9683), .B(n6109), .Y(n14813));
INVX1 mul_U8601(.A(n14813), .Y(n1451));
AND2X1 mul_U8602(.A(n9684), .B(n6110), .Y(n14815));
INVX1 mul_U8603(.A(n14815), .Y(n1452));
AND2X1 mul_U8604(.A(n9672), .B(n6111), .Y(n14817));
INVX1 mul_U8605(.A(n14817), .Y(n1453));
AND2X1 mul_U8606(.A(n9671), .B(n6112), .Y(n14819));
INVX1 mul_U8607(.A(n14819), .Y(n1454));
AND2X1 mul_U8608(.A(n9673), .B(n6113), .Y(n14821));
INVX1 mul_U8609(.A(n14821), .Y(n1455));
AND2X1 mul_U8610(.A(n9671), .B(n6114), .Y(n14823));
INVX1 mul_U8611(.A(n14823), .Y(n1456));
AND2X1 mul_U8612(.A(n9671), .B(n6115), .Y(n14825));
INVX1 mul_U8613(.A(n14825), .Y(n1457));
AND2X1 mul_U8614(.A(n9683), .B(n6116), .Y(n14827));
INVX1 mul_U8615(.A(n14827), .Y(n1458));
AND2X1 mul_U8616(.A(n9684), .B(n6117), .Y(n14829));
INVX1 mul_U8617(.A(n14829), .Y(n1459));
AND2X1 mul_U8618(.A(n9685), .B(n6118), .Y(n14831));
INVX1 mul_U8619(.A(n14831), .Y(n1460));
AND2X1 mul_U8620(.A(n9685), .B(n6119), .Y(n14833));
INVX1 mul_U8621(.A(n14833), .Y(n1461));
AND2X1 mul_U8622(.A(n9685), .B(n6120), .Y(n14835));
INVX1 mul_U8623(.A(n14835), .Y(n1462));
AND2X1 mul_U8624(.A(n9685), .B(n6121), .Y(n14837));
INVX1 mul_U8625(.A(n14837), .Y(n1463));
AND2X1 mul_U8626(.A(n9685), .B(n6122), .Y(n14839));
INVX1 mul_U8627(.A(n14839), .Y(n1464));
AND2X1 mul_U8628(.A(n9685), .B(n6123), .Y(n14841));
INVX1 mul_U8629(.A(n14841), .Y(n1465));
AND2X1 mul_U8630(.A(n9685), .B(n6124), .Y(n14843));
INVX1 mul_U8631(.A(n14843), .Y(n1466));
AND2X1 mul_U8632(.A(n9685), .B(n6125), .Y(n14845));
INVX1 mul_U8633(.A(n14845), .Y(n1467));
AND2X1 mul_U8634(.A(n9685), .B(n6126), .Y(n14847));
INVX1 mul_U8635(.A(n14847), .Y(n1468));
AND2X1 mul_U8636(.A(n9685), .B(n6127), .Y(n14849));
INVX1 mul_U8637(.A(n14849), .Y(n1469));
AND2X1 mul_U8638(.A(n9685), .B(n6128), .Y(n14851));
INVX1 mul_U8639(.A(n14851), .Y(n1470));
AND2X1 mul_U8640(.A(n9685), .B(n6129), .Y(n14853));
INVX1 mul_U8641(.A(n14853), .Y(n1471));
AND2X1 mul_U8642(.A(n9672), .B(n6130), .Y(n14855));
INVX1 mul_U8643(.A(n14855), .Y(n1472));
AND2X1 mul_U8644(.A(n9673), .B(n6131), .Y(n14857));
INVX1 mul_U8645(.A(n14857), .Y(n1473));
AND2X1 mul_U8646(.A(dpath_mulcore_x2_c2c3), .B(n6132), .Y(n14859));
INVX1 mul_U8647(.A(n14859), .Y(n1474));
AND2X1 mul_U8648(.A(n9686), .B(n6133), .Y(n14861));
INVX1 mul_U8649(.A(n14861), .Y(n1475));
AND2X1 mul_U8650(.A(n9674), .B(n6134), .Y(n14863));
INVX1 mul_U8651(.A(n14863), .Y(n1476));
AND2X1 mul_U8652(.A(n9676), .B(n6135), .Y(n14865));
INVX1 mul_U8653(.A(n14865), .Y(n1477));
AND2X1 mul_U8654(.A(n9677), .B(n6136), .Y(n14867));
INVX1 mul_U8655(.A(n14867), .Y(n1478));
AND2X1 mul_U8656(.A(n9690), .B(n6137), .Y(n14869));
INVX1 mul_U8657(.A(n14869), .Y(n1479));
AND2X1 mul_U8658(.A(n9689), .B(n6138), .Y(n14871));
INVX1 mul_U8659(.A(n14871), .Y(n1480));
AND2X1 mul_U8660(.A(n9687), .B(n6139), .Y(n14873));
INVX1 mul_U8661(.A(n14873), .Y(n1481));
AND2X1 mul_U8662(.A(n9688), .B(dpath_areg[31]), .Y(n14875));
INVX1 mul_U8663(.A(n14875), .Y(n1482));
AND2X1 mul_U8664(.A(n9673), .B(dpath_areg[30]), .Y(n14877));
INVX1 mul_U8665(.A(n14877), .Y(n1483));
AND2X1 mul_U8666(.A(n9679), .B(dpath_areg[29]), .Y(n14879));
INVX1 mul_U8667(.A(n14879), .Y(n1484));
AND2X1 mul_U8668(.A(n9671), .B(dpath_areg[28]), .Y(n14881));
INVX1 mul_U8669(.A(n14881), .Y(n1485));
AND2X1 mul_U8670(.A(n9672), .B(dpath_areg[27]), .Y(n14883));
INVX1 mul_U8671(.A(n14883), .Y(n1486));
AND2X1 mul_U8672(.A(n9673), .B(dpath_areg[26]), .Y(n14885));
INVX1 mul_U8673(.A(n14885), .Y(n1487));
AND2X1 mul_U8674(.A(dpath_mulcore_x2_c2c3), .B(dpath_areg[25]), .Y(n14887));
INVX1 mul_U8675(.A(n14887), .Y(n1488));
AND2X1 mul_U8676(.A(n9690), .B(dpath_areg[24]), .Y(n14889));
INVX1 mul_U8677(.A(n14889), .Y(n1489));
AND2X1 mul_U8678(.A(n9675), .B(dpath_areg[23]), .Y(n14891));
INVX1 mul_U8679(.A(n14891), .Y(n1490));
AND2X1 mul_U8680(.A(n9678), .B(dpath_areg[22]), .Y(n14893));
INVX1 mul_U8681(.A(n14893), .Y(n1491));
AND2X1 mul_U8682(.A(n9679), .B(dpath_areg[21]), .Y(n14895));
INVX1 mul_U8683(.A(n14895), .Y(n1492));
AND2X1 mul_U8684(.A(n9684), .B(n6075), .Y(n14898));
INVX1 mul_U8685(.A(n14898), .Y(n1493));
AND2X1 mul_U8686(.A(n9683), .B(n6076), .Y(n14900));
INVX1 mul_U8687(.A(n14900), .Y(n1494));
AND2X1 mul_U8688(.A(n9671), .B(n6077), .Y(n14902));
INVX1 mul_U8689(.A(n14902), .Y(n1495));
AND2X1 mul_U8690(.A(n9671), .B(n6078), .Y(n14904));
INVX1 mul_U8691(.A(n14904), .Y(n1496));
AND2X1 mul_U8692(.A(n9672), .B(n6079), .Y(n14906));
INVX1 mul_U8693(.A(n14906), .Y(n1497));
AND2X1 mul_U8694(.A(dpath_mulcore_x2_c2c3), .B(n6080), .Y(n14908));
INVX1 mul_U8695(.A(n14908), .Y(n1498));
AND2X1 mul_U8696(.A(n9675), .B(n6081), .Y(n14910));
INVX1 mul_U8697(.A(n14910), .Y(n1499));
AND2X1 mul_U8698(.A(n9678), .B(n6082), .Y(n14912));
INVX1 mul_U8699(.A(n14912), .Y(n1500));
AND2X1 mul_U8700(.A(n9679), .B(n6083), .Y(n14914));
INVX1 mul_U8701(.A(n14914), .Y(n1501));
AND2X1 mul_U8702(.A(n9671), .B(n6084), .Y(n14916));
INVX1 mul_U8703(.A(n14916), .Y(n1502));
AND2X1 mul_U8704(.A(n9672), .B(n6085), .Y(n14918));
INVX1 mul_U8705(.A(n14918), .Y(n1503));
AND2X1 mul_U8706(.A(dpath_mulcore_x2_c2c3), .B(n6086), .Y(n14920));
INVX1 mul_U8707(.A(n14920), .Y(n1504));
AND2X1 mul_U8708(.A(n9675), .B(dpath_areg[1]), .Y(n14922));
INVX1 mul_U8709(.A(n14922), .Y(n1505));
AND2X1 mul_U8710(.A(n9678), .B(n6089), .Y(n14924));
INVX1 mul_U8711(.A(n14924), .Y(n1506));
AND2X1 mul_U8712(.A(n9672), .B(n6090), .Y(n14926));
INVX1 mul_U8713(.A(n14926), .Y(n1507));
AND2X1 mul_U8714(.A(n9672), .B(n6091), .Y(n14928));
INVX1 mul_U8715(.A(n14928), .Y(n1508));
AND2X1 mul_U8716(.A(n9672), .B(n6092), .Y(n14930));
INVX1 mul_U8717(.A(n14930), .Y(n1509));
AND2X1 mul_U8718(.A(n9671), .B(n6093), .Y(n14932));
INVX1 mul_U8719(.A(n14932), .Y(n1510));
AND2X1 mul_U8720(.A(n9673), .B(n6094), .Y(n14934));
INVX1 mul_U8721(.A(n14934), .Y(n1511));
AND2X1 mul_U8722(.A(n9685), .B(n6095), .Y(n14936));
INVX1 mul_U8723(.A(n14936), .Y(n1512));
AND2X1 mul_U8724(.A(n9685), .B(n6096), .Y(n14938));
INVX1 mul_U8725(.A(n14938), .Y(n1513));
AND2X1 mul_U8726(.A(n9686), .B(n6097), .Y(n14940));
INVX1 mul_U8727(.A(n14940), .Y(n1514));
AND2X1 mul_U8728(.A(n9673), .B(n6098), .Y(n14942));
INVX1 mul_U8729(.A(n14942), .Y(n1515));
AND2X1 mul_U8730(.A(dpath_mulcore_x2_c2c3), .B(n6099), .Y(n14944));
INVX1 mul_U8731(.A(n14944), .Y(n1516));
AND2X1 mul_U8732(.A(n9674), .B(n6100), .Y(n14946));
INVX1 mul_U8733(.A(n14946), .Y(n1517));
AND2X1 mul_U8734(.A(n9675), .B(n6101), .Y(n14948));
INVX1 mul_U8735(.A(n14948), .Y(n1518));
AND2X1 mul_U8736(.A(n9684), .B(dpath_areg[20]), .Y(n14950));
INVX1 mul_U8737(.A(n14950), .Y(n1519));
AND2X1 mul_U8738(.A(n9684), .B(dpath_areg[19]), .Y(n14952));
INVX1 mul_U8739(.A(n14952), .Y(n1520));
AND2X1 mul_U8740(.A(n9684), .B(dpath_areg[18]), .Y(n14954));
INVX1 mul_U8741(.A(n14954), .Y(n1521));
AND2X1 mul_U8742(.A(n9684), .B(dpath_areg[17]), .Y(n14956));
INVX1 mul_U8743(.A(n14956), .Y(n1522));
AND2X1 mul_U8744(.A(n9684), .B(dpath_areg[16]), .Y(n14958));
INVX1 mul_U8745(.A(n14958), .Y(n1523));
AND2X1 mul_U8746(.A(n9684), .B(dpath_areg[5]), .Y(n14960));
INVX1 mul_U8747(.A(n14960), .Y(n1524));
AND2X1 mul_U8748(.A(n9684), .B(dpath_areg[4]), .Y(n14962));
INVX1 mul_U8749(.A(n14962), .Y(n1525));
AND2X1 mul_U8750(.A(n9684), .B(dpath_areg[3]), .Y(n14964));
INVX1 mul_U8751(.A(n14964), .Y(n1526));
AND2X1 mul_U8752(.A(n9684), .B(dpath_areg[2]), .Y(n14966));
INVX1 mul_U8753(.A(n14966), .Y(n1527));
AND2X1 mul_U8754(.A(n9684), .B(n6087), .Y(n14969));
INVX1 mul_U8755(.A(n14969), .Y(n1528));
AND2X1 mul_U8756(.A(n9684), .B(dpath_areg[15]), .Y(n14971));
INVX1 mul_U8757(.A(n14971), .Y(n1529));
AND2X1 mul_U8758(.A(n9683), .B(dpath_areg[14]), .Y(n14973));
INVX1 mul_U8759(.A(n14973), .Y(n1530));
AND2X1 mul_U8760(.A(n9683), .B(dpath_areg[13]), .Y(n14975));
INVX1 mul_U8761(.A(n14975), .Y(n1531));
AND2X1 mul_U8762(.A(n9683), .B(dpath_areg[12]), .Y(n14977));
INVX1 mul_U8763(.A(n14977), .Y(n1532));
AND2X1 mul_U8764(.A(n9683), .B(dpath_areg[11]), .Y(n14979));
INVX1 mul_U8765(.A(n14979), .Y(n1533));
AND2X1 mul_U8766(.A(n9683), .B(dpath_areg[10]), .Y(n14981));
INVX1 mul_U8767(.A(n14981), .Y(n1534));
AND2X1 mul_U8768(.A(n9683), .B(dpath_areg[9]), .Y(n14983));
INVX1 mul_U8769(.A(n14983), .Y(n1535));
AND2X1 mul_U8770(.A(n9683), .B(dpath_areg[8]), .Y(n14985));
INVX1 mul_U8771(.A(n14985), .Y(n1536));
AND2X1 mul_U8772(.A(n9683), .B(dpath_areg[7]), .Y(n14987));
INVX1 mul_U8773(.A(n14987), .Y(n1537));
AND2X1 mul_U8774(.A(n9683), .B(dpath_areg[6]), .Y(n14989));
INVX1 mul_U8775(.A(n14989), .Y(n1538));
AND2X1 mul_U8776(.A(n13756), .B(n13757), .Y(n14992));
INVX1 mul_U8777(.A(n14992), .Y(n1539));
AND2X1 mul_U8778(.A(n13758), .B(n13759), .Y(n14995));
INVX1 mul_U8779(.A(n14995), .Y(n1540));
AND2X1 mul_U8780(.A(n13760), .B(n13761), .Y(n14998));
INVX1 mul_U8781(.A(n14998), .Y(n1541));
AND2X1 mul_U8782(.A(n13762), .B(n13763), .Y(n15001));
INVX1 mul_U8783(.A(n15001), .Y(n1542));
AND2X1 mul_U8784(.A(n13764), .B(n13765), .Y(n15004));
INVX1 mul_U8785(.A(n15004), .Y(n1543));
AND2X1 mul_U8786(.A(n13766), .B(n13767), .Y(n15007));
INVX1 mul_U8787(.A(n15007), .Y(n1544));
AND2X1 mul_U8788(.A(n13768), .B(n13769), .Y(n15010));
INVX1 mul_U8789(.A(n15010), .Y(n1545));
AND2X1 mul_U8790(.A(n13770), .B(n13771), .Y(n15013));
INVX1 mul_U8791(.A(n15013), .Y(n1546));
AND2X1 mul_U8792(.A(n13772), .B(n13773), .Y(n15016));
INVX1 mul_U8793(.A(n15016), .Y(n1547));
AND2X1 mul_U8794(.A(n13774), .B(n13775), .Y(n15019));
INVX1 mul_U8795(.A(n15019), .Y(n1548));
AND2X1 mul_U8796(.A(n13776), .B(n13777), .Y(n15022));
INVX1 mul_U8797(.A(n15022), .Y(n1549));
AND2X1 mul_U8798(.A(n13778), .B(n13779), .Y(n15025));
INVX1 mul_U8799(.A(n15025), .Y(n1550));
AND2X1 mul_U8800(.A(n13780), .B(n13781), .Y(n15028));
INVX1 mul_U8801(.A(n15028), .Y(n1551));
AND2X1 mul_U8802(.A(n13782), .B(n13783), .Y(n15031));
INVX1 mul_U8803(.A(n15031), .Y(n1552));
AND2X1 mul_U8804(.A(n13784), .B(n13785), .Y(n15034));
INVX1 mul_U8805(.A(n15034), .Y(n1553));
AND2X1 mul_U8806(.A(n13786), .B(n13787), .Y(n15037));
INVX1 mul_U8807(.A(n15037), .Y(n1554));
AND2X1 mul_U8808(.A(n13788), .B(n13789), .Y(n15040));
INVX1 mul_U8809(.A(n15040), .Y(n1555));
AND2X1 mul_U8810(.A(n13790), .B(n13791), .Y(n15043));
INVX1 mul_U8811(.A(n15043), .Y(n1556));
AND2X1 mul_U8812(.A(n13792), .B(n13793), .Y(n15046));
INVX1 mul_U8813(.A(n15046), .Y(n1557));
AND2X1 mul_U8814(.A(n13794), .B(n13795), .Y(n15049));
INVX1 mul_U8815(.A(n15049), .Y(n1558));
AND2X1 mul_U8816(.A(n13796), .B(n13797), .Y(n15052));
INVX1 mul_U8817(.A(n15052), .Y(n1559));
AND2X1 mul_U8818(.A(n13798), .B(n13799), .Y(n15055));
INVX1 mul_U8819(.A(n15055), .Y(n1560));
AND2X1 mul_U8820(.A(n13800), .B(n13801), .Y(n15058));
INVX1 mul_U8821(.A(n15058), .Y(n1561));
AND2X1 mul_U8822(.A(n13802), .B(n13803), .Y(n15061));
INVX1 mul_U8823(.A(n15061), .Y(n1562));
AND2X1 mul_U8824(.A(n13804), .B(n13805), .Y(n15064));
INVX1 mul_U8825(.A(n15064), .Y(n1563));
AND2X1 mul_U8826(.A(n13806), .B(n13807), .Y(n15067));
INVX1 mul_U8827(.A(n15067), .Y(n1564));
AND2X1 mul_U8828(.A(n13808), .B(n13809), .Y(n15070));
INVX1 mul_U8829(.A(n15070), .Y(n1565));
AND2X1 mul_U8830(.A(n13810), .B(n13811), .Y(n15073));
INVX1 mul_U8831(.A(n15073), .Y(n1566));
AND2X1 mul_U8832(.A(n13812), .B(n13813), .Y(n15076));
INVX1 mul_U8833(.A(n15076), .Y(n1567));
AND2X1 mul_U8834(.A(n13814), .B(n13815), .Y(n15079));
INVX1 mul_U8835(.A(n15079), .Y(n1568));
AND2X1 mul_U8836(.A(n13816), .B(n13817), .Y(n15082));
INVX1 mul_U8837(.A(n15082), .Y(n1569));
AND2X1 mul_U8838(.A(n13818), .B(n13819), .Y(n15085));
INVX1 mul_U8839(.A(n15085), .Y(n1570));
AND2X1 mul_U8840(.A(n13820), .B(n13821), .Y(n15088));
INVX1 mul_U8841(.A(n15088), .Y(n1571));
AND2X1 mul_U8842(.A(n13822), .B(n13823), .Y(n15091));
INVX1 mul_U8843(.A(n15091), .Y(n1572));
AND2X1 mul_U8844(.A(n13824), .B(n13825), .Y(n15094));
INVX1 mul_U8845(.A(n15094), .Y(n1573));
AND2X1 mul_U8846(.A(n13826), .B(n13827), .Y(n15097));
INVX1 mul_U8847(.A(n15097), .Y(n1574));
AND2X1 mul_U8848(.A(n13828), .B(n13829), .Y(n15100));
INVX1 mul_U8849(.A(n15100), .Y(n1575));
AND2X1 mul_U8850(.A(n13830), .B(n13831), .Y(n15103));
INVX1 mul_U8851(.A(n15103), .Y(n1576));
AND2X1 mul_U8852(.A(n13832), .B(n13833), .Y(n15106));
INVX1 mul_U8853(.A(n15106), .Y(n1577));
AND2X1 mul_U8854(.A(n13834), .B(n13835), .Y(n15109));
INVX1 mul_U8855(.A(n15109), .Y(n1578));
AND2X1 mul_U8856(.A(n13836), .B(n13837), .Y(n15112));
INVX1 mul_U8857(.A(n15112), .Y(n1579));
AND2X1 mul_U8858(.A(n13838), .B(n13839), .Y(n15115));
INVX1 mul_U8859(.A(n15115), .Y(n1580));
AND2X1 mul_U8860(.A(n13840), .B(n13841), .Y(n15118));
INVX1 mul_U8861(.A(n15118), .Y(n1581));
AND2X1 mul_U8862(.A(n13842), .B(n13843), .Y(n15121));
INVX1 mul_U8863(.A(n15121), .Y(n1582));
AND2X1 mul_U8864(.A(n13844), .B(n13845), .Y(n15124));
INVX1 mul_U8865(.A(n15124), .Y(n1583));
AND2X1 mul_U8866(.A(n13846), .B(n13847), .Y(n15127));
INVX1 mul_U8867(.A(n15127), .Y(n1584));
AND2X1 mul_U8868(.A(n13848), .B(n13849), .Y(n15130));
INVX1 mul_U8869(.A(n15130), .Y(n1585));
AND2X1 mul_U8870(.A(n13850), .B(n13851), .Y(n15133));
INVX1 mul_U8871(.A(n15133), .Y(n1586));
AND2X1 mul_U8872(.A(n13852), .B(n13853), .Y(n15136));
INVX1 mul_U8873(.A(n15136), .Y(n1587));
AND2X1 mul_U8874(.A(n13854), .B(n13855), .Y(n15139));
INVX1 mul_U8875(.A(n15139), .Y(n1588));
AND2X1 mul_U8876(.A(n13856), .B(n13857), .Y(n15142));
INVX1 mul_U8877(.A(n15142), .Y(n1589));
AND2X1 mul_U8878(.A(n13858), .B(n13859), .Y(n15145));
INVX1 mul_U8879(.A(n15145), .Y(n1590));
AND2X1 mul_U8880(.A(n13860), .B(n13861), .Y(n15148));
INVX1 mul_U8881(.A(n15148), .Y(n1591));
AND2X1 mul_U8882(.A(n13862), .B(n8976), .Y(n15151));
INVX1 mul_U8883(.A(n15151), .Y(n1592));
AND2X1 mul_U8884(.A(dpath_mulcore_ary1_a0_s2[3]), .B(n8975), .Y(n15154));
INVX1 mul_U8885(.A(n15154), .Y(n1593));
AND2X1 mul_U8886(.A(dpath_mulcore_ary1_a0_s2[2]), .B(dpath_mulcore_ary1_a0_c2[1]), .Y(n15157));
INVX1 mul_U8887(.A(n15157), .Y(n1594));
AND2X1 mul_U8888(.A(dpath_mulcore_ary1_a0_s2[1]), .B(dpath_mulcore_ary1_a0_s1[7]), .Y(n15160));
INVX1 mul_U8889(.A(n15160), .Y(n1595));
AND2X1 mul_U8890(.A(dpath_mulcore_ary1_a0_s2[0]), .B(dpath_mulcore_ary1_a0_s1[6]), .Y(n15163));
INVX1 mul_U8891(.A(n15163), .Y(n1596));
AND2X1 mul_U8892(.A(n8386), .B(dpath_mulcore_ary1_a0_s1[5]), .Y(n15166));
INVX1 mul_U8893(.A(n15166), .Y(n1597));
AND2X1 mul_U8894(.A(n8387), .B(dpath_mulcore_ary1_a0_s1[4]), .Y(n15169));
INVX1 mul_U8895(.A(n15169), .Y(n1598));
AND2X1 mul_U8896(.A(n16570), .B(n16573), .Y(n15171));
INVX1 mul_U8897(.A(n15171), .Y(n1599));
AND2X1 mul_U8898(.A(n5209), .B(n4687), .Y(dpath_mulcore_a0cout[77]));
INVX1 mul_U8899(.A(dpath_mulcore_a0cout[77]), .Y(n1600));
AND2X1 mul_U8900(.A(dpath_mulcore_ary1_a0_s0[9]), .B(n8816), .Y(n15176));
INVX1 mul_U8901(.A(n15176), .Y(n1601));
AND2X1 mul_U8902(.A(dpath_mulcore_ary1_a0_s0[8]), .B(n8817), .Y(n15179));
INVX1 mul_U8903(.A(n15179), .Y(n1602));
AND2X1 mul_U8904(.A(dpath_mulcore_ary1_a0_s0[3]), .B(n8760), .Y(n15182));
INVX1 mul_U8905(.A(n15182), .Y(n1603));
AND2X1 mul_U8906(.A(n5210), .B(n4688), .Y(dpath_mulcore_a0cout[10]));
INVX1 mul_U8907(.A(dpath_mulcore_a0cout[10]), .Y(n1604));
AND2X1 mul_U8908(.A(n5211), .B(n4689), .Y(dpath_mulcore_a0cout[9]));
INVX1 mul_U8909(.A(dpath_mulcore_a0cout[9]), .Y(n1605));
AND2X1 mul_U8910(.A(n5212), .B(n4690), .Y(dpath_mulcore_a0cout[8]));
INVX1 mul_U8911(.A(dpath_mulcore_a0cout[8]), .Y(n1606));
AND2X1 mul_U8912(.A(n13752), .B(n13753), .Y(n15194));
INVX1 mul_U8913(.A(n15194), .Y(n1607));
AND2X1 mul_U8914(.A(n16572), .B(n13745), .Y(n15197));
INVX1 mul_U8915(.A(n15197), .Y(n1608));
AND2X1 mul_U8916(.A(n13746), .B(n13747), .Y(n15200));
INVX1 mul_U8917(.A(n15200), .Y(n1609));
AND2X1 mul_U8918(.A(n13748), .B(n13749), .Y(n15203));
INVX1 mul_U8919(.A(n15203), .Y(n1610));
AND2X1 mul_U8920(.A(n13750), .B(n13751), .Y(n15206));
INVX1 mul_U8921(.A(n15206), .Y(n1611));
AND2X1 mul_U8922(.A(n9425), .B(n9488), .Y(n15209));
INVX1 mul_U8923(.A(n15209), .Y(n1612));
AND2X1 mul_U8924(.A(dpath_mulcore_ary1_a0_I0_I2_net073), .B(n8940), .Y(n15212));
INVX1 mul_U8925(.A(n15212), .Y(n1613));
AND2X1 mul_U8926(.A(dpath_mulcore_ary1_a0_s0[67]), .B(n8939), .Y(n15215));
INVX1 mul_U8927(.A(n15215), .Y(n1614));
AND2X1 mul_U8928(.A(dpath_mulcore_ary1_a0_s0[66]), .B(n8938), .Y(n15218));
INVX1 mul_U8929(.A(n15218), .Y(n1615));
AND2X1 mul_U8930(.A(dpath_mulcore_ary1_a0_s0[65]), .B(n8937), .Y(n15221));
INVX1 mul_U8931(.A(n15221), .Y(n1616));
AND2X1 mul_U8932(.A(dpath_mulcore_ary1_a0_s0[64]), .B(n8765), .Y(n15224));
INVX1 mul_U8933(.A(n15224), .Y(n1617));
AND2X1 mul_U8934(.A(dpath_mulcore_ary1_a0_s0[63]), .B(n8766), .Y(n15227));
INVX1 mul_U8935(.A(n15227), .Y(n1618));
AND2X1 mul_U8936(.A(dpath_mulcore_ary1_a0_s0[62]), .B(n8767), .Y(n15230));
INVX1 mul_U8937(.A(n15230), .Y(n1619));
AND2X1 mul_U8938(.A(dpath_mulcore_ary1_a0_s0[61]), .B(n8768), .Y(n15233));
INVX1 mul_U8939(.A(n15233), .Y(n1620));
AND2X1 mul_U8940(.A(dpath_mulcore_ary1_a0_s0[60]), .B(n8769), .Y(n15236));
INVX1 mul_U8941(.A(n15236), .Y(n1621));
AND2X1 mul_U8942(.A(dpath_mulcore_ary1_a0_s0[59]), .B(n8770), .Y(n15239));
INVX1 mul_U8943(.A(n15239), .Y(n1622));
AND2X1 mul_U8944(.A(dpath_mulcore_ary1_a0_s0[58]), .B(n8771), .Y(n15242));
INVX1 mul_U8945(.A(n15242), .Y(n1623));
AND2X1 mul_U8946(.A(dpath_mulcore_ary1_a0_s0[57]), .B(n8772), .Y(n15245));
INVX1 mul_U8947(.A(n15245), .Y(n1624));
AND2X1 mul_U8948(.A(dpath_mulcore_ary1_a0_s0[56]), .B(n8773), .Y(n15248));
INVX1 mul_U8949(.A(n15248), .Y(n1625));
AND2X1 mul_U8950(.A(dpath_mulcore_ary1_a0_s0[55]), .B(n8774), .Y(n15251));
INVX1 mul_U8951(.A(n15251), .Y(n1626));
AND2X1 mul_U8952(.A(dpath_mulcore_ary1_a0_s0[54]), .B(n8775), .Y(n15254));
INVX1 mul_U8953(.A(n15254), .Y(n1627));
AND2X1 mul_U8954(.A(dpath_mulcore_ary1_a0_s0[53]), .B(n8776), .Y(n15257));
INVX1 mul_U8955(.A(n15257), .Y(n1628));
AND2X1 mul_U8956(.A(dpath_mulcore_ary1_a0_s0[52]), .B(n8777), .Y(n15260));
INVX1 mul_U8957(.A(n15260), .Y(n1629));
AND2X1 mul_U8958(.A(dpath_mulcore_ary1_a0_s0[51]), .B(n8778), .Y(n15263));
INVX1 mul_U8959(.A(n15263), .Y(n1630));
AND2X1 mul_U8960(.A(dpath_mulcore_ary1_a0_s0[50]), .B(n8779), .Y(n15266));
INVX1 mul_U8961(.A(n15266), .Y(n1631));
AND2X1 mul_U8962(.A(dpath_mulcore_ary1_a0_s0[49]), .B(n8780), .Y(n15269));
INVX1 mul_U8963(.A(n15269), .Y(n1632));
AND2X1 mul_U8964(.A(dpath_mulcore_ary1_a0_s0[48]), .B(n8781), .Y(n15272));
INVX1 mul_U8965(.A(n15272), .Y(n1633));
AND2X1 mul_U8966(.A(dpath_mulcore_ary1_a0_s0[47]), .B(n8782), .Y(n15275));
INVX1 mul_U8967(.A(n15275), .Y(n1634));
AND2X1 mul_U8968(.A(dpath_mulcore_ary1_a0_s0[46]), .B(n8783), .Y(n15278));
INVX1 mul_U8969(.A(n15278), .Y(n1635));
AND2X1 mul_U8970(.A(dpath_mulcore_ary1_a0_s0[45]), .B(n8784), .Y(n15281));
INVX1 mul_U8971(.A(n15281), .Y(n1636));
AND2X1 mul_U8972(.A(dpath_mulcore_ary1_a0_s0[44]), .B(n8785), .Y(n15284));
INVX1 mul_U8973(.A(n15284), .Y(n1637));
AND2X1 mul_U8974(.A(dpath_mulcore_ary1_a0_s0[43]), .B(n8786), .Y(n15287));
INVX1 mul_U8975(.A(n15287), .Y(n1638));
AND2X1 mul_U8976(.A(dpath_mulcore_ary1_a0_s0[42]), .B(n8787), .Y(n15290));
INVX1 mul_U8977(.A(n15290), .Y(n1639));
AND2X1 mul_U8978(.A(dpath_mulcore_ary1_a0_s0[41]), .B(n8788), .Y(n15293));
INVX1 mul_U8979(.A(n15293), .Y(n1640));
AND2X1 mul_U8980(.A(dpath_mulcore_ary1_a0_s0[40]), .B(n8789), .Y(n15296));
INVX1 mul_U8981(.A(n15296), .Y(n1641));
AND2X1 mul_U8982(.A(dpath_mulcore_ary1_a0_s0[39]), .B(n8790), .Y(n15299));
INVX1 mul_U8983(.A(n15299), .Y(n1642));
AND2X1 mul_U8984(.A(dpath_mulcore_ary1_a0_s0[38]), .B(n8791), .Y(n15302));
INVX1 mul_U8985(.A(n15302), .Y(n1643));
AND2X1 mul_U8986(.A(dpath_mulcore_ary1_a0_s0[37]), .B(n8792), .Y(n15305));
INVX1 mul_U8987(.A(n15305), .Y(n1644));
AND2X1 mul_U8988(.A(dpath_mulcore_ary1_a0_s0[36]), .B(n8793), .Y(n15308));
INVX1 mul_U8989(.A(n15308), .Y(n1645));
AND2X1 mul_U8990(.A(dpath_mulcore_ary1_a0_s0[35]), .B(n8794), .Y(n15311));
INVX1 mul_U8991(.A(n15311), .Y(n1646));
AND2X1 mul_U8992(.A(dpath_mulcore_ary1_a0_s0[34]), .B(n8795), .Y(n15314));
INVX1 mul_U8993(.A(n15314), .Y(n1647));
AND2X1 mul_U8994(.A(dpath_mulcore_ary1_a0_s0[33]), .B(n8796), .Y(n15317));
INVX1 mul_U8995(.A(n15317), .Y(n1648));
AND2X1 mul_U8996(.A(dpath_mulcore_ary1_a0_s0[32]), .B(n8797), .Y(n15320));
INVX1 mul_U8997(.A(n15320), .Y(n1649));
AND2X1 mul_U8998(.A(dpath_mulcore_ary1_a0_s0[31]), .B(n8798), .Y(n15323));
INVX1 mul_U8999(.A(n15323), .Y(n1650));
AND2X1 mul_U9000(.A(dpath_mulcore_ary1_a0_s0[30]), .B(n8799), .Y(n15326));
INVX1 mul_U9001(.A(n15326), .Y(n1651));
AND2X1 mul_U9002(.A(dpath_mulcore_ary1_a0_s0[29]), .B(n8800), .Y(n15329));
INVX1 mul_U9003(.A(n15329), .Y(n1652));
AND2X1 mul_U9004(.A(dpath_mulcore_ary1_a0_s0[28]), .B(n8801), .Y(n15332));
INVX1 mul_U9005(.A(n15332), .Y(n1653));
AND2X1 mul_U9006(.A(dpath_mulcore_ary1_a0_s0[27]), .B(n8802), .Y(n15335));
INVX1 mul_U9007(.A(n15335), .Y(n1654));
AND2X1 mul_U9008(.A(dpath_mulcore_ary1_a0_s0[26]), .B(n8803), .Y(n15338));
INVX1 mul_U9009(.A(n15338), .Y(n1655));
AND2X1 mul_U9010(.A(dpath_mulcore_ary1_a0_s0[25]), .B(n8804), .Y(n15341));
INVX1 mul_U9011(.A(n15341), .Y(n1656));
AND2X1 mul_U9012(.A(dpath_mulcore_ary1_a0_s0[24]), .B(n8805), .Y(n15344));
INVX1 mul_U9013(.A(n15344), .Y(n1657));
AND2X1 mul_U9014(.A(dpath_mulcore_ary1_a0_s0[23]), .B(n8806), .Y(n15347));
INVX1 mul_U9015(.A(n15347), .Y(n1658));
AND2X1 mul_U9016(.A(dpath_mulcore_ary1_a0_s0[22]), .B(n8807), .Y(n15350));
INVX1 mul_U9017(.A(n15350), .Y(n1659));
AND2X1 mul_U9018(.A(dpath_mulcore_ary1_a0_s0[21]), .B(n8808), .Y(n15353));
INVX1 mul_U9019(.A(n15353), .Y(n1660));
AND2X1 mul_U9020(.A(dpath_mulcore_ary1_a0_s0[20]), .B(n8809), .Y(n15356));
INVX1 mul_U9021(.A(n15356), .Y(n1661));
AND2X1 mul_U9022(.A(dpath_mulcore_ary1_a0_s0[19]), .B(n8810), .Y(n15359));
INVX1 mul_U9023(.A(n15359), .Y(n1662));
AND2X1 mul_U9024(.A(dpath_mulcore_ary1_a0_s0[18]), .B(n8811), .Y(n15362));
INVX1 mul_U9025(.A(n15362), .Y(n1663));
AND2X1 mul_U9026(.A(dpath_mulcore_ary1_a0_s0[17]), .B(n8812), .Y(n15365));
INVX1 mul_U9027(.A(n15365), .Y(n1664));
AND2X1 mul_U9028(.A(dpath_mulcore_ary1_a0_s0[16]), .B(n8813), .Y(n15368));
INVX1 mul_U9029(.A(n15368), .Y(n1665));
AND2X1 mul_U9030(.A(dpath_mulcore_ary1_a0_s0[15]), .B(n8814), .Y(n15371));
INVX1 mul_U9031(.A(n15371), .Y(n1666));
AND2X1 mul_U9032(.A(dpath_mulcore_ary1_a0_s0[14]), .B(n8815), .Y(n15374));
INVX1 mul_U9033(.A(n15374), .Y(n1667));
AND2X1 mul_U9034(.A(dpath_mulcore_ary1_a0_s0[7]), .B(n8818), .Y(n15377));
INVX1 mul_U9035(.A(n15377), .Y(n1668));
AND2X1 mul_U9036(.A(dpath_mulcore_ary1_a0_s0[6]), .B(n8819), .Y(n15380));
INVX1 mul_U9037(.A(n15380), .Y(n1669));
AND2X1 mul_U9038(.A(dpath_mulcore_ary1_a0_s0[5]), .B(n8820), .Y(n15383));
INVX1 mul_U9039(.A(n15383), .Y(n1670));
AND2X1 mul_U9040(.A(dpath_mulcore_ary1_a0_s0[4]), .B(n8759), .Y(n15386));
INVX1 mul_U9041(.A(n15386), .Y(n1671));
AND2X1 mul_U9042(.A(dpath_mulcore_ary1_a1_s2[58]), .B(n8827), .Y(n15389));
INVX1 mul_U9043(.A(n15389), .Y(n1672));
AND2X1 mul_U9044(.A(dpath_mulcore_ary1_a1_s2[57]), .B(n8828), .Y(n15392));
INVX1 mul_U9045(.A(n15392), .Y(n1673));
AND2X1 mul_U9046(.A(dpath_mulcore_ary1_a1_s2[56]), .B(n8829), .Y(n15395));
INVX1 mul_U9047(.A(n15395), .Y(n1674));
AND2X1 mul_U9048(.A(dpath_mulcore_ary1_a1_s2[55]), .B(n8830), .Y(n15398));
INVX1 mul_U9049(.A(n15398), .Y(n1675));
AND2X1 mul_U9050(.A(dpath_mulcore_ary1_a1_s2[54]), .B(n8831), .Y(n15401));
INVX1 mul_U9051(.A(n15401), .Y(n1676));
AND2X1 mul_U9052(.A(dpath_mulcore_ary1_a1_s2[53]), .B(n8832), .Y(n15404));
INVX1 mul_U9053(.A(n15404), .Y(n1677));
AND2X1 mul_U9054(.A(dpath_mulcore_ary1_a1_s2[52]), .B(n8833), .Y(n15407));
INVX1 mul_U9055(.A(n15407), .Y(n1678));
AND2X1 mul_U9056(.A(dpath_mulcore_ary1_a1_s2[51]), .B(n8834), .Y(n15410));
INVX1 mul_U9057(.A(n15410), .Y(n1679));
AND2X1 mul_U9058(.A(dpath_mulcore_ary1_a1_s2[50]), .B(n8835), .Y(n15413));
INVX1 mul_U9059(.A(n15413), .Y(n1680));
AND2X1 mul_U9060(.A(dpath_mulcore_ary1_a1_s2[49]), .B(n8836), .Y(n15416));
INVX1 mul_U9061(.A(n15416), .Y(n1681));
AND2X1 mul_U9062(.A(dpath_mulcore_ary1_a1_s2[48]), .B(n8837), .Y(n15419));
INVX1 mul_U9063(.A(n15419), .Y(n1682));
AND2X1 mul_U9064(.A(dpath_mulcore_ary1_a1_s2[47]), .B(n8838), .Y(n15422));
INVX1 mul_U9065(.A(n15422), .Y(n1683));
AND2X1 mul_U9066(.A(dpath_mulcore_ary1_a1_s2[46]), .B(n8839), .Y(n15425));
INVX1 mul_U9067(.A(n15425), .Y(n1684));
AND2X1 mul_U9068(.A(dpath_mulcore_ary1_a1_s2[45]), .B(n8840), .Y(n15428));
INVX1 mul_U9069(.A(n15428), .Y(n1685));
AND2X1 mul_U9070(.A(dpath_mulcore_ary1_a1_s2[44]), .B(n8841), .Y(n15431));
INVX1 mul_U9071(.A(n15431), .Y(n1686));
AND2X1 mul_U9072(.A(dpath_mulcore_ary1_a1_s2[43]), .B(n8842), .Y(n15434));
INVX1 mul_U9073(.A(n15434), .Y(n1687));
AND2X1 mul_U9074(.A(dpath_mulcore_ary1_a1_s2[42]), .B(n8843), .Y(n15437));
INVX1 mul_U9075(.A(n15437), .Y(n1688));
AND2X1 mul_U9076(.A(dpath_mulcore_ary1_a1_s2[41]), .B(n8844), .Y(n15440));
INVX1 mul_U9077(.A(n15440), .Y(n1689));
AND2X1 mul_U9078(.A(dpath_mulcore_ary1_a1_s2[40]), .B(n8845), .Y(n15443));
INVX1 mul_U9079(.A(n15443), .Y(n1690));
AND2X1 mul_U9080(.A(dpath_mulcore_ary1_a1_s2[39]), .B(n8846), .Y(n15446));
INVX1 mul_U9081(.A(n15446), .Y(n1691));
AND2X1 mul_U9082(.A(dpath_mulcore_ary1_a1_s2[38]), .B(n8847), .Y(n15449));
INVX1 mul_U9083(.A(n15449), .Y(n1692));
AND2X1 mul_U9084(.A(dpath_mulcore_ary1_a1_s2[37]), .B(n8848), .Y(n15452));
INVX1 mul_U9085(.A(n15452), .Y(n1693));
AND2X1 mul_U9086(.A(dpath_mulcore_ary1_a1_s2[36]), .B(n8849), .Y(n15455));
INVX1 mul_U9087(.A(n15455), .Y(n1694));
AND2X1 mul_U9088(.A(dpath_mulcore_ary1_a1_s2[35]), .B(n8850), .Y(n15458));
INVX1 mul_U9089(.A(n15458), .Y(n1695));
AND2X1 mul_U9090(.A(dpath_mulcore_ary1_a1_s2[34]), .B(n8851), .Y(n15461));
INVX1 mul_U9091(.A(n15461), .Y(n1696));
AND2X1 mul_U9092(.A(dpath_mulcore_ary1_a1_s2[33]), .B(n8852), .Y(n15464));
INVX1 mul_U9093(.A(n15464), .Y(n1697));
AND2X1 mul_U9094(.A(dpath_mulcore_ary1_a1_s2[32]), .B(n8853), .Y(n15467));
INVX1 mul_U9095(.A(n15467), .Y(n1698));
AND2X1 mul_U9096(.A(dpath_mulcore_ary1_a1_s2[31]), .B(n8854), .Y(n15470));
INVX1 mul_U9097(.A(n15470), .Y(n1699));
AND2X1 mul_U9098(.A(dpath_mulcore_ary1_a1_s2[30]), .B(n8855), .Y(n15473));
INVX1 mul_U9099(.A(n15473), .Y(n1700));
AND2X1 mul_U9100(.A(dpath_mulcore_ary1_a1_s2[29]), .B(n8856), .Y(n15476));
INVX1 mul_U9101(.A(n15476), .Y(n1701));
AND2X1 mul_U9102(.A(dpath_mulcore_ary1_a1_s2[28]), .B(n8857), .Y(n15479));
INVX1 mul_U9103(.A(n15479), .Y(n1702));
AND2X1 mul_U9104(.A(dpath_mulcore_ary1_a1_s2[27]), .B(n8858), .Y(n15482));
INVX1 mul_U9105(.A(n15482), .Y(n1703));
AND2X1 mul_U9106(.A(dpath_mulcore_ary1_a1_s2[26]), .B(n8859), .Y(n15485));
INVX1 mul_U9107(.A(n15485), .Y(n1704));
AND2X1 mul_U9108(.A(dpath_mulcore_ary1_a1_s2[25]), .B(n8860), .Y(n15488));
INVX1 mul_U9109(.A(n15488), .Y(n1705));
AND2X1 mul_U9110(.A(dpath_mulcore_ary1_a1_s2[24]), .B(n8861), .Y(n15491));
INVX1 mul_U9111(.A(n15491), .Y(n1706));
AND2X1 mul_U9112(.A(dpath_mulcore_ary1_a1_s2[23]), .B(n8862), .Y(n15494));
INVX1 mul_U9113(.A(n15494), .Y(n1707));
AND2X1 mul_U9114(.A(dpath_mulcore_ary1_a1_s2[22]), .B(n8863), .Y(n15497));
INVX1 mul_U9115(.A(n15497), .Y(n1708));
AND2X1 mul_U9116(.A(dpath_mulcore_ary1_a1_s2[21]), .B(n8864), .Y(n15500));
INVX1 mul_U9117(.A(n15500), .Y(n1709));
AND2X1 mul_U9118(.A(dpath_mulcore_ary1_a1_s2[20]), .B(n8865), .Y(n15503));
INVX1 mul_U9119(.A(n15503), .Y(n1710));
AND2X1 mul_U9120(.A(dpath_mulcore_ary1_a1_s2[19]), .B(n8866), .Y(n15506));
INVX1 mul_U9121(.A(n15506), .Y(n1711));
AND2X1 mul_U9122(.A(dpath_mulcore_ary1_a1_s2[18]), .B(n8867), .Y(n15509));
INVX1 mul_U9123(.A(n15509), .Y(n1712));
AND2X1 mul_U9124(.A(dpath_mulcore_ary1_a1_s2[17]), .B(n8868), .Y(n15512));
INVX1 mul_U9125(.A(n15512), .Y(n1713));
AND2X1 mul_U9126(.A(dpath_mulcore_ary1_a1_s2[16]), .B(n8869), .Y(n15515));
INVX1 mul_U9127(.A(n15515), .Y(n1714));
AND2X1 mul_U9128(.A(dpath_mulcore_ary1_a1_s2[15]), .B(n8870), .Y(n15518));
INVX1 mul_U9129(.A(n15518), .Y(n1715));
AND2X1 mul_U9130(.A(dpath_mulcore_ary1_a1_s2[14]), .B(n8871), .Y(n15521));
INVX1 mul_U9131(.A(n15521), .Y(n1716));
AND2X1 mul_U9132(.A(dpath_mulcore_ary1_a1_s2[13]), .B(n8872), .Y(n15524));
INVX1 mul_U9133(.A(n15524), .Y(n1717));
AND2X1 mul_U9134(.A(dpath_mulcore_ary1_a1_s2[12]), .B(n8873), .Y(n15527));
INVX1 mul_U9135(.A(n15527), .Y(n1718));
AND2X1 mul_U9136(.A(dpath_mulcore_ary1_a1_s2[11]), .B(n8874), .Y(n15530));
INVX1 mul_U9137(.A(n15530), .Y(n1719));
AND2X1 mul_U9138(.A(dpath_mulcore_ary1_a1_s2[10]), .B(n8875), .Y(n15533));
INVX1 mul_U9139(.A(n15533), .Y(n1720));
AND2X1 mul_U9140(.A(dpath_mulcore_ary1_a1_s2[9]), .B(n8876), .Y(n15536));
INVX1 mul_U9141(.A(n15536), .Y(n1721));
AND2X1 mul_U9142(.A(dpath_mulcore_ary1_a1_s2[8]), .B(n8877), .Y(n15539));
INVX1 mul_U9143(.A(n15539), .Y(n1722));
AND2X1 mul_U9144(.A(dpath_mulcore_ary1_a1_s2[7]), .B(n8878), .Y(n15542));
INVX1 mul_U9145(.A(n15542), .Y(n1723));
AND2X1 mul_U9146(.A(dpath_mulcore_ary1_a1_s2[6]), .B(n8879), .Y(n15545));
INVX1 mul_U9147(.A(n15545), .Y(n1724));
AND2X1 mul_U9148(.A(dpath_mulcore_ary1_a1_s2[5]), .B(n8880), .Y(n15548));
INVX1 mul_U9149(.A(n15548), .Y(n1725));
AND2X1 mul_U9150(.A(dpath_mulcore_ary1_a1_s2[4]), .B(n8761), .Y(n15551));
INVX1 mul_U9151(.A(n15551), .Y(n1726));
AND2X1 mul_U9152(.A(dpath_mulcore_ary1_a1_s2[3]), .B(n8762), .Y(n15554));
INVX1 mul_U9153(.A(n15554), .Y(n1727));
AND2X1 mul_U9154(.A(dpath_mulcore_ary1_a1_s2[2]), .B(dpath_mulcore_ary1_a1_c2[1]), .Y(n15557));
INVX1 mul_U9155(.A(n15557), .Y(n1728));
AND2X1 mul_U9156(.A(dpath_mulcore_ary1_a1_s2[1]), .B(dpath_mulcore_ary1_a1_s1[7]), .Y(n15560));
INVX1 mul_U9157(.A(n15560), .Y(n1729));
AND2X1 mul_U9158(.A(dpath_mulcore_ary1_a1_s2[0]), .B(dpath_mulcore_ary1_a1_s1[6]), .Y(n15563));
INVX1 mul_U9159(.A(n15563), .Y(n1730));
AND2X1 mul_U9160(.A(n8379), .B(dpath_mulcore_ary1_a1_s1[5]), .Y(n15566));
INVX1 mul_U9161(.A(n15566), .Y(n1731));
AND2X1 mul_U9162(.A(n8380), .B(dpath_mulcore_ary1_a1_s1[4]), .Y(n15569));
INVX1 mul_U9163(.A(n15569), .Y(n1732));
AND2X1 mul_U9164(.A(dpath_mulcore_ary1_a1_s2[64]), .B(n8821), .Y(n15571));
INVX1 mul_U9165(.A(n15571), .Y(n1733));
AND2X1 mul_U9166(.A(n5213), .B(n4691), .Y(dpath_mulcore_a1cout[77]));
INVX1 mul_U9167(.A(dpath_mulcore_a1cout[77]), .Y(n1734));
AND2X1 mul_U9168(.A(dpath_mulcore_ary1_a1_s0[9]), .B(n8932), .Y(n15576));
INVX1 mul_U9169(.A(n15576), .Y(n1735));
AND2X1 mul_U9170(.A(dpath_mulcore_ary1_a1_s0[8]), .B(n8933), .Y(n15579));
INVX1 mul_U9171(.A(n15579), .Y(n1736));
AND2X1 mul_U9172(.A(dpath_mulcore_ary1_a1_s0[3]), .B(n8764), .Y(n15582));
INVX1 mul_U9173(.A(n15582), .Y(n1737));
AND2X1 mul_U9174(.A(n5214), .B(n4692), .Y(dpath_mulcore_a1cout[10]));
INVX1 mul_U9175(.A(dpath_mulcore_a1cout[10]), .Y(n1738));
AND2X1 mul_U9176(.A(n5215), .B(n4693), .Y(dpath_mulcore_a1cout[9]));
INVX1 mul_U9177(.A(dpath_mulcore_a1cout[9]), .Y(n1739));
AND2X1 mul_U9178(.A(n5216), .B(n4694), .Y(dpath_mulcore_a1cout[8]));
INVX1 mul_U9179(.A(dpath_mulcore_a1cout[8]), .Y(n1740));
AND2X1 mul_U9180(.A(dpath_mulcore_ary1_a1_s2[59]), .B(n8826), .Y(n15594));
INVX1 mul_U9181(.A(n15594), .Y(n1741));
AND2X1 mul_U9182(.A(dpath_mulcore_ary1_a1_s2[63]), .B(n8822), .Y(n15597));
INVX1 mul_U9183(.A(n15597), .Y(n1742));
AND2X1 mul_U9184(.A(dpath_mulcore_ary1_a1_s2[62]), .B(n8823), .Y(n15600));
INVX1 mul_U9185(.A(n15600), .Y(n1743));
AND2X1 mul_U9186(.A(dpath_mulcore_ary1_a1_s2[61]), .B(n8824), .Y(n15603));
INVX1 mul_U9187(.A(n15603), .Y(n1744));
AND2X1 mul_U9188(.A(dpath_mulcore_ary1_a1_s2[60]), .B(n8825), .Y(n15606));
INVX1 mul_U9189(.A(n15606), .Y(n1745));
AND2X1 mul_U9190(.A(n9427), .B(n9489), .Y(n15609));
INVX1 mul_U9191(.A(n15609), .Y(n1746));
AND2X1 mul_U9192(.A(dpath_mulcore_ary1_a1_I0_I2_net073), .B(n14798), .Y(n15612));
INVX1 mul_U9193(.A(n15612), .Y(n1747));
AND2X1 mul_U9194(.A(dpath_mulcore_ary1_a1_s0[67]), .B(n8944), .Y(n15615));
INVX1 mul_U9195(.A(n15615), .Y(n1748));
AND2X1 mul_U9196(.A(dpath_mulcore_ary1_a1_s0[66]), .B(n8943), .Y(n15618));
INVX1 mul_U9197(.A(n15618), .Y(n1749));
AND2X1 mul_U9198(.A(dpath_mulcore_ary1_a1_s0[65]), .B(n8942), .Y(n15621));
INVX1 mul_U9199(.A(n15621), .Y(n1750));
AND2X1 mul_U9200(.A(dpath_mulcore_ary1_a1_s0[64]), .B(n8881), .Y(n15624));
INVX1 mul_U9201(.A(n15624), .Y(n1751));
AND2X1 mul_U9202(.A(dpath_mulcore_ary1_a1_s0[63]), .B(n8882), .Y(n15627));
INVX1 mul_U9203(.A(n15627), .Y(n1752));
AND2X1 mul_U9204(.A(dpath_mulcore_ary1_a1_s0[62]), .B(n8883), .Y(n15630));
INVX1 mul_U9205(.A(n15630), .Y(n1753));
AND2X1 mul_U9206(.A(dpath_mulcore_ary1_a1_s0[61]), .B(n8884), .Y(n15633));
INVX1 mul_U9207(.A(n15633), .Y(n1754));
AND2X1 mul_U9208(.A(dpath_mulcore_ary1_a1_s0[60]), .B(n8885), .Y(n15636));
INVX1 mul_U9209(.A(n15636), .Y(n1755));
AND2X1 mul_U9210(.A(dpath_mulcore_ary1_a1_s0[59]), .B(n8886), .Y(n15639));
INVX1 mul_U9211(.A(n15639), .Y(n1756));
AND2X1 mul_U9212(.A(dpath_mulcore_ary1_a1_s0[58]), .B(n8887), .Y(n15642));
INVX1 mul_U9213(.A(n15642), .Y(n1757));
AND2X1 mul_U9214(.A(dpath_mulcore_ary1_a1_s0[57]), .B(n8888), .Y(n15645));
INVX1 mul_U9215(.A(n15645), .Y(n1758));
AND2X1 mul_U9216(.A(dpath_mulcore_ary1_a1_s0[56]), .B(n8889), .Y(n15648));
INVX1 mul_U9217(.A(n15648), .Y(n1759));
AND2X1 mul_U9218(.A(dpath_mulcore_ary1_a1_s0[55]), .B(n8890), .Y(n15651));
INVX1 mul_U9219(.A(n15651), .Y(n1760));
AND2X1 mul_U9220(.A(dpath_mulcore_ary1_a1_s0[54]), .B(n8891), .Y(n15654));
INVX1 mul_U9221(.A(n15654), .Y(n1761));
AND2X1 mul_U9222(.A(dpath_mulcore_ary1_a1_s0[53]), .B(n8892), .Y(n15657));
INVX1 mul_U9223(.A(n15657), .Y(n1762));
AND2X1 mul_U9224(.A(dpath_mulcore_ary1_a1_s0[52]), .B(n8893), .Y(n15660));
INVX1 mul_U9225(.A(n15660), .Y(n1763));
AND2X1 mul_U9226(.A(dpath_mulcore_ary1_a1_s0[51]), .B(n8894), .Y(n15663));
INVX1 mul_U9227(.A(n15663), .Y(n1764));
AND2X1 mul_U9228(.A(dpath_mulcore_ary1_a1_s0[50]), .B(n8895), .Y(n15666));
INVX1 mul_U9229(.A(n15666), .Y(n1765));
AND2X1 mul_U9230(.A(dpath_mulcore_ary1_a1_s0[49]), .B(n8896), .Y(n15669));
INVX1 mul_U9231(.A(n15669), .Y(n1766));
AND2X1 mul_U9232(.A(dpath_mulcore_ary1_a1_s0[48]), .B(n8897), .Y(n15672));
INVX1 mul_U9233(.A(n15672), .Y(n1767));
AND2X1 mul_U9234(.A(dpath_mulcore_ary1_a1_s0[47]), .B(n8898), .Y(n15675));
INVX1 mul_U9235(.A(n15675), .Y(n1768));
AND2X1 mul_U9236(.A(dpath_mulcore_ary1_a1_s0[46]), .B(n8899), .Y(n15678));
INVX1 mul_U9237(.A(n15678), .Y(n1769));
AND2X1 mul_U9238(.A(dpath_mulcore_ary1_a1_s0[45]), .B(n8900), .Y(n15681));
INVX1 mul_U9239(.A(n15681), .Y(n1770));
AND2X1 mul_U9240(.A(dpath_mulcore_ary1_a1_s0[44]), .B(n8901), .Y(n15684));
INVX1 mul_U9241(.A(n15684), .Y(n1771));
AND2X1 mul_U9242(.A(dpath_mulcore_ary1_a1_s0[43]), .B(n8902), .Y(n15687));
INVX1 mul_U9243(.A(n15687), .Y(n1772));
AND2X1 mul_U9244(.A(dpath_mulcore_ary1_a1_s0[42]), .B(n8903), .Y(n15690));
INVX1 mul_U9245(.A(n15690), .Y(n1773));
AND2X1 mul_U9246(.A(dpath_mulcore_ary1_a1_s0[41]), .B(n8904), .Y(n15693));
INVX1 mul_U9247(.A(n15693), .Y(n1774));
AND2X1 mul_U9248(.A(dpath_mulcore_ary1_a1_s0[40]), .B(n8905), .Y(n15696));
INVX1 mul_U9249(.A(n15696), .Y(n1775));
AND2X1 mul_U9250(.A(dpath_mulcore_ary1_a1_s0[39]), .B(n8906), .Y(n15699));
INVX1 mul_U9251(.A(n15699), .Y(n1776));
AND2X1 mul_U9252(.A(dpath_mulcore_ary1_a1_s0[38]), .B(n8907), .Y(n15702));
INVX1 mul_U9253(.A(n15702), .Y(n1777));
AND2X1 mul_U9254(.A(dpath_mulcore_ary1_a1_s0[37]), .B(n8908), .Y(n15705));
INVX1 mul_U9255(.A(n15705), .Y(n1778));
AND2X1 mul_U9256(.A(dpath_mulcore_ary1_a1_s0[36]), .B(n8909), .Y(n15708));
INVX1 mul_U9257(.A(n15708), .Y(n1779));
AND2X1 mul_U9258(.A(dpath_mulcore_ary1_a1_s0[35]), .B(n8910), .Y(n15711));
INVX1 mul_U9259(.A(n15711), .Y(n1780));
AND2X1 mul_U9260(.A(dpath_mulcore_ary1_a1_s0[34]), .B(n8911), .Y(n15714));
INVX1 mul_U9261(.A(n15714), .Y(n1781));
AND2X1 mul_U9262(.A(dpath_mulcore_ary1_a1_s0[33]), .B(n8912), .Y(n15717));
INVX1 mul_U9263(.A(n15717), .Y(n1782));
AND2X1 mul_U9264(.A(dpath_mulcore_ary1_a1_s0[32]), .B(n8913), .Y(n15720));
INVX1 mul_U9265(.A(n15720), .Y(n1783));
AND2X1 mul_U9266(.A(dpath_mulcore_ary1_a1_s0[31]), .B(n8914), .Y(n15723));
INVX1 mul_U9267(.A(n15723), .Y(n1784));
AND2X1 mul_U9268(.A(dpath_mulcore_ary1_a1_s0[30]), .B(n8915), .Y(n15726));
INVX1 mul_U9269(.A(n15726), .Y(n1785));
AND2X1 mul_U9270(.A(dpath_mulcore_ary1_a1_s0[29]), .B(n8916), .Y(n15729));
INVX1 mul_U9271(.A(n15729), .Y(n1786));
AND2X1 mul_U9272(.A(dpath_mulcore_ary1_a1_s0[28]), .B(n8917), .Y(n15732));
INVX1 mul_U9273(.A(n15732), .Y(n1787));
AND2X1 mul_U9274(.A(dpath_mulcore_ary1_a1_s0[27]), .B(n8918), .Y(n15735));
INVX1 mul_U9275(.A(n15735), .Y(n1788));
AND2X1 mul_U9276(.A(dpath_mulcore_ary1_a1_s0[26]), .B(n8919), .Y(n15738));
INVX1 mul_U9277(.A(n15738), .Y(n1789));
AND2X1 mul_U9278(.A(dpath_mulcore_ary1_a1_s0[25]), .B(n8920), .Y(n15741));
INVX1 mul_U9279(.A(n15741), .Y(n1790));
AND2X1 mul_U9280(.A(dpath_mulcore_ary1_a1_s0[24]), .B(n8921), .Y(n15744));
INVX1 mul_U9281(.A(n15744), .Y(n1791));
AND2X1 mul_U9282(.A(dpath_mulcore_ary1_a1_s0[23]), .B(n8922), .Y(n15747));
INVX1 mul_U9283(.A(n15747), .Y(n1792));
AND2X1 mul_U9284(.A(dpath_mulcore_ary1_a1_s0[22]), .B(n8923), .Y(n15750));
INVX1 mul_U9285(.A(n15750), .Y(n1793));
AND2X1 mul_U9286(.A(dpath_mulcore_ary1_a1_s0[21]), .B(n8924), .Y(n15753));
INVX1 mul_U9287(.A(n15753), .Y(n1794));
AND2X1 mul_U9288(.A(dpath_mulcore_ary1_a1_s0[20]), .B(n8925), .Y(n15756));
INVX1 mul_U9289(.A(n15756), .Y(n1795));
AND2X1 mul_U9290(.A(dpath_mulcore_ary1_a1_s0[19]), .B(n8926), .Y(n15759));
INVX1 mul_U9291(.A(n15759), .Y(n1796));
AND2X1 mul_U9292(.A(dpath_mulcore_ary1_a1_s0[18]), .B(n8927), .Y(n15762));
INVX1 mul_U9293(.A(n15762), .Y(n1797));
AND2X1 mul_U9294(.A(dpath_mulcore_ary1_a1_s0[17]), .B(n8928), .Y(n15765));
INVX1 mul_U9295(.A(n15765), .Y(n1798));
AND2X1 mul_U9296(.A(dpath_mulcore_ary1_a1_s0[16]), .B(n8929), .Y(n15768));
INVX1 mul_U9297(.A(n15768), .Y(n1799));
AND2X1 mul_U9298(.A(dpath_mulcore_ary1_a1_s0[15]), .B(n8930), .Y(n15771));
INVX1 mul_U9299(.A(n15771), .Y(n1800));
AND2X1 mul_U9300(.A(dpath_mulcore_ary1_a1_s0[14]), .B(n8931), .Y(n15774));
INVX1 mul_U9301(.A(n15774), .Y(n1801));
AND2X1 mul_U9302(.A(dpath_mulcore_ary1_a1_s0[7]), .B(n8934), .Y(n15777));
INVX1 mul_U9303(.A(n15777), .Y(n1802));
AND2X1 mul_U9304(.A(dpath_mulcore_ary1_a1_s0[6]), .B(n8935), .Y(n15780));
INVX1 mul_U9305(.A(n15780), .Y(n1803));
AND2X1 mul_U9306(.A(dpath_mulcore_ary1_a1_s0[5]), .B(n8936), .Y(n15783));
INVX1 mul_U9307(.A(n15783), .Y(n1804));
AND2X1 mul_U9308(.A(dpath_mulcore_ary1_a1_s0[4]), .B(n8763), .Y(n15786));
INVX1 mul_U9309(.A(n15786), .Y(n1805));
AND2X1 mul_U9310(.A(n8385), .B(dpath_mulcore_array2_s2[82]), .Y(n15789));
INVX1 mul_U9311(.A(n15789), .Y(n1806));
AND2X1 mul_U9312(.A(n8191), .B(dpath_mulcore_array2_s3[68]), .Y(n15792));
INVX1 mul_U9313(.A(n15792), .Y(n1807));
AND2X1 mul_U9314(.A(n8192), .B(dpath_mulcore_array2_s3[67]), .Y(n15795));
INVX1 mul_U9315(.A(n15795), .Y(n1808));
AND2X1 mul_U9316(.A(n8193), .B(dpath_mulcore_array2_s3[66]), .Y(n15798));
INVX1 mul_U9317(.A(n15798), .Y(n1809));
AND2X1 mul_U9318(.A(n8194), .B(dpath_mulcore_array2_s3[65]), .Y(n15801));
INVX1 mul_U9319(.A(n15801), .Y(n1810));
AND2X1 mul_U9320(.A(n8195), .B(dpath_mulcore_array2_s3[64]), .Y(n15804));
INVX1 mul_U9321(.A(n15804), .Y(n1811));
AND2X1 mul_U9322(.A(n8196), .B(dpath_mulcore_array2_s3[63]), .Y(n15807));
INVX1 mul_U9323(.A(n15807), .Y(n1812));
AND2X1 mul_U9324(.A(n8197), .B(dpath_mulcore_array2_s3[62]), .Y(n15810));
INVX1 mul_U9325(.A(n15810), .Y(n1813));
AND2X1 mul_U9326(.A(n8198), .B(dpath_mulcore_array2_s3[61]), .Y(n15813));
INVX1 mul_U9327(.A(n15813), .Y(n1814));
AND2X1 mul_U9328(.A(n8199), .B(dpath_mulcore_array2_s3[60]), .Y(n15816));
INVX1 mul_U9329(.A(n15816), .Y(n1815));
AND2X1 mul_U9330(.A(n8200), .B(dpath_mulcore_array2_s3[59]), .Y(n15819));
INVX1 mul_U9331(.A(n15819), .Y(n1816));
AND2X1 mul_U9332(.A(n8201), .B(dpath_mulcore_array2_s3[58]), .Y(n15822));
INVX1 mul_U9333(.A(n15822), .Y(n1817));
AND2X1 mul_U9334(.A(n8202), .B(dpath_mulcore_array2_s3[57]), .Y(n15825));
INVX1 mul_U9335(.A(n15825), .Y(n1818));
AND2X1 mul_U9336(.A(n8203), .B(dpath_mulcore_array2_s3[56]), .Y(n15828));
INVX1 mul_U9337(.A(n15828), .Y(n1819));
AND2X1 mul_U9338(.A(n8204), .B(dpath_mulcore_array2_s3[55]), .Y(n15831));
INVX1 mul_U9339(.A(n15831), .Y(n1820));
AND2X1 mul_U9340(.A(n8205), .B(dpath_mulcore_array2_s3[54]), .Y(n15834));
INVX1 mul_U9341(.A(n15834), .Y(n1821));
AND2X1 mul_U9342(.A(n8206), .B(dpath_mulcore_array2_s3[53]), .Y(n15837));
INVX1 mul_U9343(.A(n15837), .Y(n1822));
AND2X1 mul_U9344(.A(n8207), .B(dpath_mulcore_array2_s3[52]), .Y(n15840));
INVX1 mul_U9345(.A(n15840), .Y(n1823));
AND2X1 mul_U9346(.A(n8208), .B(dpath_mulcore_array2_s3[51]), .Y(n15843));
INVX1 mul_U9347(.A(n15843), .Y(n1824));
AND2X1 mul_U9348(.A(n8209), .B(dpath_mulcore_array2_s3[50]), .Y(n15846));
INVX1 mul_U9349(.A(n15846), .Y(n1825));
AND2X1 mul_U9350(.A(n8210), .B(dpath_mulcore_array2_s3[49]), .Y(n15849));
INVX1 mul_U9351(.A(n15849), .Y(n1826));
AND2X1 mul_U9352(.A(n8211), .B(dpath_mulcore_array2_s3[48]), .Y(n15852));
INVX1 mul_U9353(.A(n15852), .Y(n1827));
AND2X1 mul_U9354(.A(n8212), .B(dpath_mulcore_array2_s3[47]), .Y(n15855));
INVX1 mul_U9355(.A(n15855), .Y(n1828));
AND2X1 mul_U9356(.A(n8213), .B(dpath_mulcore_array2_s3[46]), .Y(n15858));
INVX1 mul_U9357(.A(n15858), .Y(n1829));
AND2X1 mul_U9358(.A(n8214), .B(dpath_mulcore_array2_s3[45]), .Y(n15861));
INVX1 mul_U9359(.A(n15861), .Y(n1830));
AND2X1 mul_U9360(.A(n8215), .B(dpath_mulcore_array2_s3[44]), .Y(n15864));
INVX1 mul_U9361(.A(n15864), .Y(n1831));
AND2X1 mul_U9362(.A(n8216), .B(dpath_mulcore_array2_s3[43]), .Y(n15867));
INVX1 mul_U9363(.A(n15867), .Y(n1832));
AND2X1 mul_U9364(.A(n8217), .B(dpath_mulcore_array2_s3[42]), .Y(n15870));
INVX1 mul_U9365(.A(n15870), .Y(n1833));
AND2X1 mul_U9366(.A(n8218), .B(dpath_mulcore_array2_s3[41]), .Y(n15873));
INVX1 mul_U9367(.A(n15873), .Y(n1834));
AND2X1 mul_U9368(.A(n8219), .B(dpath_mulcore_array2_s3[40]), .Y(n15876));
INVX1 mul_U9369(.A(n15876), .Y(n1835));
AND2X1 mul_U9370(.A(n8220), .B(dpath_mulcore_array2_s3[39]), .Y(n15879));
INVX1 mul_U9371(.A(n15879), .Y(n1836));
AND2X1 mul_U9372(.A(n8221), .B(dpath_mulcore_array2_s3[38]), .Y(n15882));
INVX1 mul_U9373(.A(n15882), .Y(n1837));
AND2X1 mul_U9374(.A(n8222), .B(dpath_mulcore_array2_s3[37]), .Y(n15885));
INVX1 mul_U9375(.A(n15885), .Y(n1838));
AND2X1 mul_U9376(.A(n8223), .B(dpath_mulcore_array2_s3[36]), .Y(n15888));
INVX1 mul_U9377(.A(n15888), .Y(n1839));
AND2X1 mul_U9378(.A(n8224), .B(dpath_mulcore_array2_s3[35]), .Y(n15891));
INVX1 mul_U9379(.A(n15891), .Y(n1840));
AND2X1 mul_U9380(.A(n8225), .B(dpath_mulcore_array2_s3[34]), .Y(n15894));
INVX1 mul_U9381(.A(n15894), .Y(n1841));
AND2X1 mul_U9382(.A(n8226), .B(dpath_mulcore_array2_s3[33]), .Y(n15897));
INVX1 mul_U9383(.A(n15897), .Y(n1842));
AND2X1 mul_U9384(.A(n8227), .B(dpath_mulcore_array2_s3[32]), .Y(n15900));
INVX1 mul_U9385(.A(n15900), .Y(n1843));
AND2X1 mul_U9386(.A(n8228), .B(dpath_mulcore_array2_s3[31]), .Y(n15903));
INVX1 mul_U9387(.A(n15903), .Y(n1844));
AND2X1 mul_U9388(.A(n8229), .B(dpath_mulcore_array2_s3[30]), .Y(n15906));
INVX1 mul_U9389(.A(n15906), .Y(n1845));
AND2X1 mul_U9390(.A(n8230), .B(dpath_mulcore_array2_s3[29]), .Y(n15909));
INVX1 mul_U9391(.A(n15909), .Y(n1846));
AND2X1 mul_U9392(.A(n8231), .B(dpath_mulcore_array2_s3[28]), .Y(n15912));
INVX1 mul_U9393(.A(n15912), .Y(n1847));
AND2X1 mul_U9394(.A(n8232), .B(dpath_mulcore_array2_s3[27]), .Y(n15915));
INVX1 mul_U9395(.A(n15915), .Y(n1848));
AND2X1 mul_U9396(.A(n8233), .B(dpath_mulcore_array2_s3[26]), .Y(n15918));
INVX1 mul_U9397(.A(n15918), .Y(n1849));
AND2X1 mul_U9398(.A(n8234), .B(dpath_mulcore_array2_s3[25]), .Y(n15921));
INVX1 mul_U9399(.A(n15921), .Y(n1850));
AND2X1 mul_U9400(.A(n8235), .B(dpath_mulcore_array2_s3[24]), .Y(n15924));
INVX1 mul_U9401(.A(n15924), .Y(n1851));
AND2X1 mul_U9402(.A(n8236), .B(dpath_mulcore_array2_s3[23]), .Y(n15927));
INVX1 mul_U9403(.A(n15927), .Y(n1852));
AND2X1 mul_U9404(.A(n8237), .B(dpath_mulcore_array2_s3[22]), .Y(n15930));
INVX1 mul_U9405(.A(n15930), .Y(n1853));
AND2X1 mul_U9406(.A(n8238), .B(dpath_mulcore_array2_s3[21]), .Y(n15933));
INVX1 mul_U9407(.A(n15933), .Y(n1854));
AND2X1 mul_U9408(.A(n8239), .B(dpath_mulcore_array2_sc3_20__z), .Y(n15936));
INVX1 mul_U9409(.A(n15936), .Y(n1855));
AND2X1 mul_U9410(.A(n14897), .B(dpath_mulcore_array2_s2[96]), .Y(n15939));
INVX1 mul_U9411(.A(n15939), .Y(n1856));
AND2X1 mul_U9412(.A(n8240), .B(dpath_mulcore_array2_s2[95]), .Y(n15942));
INVX1 mul_U9413(.A(n15942), .Y(n1857));
AND2X1 mul_U9414(.A(n8241), .B(dpath_mulcore_array2_s2[94]), .Y(n15945));
INVX1 mul_U9415(.A(n15945), .Y(n1858));
AND2X1 mul_U9416(.A(n8242), .B(dpath_mulcore_array2_s2[93]), .Y(n15948));
INVX1 mul_U9417(.A(n15948), .Y(n1859));
AND2X1 mul_U9418(.A(n8243), .B(dpath_mulcore_array2_s2[92]), .Y(n15951));
INVX1 mul_U9419(.A(n15951), .Y(n1860));
AND2X1 mul_U9420(.A(n8244), .B(dpath_mulcore_array2_s2[91]), .Y(n15954));
INVX1 mul_U9421(.A(n15954), .Y(n1861));
AND2X1 mul_U9422(.A(n8245), .B(dpath_mulcore_array2_s2[90]), .Y(n15957));
INVX1 mul_U9423(.A(n15957), .Y(n1862));
AND2X1 mul_U9424(.A(n8246), .B(dpath_mulcore_array2_s2[89]), .Y(n15960));
INVX1 mul_U9425(.A(n15960), .Y(n1863));
AND2X1 mul_U9426(.A(n8247), .B(dpath_mulcore_array2_s2[88]), .Y(n15963));
INVX1 mul_U9427(.A(n15963), .Y(n1864));
AND2X1 mul_U9428(.A(n8248), .B(dpath_mulcore_array2_s2[87]), .Y(n15966));
INVX1 mul_U9429(.A(n15966), .Y(n1865));
AND2X1 mul_U9430(.A(n8249), .B(dpath_mulcore_array2_s2[86]), .Y(n15969));
INVX1 mul_U9431(.A(n15969), .Y(n1866));
AND2X1 mul_U9432(.A(n8250), .B(dpath_mulcore_array2_s2[85]), .Y(n15972));
INVX1 mul_U9433(.A(n15972), .Y(n1867));
AND2X1 mul_U9434(.A(n8251), .B(dpath_mulcore_array2_s2[84]), .Y(n15975));
INVX1 mul_U9435(.A(n15975), .Y(n1868));
AND2X1 mul_U9436(.A(n8252), .B(dpath_mulcore_array2_s3[81]), .Y(n15978));
INVX1 mul_U9437(.A(n15978), .Y(n1869));
AND2X1 mul_U9438(.A(n8253), .B(dpath_mulcore_array2_s3[80]), .Y(n15981));
INVX1 mul_U9439(.A(n15981), .Y(n1870));
AND2X1 mul_U9440(.A(n8254), .B(dpath_mulcore_array2_s3[79]), .Y(n15984));
INVX1 mul_U9441(.A(n15984), .Y(n1871));
AND2X1 mul_U9442(.A(n8255), .B(dpath_mulcore_array2_s3[78]), .Y(n15987));
INVX1 mul_U9443(.A(n15987), .Y(n1872));
AND2X1 mul_U9444(.A(n8256), .B(dpath_mulcore_array2_s3[77]), .Y(n15990));
INVX1 mul_U9445(.A(n15990), .Y(n1873));
AND2X1 mul_U9446(.A(n8257), .B(dpath_mulcore_array2_s3[76]), .Y(n15993));
INVX1 mul_U9447(.A(n15993), .Y(n1874));
AND2X1 mul_U9448(.A(n8258), .B(dpath_mulcore_array2_s3[75]), .Y(n15996));
INVX1 mul_U9449(.A(n15996), .Y(n1875));
AND2X1 mul_U9450(.A(n8259), .B(dpath_mulcore_array2_s3[74]), .Y(n15999));
INVX1 mul_U9451(.A(n15999), .Y(n1876));
AND2X1 mul_U9452(.A(n8260), .B(dpath_mulcore_array2_s3[73]), .Y(n16002));
INVX1 mul_U9453(.A(n16002), .Y(n1877));
AND2X1 mul_U9454(.A(n8261), .B(dpath_mulcore_array2_s3[72]), .Y(n16005));
INVX1 mul_U9455(.A(n16005), .Y(n1878));
AND2X1 mul_U9456(.A(n8262), .B(dpath_mulcore_array2_s3[71]), .Y(n16008));
INVX1 mul_U9457(.A(n16008), .Y(n1879));
AND2X1 mul_U9458(.A(n8263), .B(dpath_mulcore_array2_s3[70]), .Y(n16011));
INVX1 mul_U9459(.A(n16011), .Y(n1880));
AND2X1 mul_U9460(.A(n8264), .B(dpath_mulcore_array2_s3[69]), .Y(n16014));
INVX1 mul_U9461(.A(n16014), .Y(n1881));
AND2X1 mul_U9462(.A(n8270), .B(dpath_mulcore_array2_s2[4]), .Y(n16017));
INVX1 mul_U9463(.A(n16017), .Y(n1882));
AND2X1 mul_U9464(.A(n8271), .B(dpath_mulcore_array2_s2[3]), .Y(n16020));
INVX1 mul_U9465(.A(n16020), .Y(n1883));
AND2X1 mul_U9466(.A(n8272), .B(dpath_mulcore_array2_s2[2]), .Y(n16023));
INVX1 mul_U9467(.A(n16023), .Y(n1884));
AND2X1 mul_U9468(.A(n8273), .B(dpath_mulcore_array2_s2[1]), .Y(n16026));
INVX1 mul_U9469(.A(n16026), .Y(n1885));
AND2X1 mul_U9470(.A(n5217), .B(n4695), .Y(dpath_mulcore_pcout[97]));
INVX1 mul_U9471(.A(dpath_mulcore_pcout[97]), .Y(n1886));
AND2X1 mul_U9472(.A(dpath_mulcore_ps[51]), .B(dpath_mulcore_pc[50]), .Y(n16032));
INVX1 mul_U9473(.A(n16032), .Y(n1887));
AND2X1 mul_U9474(.A(dpath_mulcore_ps[50]), .B(dpath_mulcore_pc[49]), .Y(n16035));
INVX1 mul_U9475(.A(n16035), .Y(n1888));
AND2X1 mul_U9476(.A(dpath_mulcore_ps[49]), .B(dpath_mulcore_pc[48]), .Y(n16038));
INVX1 mul_U9477(.A(n16038), .Y(n1889));
AND2X1 mul_U9478(.A(dpath_mulcore_ps[48]), .B(dpath_mulcore_pc[47]), .Y(n16041));
INVX1 mul_U9479(.A(n16041), .Y(n1890));
AND2X1 mul_U9480(.A(n8274), .B(dpath_mulcore_array2_s2[83]), .Y(n16046));
INVX1 mul_U9481(.A(n16046), .Y(n1891));
AND2X1 mul_U9482(.A(dpath_mulcore_a1s[67]), .B(dpath_mulcore_a1c[66]), .Y(n16049));
INVX1 mul_U9483(.A(n16049), .Y(n1892));
AND2X1 mul_U9484(.A(dpath_mulcore_array2_s1[19]), .B(dpath_mulcore_a0s[19]), .Y(n16052));
INVX1 mul_U9485(.A(n16052), .Y(n1893));
AND2X1 mul_U9486(.A(dpath_mulcore_array2_s1[18]), .B(dpath_mulcore_a0s[18]), .Y(n16055));
INVX1 mul_U9487(.A(n16055), .Y(n1894));
AND2X1 mul_U9488(.A(dpath_mulcore_array2_s1[17]), .B(dpath_mulcore_a0s[17]), .Y(n16058));
INVX1 mul_U9489(.A(n16058), .Y(n1895));
AND2X1 mul_U9490(.A(dpath_mulcore_array2_s1[16]), .B(dpath_mulcore_a0s[16]), .Y(n16061));
INVX1 mul_U9491(.A(n16061), .Y(n1896));
AND2X1 mul_U9492(.A(n16043), .B(dpath_mulcore_a0s[15]), .Y(n16064));
INVX1 mul_U9493(.A(n16064), .Y(n1897));
AND2X1 mul_U9494(.A(dpath_mulcore_a1s[65]), .B(dpath_mulcore_a1c[64]), .Y(n16066));
INVX1 mul_U9495(.A(n16066), .Y(dpath_mulcore_array2_c1[81]));
AND2X1 mul_U9496(.A(dpath_mulcore_a1s[64]), .B(dpath_mulcore_a1c[63]), .Y(n16068));
INVX1 mul_U9497(.A(n16068), .Y(n1898));
AND2X1 mul_U9498(.A(dpath_mulcore_a1s[63]), .B(dpath_mulcore_a1c[62]), .Y(n16071));
INVX1 mul_U9499(.A(n16071), .Y(n1899));
AND2X1 mul_U9500(.A(dpath_mulcore_a1s[62]), .B(dpath_mulcore_a1c[61]), .Y(n16074));
INVX1 mul_U9501(.A(n16074), .Y(n1900));
AND2X1 mul_U9502(.A(dpath_mulcore_a1s[61]), .B(dpath_mulcore_a1c[60]), .Y(n16077));
INVX1 mul_U9503(.A(n16077), .Y(n1901));
AND2X1 mul_U9504(.A(dpath_mulcore_a1s[60]), .B(dpath_mulcore_a1c[59]), .Y(n16080));
INVX1 mul_U9505(.A(n16080), .Y(n1902));
AND2X1 mul_U9506(.A(dpath_mulcore_a1s[59]), .B(dpath_mulcore_a1c[58]), .Y(n16083));
INVX1 mul_U9507(.A(n16083), .Y(n1903));
AND2X1 mul_U9508(.A(dpath_mulcore_a1s[58]), .B(dpath_mulcore_a1c[57]), .Y(n16086));
INVX1 mul_U9509(.A(n16086), .Y(n1904));
AND2X1 mul_U9510(.A(dpath_mulcore_a1s[57]), .B(dpath_mulcore_a1c[56]), .Y(n16089));
INVX1 mul_U9511(.A(n16089), .Y(n1905));
AND2X1 mul_U9512(.A(dpath_mulcore_a1s[56]), .B(dpath_mulcore_a1c[55]), .Y(n16092));
INVX1 mul_U9513(.A(n16092), .Y(n1906));
AND2X1 mul_U9514(.A(dpath_mulcore_a1s[55]), .B(dpath_mulcore_a1c[54]), .Y(n16095));
INVX1 mul_U9515(.A(n16095), .Y(n1907));
AND2X1 mul_U9516(.A(dpath_mulcore_a1s[54]), .B(dpath_mulcore_a1c[53]), .Y(n16098));
INVX1 mul_U9517(.A(n16098), .Y(n1908));
AND2X1 mul_U9518(.A(dpath_mulcore_a1s[53]), .B(dpath_mulcore_a1c[52]), .Y(n16101));
INVX1 mul_U9519(.A(n16101), .Y(n1909));
AND2X1 mul_U9520(.A(dpath_mulcore_a1s[52]), .B(dpath_mulcore_a1c[51]), .Y(n16104));
INVX1 mul_U9521(.A(n16104), .Y(n1910));
AND2X1 mul_U9522(.A(dpath_mulcore_array2_s2[19]), .B(n8945), .Y(n16107));
INVX1 mul_U9523(.A(n16107), .Y(n1911));
AND2X1 mul_U9524(.A(dpath_mulcore_array2_s2[18]), .B(n8946), .Y(n16110));
INVX1 mul_U9525(.A(n16110), .Y(n1912));
AND2X1 mul_U9526(.A(dpath_mulcore_array2_s2[17]), .B(n8947), .Y(n16113));
INVX1 mul_U9527(.A(n16113), .Y(n1913));
AND2X1 mul_U9528(.A(dpath_mulcore_array2_s2[16]), .B(n16044), .Y(n16116));
INVX1 mul_U9529(.A(n16116), .Y(n1914));
AND2X1 mul_U9530(.A(dpath_mulcore_array2_s2[15]), .B(n8962), .Y(n16119));
INVX1 mul_U9531(.A(n16119), .Y(n1915));
AND2X1 mul_U9532(.A(dpath_mulcore_a1s[66]), .B(dpath_mulcore_a1c[65]), .Y(n16121));
INVX1 mul_U9533(.A(n16121), .Y(dpath_mulcore_array2_c1[82]));
AND2X1 mul_U9534(.A(n8275), .B(dpath_mulcore_array2_s2[14]), .Y(n16123));
INVX1 mul_U9535(.A(n16123), .Y(n1916));
AND2X1 mul_U9536(.A(n8276), .B(dpath_mulcore_array2_s2[13]), .Y(n16126));
INVX1 mul_U9537(.A(n16126), .Y(n1917));
AND2X1 mul_U9538(.A(n8277), .B(dpath_mulcore_array2_s2[12]), .Y(n16129));
INVX1 mul_U9539(.A(n16129), .Y(n1918));
AND2X1 mul_U9540(.A(n8278), .B(dpath_mulcore_array2_s2[11]), .Y(n16132));
INVX1 mul_U9541(.A(n16132), .Y(n1919));
AND2X1 mul_U9542(.A(n8279), .B(dpath_mulcore_array2_s2[10]), .Y(n16135));
INVX1 mul_U9543(.A(n16135), .Y(n1920));
AND2X1 mul_U9544(.A(n8280), .B(dpath_mulcore_array2_s2[9]), .Y(n16138));
INVX1 mul_U9545(.A(n16138), .Y(n1921));
AND2X1 mul_U9546(.A(n8281), .B(dpath_mulcore_array2_s2[8]), .Y(n16141));
INVX1 mul_U9547(.A(n16141), .Y(n1922));
AND2X1 mul_U9548(.A(n8282), .B(dpath_mulcore_array2_s2[7]), .Y(n16144));
INVX1 mul_U9549(.A(n16144), .Y(n1923));
AND2X1 mul_U9550(.A(n8283), .B(dpath_mulcore_array2_s2[6]), .Y(n16147));
INVX1 mul_U9551(.A(n16147), .Y(n1924));
AND2X1 mul_U9552(.A(n8284), .B(dpath_mulcore_array2_s2[5]), .Y(n16150));
INVX1 mul_U9553(.A(n16150), .Y(n1925));
AND2X1 mul_U9554(.A(dpath_mulcore_a0s[67]), .B(n8973), .Y(n16153));
INVX1 mul_U9555(.A(n16153), .Y(n1926));
AND2X1 mul_U9556(.A(dpath_mulcore_ps[46]), .B(dpath_mulcore_pc[45]), .Y(n16156));
INVX1 mul_U9557(.A(n16156), .Y(n1927));
AND2X1 mul_U9558(.A(dpath_mulcore_ps[45]), .B(dpath_mulcore_pc[44]), .Y(n16159));
INVX1 mul_U9559(.A(n16159), .Y(n1928));
AND2X1 mul_U9560(.A(dpath_mulcore_ps[44]), .B(dpath_mulcore_pc[43]), .Y(n16162));
INVX1 mul_U9561(.A(n16162), .Y(n1929));
AND2X1 mul_U9562(.A(dpath_mulcore_ps[43]), .B(dpath_mulcore_pc[42]), .Y(n16165));
INVX1 mul_U9563(.A(n16165), .Y(n1930));
AND2X1 mul_U9564(.A(dpath_mulcore_ps[42]), .B(dpath_mulcore_pc[41]), .Y(n16168));
INVX1 mul_U9565(.A(n16168), .Y(n1931));
AND2X1 mul_U9566(.A(dpath_mulcore_ps[41]), .B(dpath_mulcore_pc[40]), .Y(n16171));
INVX1 mul_U9567(.A(n16171), .Y(n1932));
AND2X1 mul_U9568(.A(dpath_mulcore_ps[40]), .B(dpath_mulcore_pc[39]), .Y(n16174));
INVX1 mul_U9569(.A(n16174), .Y(n1933));
AND2X1 mul_U9570(.A(dpath_mulcore_ps[39]), .B(dpath_mulcore_pc[38]), .Y(n16177));
INVX1 mul_U9571(.A(n16177), .Y(n1934));
AND2X1 mul_U9572(.A(dpath_mulcore_ps[38]), .B(dpath_mulcore_pc[37]), .Y(n16180));
INVX1 mul_U9573(.A(n16180), .Y(n1935));
AND2X1 mul_U9574(.A(dpath_mulcore_ps[37]), .B(dpath_mulcore_pc[36]), .Y(n16183));
INVX1 mul_U9575(.A(n16183), .Y(n1936));
AND2X1 mul_U9576(.A(dpath_mulcore_array2_s1[14]), .B(n8963), .Y(n16186));
INVX1 mul_U9577(.A(n16186), .Y(n1937));
AND2X1 mul_U9578(.A(dpath_mulcore_array2_s1[13]), .B(n8964), .Y(n16189));
INVX1 mul_U9579(.A(n16189), .Y(n1938));
AND2X1 mul_U9580(.A(dpath_mulcore_array2_s1[12]), .B(n8965), .Y(n16192));
INVX1 mul_U9581(.A(n16192), .Y(n1939));
AND2X1 mul_U9582(.A(dpath_mulcore_array2_s1[11]), .B(n8966), .Y(n16195));
INVX1 mul_U9583(.A(n16195), .Y(n1940));
AND2X1 mul_U9584(.A(dpath_mulcore_array2_s1[10]), .B(n8967), .Y(n16198));
INVX1 mul_U9585(.A(n16198), .Y(n1941));
AND2X1 mul_U9586(.A(dpath_mulcore_array2_s1[9]), .B(n8968), .Y(n16201));
INVX1 mul_U9587(.A(n16201), .Y(n1942));
AND2X1 mul_U9588(.A(dpath_mulcore_array2_s1[8]), .B(n8969), .Y(n16204));
INVX1 mul_U9589(.A(n16204), .Y(n1943));
AND2X1 mul_U9590(.A(dpath_mulcore_array2_s1[7]), .B(n8970), .Y(n16207));
INVX1 mul_U9591(.A(n16207), .Y(n1944));
AND2X1 mul_U9592(.A(dpath_mulcore_array2_s1[6]), .B(n8971), .Y(n16210));
INVX1 mul_U9593(.A(n16210), .Y(n1945));
AND2X1 mul_U9594(.A(dpath_mulcore_array2_s1[5]), .B(n8972), .Y(n16213));
INVX1 mul_U9595(.A(n16213), .Y(n1946));
AND2X1 mul_U9596(.A(dpath_mulcore_array2_s1[82]), .B(n8948), .Y(n16216));
INVX1 mul_U9597(.A(n16216), .Y(n1947));
AND2X1 mul_U9598(.A(dpath_mulcore_ps[36]), .B(dpath_mulcore_pc[35]), .Y(n16219));
INVX1 mul_U9599(.A(n16219), .Y(n1948));
AND2X1 mul_U9600(.A(dpath_mulcore_ps[35]), .B(dpath_mulcore_pc[34]), .Y(n16222));
INVX1 mul_U9601(.A(n16222), .Y(n1949));
AND2X1 mul_U9602(.A(dpath_mulcore_ps[34]), .B(dpath_mulcore_pc[33]), .Y(n16225));
INVX1 mul_U9603(.A(n16225), .Y(n1950));
AND2X1 mul_U9604(.A(dpath_mulcore_ps[33]), .B(dpath_mulcore_pc[32]), .Y(n16228));
INVX1 mul_U9605(.A(n16228), .Y(n1951));
AND2X1 mul_U9606(.A(dpath_mulcore_a1c[49]), .B(dpath_mulcore_a0s[66]), .Y(n16231));
INVX1 mul_U9607(.A(n16231), .Y(n1952));
AND2X1 mul_U9608(.A(dpath_mulcore_a1c[48]), .B(dpath_mulcore_a0s[65]), .Y(n16234));
INVX1 mul_U9609(.A(n16234), .Y(n1953));
AND2X1 mul_U9610(.A(dpath_mulcore_a1c[47]), .B(dpath_mulcore_a0s[64]), .Y(n16237));
INVX1 mul_U9611(.A(n16237), .Y(n1954));
AND2X1 mul_U9612(.A(dpath_mulcore_a1c[46]), .B(dpath_mulcore_a0s[63]), .Y(n16240));
INVX1 mul_U9613(.A(n16240), .Y(n1955));
AND2X1 mul_U9614(.A(dpath_mulcore_a1c[45]), .B(dpath_mulcore_a0s[62]), .Y(n16243));
INVX1 mul_U9615(.A(n16243), .Y(n1956));
AND2X1 mul_U9616(.A(dpath_mulcore_a1c[44]), .B(dpath_mulcore_a0s[61]), .Y(n16246));
INVX1 mul_U9617(.A(n16246), .Y(n1957));
AND2X1 mul_U9618(.A(dpath_mulcore_a1c[43]), .B(dpath_mulcore_a0s[60]), .Y(n16249));
INVX1 mul_U9619(.A(n16249), .Y(n1958));
AND2X1 mul_U9620(.A(dpath_mulcore_a1c[42]), .B(dpath_mulcore_a0s[59]), .Y(n16252));
INVX1 mul_U9621(.A(n16252), .Y(n1959));
AND2X1 mul_U9622(.A(dpath_mulcore_a1c[41]), .B(dpath_mulcore_a0s[58]), .Y(n16255));
INVX1 mul_U9623(.A(n16255), .Y(n1960));
AND2X1 mul_U9624(.A(dpath_mulcore_a1c[40]), .B(dpath_mulcore_a0s[57]), .Y(n16258));
INVX1 mul_U9625(.A(n16258), .Y(n1961));
AND2X1 mul_U9626(.A(dpath_mulcore_a1c[39]), .B(dpath_mulcore_a0s[56]), .Y(n16261));
INVX1 mul_U9627(.A(n16261), .Y(n1962));
AND2X1 mul_U9628(.A(dpath_mulcore_a1c[38]), .B(dpath_mulcore_a0s[55]), .Y(n16264));
INVX1 mul_U9629(.A(n16264), .Y(n1963));
AND2X1 mul_U9630(.A(dpath_mulcore_a1c[37]), .B(dpath_mulcore_a0s[54]), .Y(n16267));
INVX1 mul_U9631(.A(n16267), .Y(n1964));
AND2X1 mul_U9632(.A(dpath_mulcore_a1c[36]), .B(dpath_mulcore_a0s[53]), .Y(n16270));
INVX1 mul_U9633(.A(n16270), .Y(n1965));
AND2X1 mul_U9634(.A(dpath_mulcore_a1c[35]), .B(dpath_mulcore_a0s[52]), .Y(n16273));
INVX1 mul_U9635(.A(n16273), .Y(n1966));
AND2X1 mul_U9636(.A(dpath_mulcore_a1c[34]), .B(dpath_mulcore_a0s[51]), .Y(n16276));
INVX1 mul_U9637(.A(n16276), .Y(n1967));
AND2X1 mul_U9638(.A(dpath_mulcore_a1c[33]), .B(dpath_mulcore_a0s[50]), .Y(n16279));
INVX1 mul_U9639(.A(n16279), .Y(n1968));
AND2X1 mul_U9640(.A(dpath_mulcore_a1c[32]), .B(dpath_mulcore_a0s[49]), .Y(n16282));
INVX1 mul_U9641(.A(n16282), .Y(n1969));
AND2X1 mul_U9642(.A(dpath_mulcore_a1c[31]), .B(dpath_mulcore_a0s[48]), .Y(n16285));
INVX1 mul_U9643(.A(n16285), .Y(n1970));
AND2X1 mul_U9644(.A(dpath_mulcore_a1c[30]), .B(dpath_mulcore_a0s[47]), .Y(n16288));
INVX1 mul_U9645(.A(n16288), .Y(n1971));
AND2X1 mul_U9646(.A(dpath_mulcore_a1c[29]), .B(dpath_mulcore_a0s[46]), .Y(n16291));
INVX1 mul_U9647(.A(n16291), .Y(n1972));
AND2X1 mul_U9648(.A(dpath_mulcore_a1c[28]), .B(dpath_mulcore_a0s[45]), .Y(n16294));
INVX1 mul_U9649(.A(n16294), .Y(n1973));
AND2X1 mul_U9650(.A(dpath_mulcore_a1c[27]), .B(dpath_mulcore_a0s[44]), .Y(n16297));
INVX1 mul_U9651(.A(n16297), .Y(n1974));
AND2X1 mul_U9652(.A(dpath_mulcore_a1c[26]), .B(dpath_mulcore_a0s[43]), .Y(n16300));
INVX1 mul_U9653(.A(n16300), .Y(n1975));
AND2X1 mul_U9654(.A(dpath_mulcore_a1c[25]), .B(dpath_mulcore_a0s[42]), .Y(n16303));
INVX1 mul_U9655(.A(n16303), .Y(n1976));
AND2X1 mul_U9656(.A(dpath_mulcore_a1c[24]), .B(dpath_mulcore_a0s[41]), .Y(n16306));
INVX1 mul_U9657(.A(n16306), .Y(n1977));
AND2X1 mul_U9658(.A(dpath_mulcore_a1c[23]), .B(dpath_mulcore_a0s[40]), .Y(n16309));
INVX1 mul_U9659(.A(n16309), .Y(n1978));
AND2X1 mul_U9660(.A(dpath_mulcore_a1c[22]), .B(dpath_mulcore_a0s[39]), .Y(n16312));
INVX1 mul_U9661(.A(n16312), .Y(n1979));
AND2X1 mul_U9662(.A(dpath_mulcore_a1c[21]), .B(dpath_mulcore_a0s[38]), .Y(n16315));
INVX1 mul_U9663(.A(n16315), .Y(n1980));
AND2X1 mul_U9664(.A(dpath_mulcore_a1c[20]), .B(dpath_mulcore_a0s[37]), .Y(n16318));
INVX1 mul_U9665(.A(n16318), .Y(n1981));
AND2X1 mul_U9666(.A(dpath_mulcore_a1c[19]), .B(dpath_mulcore_a0s[36]), .Y(n16321));
INVX1 mul_U9667(.A(n16321), .Y(n1982));
AND2X1 mul_U9668(.A(dpath_mulcore_a1c[18]), .B(dpath_mulcore_a0s[35]), .Y(n16324));
INVX1 mul_U9669(.A(n16324), .Y(n1983));
AND2X1 mul_U9670(.A(dpath_mulcore_a1c[17]), .B(dpath_mulcore_a0s[34]), .Y(n16327));
INVX1 mul_U9671(.A(n16327), .Y(n1984));
AND2X1 mul_U9672(.A(dpath_mulcore_a1c[16]), .B(dpath_mulcore_a0s[33]), .Y(n16330));
INVX1 mul_U9673(.A(n16330), .Y(n1985));
AND2X1 mul_U9674(.A(dpath_mulcore_a1c[15]), .B(dpath_mulcore_a0s[32]), .Y(n16333));
INVX1 mul_U9675(.A(n16333), .Y(n1986));
AND2X1 mul_U9676(.A(dpath_mulcore_a1c[14]), .B(dpath_mulcore_a0s[31]), .Y(n16336));
INVX1 mul_U9677(.A(n16336), .Y(n1987));
AND2X1 mul_U9678(.A(dpath_mulcore_a1c[13]), .B(dpath_mulcore_a0s[30]), .Y(n16339));
INVX1 mul_U9679(.A(n16339), .Y(n1988));
AND2X1 mul_U9680(.A(dpath_mulcore_a1c[12]), .B(dpath_mulcore_a0s[29]), .Y(n16342));
INVX1 mul_U9681(.A(n16342), .Y(n1989));
AND2X1 mul_U9682(.A(dpath_mulcore_a1c[11]), .B(dpath_mulcore_a0s[28]), .Y(n16345));
INVX1 mul_U9683(.A(n16345), .Y(n1990));
AND2X1 mul_U9684(.A(dpath_mulcore_a1c[10]), .B(dpath_mulcore_a0s[27]), .Y(n16348));
INVX1 mul_U9685(.A(n16348), .Y(n1991));
AND2X1 mul_U9686(.A(dpath_mulcore_a1c[9]), .B(dpath_mulcore_a0s[26]), .Y(n16351));
INVX1 mul_U9687(.A(n16351), .Y(n1992));
AND2X1 mul_U9688(.A(dpath_mulcore_a1c[8]), .B(dpath_mulcore_a0s[25]), .Y(n16354));
INVX1 mul_U9689(.A(n16354), .Y(n1993));
AND2X1 mul_U9690(.A(dpath_mulcore_a1c[7]), .B(dpath_mulcore_a0s[24]), .Y(n16357));
INVX1 mul_U9691(.A(n16357), .Y(n1994));
AND2X1 mul_U9692(.A(dpath_mulcore_a1c[6]), .B(dpath_mulcore_a0s[23]), .Y(n16360));
INVX1 mul_U9693(.A(n16360), .Y(n1995));
AND2X1 mul_U9694(.A(dpath_mulcore_a1c[5]), .B(dpath_mulcore_a0s[22]), .Y(n16363));
INVX1 mul_U9695(.A(n16363), .Y(n1996));
AND2X1 mul_U9696(.A(dpath_mulcore_a1c[4]), .B(dpath_mulcore_a0s[21]), .Y(n16366));
INVX1 mul_U9697(.A(n16366), .Y(n1997));
AND2X1 mul_U9698(.A(dpath_mulcore_ps[98]), .B(dpath_mulcore_pc[97]), .Y(n16370));
INVX1 mul_U9699(.A(n16370), .Y(n1998));
AND2X1 mul_U9700(.A(dpath_mulcore_ps[97]), .B(dpath_mulcore_pc[96]), .Y(n16373));
INVX1 mul_U9701(.A(n16373), .Y(n1999));
AND2X1 mul_U9702(.A(dpath_mulcore_ps[96]), .B(dpath_mulcore_pc[95]), .Y(n16376));
INVX1 mul_U9703(.A(n16376), .Y(n2000));
AND2X1 mul_U9704(.A(dpath_mulcore_ps[95]), .B(dpath_mulcore_pc[94]), .Y(n16379));
INVX1 mul_U9705(.A(n16379), .Y(n2001));
AND2X1 mul_U9706(.A(dpath_mulcore_ps[94]), .B(dpath_mulcore_pc[93]), .Y(n16382));
INVX1 mul_U9707(.A(n16382), .Y(n2002));
AND2X1 mul_U9708(.A(dpath_mulcore_ps[93]), .B(dpath_mulcore_pc[92]), .Y(n16385));
INVX1 mul_U9709(.A(n16385), .Y(n2003));
AND2X1 mul_U9710(.A(dpath_mulcore_ps[92]), .B(dpath_mulcore_pc[91]), .Y(n16388));
INVX1 mul_U9711(.A(n16388), .Y(n2004));
AND2X1 mul_U9712(.A(dpath_mulcore_ps[91]), .B(dpath_mulcore_pc[90]), .Y(n16391));
INVX1 mul_U9713(.A(n16391), .Y(n2005));
AND2X1 mul_U9714(.A(dpath_mulcore_ps[90]), .B(dpath_mulcore_pc[89]), .Y(n16394));
INVX1 mul_U9715(.A(n16394), .Y(n2006));
AND2X1 mul_U9716(.A(dpath_mulcore_ps[89]), .B(dpath_mulcore_pc[88]), .Y(n16397));
INVX1 mul_U9717(.A(n16397), .Y(n2007));
AND2X1 mul_U9718(.A(dpath_mulcore_ps[88]), .B(dpath_mulcore_pc[87]), .Y(n16400));
INVX1 mul_U9719(.A(n16400), .Y(n2008));
AND2X1 mul_U9720(.A(dpath_mulcore_ps[87]), .B(dpath_mulcore_pc[86]), .Y(n16403));
INVX1 mul_U9721(.A(n16403), .Y(n2009));
AND2X1 mul_U9722(.A(dpath_mulcore_ps[86]), .B(dpath_mulcore_pc[85]), .Y(n16406));
INVX1 mul_U9723(.A(n16406), .Y(n2010));
AND2X1 mul_U9724(.A(dpath_mulcore_ps[85]), .B(dpath_mulcore_pc[84]), .Y(n16409));
INVX1 mul_U9725(.A(n16409), .Y(n2011));
AND2X1 mul_U9726(.A(dpath_mulcore_ps[84]), .B(dpath_mulcore_pc[83]), .Y(n16412));
INVX1 mul_U9727(.A(n16412), .Y(n2012));
AND2X1 mul_U9728(.A(dpath_mulcore_ps[83]), .B(dpath_mulcore_pc[82]), .Y(n16415));
INVX1 mul_U9729(.A(n16415), .Y(n2013));
AND2X1 mul_U9730(.A(dpath_mulcore_ps[82]), .B(dpath_mulcore_pc[81]), .Y(n16418));
INVX1 mul_U9731(.A(n16418), .Y(n2014));
AND2X1 mul_U9732(.A(dpath_mulcore_ps[81]), .B(dpath_mulcore_pc[80]), .Y(n16421));
INVX1 mul_U9733(.A(n16421), .Y(n2015));
AND2X1 mul_U9734(.A(dpath_mulcore_ps[80]), .B(dpath_mulcore_pc[79]), .Y(n16424));
INVX1 mul_U9735(.A(n16424), .Y(n2016));
AND2X1 mul_U9736(.A(dpath_mulcore_ps[79]), .B(dpath_mulcore_pc[78]), .Y(n16427));
INVX1 mul_U9737(.A(n16427), .Y(n2017));
AND2X1 mul_U9738(.A(dpath_mulcore_ps[78]), .B(dpath_mulcore_pc[77]), .Y(n16430));
INVX1 mul_U9739(.A(n16430), .Y(n2018));
AND2X1 mul_U9740(.A(dpath_mulcore_ps[77]), .B(dpath_mulcore_pc[76]), .Y(n16433));
INVX1 mul_U9741(.A(n16433), .Y(n2019));
AND2X1 mul_U9742(.A(dpath_mulcore_ps[76]), .B(dpath_mulcore_pc[75]), .Y(n16436));
INVX1 mul_U9743(.A(n16436), .Y(n2020));
AND2X1 mul_U9744(.A(dpath_mulcore_ps[75]), .B(dpath_mulcore_pc[74]), .Y(n16439));
INVX1 mul_U9745(.A(n16439), .Y(n2021));
AND2X1 mul_U9746(.A(dpath_mulcore_ps[74]), .B(dpath_mulcore_pc[73]), .Y(n16442));
INVX1 mul_U9747(.A(n16442), .Y(n2022));
AND2X1 mul_U9748(.A(dpath_mulcore_ps[73]), .B(dpath_mulcore_pc[72]), .Y(n16445));
INVX1 mul_U9749(.A(n16445), .Y(n2023));
AND2X1 mul_U9750(.A(dpath_mulcore_ps[72]), .B(dpath_mulcore_pc[71]), .Y(n16448));
INVX1 mul_U9751(.A(n16448), .Y(n2024));
AND2X1 mul_U9752(.A(dpath_mulcore_ps[71]), .B(dpath_mulcore_pc[70]), .Y(n16451));
INVX1 mul_U9753(.A(n16451), .Y(n2025));
AND2X1 mul_U9754(.A(dpath_mulcore_ps[70]), .B(dpath_mulcore_pc[69]), .Y(n16454));
INVX1 mul_U9755(.A(n16454), .Y(n2026));
AND2X1 mul_U9756(.A(dpath_mulcore_ps[69]), .B(dpath_mulcore_pc[68]), .Y(n16457));
INVX1 mul_U9757(.A(n16457), .Y(n2027));
AND2X1 mul_U9758(.A(dpath_mulcore_ps[68]), .B(dpath_mulcore_pc[67]), .Y(n16460));
INVX1 mul_U9759(.A(n16460), .Y(n2028));
AND2X1 mul_U9760(.A(dpath_mulcore_ps[67]), .B(dpath_mulcore_pc[66]), .Y(n16463));
INVX1 mul_U9761(.A(n16463), .Y(n2029));
AND2X1 mul_U9762(.A(dpath_mulcore_ps[66]), .B(dpath_mulcore_pc[65]), .Y(n16466));
INVX1 mul_U9763(.A(n16466), .Y(n2030));
AND2X1 mul_U9764(.A(dpath_mulcore_ps[65]), .B(dpath_mulcore_pc[64]), .Y(n16469));
INVX1 mul_U9765(.A(n16469), .Y(n2031));
AND2X1 mul_U9766(.A(dpath_mulcore_ps[64]), .B(dpath_mulcore_pc[63]), .Y(n16472));
INVX1 mul_U9767(.A(n16472), .Y(n2032));
AND2X1 mul_U9768(.A(dpath_mulcore_ps[63]), .B(dpath_mulcore_pc[62]), .Y(n16475));
INVX1 mul_U9769(.A(n16475), .Y(n2033));
AND2X1 mul_U9770(.A(dpath_mulcore_ps[62]), .B(dpath_mulcore_pc[61]), .Y(n16478));
INVX1 mul_U9771(.A(n16478), .Y(n2034));
AND2X1 mul_U9772(.A(dpath_mulcore_ps[61]), .B(dpath_mulcore_pc[60]), .Y(n16481));
INVX1 mul_U9773(.A(n16481), .Y(n2035));
AND2X1 mul_U9774(.A(dpath_mulcore_ps[60]), .B(dpath_mulcore_pc[59]), .Y(n16484));
INVX1 mul_U9775(.A(n16484), .Y(n2036));
AND2X1 mul_U9776(.A(dpath_mulcore_ps[59]), .B(dpath_mulcore_pc[58]), .Y(n16487));
INVX1 mul_U9777(.A(n16487), .Y(n2037));
AND2X1 mul_U9778(.A(dpath_mulcore_ps[58]), .B(dpath_mulcore_pc[57]), .Y(n16490));
INVX1 mul_U9779(.A(n16490), .Y(n2038));
AND2X1 mul_U9780(.A(dpath_mulcore_ps[57]), .B(dpath_mulcore_pc[56]), .Y(n16493));
INVX1 mul_U9781(.A(n16493), .Y(n2039));
AND2X1 mul_U9782(.A(dpath_mulcore_ps[56]), .B(dpath_mulcore_pc[55]), .Y(n16496));
INVX1 mul_U9783(.A(n16496), .Y(n2040));
AND2X1 mul_U9784(.A(dpath_mulcore_ps[55]), .B(dpath_mulcore_pc[54]), .Y(n16499));
INVX1 mul_U9785(.A(n16499), .Y(n2041));
AND2X1 mul_U9786(.A(dpath_mulcore_ps[54]), .B(dpath_mulcore_pc[53]), .Y(n16502));
INVX1 mul_U9787(.A(n16502), .Y(n2042));
AND2X1 mul_U9788(.A(dpath_mulcore_ps[53]), .B(dpath_mulcore_pc[52]), .Y(n16505));
INVX1 mul_U9789(.A(n16505), .Y(n2043));
AND2X1 mul_U9790(.A(dpath_mulcore_ps[52]), .B(dpath_mulcore_pc[51]), .Y(n16508));
INVX1 mul_U9791(.A(n16508), .Y(n2044));
AND2X1 mul_U9792(.A(dpath_mulcore_array2_s1[81]), .B(n8949), .Y(n16510));
INVX1 mul_U9793(.A(n16510), .Y(dpath_mulcore_array2_c2[81]));
AND2X1 mul_U9794(.A(dpath_mulcore_array2_s1[80]), .B(n8950), .Y(n16512));
INVX1 mul_U9795(.A(n16512), .Y(n2045));
AND2X1 mul_U9796(.A(dpath_mulcore_array2_s1[79]), .B(n8951), .Y(n16515));
INVX1 mul_U9797(.A(n16515), .Y(n2046));
AND2X1 mul_U9798(.A(dpath_mulcore_array2_s1[78]), .B(n8952), .Y(n16518));
INVX1 mul_U9799(.A(n16518), .Y(n2047));
AND2X1 mul_U9800(.A(dpath_mulcore_array2_s1[77]), .B(n8953), .Y(n16521));
INVX1 mul_U9801(.A(n16521), .Y(n2048));
AND2X1 mul_U9802(.A(dpath_mulcore_array2_s1[76]), .B(n8954), .Y(n16524));
INVX1 mul_U9803(.A(n16524), .Y(n2049));
AND2X1 mul_U9804(.A(dpath_mulcore_array2_s1[75]), .B(n8955), .Y(n16527));
INVX1 mul_U9805(.A(n16527), .Y(n2050));
AND2X1 mul_U9806(.A(dpath_mulcore_array2_s1[74]), .B(n8956), .Y(n16530));
INVX1 mul_U9807(.A(n16530), .Y(n2051));
AND2X1 mul_U9808(.A(dpath_mulcore_array2_s1[73]), .B(n8957), .Y(n16533));
INVX1 mul_U9809(.A(n16533), .Y(n2052));
AND2X1 mul_U9810(.A(dpath_mulcore_array2_s1[72]), .B(n8958), .Y(n16536));
INVX1 mul_U9811(.A(n16536), .Y(n2053));
AND2X1 mul_U9812(.A(dpath_mulcore_array2_s1[71]), .B(n8959), .Y(n16539));
INVX1 mul_U9813(.A(n16539), .Y(n2054));
AND2X1 mul_U9814(.A(dpath_mulcore_array2_s1[70]), .B(n8960), .Y(n16542));
INVX1 mul_U9815(.A(n16542), .Y(n2055));
AND2X1 mul_U9816(.A(dpath_mulcore_array2_s1[69]), .B(n8961), .Y(n16545));
INVX1 mul_U9817(.A(n16545), .Y(n2056));
AND2X1 mul_U9818(.A(dpath_mulcore_array2_s1[68]), .B(n8974), .Y(n16548));
INVX1 mul_U9819(.A(n16548), .Y(n2057));
AND2X1 mul_U9820(.A(n8265), .B(dpath_mulcore_array2_s3[19]), .Y(n16551));
INVX1 mul_U9821(.A(n16551), .Y(n2058));
AND2X1 mul_U9822(.A(n8266), .B(dpath_mulcore_array2_s3[18]), .Y(n16554));
INVX1 mul_U9823(.A(n16554), .Y(n2059));
AND2X1 mul_U9824(.A(n8267), .B(dpath_mulcore_array2_s3[17]), .Y(n16557));
INVX1 mul_U9825(.A(n16557), .Y(n2060));
AND2X1 mul_U9826(.A(n8268), .B(dpath_mulcore_array2_s3[16]), .Y(n16560));
INVX1 mul_U9827(.A(n16560), .Y(n2061));
AND2X1 mul_U9828(.A(dpath_mulcore_ps[32]), .B(dpath_mulcore_pc[31]), .Y(n16565));
INVX1 mul_U9829(.A(n16565), .Y(n2062));
AND2X1 mul_U9830(.A(n7480), .B(n9853), .Y(n16575));
INVX1 mul_U9831(.A(n16575), .Y(n2063));
AND2X1 mul_U9832(.A(n7479), .B(n8448), .Y(n16578));
INVX1 mul_U9833(.A(n16578), .Y(n2064));
AND2X1 mul_U9834(.A(n7484), .B(n9475), .Y(n16583));
INVX1 mul_U9835(.A(n16583), .Y(n2065));
AND2X1 mul_U9836(.A(n7485), .B(n8754), .Y(n16586));
INVX1 mul_U9837(.A(n16586), .Y(n2066));
AND2X1 mul_U9838(.A(n5218), .B(n4696), .Y(dpath_mulcore_a0cout[75]));
INVX1 mul_U9839(.A(dpath_mulcore_a0cout[75]), .Y(n2067));
AND2X1 mul_U9840(.A(n5219), .B(n4697), .Y(dpath_mulcore_a0cout[74]));
INVX1 mul_U9841(.A(dpath_mulcore_a0cout[74]), .Y(n2068));
AND2X1 mul_U9842(.A(n5220), .B(n4698), .Y(dpath_mulcore_a0cout[73]));
INVX1 mul_U9843(.A(dpath_mulcore_a0cout[73]), .Y(n2069));
AND2X1 mul_U9844(.A(n5221), .B(n4699), .Y(dpath_mulcore_a0cout[72]));
INVX1 mul_U9845(.A(dpath_mulcore_a0cout[72]), .Y(n2070));
AND2X1 mul_U9846(.A(n5222), .B(n4700), .Y(dpath_mulcore_a0cout[76]));
INVX1 mul_U9847(.A(dpath_mulcore_a0cout[76]), .Y(n2071));
AND2X1 mul_U9848(.A(dpath_mulcore_ary1_a0_s_2[70]), .B(n9313), .Y(n16606));
INVX1 mul_U9849(.A(n16606), .Y(n2072));
AND2X1 mul_U9850(.A(n5223), .B(n4701), .Y(dpath_mulcore_a0cout[70]));
INVX1 mul_U9851(.A(dpath_mulcore_a0cout[70]), .Y(n2073));
AND2X1 mul_U9852(.A(dpath_mulcore_ary1_a0_s_2[69]), .B(n9314), .Y(n16613));
INVX1 mul_U9853(.A(n16613), .Y(n2074));
AND2X1 mul_U9854(.A(n5224), .B(n4702), .Y(dpath_mulcore_a0cout[69]));
INVX1 mul_U9855(.A(dpath_mulcore_a0cout[69]), .Y(n2075));
AND2X1 mul_U9856(.A(dpath_mulcore_ary1_a0_s_2[68]), .B(n9315), .Y(n16620));
INVX1 mul_U9857(.A(n16620), .Y(n2076));
AND2X1 mul_U9858(.A(n5225), .B(n4703), .Y(dpath_mulcore_a0cout[68]));
INVX1 mul_U9859(.A(dpath_mulcore_a0cout[68]), .Y(n2077));
AND2X1 mul_U9860(.A(dpath_mulcore_ary1_a0_s_2[67]), .B(n9316), .Y(n16627));
INVX1 mul_U9861(.A(n16627), .Y(n2078));
AND2X1 mul_U9862(.A(n5226), .B(n4704), .Y(dpath_mulcore_a0cout[67]));
INVX1 mul_U9863(.A(dpath_mulcore_a0cout[67]), .Y(n2079));
AND2X1 mul_U9864(.A(dpath_mulcore_ary1_a0_s_2[66]), .B(n9317), .Y(n16634));
INVX1 mul_U9865(.A(n16634), .Y(n2080));
AND2X1 mul_U9866(.A(n5227), .B(n4705), .Y(dpath_mulcore_a0cout[66]));
INVX1 mul_U9867(.A(dpath_mulcore_a0cout[66]), .Y(n2081));
AND2X1 mul_U9868(.A(dpath_mulcore_ary1_a0_s_2[65]), .B(n9318), .Y(n16641));
INVX1 mul_U9869(.A(n16641), .Y(n2082));
AND2X1 mul_U9870(.A(n5228), .B(n4706), .Y(dpath_mulcore_a0cout[65]));
INVX1 mul_U9871(.A(dpath_mulcore_a0cout[65]), .Y(n2083));
AND2X1 mul_U9872(.A(dpath_mulcore_ary1_a0_s_2[64]), .B(n9319), .Y(n16648));
INVX1 mul_U9873(.A(n16648), .Y(n2084));
AND2X1 mul_U9874(.A(n5229), .B(n4707), .Y(dpath_mulcore_a0cout[64]));
INVX1 mul_U9875(.A(dpath_mulcore_a0cout[64]), .Y(n2085));
AND2X1 mul_U9876(.A(dpath_mulcore_ary1_a0_s_2[63]), .B(n9320), .Y(n16655));
INVX1 mul_U9877(.A(n16655), .Y(n2086));
AND2X1 mul_U9878(.A(n5230), .B(n4708), .Y(dpath_mulcore_a0cout[63]));
INVX1 mul_U9879(.A(dpath_mulcore_a0cout[63]), .Y(n2087));
AND2X1 mul_U9880(.A(dpath_mulcore_ary1_a0_s_2[62]), .B(n9321), .Y(n16662));
INVX1 mul_U9881(.A(n16662), .Y(n2088));
AND2X1 mul_U9882(.A(n5231), .B(n4709), .Y(dpath_mulcore_a0cout[62]));
INVX1 mul_U9883(.A(dpath_mulcore_a0cout[62]), .Y(n2089));
AND2X1 mul_U9884(.A(dpath_mulcore_ary1_a0_s_2[61]), .B(n9322), .Y(n16669));
INVX1 mul_U9885(.A(n16669), .Y(n2090));
AND2X1 mul_U9886(.A(n5232), .B(n4710), .Y(dpath_mulcore_a0cout[61]));
INVX1 mul_U9887(.A(dpath_mulcore_a0cout[61]), .Y(n2091));
AND2X1 mul_U9888(.A(dpath_mulcore_ary1_a0_s_2[60]), .B(n9323), .Y(n16676));
INVX1 mul_U9889(.A(n16676), .Y(n2092));
AND2X1 mul_U9890(.A(n5233), .B(n4711), .Y(dpath_mulcore_a0cout[60]));
INVX1 mul_U9891(.A(dpath_mulcore_a0cout[60]), .Y(n2093));
AND2X1 mul_U9892(.A(dpath_mulcore_ary1_a0_s_2[59]), .B(n9324), .Y(n16683));
INVX1 mul_U9893(.A(n16683), .Y(n2094));
AND2X1 mul_U9894(.A(n5234), .B(n4712), .Y(dpath_mulcore_a0cout[59]));
INVX1 mul_U9895(.A(dpath_mulcore_a0cout[59]), .Y(n2095));
AND2X1 mul_U9896(.A(dpath_mulcore_ary1_a0_s_2[58]), .B(n9325), .Y(n16690));
INVX1 mul_U9897(.A(n16690), .Y(n2096));
AND2X1 mul_U9898(.A(n5235), .B(n4713), .Y(dpath_mulcore_a0cout[58]));
INVX1 mul_U9899(.A(dpath_mulcore_a0cout[58]), .Y(n2097));
AND2X1 mul_U9900(.A(dpath_mulcore_ary1_a0_s_2[57]), .B(n9326), .Y(n16697));
INVX1 mul_U9901(.A(n16697), .Y(n2098));
AND2X1 mul_U9902(.A(n5236), .B(n4714), .Y(dpath_mulcore_a0cout[57]));
INVX1 mul_U9903(.A(dpath_mulcore_a0cout[57]), .Y(n2099));
AND2X1 mul_U9904(.A(dpath_mulcore_ary1_a0_s_2[56]), .B(n9327), .Y(n16704));
INVX1 mul_U9905(.A(n16704), .Y(n2100));
AND2X1 mul_U9906(.A(n5237), .B(n4715), .Y(dpath_mulcore_a0cout[56]));
INVX1 mul_U9907(.A(dpath_mulcore_a0cout[56]), .Y(n2101));
AND2X1 mul_U9908(.A(dpath_mulcore_ary1_a0_s_2[55]), .B(n9328), .Y(n16711));
INVX1 mul_U9909(.A(n16711), .Y(n2102));
AND2X1 mul_U9910(.A(n5238), .B(n4716), .Y(dpath_mulcore_a0cout[55]));
INVX1 mul_U9911(.A(dpath_mulcore_a0cout[55]), .Y(n2103));
AND2X1 mul_U9912(.A(dpath_mulcore_ary1_a0_s_2[54]), .B(n9329), .Y(n16718));
INVX1 mul_U9913(.A(n16718), .Y(n2104));
AND2X1 mul_U9914(.A(n5239), .B(n4717), .Y(dpath_mulcore_a0cout[54]));
INVX1 mul_U9915(.A(dpath_mulcore_a0cout[54]), .Y(n2105));
AND2X1 mul_U9916(.A(dpath_mulcore_ary1_a0_s_2[53]), .B(n9330), .Y(n16725));
INVX1 mul_U9917(.A(n16725), .Y(n2106));
AND2X1 mul_U9918(.A(n5240), .B(n4718), .Y(dpath_mulcore_a0cout[53]));
INVX1 mul_U9919(.A(dpath_mulcore_a0cout[53]), .Y(n2107));
AND2X1 mul_U9920(.A(dpath_mulcore_ary1_a0_s_2[52]), .B(n9331), .Y(n16732));
INVX1 mul_U9921(.A(n16732), .Y(n2108));
AND2X1 mul_U9922(.A(n5241), .B(n4719), .Y(dpath_mulcore_a0cout[52]));
INVX1 mul_U9923(.A(dpath_mulcore_a0cout[52]), .Y(n2109));
AND2X1 mul_U9924(.A(dpath_mulcore_ary1_a0_s_2[51]), .B(n9332), .Y(n16739));
INVX1 mul_U9925(.A(n16739), .Y(n2110));
AND2X1 mul_U9926(.A(n5242), .B(n4720), .Y(dpath_mulcore_a0cout[51]));
INVX1 mul_U9927(.A(dpath_mulcore_a0cout[51]), .Y(n2111));
AND2X1 mul_U9928(.A(dpath_mulcore_ary1_a0_s_2[50]), .B(n9333), .Y(n16746));
INVX1 mul_U9929(.A(n16746), .Y(n2112));
AND2X1 mul_U9930(.A(n5243), .B(n4721), .Y(dpath_mulcore_a0cout[50]));
INVX1 mul_U9931(.A(dpath_mulcore_a0cout[50]), .Y(n2113));
AND2X1 mul_U9932(.A(dpath_mulcore_ary1_a0_s_2[49]), .B(n9334), .Y(n16753));
INVX1 mul_U9933(.A(n16753), .Y(n2114));
AND2X1 mul_U9934(.A(n5244), .B(n4722), .Y(dpath_mulcore_a0cout[49]));
INVX1 mul_U9935(.A(dpath_mulcore_a0cout[49]), .Y(n2115));
AND2X1 mul_U9936(.A(dpath_mulcore_ary1_a0_s_2[48]), .B(n9335), .Y(n16760));
INVX1 mul_U9937(.A(n16760), .Y(n2116));
AND2X1 mul_U9938(.A(n5245), .B(n4723), .Y(dpath_mulcore_a0cout[48]));
INVX1 mul_U9939(.A(dpath_mulcore_a0cout[48]), .Y(n2117));
AND2X1 mul_U9940(.A(dpath_mulcore_ary1_a0_s_2[47]), .B(n9336), .Y(n16767));
INVX1 mul_U9941(.A(n16767), .Y(n2118));
AND2X1 mul_U9942(.A(n5246), .B(n4724), .Y(dpath_mulcore_a0cout[47]));
INVX1 mul_U9943(.A(dpath_mulcore_a0cout[47]), .Y(n2119));
AND2X1 mul_U9944(.A(dpath_mulcore_ary1_a0_s_2[46]), .B(n9337), .Y(n16774));
INVX1 mul_U9945(.A(n16774), .Y(n2120));
AND2X1 mul_U9946(.A(n5247), .B(n4725), .Y(dpath_mulcore_a0cout[46]));
INVX1 mul_U9947(.A(dpath_mulcore_a0cout[46]), .Y(n2121));
AND2X1 mul_U9948(.A(dpath_mulcore_ary1_a0_s_2[45]), .B(n9338), .Y(n16781));
INVX1 mul_U9949(.A(n16781), .Y(n2122));
AND2X1 mul_U9950(.A(n5248), .B(n4726), .Y(dpath_mulcore_a0cout[45]));
INVX1 mul_U9951(.A(dpath_mulcore_a0cout[45]), .Y(n2123));
AND2X1 mul_U9952(.A(dpath_mulcore_ary1_a0_s_2[44]), .B(n9339), .Y(n16788));
INVX1 mul_U9953(.A(n16788), .Y(n2124));
AND2X1 mul_U9954(.A(n5249), .B(n4727), .Y(dpath_mulcore_a0cout[44]));
INVX1 mul_U9955(.A(dpath_mulcore_a0cout[44]), .Y(n2125));
AND2X1 mul_U9956(.A(dpath_mulcore_ary1_a0_s_2[43]), .B(n9340), .Y(n16795));
INVX1 mul_U9957(.A(n16795), .Y(n2126));
AND2X1 mul_U9958(.A(n5250), .B(n4728), .Y(dpath_mulcore_a0cout[43]));
INVX1 mul_U9959(.A(dpath_mulcore_a0cout[43]), .Y(n2127));
AND2X1 mul_U9960(.A(dpath_mulcore_ary1_a0_s_2[42]), .B(n9341), .Y(n16802));
INVX1 mul_U9961(.A(n16802), .Y(n2128));
AND2X1 mul_U9962(.A(n5251), .B(n4729), .Y(dpath_mulcore_a0cout[42]));
INVX1 mul_U9963(.A(dpath_mulcore_a0cout[42]), .Y(n2129));
AND2X1 mul_U9964(.A(dpath_mulcore_ary1_a0_s_2[41]), .B(n9342), .Y(n16809));
INVX1 mul_U9965(.A(n16809), .Y(n2130));
AND2X1 mul_U9966(.A(n5252), .B(n4730), .Y(dpath_mulcore_a0cout[41]));
INVX1 mul_U9967(.A(dpath_mulcore_a0cout[41]), .Y(n2131));
AND2X1 mul_U9968(.A(dpath_mulcore_ary1_a0_s_2[40]), .B(n9343), .Y(n16816));
INVX1 mul_U9969(.A(n16816), .Y(n2132));
AND2X1 mul_U9970(.A(n5253), .B(n4731), .Y(dpath_mulcore_a0cout[40]));
INVX1 mul_U9971(.A(dpath_mulcore_a0cout[40]), .Y(n2133));
AND2X1 mul_U9972(.A(dpath_mulcore_ary1_a0_s_2[39]), .B(n9344), .Y(n16823));
INVX1 mul_U9973(.A(n16823), .Y(n2134));
AND2X1 mul_U9974(.A(n5254), .B(n4732), .Y(dpath_mulcore_a0cout[39]));
INVX1 mul_U9975(.A(dpath_mulcore_a0cout[39]), .Y(n2135));
AND2X1 mul_U9976(.A(dpath_mulcore_ary1_a0_s_2[38]), .B(n9345), .Y(n16830));
INVX1 mul_U9977(.A(n16830), .Y(n2136));
AND2X1 mul_U9978(.A(n5255), .B(n4733), .Y(dpath_mulcore_a0cout[38]));
INVX1 mul_U9979(.A(dpath_mulcore_a0cout[38]), .Y(n2137));
AND2X1 mul_U9980(.A(dpath_mulcore_ary1_a0_s_2[37]), .B(n9346), .Y(n16837));
INVX1 mul_U9981(.A(n16837), .Y(n2138));
AND2X1 mul_U9982(.A(n5256), .B(n4734), .Y(dpath_mulcore_a0cout[37]));
INVX1 mul_U9983(.A(dpath_mulcore_a0cout[37]), .Y(n2139));
AND2X1 mul_U9984(.A(dpath_mulcore_ary1_a0_s_2[36]), .B(n9347), .Y(n16844));
INVX1 mul_U9985(.A(n16844), .Y(n2140));
AND2X1 mul_U9986(.A(n5257), .B(n4735), .Y(dpath_mulcore_a0cout[36]));
INVX1 mul_U9987(.A(dpath_mulcore_a0cout[36]), .Y(n2141));
AND2X1 mul_U9988(.A(dpath_mulcore_ary1_a0_s_2[35]), .B(n9348), .Y(n16851));
INVX1 mul_U9989(.A(n16851), .Y(n2142));
AND2X1 mul_U9990(.A(n5258), .B(n4736), .Y(dpath_mulcore_a0cout[35]));
INVX1 mul_U9991(.A(dpath_mulcore_a0cout[35]), .Y(n2143));
AND2X1 mul_U9992(.A(dpath_mulcore_ary1_a0_s_2[34]), .B(n9349), .Y(n16858));
INVX1 mul_U9993(.A(n16858), .Y(n2144));
AND2X1 mul_U9994(.A(n5259), .B(n4737), .Y(dpath_mulcore_a0cout[34]));
INVX1 mul_U9995(.A(dpath_mulcore_a0cout[34]), .Y(n2145));
AND2X1 mul_U9996(.A(dpath_mulcore_ary1_a0_s_2[33]), .B(n9350), .Y(n16865));
INVX1 mul_U9997(.A(n16865), .Y(n2146));
AND2X1 mul_U9998(.A(n5260), .B(n4738), .Y(dpath_mulcore_a0cout[33]));
INVX1 mul_U9999(.A(dpath_mulcore_a0cout[33]), .Y(n2147));
AND2X1 mul_U10000(.A(dpath_mulcore_ary1_a0_s_2[32]), .B(n9351), .Y(n16872));
INVX1 mul_U10001(.A(n16872), .Y(n2148));
AND2X1 mul_U10002(.A(n5261), .B(n4739), .Y(dpath_mulcore_a0cout[32]));
INVX1 mul_U10003(.A(dpath_mulcore_a0cout[32]), .Y(n2149));
AND2X1 mul_U10004(.A(dpath_mulcore_ary1_a0_s_2[31]), .B(n9352), .Y(n16879));
INVX1 mul_U10005(.A(n16879), .Y(n2150));
AND2X1 mul_U10006(.A(n5262), .B(n4740), .Y(dpath_mulcore_a0cout[31]));
INVX1 mul_U10007(.A(dpath_mulcore_a0cout[31]), .Y(n2151));
AND2X1 mul_U10008(.A(dpath_mulcore_ary1_a0_s_2[30]), .B(n9353), .Y(n16886));
INVX1 mul_U10009(.A(n16886), .Y(n2152));
AND2X1 mul_U10010(.A(n5263), .B(n4741), .Y(dpath_mulcore_a0cout[30]));
INVX1 mul_U10011(.A(dpath_mulcore_a0cout[30]), .Y(n2153));
AND2X1 mul_U10012(.A(dpath_mulcore_ary1_a0_s_2[29]), .B(n9354), .Y(n16893));
INVX1 mul_U10013(.A(n16893), .Y(n2154));
AND2X1 mul_U10014(.A(n5264), .B(n4742), .Y(dpath_mulcore_a0cout[29]));
INVX1 mul_U10015(.A(dpath_mulcore_a0cout[29]), .Y(n2155));
AND2X1 mul_U10016(.A(dpath_mulcore_ary1_a0_s_2[28]), .B(n9355), .Y(n16900));
INVX1 mul_U10017(.A(n16900), .Y(n2156));
AND2X1 mul_U10018(.A(n5265), .B(n4743), .Y(dpath_mulcore_a0cout[28]));
INVX1 mul_U10019(.A(dpath_mulcore_a0cout[28]), .Y(n2157));
AND2X1 mul_U10020(.A(dpath_mulcore_ary1_a0_s_2[27]), .B(n9356), .Y(n16907));
INVX1 mul_U10021(.A(n16907), .Y(n2158));
AND2X1 mul_U10022(.A(n5266), .B(n4744), .Y(dpath_mulcore_a0cout[27]));
INVX1 mul_U10023(.A(dpath_mulcore_a0cout[27]), .Y(n2159));
AND2X1 mul_U10024(.A(dpath_mulcore_ary1_a0_s_2[26]), .B(n9357), .Y(n16914));
INVX1 mul_U10025(.A(n16914), .Y(n2160));
AND2X1 mul_U10026(.A(n5267), .B(n4745), .Y(dpath_mulcore_a0cout[26]));
INVX1 mul_U10027(.A(dpath_mulcore_a0cout[26]), .Y(n2161));
AND2X1 mul_U10028(.A(dpath_mulcore_ary1_a0_s_2[25]), .B(n9358), .Y(n16921));
INVX1 mul_U10029(.A(n16921), .Y(n2162));
AND2X1 mul_U10030(.A(n5268), .B(n4746), .Y(dpath_mulcore_a0cout[25]));
INVX1 mul_U10031(.A(dpath_mulcore_a0cout[25]), .Y(n2163));
AND2X1 mul_U10032(.A(dpath_mulcore_ary1_a0_s_2[24]), .B(n9359), .Y(n16928));
INVX1 mul_U10033(.A(n16928), .Y(n2164));
AND2X1 mul_U10034(.A(n5269), .B(n4747), .Y(dpath_mulcore_a0cout[24]));
INVX1 mul_U10035(.A(dpath_mulcore_a0cout[24]), .Y(n2165));
AND2X1 mul_U10036(.A(dpath_mulcore_ary1_a0_s_2[23]), .B(n9360), .Y(n16935));
INVX1 mul_U10037(.A(n16935), .Y(n2166));
AND2X1 mul_U10038(.A(n5270), .B(n4748), .Y(dpath_mulcore_a0cout[23]));
INVX1 mul_U10039(.A(dpath_mulcore_a0cout[23]), .Y(n2167));
AND2X1 mul_U10040(.A(dpath_mulcore_ary1_a0_s_2[22]), .B(n9361), .Y(n16942));
INVX1 mul_U10041(.A(n16942), .Y(n2168));
AND2X1 mul_U10042(.A(n5271), .B(n4749), .Y(dpath_mulcore_a0cout[22]));
INVX1 mul_U10043(.A(dpath_mulcore_a0cout[22]), .Y(n2169));
AND2X1 mul_U10044(.A(dpath_mulcore_ary1_a0_s_2[21]), .B(n9362), .Y(n16949));
INVX1 mul_U10045(.A(n16949), .Y(n2170));
AND2X1 mul_U10046(.A(n5272), .B(n4750), .Y(dpath_mulcore_a0cout[21]));
INVX1 mul_U10047(.A(dpath_mulcore_a0cout[21]), .Y(n2171));
AND2X1 mul_U10048(.A(dpath_mulcore_ary1_a0_s_2[20]), .B(n9363), .Y(n16956));
INVX1 mul_U10049(.A(n16956), .Y(n2172));
AND2X1 mul_U10050(.A(n5273), .B(n4751), .Y(dpath_mulcore_a0cout[20]));
INVX1 mul_U10051(.A(dpath_mulcore_a0cout[20]), .Y(n2173));
AND2X1 mul_U10052(.A(dpath_mulcore_ary1_a0_s_2[19]), .B(n9364), .Y(n16963));
INVX1 mul_U10053(.A(n16963), .Y(n2174));
AND2X1 mul_U10054(.A(n5274), .B(n4752), .Y(dpath_mulcore_a0cout[19]));
INVX1 mul_U10055(.A(dpath_mulcore_a0cout[19]), .Y(n2175));
AND2X1 mul_U10056(.A(dpath_mulcore_ary1_a0_s_2[18]), .B(n9365), .Y(n16970));
INVX1 mul_U10057(.A(n16970), .Y(n2176));
AND2X1 mul_U10058(.A(n5275), .B(n4753), .Y(dpath_mulcore_a0cout[18]));
INVX1 mul_U10059(.A(dpath_mulcore_a0cout[18]), .Y(n2177));
AND2X1 mul_U10060(.A(dpath_mulcore_ary1_a0_s_2[17]), .B(n9366), .Y(n16977));
INVX1 mul_U10061(.A(n16977), .Y(n2178));
AND2X1 mul_U10062(.A(n5276), .B(n4754), .Y(dpath_mulcore_a0cout[17]));
INVX1 mul_U10063(.A(dpath_mulcore_a0cout[17]), .Y(n2179));
AND2X1 mul_U10064(.A(dpath_mulcore_ary1_a0_s_2[16]), .B(n9367), .Y(n16984));
INVX1 mul_U10065(.A(n16984), .Y(n2180));
AND2X1 mul_U10066(.A(n5277), .B(n4755), .Y(dpath_mulcore_a0cout[16]));
INVX1 mul_U10067(.A(dpath_mulcore_a0cout[16]), .Y(n2181));
AND2X1 mul_U10068(.A(dpath_mulcore_ary1_a0_s_2[15]), .B(n9368), .Y(n16991));
INVX1 mul_U10069(.A(n16991), .Y(n2182));
AND2X1 mul_U10070(.A(n5278), .B(n4756), .Y(dpath_mulcore_a0cout[15]));
INVX1 mul_U10071(.A(dpath_mulcore_a0cout[15]), .Y(n2183));
AND2X1 mul_U10072(.A(dpath_mulcore_ary1_a0_s_2[14]), .B(dpath_mulcore_ary1_a0_c_1[13]), .Y(n16998));
INVX1 mul_U10073(.A(n16998), .Y(n2184));
AND2X1 mul_U10074(.A(n5279), .B(n4757), .Y(dpath_mulcore_a0cout[14]));
INVX1 mul_U10075(.A(dpath_mulcore_a0cout[14]), .Y(n2185));
AND2X1 mul_U10076(.A(dpath_mulcore_ary1_a0_s_2[13]), .B(dpath_mulcore_ary1_a0_c_1[12]), .Y(n17005));
INVX1 mul_U10077(.A(n17005), .Y(n2186));
AND2X1 mul_U10078(.A(n5280), .B(n4758), .Y(dpath_mulcore_a0cout[13]));
INVX1 mul_U10079(.A(dpath_mulcore_a0cout[13]), .Y(n2187));
AND2X1 mul_U10080(.A(dpath_mulcore_ary1_a0_s_2[12]), .B(dpath_mulcore_ary1_a0_c_1[11]), .Y(n17012));
INVX1 mul_U10081(.A(n17012), .Y(n2188));
AND2X1 mul_U10082(.A(n5281), .B(n4759), .Y(dpath_mulcore_a0cout[12]));
INVX1 mul_U10083(.A(dpath_mulcore_a0cout[12]), .Y(n2189));
AND2X1 mul_U10084(.A(dpath_mulcore_ary1_a0_s_2[11]), .B(dpath_mulcore_ary1_a0_c_1[10]), .Y(n17019));
INVX1 mul_U10085(.A(n17019), .Y(n2190));
AND2X1 mul_U10086(.A(dpath_mulcore_ary1_a1_s_2[71]), .B(dpath_mulcore_ary1_a1_s1[64]), .Y(n17025));
INVX1 mul_U10087(.A(n17025), .Y(n2191));
AND2X1 mul_U10088(.A(n5282), .B(n4760), .Y(dpath_mulcore_a1cout[71]));
INVX1 mul_U10089(.A(dpath_mulcore_a1cout[71]), .Y(n2192));
AND2X1 mul_U10090(.A(n5283), .B(n4761), .Y(dpath_mulcore_a1cout[75]));
INVX1 mul_U10091(.A(dpath_mulcore_a1cout[75]), .Y(n2193));
AND2X1 mul_U10092(.A(n5284), .B(n4762), .Y(dpath_mulcore_a1cout[74]));
INVX1 mul_U10093(.A(dpath_mulcore_a1cout[74]), .Y(n2194));
AND2X1 mul_U10094(.A(n5285), .B(n4763), .Y(dpath_mulcore_a1cout[73]));
INVX1 mul_U10095(.A(dpath_mulcore_a1cout[73]), .Y(n2195));
AND2X1 mul_U10096(.A(n5286), .B(n4764), .Y(dpath_mulcore_a1cout[72]));
INVX1 mul_U10097(.A(dpath_mulcore_a1cout[72]), .Y(n2196));
AND2X1 mul_U10098(.A(n5287), .B(n4765), .Y(dpath_mulcore_a1cout[76]));
INVX1 mul_U10099(.A(dpath_mulcore_a1cout[76]), .Y(n2197));
AND2X1 mul_U10100(.A(dpath_mulcore_ary1_a1_s_2[70]), .B(n9369), .Y(n17050));
INVX1 mul_U10101(.A(n17050), .Y(n2198));
AND2X1 mul_U10102(.A(n5288), .B(n4766), .Y(dpath_mulcore_a1cout[70]));
INVX1 mul_U10103(.A(dpath_mulcore_a1cout[70]), .Y(n2199));
AND2X1 mul_U10104(.A(dpath_mulcore_ary1_a1_s_2[69]), .B(n9370), .Y(n17057));
INVX1 mul_U10105(.A(n17057), .Y(n2200));
AND2X1 mul_U10106(.A(n5289), .B(n4767), .Y(dpath_mulcore_a1cout[69]));
INVX1 mul_U10107(.A(dpath_mulcore_a1cout[69]), .Y(n2201));
AND2X1 mul_U10108(.A(dpath_mulcore_ary1_a1_s_2[68]), .B(n9371), .Y(n17064));
INVX1 mul_U10109(.A(n17064), .Y(n2202));
AND2X1 mul_U10110(.A(n5290), .B(n4768), .Y(dpath_mulcore_a1cout[68]));
INVX1 mul_U10111(.A(dpath_mulcore_a1cout[68]), .Y(n2203));
AND2X1 mul_U10112(.A(dpath_mulcore_ary1_a1_s_2[67]), .B(n9372), .Y(n17071));
INVX1 mul_U10113(.A(n17071), .Y(n2204));
AND2X1 mul_U10114(.A(n5291), .B(n4769), .Y(dpath_mulcore_a1cout[67]));
INVX1 mul_U10115(.A(dpath_mulcore_a1cout[67]), .Y(n2205));
AND2X1 mul_U10116(.A(dpath_mulcore_ary1_a1_s_2[66]), .B(n9373), .Y(n17078));
INVX1 mul_U10117(.A(n17078), .Y(n2206));
AND2X1 mul_U10118(.A(n5292), .B(n4770), .Y(dpath_mulcore_a1cout[66]));
INVX1 mul_U10119(.A(dpath_mulcore_a1cout[66]), .Y(n2207));
AND2X1 mul_U10120(.A(dpath_mulcore_ary1_a1_s_2[65]), .B(n9374), .Y(n17085));
INVX1 mul_U10121(.A(n17085), .Y(n2208));
AND2X1 mul_U10122(.A(n5293), .B(n4771), .Y(dpath_mulcore_a1cout[65]));
INVX1 mul_U10123(.A(dpath_mulcore_a1cout[65]), .Y(n2209));
AND2X1 mul_U10124(.A(dpath_mulcore_ary1_a1_s_2[64]), .B(n9375), .Y(n17092));
INVX1 mul_U10125(.A(n17092), .Y(n2210));
AND2X1 mul_U10126(.A(n5294), .B(n4772), .Y(dpath_mulcore_a1cout[64]));
INVX1 mul_U10127(.A(dpath_mulcore_a1cout[64]), .Y(n2211));
AND2X1 mul_U10128(.A(dpath_mulcore_ary1_a1_s_2[63]), .B(n9376), .Y(n17099));
INVX1 mul_U10129(.A(n17099), .Y(n2212));
AND2X1 mul_U10130(.A(n5295), .B(n4773), .Y(dpath_mulcore_a1cout[63]));
INVX1 mul_U10131(.A(dpath_mulcore_a1cout[63]), .Y(n2213));
AND2X1 mul_U10132(.A(dpath_mulcore_ary1_a1_s_2[62]), .B(n9377), .Y(n17106));
INVX1 mul_U10133(.A(n17106), .Y(n2214));
AND2X1 mul_U10134(.A(n5296), .B(n4774), .Y(dpath_mulcore_a1cout[62]));
INVX1 mul_U10135(.A(dpath_mulcore_a1cout[62]), .Y(n2215));
AND2X1 mul_U10136(.A(dpath_mulcore_ary1_a1_s_2[61]), .B(n9378), .Y(n17113));
INVX1 mul_U10137(.A(n17113), .Y(n2216));
AND2X1 mul_U10138(.A(n5297), .B(n4775), .Y(dpath_mulcore_a1cout[61]));
INVX1 mul_U10139(.A(dpath_mulcore_a1cout[61]), .Y(n2217));
AND2X1 mul_U10140(.A(dpath_mulcore_ary1_a1_s_2[60]), .B(n9379), .Y(n17120));
INVX1 mul_U10141(.A(n17120), .Y(n2218));
AND2X1 mul_U10142(.A(n5298), .B(n4776), .Y(dpath_mulcore_a1cout[60]));
INVX1 mul_U10143(.A(dpath_mulcore_a1cout[60]), .Y(n2219));
AND2X1 mul_U10144(.A(dpath_mulcore_ary1_a1_s_2[59]), .B(n9380), .Y(n17127));
INVX1 mul_U10145(.A(n17127), .Y(n2220));
AND2X1 mul_U10146(.A(n5299), .B(n4777), .Y(dpath_mulcore_a1cout[59]));
INVX1 mul_U10147(.A(dpath_mulcore_a1cout[59]), .Y(n2221));
AND2X1 mul_U10148(.A(dpath_mulcore_ary1_a1_s_2[58]), .B(n9381), .Y(n17134));
INVX1 mul_U10149(.A(n17134), .Y(n2222));
AND2X1 mul_U10150(.A(n5300), .B(n4778), .Y(dpath_mulcore_a1cout[58]));
INVX1 mul_U10151(.A(dpath_mulcore_a1cout[58]), .Y(n2223));
AND2X1 mul_U10152(.A(dpath_mulcore_ary1_a1_s_2[57]), .B(n9382), .Y(n17141));
INVX1 mul_U10153(.A(n17141), .Y(n2224));
AND2X1 mul_U10154(.A(n5301), .B(n4779), .Y(dpath_mulcore_a1cout[57]));
INVX1 mul_U10155(.A(dpath_mulcore_a1cout[57]), .Y(n2225));
AND2X1 mul_U10156(.A(dpath_mulcore_ary1_a1_s_2[56]), .B(n9383), .Y(n17148));
INVX1 mul_U10157(.A(n17148), .Y(n2226));
AND2X1 mul_U10158(.A(n5302), .B(n4780), .Y(dpath_mulcore_a1cout[56]));
INVX1 mul_U10159(.A(dpath_mulcore_a1cout[56]), .Y(n2227));
AND2X1 mul_U10160(.A(dpath_mulcore_ary1_a1_s_2[55]), .B(n9384), .Y(n17155));
INVX1 mul_U10161(.A(n17155), .Y(n2228));
AND2X1 mul_U10162(.A(n5303), .B(n4781), .Y(dpath_mulcore_a1cout[55]));
INVX1 mul_U10163(.A(dpath_mulcore_a1cout[55]), .Y(n2229));
AND2X1 mul_U10164(.A(dpath_mulcore_ary1_a1_s_2[54]), .B(n9385), .Y(n17162));
INVX1 mul_U10165(.A(n17162), .Y(n2230));
AND2X1 mul_U10166(.A(n5304), .B(n4782), .Y(dpath_mulcore_a1cout[54]));
INVX1 mul_U10167(.A(dpath_mulcore_a1cout[54]), .Y(n2231));
AND2X1 mul_U10168(.A(dpath_mulcore_ary1_a1_s_2[53]), .B(n9386), .Y(n17169));
INVX1 mul_U10169(.A(n17169), .Y(n2232));
AND2X1 mul_U10170(.A(n5305), .B(n4783), .Y(dpath_mulcore_a1cout[53]));
INVX1 mul_U10171(.A(dpath_mulcore_a1cout[53]), .Y(n2233));
AND2X1 mul_U10172(.A(dpath_mulcore_ary1_a1_s_2[52]), .B(n9387), .Y(n17176));
INVX1 mul_U10173(.A(n17176), .Y(n2234));
AND2X1 mul_U10174(.A(n5306), .B(n4784), .Y(dpath_mulcore_a1cout[52]));
INVX1 mul_U10175(.A(dpath_mulcore_a1cout[52]), .Y(n2235));
AND2X1 mul_U10176(.A(dpath_mulcore_ary1_a1_s_2[51]), .B(n9388), .Y(n17183));
INVX1 mul_U10177(.A(n17183), .Y(n2236));
AND2X1 mul_U10178(.A(n5307), .B(n4785), .Y(dpath_mulcore_a1cout[51]));
INVX1 mul_U10179(.A(dpath_mulcore_a1cout[51]), .Y(n2237));
AND2X1 mul_U10180(.A(dpath_mulcore_ary1_a1_s_2[50]), .B(n9389), .Y(n17190));
INVX1 mul_U10181(.A(n17190), .Y(n2238));
AND2X1 mul_U10182(.A(n5308), .B(n4786), .Y(dpath_mulcore_a1cout[50]));
INVX1 mul_U10183(.A(dpath_mulcore_a1cout[50]), .Y(n2239));
AND2X1 mul_U10184(.A(dpath_mulcore_ary1_a1_s_2[49]), .B(n9390), .Y(n17197));
INVX1 mul_U10185(.A(n17197), .Y(n2240));
AND2X1 mul_U10186(.A(n5309), .B(n4787), .Y(dpath_mulcore_a1cout[49]));
INVX1 mul_U10187(.A(dpath_mulcore_a1cout[49]), .Y(n2241));
AND2X1 mul_U10188(.A(dpath_mulcore_ary1_a1_s_2[48]), .B(n9391), .Y(n17204));
INVX1 mul_U10189(.A(n17204), .Y(n2242));
AND2X1 mul_U10190(.A(n5310), .B(n4788), .Y(dpath_mulcore_a1cout[48]));
INVX1 mul_U10191(.A(dpath_mulcore_a1cout[48]), .Y(n2243));
AND2X1 mul_U10192(.A(dpath_mulcore_ary1_a1_s_2[47]), .B(n9392), .Y(n17211));
INVX1 mul_U10193(.A(n17211), .Y(n2244));
AND2X1 mul_U10194(.A(n5311), .B(n4789), .Y(dpath_mulcore_a1cout[47]));
INVX1 mul_U10195(.A(dpath_mulcore_a1cout[47]), .Y(n2245));
AND2X1 mul_U10196(.A(dpath_mulcore_ary1_a1_s_2[46]), .B(n9393), .Y(n17218));
INVX1 mul_U10197(.A(n17218), .Y(n2246));
AND2X1 mul_U10198(.A(n5312), .B(n4790), .Y(dpath_mulcore_a1cout[46]));
INVX1 mul_U10199(.A(dpath_mulcore_a1cout[46]), .Y(n2247));
AND2X1 mul_U10200(.A(dpath_mulcore_ary1_a1_s_2[45]), .B(n9394), .Y(n17225));
INVX1 mul_U10201(.A(n17225), .Y(n2248));
AND2X1 mul_U10202(.A(n5313), .B(n4791), .Y(dpath_mulcore_a1cout[45]));
INVX1 mul_U10203(.A(dpath_mulcore_a1cout[45]), .Y(n2249));
AND2X1 mul_U10204(.A(dpath_mulcore_ary1_a1_s_2[44]), .B(n9395), .Y(n17232));
INVX1 mul_U10205(.A(n17232), .Y(n2250));
AND2X1 mul_U10206(.A(n5314), .B(n4792), .Y(dpath_mulcore_a1cout[44]));
INVX1 mul_U10207(.A(dpath_mulcore_a1cout[44]), .Y(n2251));
AND2X1 mul_U10208(.A(dpath_mulcore_ary1_a1_s_2[43]), .B(n9396), .Y(n17239));
INVX1 mul_U10209(.A(n17239), .Y(n2252));
AND2X1 mul_U10210(.A(n5315), .B(n4793), .Y(dpath_mulcore_a1cout[43]));
INVX1 mul_U10211(.A(dpath_mulcore_a1cout[43]), .Y(n2253));
AND2X1 mul_U10212(.A(dpath_mulcore_ary1_a1_s_2[42]), .B(n9397), .Y(n17246));
INVX1 mul_U10213(.A(n17246), .Y(n2254));
AND2X1 mul_U10214(.A(n5316), .B(n4794), .Y(dpath_mulcore_a1cout[42]));
INVX1 mul_U10215(.A(dpath_mulcore_a1cout[42]), .Y(n2255));
AND2X1 mul_U10216(.A(dpath_mulcore_ary1_a1_s_2[41]), .B(n9398), .Y(n17253));
INVX1 mul_U10217(.A(n17253), .Y(n2256));
AND2X1 mul_U10218(.A(n5317), .B(n4795), .Y(dpath_mulcore_a1cout[41]));
INVX1 mul_U10219(.A(dpath_mulcore_a1cout[41]), .Y(n2257));
AND2X1 mul_U10220(.A(dpath_mulcore_ary1_a1_s_2[40]), .B(n9399), .Y(n17260));
INVX1 mul_U10221(.A(n17260), .Y(n2258));
AND2X1 mul_U10222(.A(n5318), .B(n4796), .Y(dpath_mulcore_a1cout[40]));
INVX1 mul_U10223(.A(dpath_mulcore_a1cout[40]), .Y(n2259));
AND2X1 mul_U10224(.A(dpath_mulcore_ary1_a1_s_2[39]), .B(n9400), .Y(n17267));
INVX1 mul_U10225(.A(n17267), .Y(n2260));
AND2X1 mul_U10226(.A(n5319), .B(n4797), .Y(dpath_mulcore_a1cout[39]));
INVX1 mul_U10227(.A(dpath_mulcore_a1cout[39]), .Y(n2261));
AND2X1 mul_U10228(.A(dpath_mulcore_ary1_a1_s_2[38]), .B(n9401), .Y(n17274));
INVX1 mul_U10229(.A(n17274), .Y(n2262));
AND2X1 mul_U10230(.A(n5320), .B(n4798), .Y(dpath_mulcore_a1cout[38]));
INVX1 mul_U10231(.A(dpath_mulcore_a1cout[38]), .Y(n2263));
AND2X1 mul_U10232(.A(dpath_mulcore_ary1_a1_s_2[37]), .B(n9402), .Y(n17281));
INVX1 mul_U10233(.A(n17281), .Y(n2264));
AND2X1 mul_U10234(.A(n5321), .B(n4799), .Y(dpath_mulcore_a1cout[37]));
INVX1 mul_U10235(.A(dpath_mulcore_a1cout[37]), .Y(n2265));
AND2X1 mul_U10236(.A(dpath_mulcore_ary1_a1_s_2[36]), .B(n9403), .Y(n17288));
INVX1 mul_U10237(.A(n17288), .Y(n2266));
AND2X1 mul_U10238(.A(n5322), .B(n4800), .Y(dpath_mulcore_a1cout[36]));
INVX1 mul_U10239(.A(dpath_mulcore_a1cout[36]), .Y(n2267));
AND2X1 mul_U10240(.A(dpath_mulcore_ary1_a1_s_2[35]), .B(n9404), .Y(n17295));
INVX1 mul_U10241(.A(n17295), .Y(n2268));
AND2X1 mul_U10242(.A(n5323), .B(n4801), .Y(dpath_mulcore_a1cout[35]));
INVX1 mul_U10243(.A(dpath_mulcore_a1cout[35]), .Y(n2269));
AND2X1 mul_U10244(.A(dpath_mulcore_ary1_a1_s_2[34]), .B(n9405), .Y(n17302));
INVX1 mul_U10245(.A(n17302), .Y(n2270));
AND2X1 mul_U10246(.A(n5324), .B(n4802), .Y(dpath_mulcore_a1cout[34]));
INVX1 mul_U10247(.A(dpath_mulcore_a1cout[34]), .Y(n2271));
AND2X1 mul_U10248(.A(dpath_mulcore_ary1_a1_s_2[33]), .B(n9406), .Y(n17309));
INVX1 mul_U10249(.A(n17309), .Y(n2272));
AND2X1 mul_U10250(.A(n5325), .B(n4803), .Y(dpath_mulcore_a1cout[33]));
INVX1 mul_U10251(.A(dpath_mulcore_a1cout[33]), .Y(n2273));
AND2X1 mul_U10252(.A(dpath_mulcore_ary1_a1_s_2[32]), .B(n9407), .Y(n17316));
INVX1 mul_U10253(.A(n17316), .Y(n2274));
AND2X1 mul_U10254(.A(n5326), .B(n4804), .Y(dpath_mulcore_a1cout[32]));
INVX1 mul_U10255(.A(dpath_mulcore_a1cout[32]), .Y(n2275));
AND2X1 mul_U10256(.A(dpath_mulcore_ary1_a1_s_2[31]), .B(n9408), .Y(n17323));
INVX1 mul_U10257(.A(n17323), .Y(n2276));
AND2X1 mul_U10258(.A(n5327), .B(n4805), .Y(dpath_mulcore_a1cout[31]));
INVX1 mul_U10259(.A(dpath_mulcore_a1cout[31]), .Y(n2277));
AND2X1 mul_U10260(.A(dpath_mulcore_ary1_a1_s_2[30]), .B(n9409), .Y(n17330));
INVX1 mul_U10261(.A(n17330), .Y(n2278));
AND2X1 mul_U10262(.A(n5328), .B(n4806), .Y(dpath_mulcore_a1cout[30]));
INVX1 mul_U10263(.A(dpath_mulcore_a1cout[30]), .Y(n2279));
AND2X1 mul_U10264(.A(dpath_mulcore_ary1_a1_s_2[29]), .B(n9410), .Y(n17337));
INVX1 mul_U10265(.A(n17337), .Y(n2280));
AND2X1 mul_U10266(.A(n5329), .B(n4807), .Y(dpath_mulcore_a1cout[29]));
INVX1 mul_U10267(.A(dpath_mulcore_a1cout[29]), .Y(n2281));
AND2X1 mul_U10268(.A(dpath_mulcore_ary1_a1_s_2[28]), .B(n9411), .Y(n17344));
INVX1 mul_U10269(.A(n17344), .Y(n2282));
AND2X1 mul_U10270(.A(n5330), .B(n4808), .Y(dpath_mulcore_a1cout[28]));
INVX1 mul_U10271(.A(dpath_mulcore_a1cout[28]), .Y(n2283));
AND2X1 mul_U10272(.A(dpath_mulcore_ary1_a1_s_2[27]), .B(n9412), .Y(n17351));
INVX1 mul_U10273(.A(n17351), .Y(n2284));
AND2X1 mul_U10274(.A(n5331), .B(n4809), .Y(dpath_mulcore_a1cout[27]));
INVX1 mul_U10275(.A(dpath_mulcore_a1cout[27]), .Y(n2285));
AND2X1 mul_U10276(.A(dpath_mulcore_ary1_a1_s_2[26]), .B(n9413), .Y(n17358));
INVX1 mul_U10277(.A(n17358), .Y(n2286));
AND2X1 mul_U10278(.A(n5332), .B(n4810), .Y(dpath_mulcore_a1cout[26]));
INVX1 mul_U10279(.A(dpath_mulcore_a1cout[26]), .Y(n2287));
AND2X1 mul_U10280(.A(dpath_mulcore_ary1_a1_s_2[25]), .B(n9414), .Y(n17365));
INVX1 mul_U10281(.A(n17365), .Y(n2288));
AND2X1 mul_U10282(.A(n5333), .B(n4811), .Y(dpath_mulcore_a1cout[25]));
INVX1 mul_U10283(.A(dpath_mulcore_a1cout[25]), .Y(n2289));
AND2X1 mul_U10284(.A(dpath_mulcore_ary1_a1_s_2[24]), .B(n9415), .Y(n17372));
INVX1 mul_U10285(.A(n17372), .Y(n2290));
AND2X1 mul_U10286(.A(n5334), .B(n4812), .Y(dpath_mulcore_a1cout[24]));
INVX1 mul_U10287(.A(dpath_mulcore_a1cout[24]), .Y(n2291));
AND2X1 mul_U10288(.A(dpath_mulcore_ary1_a1_s_2[23]), .B(n9416), .Y(n17379));
INVX1 mul_U10289(.A(n17379), .Y(n2292));
AND2X1 mul_U10290(.A(n5335), .B(n4813), .Y(dpath_mulcore_a1cout[23]));
INVX1 mul_U10291(.A(dpath_mulcore_a1cout[23]), .Y(n2293));
AND2X1 mul_U10292(.A(dpath_mulcore_ary1_a1_s_2[22]), .B(n9417), .Y(n17386));
INVX1 mul_U10293(.A(n17386), .Y(n2294));
AND2X1 mul_U10294(.A(n5336), .B(n4814), .Y(dpath_mulcore_a1cout[22]));
INVX1 mul_U10295(.A(dpath_mulcore_a1cout[22]), .Y(n2295));
AND2X1 mul_U10296(.A(dpath_mulcore_ary1_a1_s_2[21]), .B(n9418), .Y(n17393));
INVX1 mul_U10297(.A(n17393), .Y(n2296));
AND2X1 mul_U10298(.A(n5337), .B(n4815), .Y(dpath_mulcore_a1cout[21]));
INVX1 mul_U10299(.A(dpath_mulcore_a1cout[21]), .Y(n2297));
AND2X1 mul_U10300(.A(dpath_mulcore_ary1_a1_s_2[20]), .B(n9419), .Y(n17400));
INVX1 mul_U10301(.A(n17400), .Y(n2298));
AND2X1 mul_U10302(.A(n5338), .B(n4816), .Y(dpath_mulcore_a1cout[20]));
INVX1 mul_U10303(.A(dpath_mulcore_a1cout[20]), .Y(n2299));
AND2X1 mul_U10304(.A(dpath_mulcore_ary1_a1_s_2[19]), .B(n9420), .Y(n17407));
INVX1 mul_U10305(.A(n17407), .Y(n2300));
AND2X1 mul_U10306(.A(n5339), .B(n4817), .Y(dpath_mulcore_a1cout[19]));
INVX1 mul_U10307(.A(dpath_mulcore_a1cout[19]), .Y(n2301));
AND2X1 mul_U10308(.A(dpath_mulcore_ary1_a1_s_2[18]), .B(n9421), .Y(n17414));
INVX1 mul_U10309(.A(n17414), .Y(n2302));
AND2X1 mul_U10310(.A(n5340), .B(n4818), .Y(dpath_mulcore_a1cout[18]));
INVX1 mul_U10311(.A(dpath_mulcore_a1cout[18]), .Y(n2303));
AND2X1 mul_U10312(.A(dpath_mulcore_ary1_a1_s_2[17]), .B(n9422), .Y(n17421));
INVX1 mul_U10313(.A(n17421), .Y(n2304));
AND2X1 mul_U10314(.A(n5341), .B(n4819), .Y(dpath_mulcore_a1cout[17]));
INVX1 mul_U10315(.A(dpath_mulcore_a1cout[17]), .Y(n2305));
AND2X1 mul_U10316(.A(dpath_mulcore_ary1_a1_s_2[16]), .B(n9423), .Y(n17428));
INVX1 mul_U10317(.A(n17428), .Y(n2306));
AND2X1 mul_U10318(.A(n5342), .B(n4820), .Y(dpath_mulcore_a1cout[16]));
INVX1 mul_U10319(.A(dpath_mulcore_a1cout[16]), .Y(n2307));
AND2X1 mul_U10320(.A(dpath_mulcore_ary1_a1_s_2[15]), .B(n9424), .Y(n17435));
INVX1 mul_U10321(.A(n17435), .Y(n2308));
AND2X1 mul_U10322(.A(n5343), .B(n4821), .Y(dpath_mulcore_a1cout[15]));
INVX1 mul_U10323(.A(dpath_mulcore_a1cout[15]), .Y(n2309));
AND2X1 mul_U10324(.A(dpath_mulcore_ary1_a1_s_2[14]), .B(dpath_mulcore_ary1_a1_c_1[13]), .Y(n17442));
INVX1 mul_U10325(.A(n17442), .Y(n2310));
AND2X1 mul_U10326(.A(n5344), .B(n4822), .Y(dpath_mulcore_a1cout[14]));
INVX1 mul_U10327(.A(dpath_mulcore_a1cout[14]), .Y(n2311));
AND2X1 mul_U10328(.A(dpath_mulcore_ary1_a1_s_2[13]), .B(dpath_mulcore_ary1_a1_c_1[12]), .Y(n17449));
INVX1 mul_U10329(.A(n17449), .Y(n2312));
AND2X1 mul_U10330(.A(n5345), .B(n4823), .Y(dpath_mulcore_a1cout[13]));
INVX1 mul_U10331(.A(dpath_mulcore_a1cout[13]), .Y(n2313));
AND2X1 mul_U10332(.A(dpath_mulcore_ary1_a1_s_2[12]), .B(dpath_mulcore_ary1_a1_c_1[11]), .Y(n17456));
INVX1 mul_U10333(.A(n17456), .Y(n2314));
AND2X1 mul_U10334(.A(n5346), .B(n4824), .Y(dpath_mulcore_a1cout[12]));
INVX1 mul_U10335(.A(dpath_mulcore_a1cout[12]), .Y(n2315));
AND2X1 mul_U10336(.A(dpath_mulcore_ary1_a1_s_2[11]), .B(dpath_mulcore_ary1_a1_c_1[10]), .Y(n17463));
INVX1 mul_U10337(.A(n17463), .Y(n2316));
AND2X1 mul_U10338(.A(dpath_mulcore_array2_sc3_68__z), .B(n17471), .Y(n17469));
INVX1 mul_U10339(.A(n17469), .Y(n2317));
AND2X1 mul_U10340(.A(dpath_mulcore_array2_sc3_67__z), .B(n7348), .Y(n17472));
INVX1 mul_U10341(.A(n17472), .Y(n2318));
AND2X1 mul_U10342(.A(n9429), .B(dpath_mulcore_array2_s1[66]), .Y(n17475));
INVX1 mul_U10343(.A(n17475), .Y(n2319));
AND2X1 mul_U10344(.A(dpath_mulcore_array2_sc3_66__z), .B(n7349), .Y(n17478));
INVX1 mul_U10345(.A(n17478), .Y(n2320));
AND2X1 mul_U10346(.A(n9430), .B(dpath_mulcore_array2_s1[65]), .Y(n17482));
INVX1 mul_U10347(.A(n17482), .Y(n2321));
AND2X1 mul_U10348(.A(dpath_mulcore_array2_sc3_65__z), .B(n7350), .Y(n17485));
INVX1 mul_U10349(.A(n17485), .Y(n2322));
AND2X1 mul_U10350(.A(n9431), .B(dpath_mulcore_array2_s1[64]), .Y(n17489));
INVX1 mul_U10351(.A(n17489), .Y(n2323));
AND2X1 mul_U10352(.A(dpath_mulcore_array2_sc3_64__z), .B(n7351), .Y(n17492));
INVX1 mul_U10353(.A(n17492), .Y(n2324));
AND2X1 mul_U10354(.A(n9432), .B(dpath_mulcore_array2_s1[63]), .Y(n17496));
INVX1 mul_U10355(.A(n17496), .Y(n2325));
AND2X1 mul_U10356(.A(dpath_mulcore_array2_sc3_63__z), .B(n7352), .Y(n17499));
INVX1 mul_U10357(.A(n17499), .Y(n2326));
AND2X1 mul_U10358(.A(n9433), .B(dpath_mulcore_array2_s1[62]), .Y(n17503));
INVX1 mul_U10359(.A(n17503), .Y(n2327));
AND2X1 mul_U10360(.A(dpath_mulcore_array2_sc3_62__z), .B(n7353), .Y(n17506));
INVX1 mul_U10361(.A(n17506), .Y(n2328));
AND2X1 mul_U10362(.A(n9434), .B(dpath_mulcore_array2_s1[61]), .Y(n17510));
INVX1 mul_U10363(.A(n17510), .Y(n2329));
AND2X1 mul_U10364(.A(dpath_mulcore_array2_sc3_61__z), .B(n7354), .Y(n17513));
INVX1 mul_U10365(.A(n17513), .Y(n2330));
AND2X1 mul_U10366(.A(n9435), .B(dpath_mulcore_array2_s1[60]), .Y(n17517));
INVX1 mul_U10367(.A(n17517), .Y(n2331));
AND2X1 mul_U10368(.A(dpath_mulcore_array2_sc3_60__z), .B(n7355), .Y(n17520));
INVX1 mul_U10369(.A(n17520), .Y(n2332));
AND2X1 mul_U10370(.A(n9436), .B(dpath_mulcore_array2_s1[59]), .Y(n17524));
INVX1 mul_U10371(.A(n17524), .Y(n2333));
AND2X1 mul_U10372(.A(dpath_mulcore_array2_sc3_59__z), .B(n7356), .Y(n17527));
INVX1 mul_U10373(.A(n17527), .Y(n2334));
AND2X1 mul_U10374(.A(n9437), .B(dpath_mulcore_array2_s1[58]), .Y(n17531));
INVX1 mul_U10375(.A(n17531), .Y(n2335));
AND2X1 mul_U10376(.A(dpath_mulcore_array2_sc3_58__z), .B(n7357), .Y(n17534));
INVX1 mul_U10377(.A(n17534), .Y(n2336));
AND2X1 mul_U10378(.A(n9438), .B(dpath_mulcore_array2_s1[57]), .Y(n17538));
INVX1 mul_U10379(.A(n17538), .Y(n2337));
AND2X1 mul_U10380(.A(dpath_mulcore_array2_sc3_57__z), .B(n7358), .Y(n17541));
INVX1 mul_U10381(.A(n17541), .Y(n2338));
AND2X1 mul_U10382(.A(n9439), .B(dpath_mulcore_array2_s1[56]), .Y(n17545));
INVX1 mul_U10383(.A(n17545), .Y(n2339));
AND2X1 mul_U10384(.A(dpath_mulcore_array2_sc3_56__z), .B(n7359), .Y(n17548));
INVX1 mul_U10385(.A(n17548), .Y(n2340));
AND2X1 mul_U10386(.A(n9440), .B(dpath_mulcore_array2_s1[55]), .Y(n17552));
INVX1 mul_U10387(.A(n17552), .Y(n2341));
AND2X1 mul_U10388(.A(dpath_mulcore_array2_sc3_55__z), .B(n7360), .Y(n17555));
INVX1 mul_U10389(.A(n17555), .Y(n2342));
AND2X1 mul_U10390(.A(n9441), .B(dpath_mulcore_array2_s1[54]), .Y(n17559));
INVX1 mul_U10391(.A(n17559), .Y(n2343));
AND2X1 mul_U10392(.A(dpath_mulcore_array2_sc3_54__z), .B(n7361), .Y(n17562));
INVX1 mul_U10393(.A(n17562), .Y(n2344));
AND2X1 mul_U10394(.A(n9442), .B(dpath_mulcore_array2_s1[53]), .Y(n17566));
INVX1 mul_U10395(.A(n17566), .Y(n2345));
AND2X1 mul_U10396(.A(dpath_mulcore_array2_sc3_53__z), .B(n7362), .Y(n17569));
INVX1 mul_U10397(.A(n17569), .Y(n2346));
AND2X1 mul_U10398(.A(n9443), .B(dpath_mulcore_array2_s1[52]), .Y(n17573));
INVX1 mul_U10399(.A(n17573), .Y(n2347));
AND2X1 mul_U10400(.A(dpath_mulcore_array2_sc3_52__z), .B(n7363), .Y(n17576));
INVX1 mul_U10401(.A(n17576), .Y(n2348));
AND2X1 mul_U10402(.A(n9444), .B(dpath_mulcore_array2_s1[51]), .Y(n17580));
INVX1 mul_U10403(.A(n17580), .Y(n2349));
AND2X1 mul_U10404(.A(dpath_mulcore_array2_sc3_51__z), .B(n7364), .Y(n17583));
INVX1 mul_U10405(.A(n17583), .Y(n2350));
AND2X1 mul_U10406(.A(n9445), .B(dpath_mulcore_array2_s1[50]), .Y(n17587));
INVX1 mul_U10407(.A(n17587), .Y(n2351));
AND2X1 mul_U10408(.A(dpath_mulcore_array2_sc3_50__z), .B(n7365), .Y(n17590));
INVX1 mul_U10409(.A(n17590), .Y(n2352));
AND2X1 mul_U10410(.A(n9446), .B(dpath_mulcore_array2_s1[49]), .Y(n17594));
INVX1 mul_U10411(.A(n17594), .Y(n2353));
AND2X1 mul_U10412(.A(dpath_mulcore_array2_sc3_49__z), .B(n7366), .Y(n17597));
INVX1 mul_U10413(.A(n17597), .Y(n2354));
AND2X1 mul_U10414(.A(n9447), .B(dpath_mulcore_array2_s1[48]), .Y(n17601));
INVX1 mul_U10415(.A(n17601), .Y(n2355));
AND2X1 mul_U10416(.A(dpath_mulcore_array2_sc3_48__z), .B(n7367), .Y(n17604));
INVX1 mul_U10417(.A(n17604), .Y(n2356));
AND2X1 mul_U10418(.A(n9448), .B(dpath_mulcore_array2_s1[47]), .Y(n17608));
INVX1 mul_U10419(.A(n17608), .Y(n2357));
AND2X1 mul_U10420(.A(dpath_mulcore_array2_sc3_47__z), .B(n7368), .Y(n17611));
INVX1 mul_U10421(.A(n17611), .Y(n2358));
AND2X1 mul_U10422(.A(n9449), .B(dpath_mulcore_array2_s1[46]), .Y(n17615));
INVX1 mul_U10423(.A(n17615), .Y(n2359));
AND2X1 mul_U10424(.A(dpath_mulcore_array2_sc3_46__z), .B(n7369), .Y(n17618));
INVX1 mul_U10425(.A(n17618), .Y(n2360));
AND2X1 mul_U10426(.A(n9450), .B(dpath_mulcore_array2_s1[45]), .Y(n17622));
INVX1 mul_U10427(.A(n17622), .Y(n2361));
AND2X1 mul_U10428(.A(dpath_mulcore_array2_sc3_45__z), .B(n7370), .Y(n17625));
INVX1 mul_U10429(.A(n17625), .Y(n2362));
AND2X1 mul_U10430(.A(n9451), .B(dpath_mulcore_array2_s1[44]), .Y(n17629));
INVX1 mul_U10431(.A(n17629), .Y(n2363));
AND2X1 mul_U10432(.A(dpath_mulcore_array2_sc3_44__z), .B(n7371), .Y(n17632));
INVX1 mul_U10433(.A(n17632), .Y(n2364));
AND2X1 mul_U10434(.A(n9452), .B(dpath_mulcore_array2_s1[43]), .Y(n17636));
INVX1 mul_U10435(.A(n17636), .Y(n2365));
AND2X1 mul_U10436(.A(dpath_mulcore_array2_sc3_43__z), .B(n7372), .Y(n17639));
INVX1 mul_U10437(.A(n17639), .Y(n2366));
AND2X1 mul_U10438(.A(n9453), .B(dpath_mulcore_array2_s1[42]), .Y(n17643));
INVX1 mul_U10439(.A(n17643), .Y(n2367));
AND2X1 mul_U10440(.A(dpath_mulcore_array2_sc3_42__z), .B(n7373), .Y(n17646));
INVX1 mul_U10441(.A(n17646), .Y(n2368));
AND2X1 mul_U10442(.A(n9454), .B(dpath_mulcore_array2_s1[41]), .Y(n17650));
INVX1 mul_U10443(.A(n17650), .Y(n2369));
AND2X1 mul_U10444(.A(dpath_mulcore_array2_sc3_41__z), .B(n7374), .Y(n17653));
INVX1 mul_U10445(.A(n17653), .Y(n2370));
AND2X1 mul_U10446(.A(n9455), .B(dpath_mulcore_array2_s1[40]), .Y(n17657));
INVX1 mul_U10447(.A(n17657), .Y(n2371));
AND2X1 mul_U10448(.A(dpath_mulcore_array2_sc3_40__z), .B(n7375), .Y(n17660));
INVX1 mul_U10449(.A(n17660), .Y(n2372));
AND2X1 mul_U10450(.A(n9456), .B(dpath_mulcore_array2_s1[39]), .Y(n17664));
INVX1 mul_U10451(.A(n17664), .Y(n2373));
AND2X1 mul_U10452(.A(dpath_mulcore_array2_sc3_39__z), .B(n7376), .Y(n17667));
INVX1 mul_U10453(.A(n17667), .Y(n2374));
AND2X1 mul_U10454(.A(n9457), .B(dpath_mulcore_array2_s1[38]), .Y(n17671));
INVX1 mul_U10455(.A(n17671), .Y(n2375));
AND2X1 mul_U10456(.A(dpath_mulcore_array2_sc3_38__z), .B(n7377), .Y(n17674));
INVX1 mul_U10457(.A(n17674), .Y(n2376));
AND2X1 mul_U10458(.A(n9458), .B(dpath_mulcore_array2_s1[37]), .Y(n17678));
INVX1 mul_U10459(.A(n17678), .Y(n2377));
AND2X1 mul_U10460(.A(dpath_mulcore_array2_sc3_37__z), .B(n7378), .Y(n17681));
INVX1 mul_U10461(.A(n17681), .Y(n2378));
AND2X1 mul_U10462(.A(n9459), .B(dpath_mulcore_array2_s1[36]), .Y(n17685));
INVX1 mul_U10463(.A(n17685), .Y(n2379));
AND2X1 mul_U10464(.A(dpath_mulcore_array2_sc3_36__z), .B(n7379), .Y(n17688));
INVX1 mul_U10465(.A(n17688), .Y(n2380));
AND2X1 mul_U10466(.A(n9460), .B(dpath_mulcore_array2_s1[35]), .Y(n17692));
INVX1 mul_U10467(.A(n17692), .Y(n2381));
AND2X1 mul_U10468(.A(dpath_mulcore_array2_sc3_35__z), .B(n7380), .Y(n17695));
INVX1 mul_U10469(.A(n17695), .Y(n2382));
AND2X1 mul_U10470(.A(n9461), .B(dpath_mulcore_array2_s1[34]), .Y(n17699));
INVX1 mul_U10471(.A(n17699), .Y(n2383));
AND2X1 mul_U10472(.A(dpath_mulcore_array2_sc3_34__z), .B(n7381), .Y(n17702));
INVX1 mul_U10473(.A(n17702), .Y(n2384));
AND2X1 mul_U10474(.A(n9462), .B(dpath_mulcore_array2_s1[33]), .Y(n17706));
INVX1 mul_U10475(.A(n17706), .Y(n2385));
AND2X1 mul_U10476(.A(dpath_mulcore_array2_sc3_33__z), .B(n7382), .Y(n17709));
INVX1 mul_U10477(.A(n17709), .Y(n2386));
AND2X1 mul_U10478(.A(n9463), .B(dpath_mulcore_array2_s1[32]), .Y(n17713));
INVX1 mul_U10479(.A(n17713), .Y(n2387));
AND2X1 mul_U10480(.A(dpath_mulcore_array2_sc3_32__z), .B(n7383), .Y(n17716));
INVX1 mul_U10481(.A(n17716), .Y(n2388));
AND2X1 mul_U10482(.A(n9464), .B(dpath_mulcore_array2_s1[31]), .Y(n17720));
INVX1 mul_U10483(.A(n17720), .Y(n2389));
AND2X1 mul_U10484(.A(dpath_mulcore_array2_sc3_31__z), .B(n7384), .Y(n17723));
INVX1 mul_U10485(.A(n17723), .Y(n2390));
AND2X1 mul_U10486(.A(n9465), .B(dpath_mulcore_array2_s1[30]), .Y(n17727));
INVX1 mul_U10487(.A(n17727), .Y(n2391));
AND2X1 mul_U10488(.A(dpath_mulcore_array2_sc3_30__z), .B(n7385), .Y(n17730));
INVX1 mul_U10489(.A(n17730), .Y(n2392));
AND2X1 mul_U10490(.A(n9466), .B(dpath_mulcore_array2_s1[29]), .Y(n17734));
INVX1 mul_U10491(.A(n17734), .Y(n2393));
AND2X1 mul_U10492(.A(dpath_mulcore_array2_sc3_29__z), .B(n7386), .Y(n17737));
INVX1 mul_U10493(.A(n17737), .Y(n2394));
AND2X1 mul_U10494(.A(n9467), .B(dpath_mulcore_array2_s1[28]), .Y(n17741));
INVX1 mul_U10495(.A(n17741), .Y(n2395));
AND2X1 mul_U10496(.A(dpath_mulcore_array2_sc3_28__z), .B(n7387), .Y(n17744));
INVX1 mul_U10497(.A(n17744), .Y(n2396));
AND2X1 mul_U10498(.A(n9468), .B(dpath_mulcore_array2_s1[27]), .Y(n17748));
INVX1 mul_U10499(.A(n17748), .Y(n2397));
AND2X1 mul_U10500(.A(dpath_mulcore_array2_sc3_27__z), .B(n7388), .Y(n17751));
INVX1 mul_U10501(.A(n17751), .Y(n2398));
AND2X1 mul_U10502(.A(n9469), .B(dpath_mulcore_array2_s1[26]), .Y(n17755));
INVX1 mul_U10503(.A(n17755), .Y(n2399));
AND2X1 mul_U10504(.A(dpath_mulcore_array2_sc3_26__z), .B(n7389), .Y(n17758));
INVX1 mul_U10505(.A(n17758), .Y(n2400));
AND2X1 mul_U10506(.A(n9470), .B(dpath_mulcore_array2_s1[25]), .Y(n17762));
INVX1 mul_U10507(.A(n17762), .Y(n2401));
AND2X1 mul_U10508(.A(dpath_mulcore_array2_sc3_25__z), .B(n7390), .Y(n17765));
INVX1 mul_U10509(.A(n17765), .Y(n2402));
AND2X1 mul_U10510(.A(n9471), .B(dpath_mulcore_array2_s1[24]), .Y(n17769));
INVX1 mul_U10511(.A(n17769), .Y(n2403));
AND2X1 mul_U10512(.A(dpath_mulcore_array2_sc3_24__z), .B(n7391), .Y(n17772));
INVX1 mul_U10513(.A(n17772), .Y(n2404));
AND2X1 mul_U10514(.A(n9472), .B(dpath_mulcore_array2_s1[23]), .Y(n17776));
INVX1 mul_U10515(.A(n17776), .Y(n2405));
AND2X1 mul_U10516(.A(dpath_mulcore_array2_sc3_23__z), .B(n7392), .Y(n17779));
INVX1 mul_U10517(.A(n17779), .Y(n2406));
AND2X1 mul_U10518(.A(n9473), .B(dpath_mulcore_array2_s1[22]), .Y(n17783));
INVX1 mul_U10519(.A(n17783), .Y(n2407));
AND2X1 mul_U10520(.A(dpath_mulcore_array2_sc3_22__z), .B(n7393), .Y(n17786));
INVX1 mul_U10521(.A(n17786), .Y(n2408));
AND2X1 mul_U10522(.A(n16368), .B(dpath_mulcore_array2_s1[21]), .Y(n17790));
INVX1 mul_U10523(.A(n17790), .Y(n2409));
AND2X1 mul_U10524(.A(dpath_mulcore_array2_sc3_21__z), .B(n7394), .Y(n17793));
INVX1 mul_U10525(.A(n17793), .Y(n2410));
AND2X1 mul_U10526(.A(n9428), .B(dpath_mulcore_array2_s1[20]), .Y(n17797));
INVX1 mul_U10527(.A(n17797), .Y(n2411));
AND2X1 mul_U10528(.A(n5347), .B(n4825), .Y(dpath_mulcore_booth_b1_outmx[2]));
INVX1 mul_U10529(.A(dpath_mulcore_booth_b1_outmx[2]), .Y(n2412));
AND2X1 mul_U10530(.A(n5348), .B(n4826), .Y(dpath_mulcore_booth_b1_outmx[1]));
INVX1 mul_U10531(.A(dpath_mulcore_booth_b1_outmx[1]), .Y(n2413));
AND2X1 mul_U10532(.A(n5349), .B(n4827), .Y(dpath_mulcore_booth_b1_outmx[0]));
INVX1 mul_U10533(.A(dpath_mulcore_booth_b1_outmx[0]), .Y(n2414));
AND2X1 mul_U10534(.A(n5350), .B(n4828), .Y(dpath_mulcore_booth_b2_outmx[2]));
INVX1 mul_U10535(.A(dpath_mulcore_booth_b2_outmx[2]), .Y(n2415));
AND2X1 mul_U10536(.A(n5351), .B(n4829), .Y(dpath_mulcore_booth_b2_outmx[1]));
INVX1 mul_U10537(.A(dpath_mulcore_booth_b2_outmx[1]), .Y(n2416));
AND2X1 mul_U10538(.A(n5352), .B(n4830), .Y(dpath_mulcore_booth_b2_outmx[0]));
INVX1 mul_U10539(.A(dpath_mulcore_booth_b2_outmx[0]), .Y(n2417));
AND2X1 mul_U10540(.A(n5353), .B(n4831), .Y(dpath_mulcore_booth_b3_outmx[2]));
INVX1 mul_U10541(.A(dpath_mulcore_booth_b3_outmx[2]), .Y(n2418));
AND2X1 mul_U10542(.A(n5354), .B(n4832), .Y(dpath_mulcore_booth_b3_outmx[1]));
INVX1 mul_U10543(.A(dpath_mulcore_booth_b3_outmx[1]), .Y(n2419));
AND2X1 mul_U10544(.A(n5355), .B(n4833), .Y(dpath_mulcore_booth_b3_outmx[0]));
INVX1 mul_U10545(.A(dpath_mulcore_booth_b3_outmx[0]), .Y(n2420));
AND2X1 mul_U10546(.A(n5356), .B(n4834), .Y(dpath_mulcore_booth_b4_outmx[2]));
INVX1 mul_U10547(.A(dpath_mulcore_booth_b4_outmx[2]), .Y(n2421));
AND2X1 mul_U10548(.A(n5357), .B(n4835), .Y(dpath_mulcore_booth_b4_outmx[1]));
INVX1 mul_U10549(.A(dpath_mulcore_booth_b4_outmx[1]), .Y(n2422));
AND2X1 mul_U10550(.A(n5358), .B(n4836), .Y(dpath_mulcore_booth_b4_outmx[0]));
INVX1 mul_U10551(.A(dpath_mulcore_booth_b4_outmx[0]), .Y(n2423));
AND2X1 mul_U10552(.A(n5359), .B(n4837), .Y(dpath_mulcore_booth_b5_outmx[2]));
INVX1 mul_U10553(.A(dpath_mulcore_booth_b5_outmx[2]), .Y(n2424));
AND2X1 mul_U10554(.A(n5360), .B(n4838), .Y(dpath_mulcore_booth_b5_outmx[1]));
INVX1 mul_U10555(.A(dpath_mulcore_booth_b5_outmx[1]), .Y(n2425));
AND2X1 mul_U10556(.A(n5361), .B(n4839), .Y(dpath_mulcore_booth_b5_outmx[0]));
INVX1 mul_U10557(.A(dpath_mulcore_booth_b5_outmx[0]), .Y(n2426));
AND2X1 mul_U10558(.A(n5362), .B(n4840), .Y(dpath_mulcore_booth_b6_outmx[2]));
INVX1 mul_U10559(.A(dpath_mulcore_booth_b6_outmx[2]), .Y(n2427));
AND2X1 mul_U10560(.A(n5363), .B(n4841), .Y(dpath_mulcore_booth_b6_outmx[1]));
INVX1 mul_U10561(.A(dpath_mulcore_booth_b6_outmx[1]), .Y(n2428));
AND2X1 mul_U10562(.A(n5364), .B(n4842), .Y(dpath_mulcore_booth_b6_outmx[0]));
INVX1 mul_U10563(.A(dpath_mulcore_booth_b6_outmx[0]), .Y(n2429));
AND2X1 mul_U10564(.A(n5365), .B(n4843), .Y(dpath_mulcore_booth_b7_outmx[2]));
INVX1 mul_U10565(.A(dpath_mulcore_booth_b7_outmx[2]), .Y(n2430));
AND2X1 mul_U10566(.A(n5366), .B(n4844), .Y(dpath_mulcore_booth_b7_outmx[1]));
INVX1 mul_U10567(.A(dpath_mulcore_booth_b7_outmx[1]), .Y(n2431));
AND2X1 mul_U10568(.A(n5367), .B(n4845), .Y(dpath_mulcore_booth_b7_outmx[0]));
INVX1 mul_U10569(.A(dpath_mulcore_booth_b7_outmx[0]), .Y(n2432));
AND2X1 mul_U10570(.A(n5368), .B(n4846), .Y(dpath_mulcore_booth_b8_outmx[2]));
INVX1 mul_U10571(.A(dpath_mulcore_booth_b8_outmx[2]), .Y(n2433));
AND2X1 mul_U10572(.A(n5369), .B(n4847), .Y(dpath_mulcore_booth_b8_outmx[1]));
INVX1 mul_U10573(.A(dpath_mulcore_booth_b8_outmx[1]), .Y(n2434));
AND2X1 mul_U10574(.A(n5370), .B(n4848), .Y(dpath_mulcore_booth_b8_outmx[0]));
INVX1 mul_U10575(.A(dpath_mulcore_booth_b8_outmx[0]), .Y(n2435));
AND2X1 mul_U10576(.A(n5371), .B(n4849), .Y(dpath_mulcore_booth_b9_outmx[2]));
INVX1 mul_U10577(.A(dpath_mulcore_booth_b9_outmx[2]), .Y(n2436));
AND2X1 mul_U10578(.A(n5372), .B(n4850), .Y(dpath_mulcore_booth_b9_outmx[1]));
INVX1 mul_U10579(.A(dpath_mulcore_booth_b9_outmx[1]), .Y(n2437));
AND2X1 mul_U10580(.A(n5373), .B(n4851), .Y(dpath_mulcore_booth_b9_outmx[0]));
INVX1 mul_U10581(.A(dpath_mulcore_booth_b9_outmx[0]), .Y(n2438));
AND2X1 mul_U10582(.A(n5374), .B(n4852), .Y(dpath_mulcore_booth_b10_outmx[2]));
INVX1 mul_U10583(.A(dpath_mulcore_booth_b10_outmx[2]), .Y(n2439));
AND2X1 mul_U10584(.A(n5375), .B(n4853), .Y(dpath_mulcore_booth_b10_outmx[1]));
INVX1 mul_U10585(.A(dpath_mulcore_booth_b10_outmx[1]), .Y(n2440));
AND2X1 mul_U10586(.A(n5376), .B(n4854), .Y(dpath_mulcore_booth_b10_outmx[0]));
INVX1 mul_U10587(.A(dpath_mulcore_booth_b10_outmx[0]), .Y(n2441));
AND2X1 mul_U10588(.A(n5377), .B(n4855), .Y(dpath_mulcore_booth_b11_outmx[2]));
INVX1 mul_U10589(.A(dpath_mulcore_booth_b11_outmx[2]), .Y(n2442));
AND2X1 mul_U10590(.A(n5378), .B(n4856), .Y(dpath_mulcore_booth_b11_outmx[1]));
INVX1 mul_U10591(.A(dpath_mulcore_booth_b11_outmx[1]), .Y(n2443));
AND2X1 mul_U10592(.A(n5379), .B(n4857), .Y(dpath_mulcore_booth_b11_outmx[0]));
INVX1 mul_U10593(.A(dpath_mulcore_booth_b11_outmx[0]), .Y(n2444));
AND2X1 mul_U10594(.A(n5380), .B(n4858), .Y(dpath_mulcore_booth_b12_outmx[2]));
INVX1 mul_U10595(.A(dpath_mulcore_booth_b12_outmx[2]), .Y(n2445));
AND2X1 mul_U10596(.A(n5381), .B(n4859), .Y(dpath_mulcore_booth_b12_outmx[1]));
INVX1 mul_U10597(.A(dpath_mulcore_booth_b12_outmx[1]), .Y(n2446));
AND2X1 mul_U10598(.A(n5382), .B(n4860), .Y(dpath_mulcore_booth_b12_outmx[0]));
INVX1 mul_U10599(.A(dpath_mulcore_booth_b12_outmx[0]), .Y(n2447));
AND2X1 mul_U10600(.A(n5383), .B(n4861), .Y(dpath_mulcore_booth_b13_outmx[2]));
INVX1 mul_U10601(.A(dpath_mulcore_booth_b13_outmx[2]), .Y(n2448));
AND2X1 mul_U10602(.A(n5384), .B(n4862), .Y(dpath_mulcore_booth_b13_outmx[1]));
INVX1 mul_U10603(.A(dpath_mulcore_booth_b13_outmx[1]), .Y(n2449));
AND2X1 mul_U10604(.A(n5385), .B(n4863), .Y(dpath_mulcore_booth_b13_outmx[0]));
INVX1 mul_U10605(.A(dpath_mulcore_booth_b13_outmx[0]), .Y(n2450));
AND2X1 mul_U10606(.A(n5386), .B(n4864), .Y(dpath_mulcore_booth_b14_outmx[2]));
INVX1 mul_U10607(.A(dpath_mulcore_booth_b14_outmx[2]), .Y(n2451));
AND2X1 mul_U10608(.A(n5387), .B(n4865), .Y(dpath_mulcore_booth_b14_outmx[1]));
INVX1 mul_U10609(.A(dpath_mulcore_booth_b14_outmx[1]), .Y(n2452));
AND2X1 mul_U10610(.A(n5388), .B(n4866), .Y(dpath_mulcore_booth_b14_outmx[0]));
INVX1 mul_U10611(.A(dpath_mulcore_booth_b14_outmx[0]), .Y(n2453));
AND2X1 mul_U10612(.A(n6064), .B(n4867), .Y(dpath_mulcore_booth_b15_outmx[2]));
INVX1 mul_U10613(.A(dpath_mulcore_booth_b15_outmx[2]), .Y(n2454));
AND2X1 mul_U10614(.A(n5389), .B(n4868), .Y(dpath_mulcore_booth_b15_outmx[1]));
INVX1 mul_U10615(.A(dpath_mulcore_booth_b15_outmx[1]), .Y(n2455));
AND2X1 mul_U10616(.A(n5390), .B(n4869), .Y(dpath_mulcore_booth_b15_outmx[0]));
INVX1 mul_U10617(.A(dpath_mulcore_booth_b15_outmx[0]), .Y(n2456));
AND2X1 mul_U10618(.A(dpath_mulcore_booth_b13_in0[2]), .B(n9805), .Y(n17957));
INVX1 mul_U10619(.A(n17957), .Y(n2457));
AND2X1 mul_U10620(.A(dpath_mulcore_booth_b12_in0[2]), .B(n9803), .Y(n17961));
INVX1 mul_U10621(.A(n17961), .Y(n2458));
AND2X1 mul_U10622(.A(dpath_mulcore_booth_b11_in0[2]), .B(n9801), .Y(n17965));
INVX1 mul_U10623(.A(n17965), .Y(n2459));
AND2X1 mul_U10624(.A(dpath_mulcore_booth_b10_in0[2]), .B(n9799), .Y(n17969));
INVX1 mul_U10625(.A(n17969), .Y(n2460));
AND2X1 mul_U10626(.A(dpath_mulcore_booth_b9_in0[2]), .B(n9797), .Y(n17973));
INVX1 mul_U10627(.A(n17973), .Y(n2461));
AND2X1 mul_U10628(.A(dpath_mulcore_booth_b8_in0[2]), .B(n9794), .Y(n17977));
INVX1 mul_U10629(.A(n17977), .Y(n2462));
AND2X1 mul_U10630(.A(n18011), .B(n4870), .Y(dpath_mulcore_booth_b0_in1[1]));
INVX1 mul_U10631(.A(dpath_mulcore_booth_b0_in1[1]), .Y(n2463));
AND2X1 mul_U10632(.A(dpath_mulcore_booth_b5_in1[2]), .B(n10094), .Y(n18021));
INVX1 mul_U10633(.A(n18021), .Y(n2464));
AND2X1 mul_U10634(.A(dpath_mulcore_booth_b4_in1[2]), .B(n10092), .Y(n18025));
INVX1 mul_U10635(.A(n18025), .Y(n2465));
AND2X1 mul_U10636(.A(dpath_mulcore_booth_b3_in1[2]), .B(n10090), .Y(n18029));
INVX1 mul_U10637(.A(n18029), .Y(n2466));
AND2X1 mul_U10638(.A(dpath_mulcore_booth_b2_in1[2]), .B(n10088), .Y(n18033));
INVX1 mul_U10639(.A(n18033), .Y(n2467));
AND2X1 mul_U10640(.A(dpath_mulcore_booth_b1_in1[2]), .B(n10086), .Y(n18037));
INVX1 mul_U10641(.A(n18037), .Y(n2468));
AND2X1 mul_U10642(.A(dpath_mulcore_booth_b0_in1[2]), .B(n10084), .Y(n18041));
INVX1 mul_U10643(.A(n18041), .Y(n2469));
AND2X1 mul_U10644(.A(n5441), .B(n4871), .Y(dpath_mulcore_booth_b0_in1[0]));
INVX1 mul_U10645(.A(dpath_mulcore_booth_b0_in1[0]), .Y(n2470));
AND2X1 mul_U10646(.A(dpath_mulcore_booth_b13_in1[2]), .B(n10108), .Y(n18085));
INVX1 mul_U10647(.A(n18085), .Y(n2471));
AND2X1 mul_U10648(.A(dpath_mulcore_booth_b12_in1[2]), .B(n10106), .Y(n18089));
INVX1 mul_U10649(.A(n18089), .Y(n2472));
AND2X1 mul_U10650(.A(dpath_mulcore_booth_b11_in1[2]), .B(n10104), .Y(n18093));
INVX1 mul_U10651(.A(n18093), .Y(n2473));
AND2X1 mul_U10652(.A(dpath_mulcore_booth_b10_in1[2]), .B(n10102), .Y(n18097));
INVX1 mul_U10653(.A(n18097), .Y(n2474));
AND2X1 mul_U10654(.A(dpath_mulcore_booth_b9_in1[2]), .B(n10100), .Y(n18101));
INVX1 mul_U10655(.A(n18101), .Y(n2475));
AND2X1 mul_U10656(.A(dpath_mulcore_booth_b8_in1[2]), .B(n10098), .Y(n18105));
INVX1 mul_U10657(.A(n18105), .Y(n2476));
AND2X1 mul_U10658(.A(dpath_mulcore_ary1_a0_I2_p0_l[63]), .B(dpath_mulcore_b6[0]), .Y(dpath_mulcore_ary1_a0_I2_I2_p0_64__n2));
INVX1 mul_U10659(.A(dpath_mulcore_ary1_a0_I2_I2_p0_64__n2), .Y(n2477));
AND2X1 mul_U10660(.A(n9683), .B(n6088), .Y(dpath_mulcore_array2_sh_82__n2));
INVX1 mul_U10661(.A(dpath_mulcore_array2_sh_82__n2), .Y(n2478));
AND2X1 mul_U10662(.A(n13754), .B(n13755), .Y(dpath_mulcore_ary1_a0_sc2_2_70__n2));
INVX1 mul_U10663(.A(dpath_mulcore_ary1_a0_sc2_2_70__n2), .Y(n2479));
AND2X1 mul_U10664(.A(dpath_mulcore_ary1_a0_s_2[71]), .B(dpath_mulcore_ary1_a0_s1[64]), .Y(dpath_mulcore_ary1_a0_sc3_71__n2));
INVX1 mul_U10665(.A(dpath_mulcore_ary1_a0_sc3_71__n2), .Y(n2480));
AND2X1 mul_U10666(.A(n5470), .B(n4872), .Y(dpath_mulcore_a0cout[71]));
INVX1 mul_U10667(.A(dpath_mulcore_a0cout[71]), .Y(n2481));
AND2X1 mul_U10668(.A(n5471), .B(n4873), .Y(dpath_mulcore_booth_b0_outmx[2]));
INVX1 mul_U10669(.A(dpath_mulcore_booth_b0_outmx[2]), .Y(n2482));
AND2X1 mul_U10670(.A(n5472), .B(n4874), .Y(dpath_mulcore_booth_b0_outmx[1]));
INVX1 mul_U10671(.A(dpath_mulcore_booth_b0_outmx[1]), .Y(n2483));
AND2X1 mul_U10672(.A(n5473), .B(n4875), .Y(dpath_mulcore_booth_b0_outmx[0]));
INVX1 mul_U10673(.A(dpath_mulcore_booth_b0_outmx[0]), .Y(n2484));
AND2X1 mul_U10674(.A(dpath_mulcore_booth_b5_in0[2]), .B(n9790), .Y(dpath_mulcore_booth_encode0_a_n25));
INVX1 mul_U10675(.A(dpath_mulcore_booth_encode0_a_n25), .Y(n2485));
AND2X1 mul_U10676(.A(dpath_mulcore_booth_b4_in0[2]), .B(n9788), .Y(dpath_mulcore_booth_encode0_a_n29));
INVX1 mul_U10677(.A(dpath_mulcore_booth_encode0_a_n29), .Y(n2486));
AND2X1 mul_U10678(.A(dpath_mulcore_booth_b3_in0[2]), .B(n9813), .Y(dpath_mulcore_booth_encode0_a_n33));
INVX1 mul_U10679(.A(dpath_mulcore_booth_encode0_a_n33), .Y(n2487));
AND2X1 mul_U10680(.A(dpath_mulcore_booth_b2_in0[2]), .B(n9811), .Y(dpath_mulcore_booth_encode0_a_n37));
INVX1 mul_U10681(.A(dpath_mulcore_booth_encode0_a_n37), .Y(n2488));
AND2X1 mul_U10682(.A(dpath_mulcore_booth_b1_in0[2]), .B(n9809), .Y(dpath_mulcore_booth_encode0_a_n41));
INVX1 mul_U10683(.A(dpath_mulcore_booth_encode0_a_n41), .Y(n2489));
AND2X1 mul_U10684(.A(dpath_mulcore_booth_b0_in0[2]), .B(n9807), .Y(dpath_mulcore_booth_encode0_a_n45));
INVX1 mul_U10685(.A(dpath_mulcore_booth_encode0_a_n45), .Y(n2490));
AND2X1 mul_U10686(.A(n5498), .B(n4876), .Y(dpath_mulcore_ary2_sum[9]));
INVX1 mul_U10687(.A(dpath_mulcore_ary2_sum[9]), .Y(n2491));
AND2X1 mul_U10688(.A(n5499), .B(n4877), .Y(dpath_mulcore_ary2_sum[97]));
INVX1 mul_U10689(.A(dpath_mulcore_ary2_sum[97]), .Y(n2492));
AND2X1 mul_U10690(.A(n5500), .B(n4878), .Y(dpath_mulcore_ary2_sum[96]));
INVX1 mul_U10691(.A(dpath_mulcore_ary2_sum[96]), .Y(n2493));
AND2X1 mul_U10692(.A(n5501), .B(n4879), .Y(dpath_mulcore_ary2_sum[95]));
INVX1 mul_U10693(.A(dpath_mulcore_ary2_sum[95]), .Y(n2494));
AND2X1 mul_U10694(.A(n5502), .B(n4880), .Y(dpath_mulcore_ary2_sum[94]));
INVX1 mul_U10695(.A(dpath_mulcore_ary2_sum[94]), .Y(n2495));
AND2X1 mul_U10696(.A(n5503), .B(n4881), .Y(dpath_mulcore_ary2_sum[93]));
INVX1 mul_U10697(.A(dpath_mulcore_ary2_sum[93]), .Y(n2496));
AND2X1 mul_U10698(.A(n5504), .B(n4882), .Y(dpath_mulcore_ary2_sum[92]));
INVX1 mul_U10699(.A(dpath_mulcore_ary2_sum[92]), .Y(n2497));
AND2X1 mul_U10700(.A(n5505), .B(n4883), .Y(dpath_mulcore_ary2_sum[91]));
INVX1 mul_U10701(.A(dpath_mulcore_ary2_sum[91]), .Y(n2498));
AND2X1 mul_U10702(.A(n5506), .B(n4884), .Y(dpath_mulcore_ary2_sum[90]));
INVX1 mul_U10703(.A(dpath_mulcore_ary2_sum[90]), .Y(n2499));
AND2X1 mul_U10704(.A(n5507), .B(n4885), .Y(dpath_mulcore_ary2_sum[8]));
INVX1 mul_U10705(.A(dpath_mulcore_ary2_sum[8]), .Y(n2500));
AND2X1 mul_U10706(.A(n5508), .B(n4886), .Y(dpath_mulcore_ary2_sum[89]));
INVX1 mul_U10707(.A(dpath_mulcore_ary2_sum[89]), .Y(n2501));
AND2X1 mul_U10708(.A(n5509), .B(n4887), .Y(dpath_mulcore_ary2_sum[88]));
INVX1 mul_U10709(.A(dpath_mulcore_ary2_sum[88]), .Y(n2502));
AND2X1 mul_U10710(.A(n5510), .B(n4888), .Y(dpath_mulcore_ary2_sum[87]));
INVX1 mul_U10711(.A(dpath_mulcore_ary2_sum[87]), .Y(n2503));
AND2X1 mul_U10712(.A(n5511), .B(n4889), .Y(dpath_mulcore_ary2_sum[86]));
INVX1 mul_U10713(.A(dpath_mulcore_ary2_sum[86]), .Y(n2504));
AND2X1 mul_U10714(.A(n5512), .B(n4890), .Y(dpath_mulcore_ary2_sum[85]));
INVX1 mul_U10715(.A(dpath_mulcore_ary2_sum[85]), .Y(n2505));
AND2X1 mul_U10716(.A(n5513), .B(n4891), .Y(dpath_mulcore_ary2_sum[84]));
INVX1 mul_U10717(.A(dpath_mulcore_ary2_sum[84]), .Y(n2506));
AND2X1 mul_U10718(.A(n5514), .B(n4892), .Y(dpath_mulcore_ary2_sum[83]));
INVX1 mul_U10719(.A(dpath_mulcore_ary2_sum[83]), .Y(n2507));
AND2X1 mul_U10720(.A(n5515), .B(n4893), .Y(dpath_mulcore_ary2_sum[82]));
INVX1 mul_U10721(.A(dpath_mulcore_ary2_sum[82]), .Y(n2508));
AND2X1 mul_U10722(.A(n5516), .B(n4894), .Y(dpath_mulcore_ary2_sum[81]));
INVX1 mul_U10723(.A(dpath_mulcore_ary2_sum[81]), .Y(n2509));
AND2X1 mul_U10724(.A(n5517), .B(n4895), .Y(dpath_mulcore_ary2_sum[80]));
INVX1 mul_U10725(.A(dpath_mulcore_ary2_sum[80]), .Y(n2510));
AND2X1 mul_U10726(.A(n5518), .B(n4896), .Y(dpath_mulcore_ary2_sum[7]));
INVX1 mul_U10727(.A(dpath_mulcore_ary2_sum[7]), .Y(n2511));
AND2X1 mul_U10728(.A(n5519), .B(n4897), .Y(dpath_mulcore_ary2_sum[79]));
INVX1 mul_U10729(.A(dpath_mulcore_ary2_sum[79]), .Y(n2512));
AND2X1 mul_U10730(.A(n5520), .B(n4898), .Y(dpath_mulcore_ary2_sum[78]));
INVX1 mul_U10731(.A(dpath_mulcore_ary2_sum[78]), .Y(n2513));
AND2X1 mul_U10732(.A(n5521), .B(n4899), .Y(dpath_mulcore_ary2_sum[77]));
INVX1 mul_U10733(.A(dpath_mulcore_ary2_sum[77]), .Y(n2514));
AND2X1 mul_U10734(.A(n5522), .B(n4900), .Y(dpath_mulcore_ary2_sum[76]));
INVX1 mul_U10735(.A(dpath_mulcore_ary2_sum[76]), .Y(n2515));
AND2X1 mul_U10736(.A(n5523), .B(n4901), .Y(dpath_mulcore_ary2_sum[75]));
INVX1 mul_U10737(.A(dpath_mulcore_ary2_sum[75]), .Y(n2516));
AND2X1 mul_U10738(.A(n5524), .B(n4902), .Y(dpath_mulcore_ary2_sum[74]));
INVX1 mul_U10739(.A(dpath_mulcore_ary2_sum[74]), .Y(n2517));
AND2X1 mul_U10740(.A(n5525), .B(n4903), .Y(dpath_mulcore_ary2_sum[73]));
INVX1 mul_U10741(.A(dpath_mulcore_ary2_sum[73]), .Y(n2518));
AND2X1 mul_U10742(.A(n5526), .B(n4904), .Y(dpath_mulcore_ary2_sum[72]));
INVX1 mul_U10743(.A(dpath_mulcore_ary2_sum[72]), .Y(n2519));
AND2X1 mul_U10744(.A(n5527), .B(n4905), .Y(dpath_mulcore_ary2_sum[71]));
INVX1 mul_U10745(.A(dpath_mulcore_ary2_sum[71]), .Y(n2520));
AND2X1 mul_U10746(.A(n5528), .B(n4906), .Y(dpath_mulcore_ary2_sum[70]));
INVX1 mul_U10747(.A(dpath_mulcore_ary2_sum[70]), .Y(n2521));
AND2X1 mul_U10748(.A(n5529), .B(n4907), .Y(dpath_mulcore_ary2_sum[6]));
INVX1 mul_U10749(.A(dpath_mulcore_ary2_sum[6]), .Y(n2522));
AND2X1 mul_U10750(.A(n5530), .B(n4908), .Y(dpath_mulcore_ary2_sum[69]));
INVX1 mul_U10751(.A(dpath_mulcore_ary2_sum[69]), .Y(n2523));
AND2X1 mul_U10752(.A(n5531), .B(n4909), .Y(dpath_mulcore_ary2_sum[68]));
INVX1 mul_U10753(.A(dpath_mulcore_ary2_sum[68]), .Y(n2524));
AND2X1 mul_U10754(.A(n5532), .B(n4910), .Y(dpath_mulcore_ary2_sum[67]));
INVX1 mul_U10755(.A(dpath_mulcore_ary2_sum[67]), .Y(n2525));
AND2X1 mul_U10756(.A(n5533), .B(n4911), .Y(dpath_mulcore_ary2_sum[66]));
INVX1 mul_U10757(.A(dpath_mulcore_ary2_sum[66]), .Y(n2526));
AND2X1 mul_U10758(.A(n5534), .B(n4912), .Y(dpath_mulcore_ary2_sum[65]));
INVX1 mul_U10759(.A(dpath_mulcore_ary2_sum[65]), .Y(n2527));
AND2X1 mul_U10760(.A(n5535), .B(n4913), .Y(dpath_mulcore_ary2_sum[64]));
INVX1 mul_U10761(.A(dpath_mulcore_ary2_sum[64]), .Y(n2528));
AND2X1 mul_U10762(.A(n5536), .B(n4914), .Y(dpath_mulcore_ary2_sum[63]));
INVX1 mul_U10763(.A(dpath_mulcore_ary2_sum[63]), .Y(n2529));
AND2X1 mul_U10764(.A(n5537), .B(n4915), .Y(dpath_mulcore_ary2_sum[62]));
INVX1 mul_U10765(.A(dpath_mulcore_ary2_sum[62]), .Y(n2530));
AND2X1 mul_U10766(.A(n5538), .B(n4916), .Y(dpath_mulcore_ary2_sum[61]));
INVX1 mul_U10767(.A(dpath_mulcore_ary2_sum[61]), .Y(n2531));
AND2X1 mul_U10768(.A(n5539), .B(n4917), .Y(dpath_mulcore_ary2_sum[60]));
INVX1 mul_U10769(.A(dpath_mulcore_ary2_sum[60]), .Y(n2532));
AND2X1 mul_U10770(.A(n5540), .B(n4918), .Y(dpath_mulcore_ary2_sum[5]));
INVX1 mul_U10771(.A(dpath_mulcore_ary2_sum[5]), .Y(n2533));
AND2X1 mul_U10772(.A(n5541), .B(n4919), .Y(dpath_mulcore_ary2_sum[59]));
INVX1 mul_U10773(.A(dpath_mulcore_ary2_sum[59]), .Y(n2534));
AND2X1 mul_U10774(.A(n5542), .B(n4920), .Y(dpath_mulcore_ary2_sum[58]));
INVX1 mul_U10775(.A(dpath_mulcore_ary2_sum[58]), .Y(n2535));
AND2X1 mul_U10776(.A(n5543), .B(n4921), .Y(dpath_mulcore_ary2_sum[57]));
INVX1 mul_U10777(.A(dpath_mulcore_ary2_sum[57]), .Y(n2536));
AND2X1 mul_U10778(.A(n5544), .B(n4922), .Y(dpath_mulcore_ary2_sum[56]));
INVX1 mul_U10779(.A(dpath_mulcore_ary2_sum[56]), .Y(n2537));
AND2X1 mul_U10780(.A(n5545), .B(n4923), .Y(dpath_mulcore_ary2_sum[55]));
INVX1 mul_U10781(.A(dpath_mulcore_ary2_sum[55]), .Y(n2538));
AND2X1 mul_U10782(.A(n5546), .B(n4924), .Y(dpath_mulcore_ary2_sum[54]));
INVX1 mul_U10783(.A(dpath_mulcore_ary2_sum[54]), .Y(n2539));
AND2X1 mul_U10784(.A(n5547), .B(n4925), .Y(dpath_mulcore_ary2_sum[53]));
INVX1 mul_U10785(.A(dpath_mulcore_ary2_sum[53]), .Y(n2540));
AND2X1 mul_U10786(.A(n5548), .B(n4926), .Y(dpath_mulcore_ary2_sum[52]));
INVX1 mul_U10787(.A(dpath_mulcore_ary2_sum[52]), .Y(n2541));
AND2X1 mul_U10788(.A(n5549), .B(n4927), .Y(dpath_mulcore_ary2_sum[51]));
INVX1 mul_U10789(.A(dpath_mulcore_ary2_sum[51]), .Y(n2542));
AND2X1 mul_U10790(.A(n5550), .B(n4928), .Y(dpath_mulcore_ary2_sum[50]));
INVX1 mul_U10791(.A(dpath_mulcore_ary2_sum[50]), .Y(n2543));
AND2X1 mul_U10792(.A(n5551), .B(n4929), .Y(dpath_mulcore_ary2_sum[4]));
INVX1 mul_U10793(.A(dpath_mulcore_ary2_sum[4]), .Y(n2544));
AND2X1 mul_U10794(.A(n5552), .B(n4930), .Y(dpath_mulcore_ary2_sum[49]));
INVX1 mul_U10795(.A(dpath_mulcore_ary2_sum[49]), .Y(n2545));
AND2X1 mul_U10796(.A(n5553), .B(n4931), .Y(dpath_mulcore_ary2_sum[48]));
INVX1 mul_U10797(.A(dpath_mulcore_ary2_sum[48]), .Y(n2546));
AND2X1 mul_U10798(.A(n5554), .B(n4932), .Y(dpath_mulcore_ary2_sum[47]));
INVX1 mul_U10799(.A(dpath_mulcore_ary2_sum[47]), .Y(n2547));
AND2X1 mul_U10800(.A(n5555), .B(n4933), .Y(dpath_mulcore_ary2_sum[46]));
INVX1 mul_U10801(.A(dpath_mulcore_ary2_sum[46]), .Y(n2548));
AND2X1 mul_U10802(.A(n5556), .B(n4934), .Y(dpath_mulcore_ary2_sum[45]));
INVX1 mul_U10803(.A(dpath_mulcore_ary2_sum[45]), .Y(n2549));
AND2X1 mul_U10804(.A(n5557), .B(n4935), .Y(dpath_mulcore_ary2_sum[44]));
INVX1 mul_U10805(.A(dpath_mulcore_ary2_sum[44]), .Y(n2550));
AND2X1 mul_U10806(.A(n5558), .B(n4936), .Y(dpath_mulcore_ary2_sum[43]));
INVX1 mul_U10807(.A(dpath_mulcore_ary2_sum[43]), .Y(n2551));
AND2X1 mul_U10808(.A(n5559), .B(n4937), .Y(dpath_mulcore_ary2_sum[42]));
INVX1 mul_U10809(.A(dpath_mulcore_ary2_sum[42]), .Y(n2552));
AND2X1 mul_U10810(.A(n5560), .B(n4938), .Y(dpath_mulcore_ary2_sum[41]));
INVX1 mul_U10811(.A(dpath_mulcore_ary2_sum[41]), .Y(n2553));
AND2X1 mul_U10812(.A(n5561), .B(n4939), .Y(dpath_mulcore_ary2_sum[40]));
INVX1 mul_U10813(.A(dpath_mulcore_ary2_sum[40]), .Y(n2554));
AND2X1 mul_U10814(.A(n5562), .B(n4940), .Y(dpath_mulcore_ary2_sum[3]));
INVX1 mul_U10815(.A(dpath_mulcore_ary2_sum[3]), .Y(n2555));
AND2X1 mul_U10816(.A(n5563), .B(n4941), .Y(dpath_mulcore_ary2_sum[39]));
INVX1 mul_U10817(.A(dpath_mulcore_ary2_sum[39]), .Y(n2556));
AND2X1 mul_U10818(.A(n5564), .B(n4942), .Y(dpath_mulcore_ary2_sum[38]));
INVX1 mul_U10819(.A(dpath_mulcore_ary2_sum[38]), .Y(n2557));
AND2X1 mul_U10820(.A(n5565), .B(n4943), .Y(dpath_mulcore_ary2_sum[37]));
INVX1 mul_U10821(.A(dpath_mulcore_ary2_sum[37]), .Y(n2558));
AND2X1 mul_U10822(.A(n5566), .B(n4944), .Y(dpath_mulcore_ary2_sum[36]));
INVX1 mul_U10823(.A(dpath_mulcore_ary2_sum[36]), .Y(n2559));
AND2X1 mul_U10824(.A(n5567), .B(n4945), .Y(dpath_mulcore_ary2_sum[35]));
INVX1 mul_U10825(.A(dpath_mulcore_ary2_sum[35]), .Y(n2560));
AND2X1 mul_U10826(.A(n5568), .B(n4946), .Y(dpath_mulcore_ary2_sum[34]));
INVX1 mul_U10827(.A(dpath_mulcore_ary2_sum[34]), .Y(n2561));
AND2X1 mul_U10828(.A(n5569), .B(n4947), .Y(dpath_mulcore_ary2_sum[33]));
INVX1 mul_U10829(.A(dpath_mulcore_ary2_sum[33]), .Y(n2562));
AND2X1 mul_U10830(.A(n5570), .B(n4948), .Y(dpath_mulcore_ary2_sum[32]));
INVX1 mul_U10831(.A(dpath_mulcore_ary2_sum[32]), .Y(n2563));
AND2X1 mul_U10832(.A(n5571), .B(n4949), .Y(dpath_mulcore_ary2_sum[31]));
INVX1 mul_U10833(.A(dpath_mulcore_ary2_sum[31]), .Y(n2564));
AND2X1 mul_U10834(.A(n5572), .B(n4950), .Y(dpath_mulcore_ary2_sum[30]));
INVX1 mul_U10835(.A(dpath_mulcore_ary2_sum[30]), .Y(n2565));
AND2X1 mul_U10836(.A(n5573), .B(n4951), .Y(dpath_mulcore_ary2_sum[2]));
INVX1 mul_U10837(.A(dpath_mulcore_ary2_sum[2]), .Y(n2566));
AND2X1 mul_U10838(.A(n5574), .B(n4952), .Y(dpath_mulcore_ary2_sum[29]));
INVX1 mul_U10839(.A(dpath_mulcore_ary2_sum[29]), .Y(n2567));
AND2X1 mul_U10840(.A(n5575), .B(n4953), .Y(dpath_mulcore_ary2_sum[28]));
INVX1 mul_U10841(.A(dpath_mulcore_ary2_sum[28]), .Y(n2568));
AND2X1 mul_U10842(.A(n5576), .B(n4954), .Y(dpath_mulcore_ary2_sum[27]));
INVX1 mul_U10843(.A(dpath_mulcore_ary2_sum[27]), .Y(n2569));
AND2X1 mul_U10844(.A(n5577), .B(n4955), .Y(dpath_mulcore_ary2_sum[26]));
INVX1 mul_U10845(.A(dpath_mulcore_ary2_sum[26]), .Y(n2570));
AND2X1 mul_U10846(.A(n5578), .B(n4956), .Y(dpath_mulcore_ary2_sum[25]));
INVX1 mul_U10847(.A(dpath_mulcore_ary2_sum[25]), .Y(n2571));
AND2X1 mul_U10848(.A(n5579), .B(n4957), .Y(dpath_mulcore_ary2_sum[24]));
INVX1 mul_U10849(.A(dpath_mulcore_ary2_sum[24]), .Y(n2572));
AND2X1 mul_U10850(.A(n5580), .B(n4958), .Y(dpath_mulcore_ary2_sum[23]));
INVX1 mul_U10851(.A(dpath_mulcore_ary2_sum[23]), .Y(n2573));
AND2X1 mul_U10852(.A(n5581), .B(n4959), .Y(dpath_mulcore_ary2_sum[22]));
INVX1 mul_U10853(.A(dpath_mulcore_ary2_sum[22]), .Y(n2574));
AND2X1 mul_U10854(.A(n5582), .B(n4960), .Y(dpath_mulcore_ary2_sum[21]));
INVX1 mul_U10855(.A(dpath_mulcore_ary2_sum[21]), .Y(n2575));
AND2X1 mul_U10856(.A(n5583), .B(n4961), .Y(dpath_mulcore_ary2_sum[20]));
INVX1 mul_U10857(.A(dpath_mulcore_ary2_sum[20]), .Y(n2576));
AND2X1 mul_U10858(.A(n5584), .B(n4962), .Y(dpath_mulcore_ary2_sum[1]));
INVX1 mul_U10859(.A(dpath_mulcore_ary2_sum[1]), .Y(n2577));
AND2X1 mul_U10860(.A(n5585), .B(n4963), .Y(dpath_mulcore_ary2_sum[19]));
INVX1 mul_U10861(.A(dpath_mulcore_ary2_sum[19]), .Y(n2578));
AND2X1 mul_U10862(.A(n5586), .B(n4964), .Y(dpath_mulcore_ary2_sum[18]));
INVX1 mul_U10863(.A(dpath_mulcore_ary2_sum[18]), .Y(n2579));
AND2X1 mul_U10864(.A(n5587), .B(n4965), .Y(dpath_mulcore_ary2_sum[17]));
INVX1 mul_U10865(.A(dpath_mulcore_ary2_sum[17]), .Y(n2580));
AND2X1 mul_U10866(.A(n5588), .B(n4966), .Y(dpath_mulcore_ary2_sum[16]));
INVX1 mul_U10867(.A(dpath_mulcore_ary2_sum[16]), .Y(n2581));
AND2X1 mul_U10868(.A(n5589), .B(n4967), .Y(dpath_mulcore_ary2_sum[15]));
INVX1 mul_U10869(.A(dpath_mulcore_ary2_sum[15]), .Y(n2582));
AND2X1 mul_U10870(.A(n5590), .B(n4968), .Y(dpath_mulcore_ary2_sum[14]));
INVX1 mul_U10871(.A(dpath_mulcore_ary2_sum[14]), .Y(n2583));
AND2X1 mul_U10872(.A(n5591), .B(n4969), .Y(dpath_mulcore_ary2_sum[13]));
INVX1 mul_U10873(.A(dpath_mulcore_ary2_sum[13]), .Y(n2584));
AND2X1 mul_U10874(.A(n5592), .B(n4970), .Y(dpath_mulcore_ary2_sum[12]));
INVX1 mul_U10875(.A(dpath_mulcore_ary2_sum[12]), .Y(n2585));
AND2X1 mul_U10876(.A(n5593), .B(n4971), .Y(dpath_mulcore_ary2_sum[11]));
INVX1 mul_U10877(.A(dpath_mulcore_ary2_sum[11]), .Y(n2586));
AND2X1 mul_U10878(.A(n5594), .B(n4972), .Y(dpath_mulcore_ary2_sum[10]));
INVX1 mul_U10879(.A(dpath_mulcore_ary2_sum[10]), .Y(n2587));
AND2X1 mul_U10880(.A(n5595), .B(n4973), .Y(dpath_mulcore_ary2_sum[0]));
INVX1 mul_U10881(.A(dpath_mulcore_ary2_sum[0]), .Y(n2588));
AND2X1 mul_U10882(.A(n5596), .B(n4974), .Y(dpath_mulcore_ary2_cout[9]));
INVX1 mul_U10883(.A(dpath_mulcore_ary2_cout[9]), .Y(n2589));
AND2X1 mul_U10884(.A(n5597), .B(n4975), .Y(dpath_mulcore_ary2_cout[96]));
INVX1 mul_U10885(.A(dpath_mulcore_ary2_cout[96]), .Y(n2590));
AND2X1 mul_U10886(.A(n5598), .B(n4976), .Y(dpath_mulcore_ary2_cout[95]));
INVX1 mul_U10887(.A(dpath_mulcore_ary2_cout[95]), .Y(n2591));
AND2X1 mul_U10888(.A(n5599), .B(n4977), .Y(dpath_mulcore_ary2_cout[94]));
INVX1 mul_U10889(.A(dpath_mulcore_ary2_cout[94]), .Y(n2592));
AND2X1 mul_U10890(.A(n5600), .B(n4978), .Y(dpath_mulcore_ary2_cout[93]));
INVX1 mul_U10891(.A(dpath_mulcore_ary2_cout[93]), .Y(n2593));
AND2X1 mul_U10892(.A(n5601), .B(n4979), .Y(dpath_mulcore_ary2_cout[92]));
INVX1 mul_U10893(.A(dpath_mulcore_ary2_cout[92]), .Y(n2594));
AND2X1 mul_U10894(.A(n5602), .B(n4980), .Y(dpath_mulcore_ary2_cout[91]));
INVX1 mul_U10895(.A(dpath_mulcore_ary2_cout[91]), .Y(n2595));
AND2X1 mul_U10896(.A(n5603), .B(n4981), .Y(dpath_mulcore_ary2_cout[90]));
INVX1 mul_U10897(.A(dpath_mulcore_ary2_cout[90]), .Y(n2596));
AND2X1 mul_U10898(.A(n5604), .B(n4982), .Y(dpath_mulcore_ary2_cout[8]));
INVX1 mul_U10899(.A(dpath_mulcore_ary2_cout[8]), .Y(n2597));
AND2X1 mul_U10900(.A(n5605), .B(n4983), .Y(dpath_mulcore_ary2_cout[89]));
INVX1 mul_U10901(.A(dpath_mulcore_ary2_cout[89]), .Y(n2598));
AND2X1 mul_U10902(.A(n5606), .B(n4984), .Y(dpath_mulcore_ary2_cout[88]));
INVX1 mul_U10903(.A(dpath_mulcore_ary2_cout[88]), .Y(n2599));
AND2X1 mul_U10904(.A(n5607), .B(n4985), .Y(dpath_mulcore_ary2_cout[87]));
INVX1 mul_U10905(.A(dpath_mulcore_ary2_cout[87]), .Y(n2600));
AND2X1 mul_U10906(.A(n5608), .B(n4986), .Y(dpath_mulcore_ary2_cout[86]));
INVX1 mul_U10907(.A(dpath_mulcore_ary2_cout[86]), .Y(n2601));
AND2X1 mul_U10908(.A(n5609), .B(n4987), .Y(dpath_mulcore_ary2_cout[85]));
INVX1 mul_U10909(.A(dpath_mulcore_ary2_cout[85]), .Y(n2602));
AND2X1 mul_U10910(.A(n5610), .B(n4988), .Y(dpath_mulcore_ary2_cout[84]));
INVX1 mul_U10911(.A(dpath_mulcore_ary2_cout[84]), .Y(n2603));
AND2X1 mul_U10912(.A(n5611), .B(n4989), .Y(dpath_mulcore_ary2_cout[83]));
INVX1 mul_U10913(.A(dpath_mulcore_ary2_cout[83]), .Y(n2604));
AND2X1 mul_U10914(.A(n5612), .B(n4990), .Y(dpath_mulcore_ary2_cout[82]));
INVX1 mul_U10915(.A(dpath_mulcore_ary2_cout[82]), .Y(n2605));
AND2X1 mul_U10916(.A(n5613), .B(n4991), .Y(dpath_mulcore_ary2_cout[81]));
INVX1 mul_U10917(.A(dpath_mulcore_ary2_cout[81]), .Y(n2606));
AND2X1 mul_U10918(.A(n5614), .B(n4992), .Y(dpath_mulcore_ary2_cout[80]));
INVX1 mul_U10919(.A(dpath_mulcore_ary2_cout[80]), .Y(n2607));
AND2X1 mul_U10920(.A(n5615), .B(n4993), .Y(dpath_mulcore_ary2_cout[7]));
INVX1 mul_U10921(.A(dpath_mulcore_ary2_cout[7]), .Y(n2608));
AND2X1 mul_U10922(.A(n5616), .B(n4994), .Y(dpath_mulcore_ary2_cout[79]));
INVX1 mul_U10923(.A(dpath_mulcore_ary2_cout[79]), .Y(n2609));
AND2X1 mul_U10924(.A(n5617), .B(n4995), .Y(dpath_mulcore_ary2_cout[78]));
INVX1 mul_U10925(.A(dpath_mulcore_ary2_cout[78]), .Y(n2610));
AND2X1 mul_U10926(.A(n5618), .B(n4996), .Y(dpath_mulcore_ary2_cout[77]));
INVX1 mul_U10927(.A(dpath_mulcore_ary2_cout[77]), .Y(n2611));
AND2X1 mul_U10928(.A(n5619), .B(n4997), .Y(dpath_mulcore_ary2_cout[76]));
INVX1 mul_U10929(.A(dpath_mulcore_ary2_cout[76]), .Y(n2612));
AND2X1 mul_U10930(.A(n5620), .B(n4998), .Y(dpath_mulcore_ary2_cout[75]));
INVX1 mul_U10931(.A(dpath_mulcore_ary2_cout[75]), .Y(n2613));
AND2X1 mul_U10932(.A(n5621), .B(n4999), .Y(dpath_mulcore_ary2_cout[74]));
INVX1 mul_U10933(.A(dpath_mulcore_ary2_cout[74]), .Y(n2614));
AND2X1 mul_U10934(.A(n5622), .B(n5000), .Y(dpath_mulcore_ary2_cout[73]));
INVX1 mul_U10935(.A(dpath_mulcore_ary2_cout[73]), .Y(n2615));
AND2X1 mul_U10936(.A(n5623), .B(n5001), .Y(dpath_mulcore_ary2_cout[72]));
INVX1 mul_U10937(.A(dpath_mulcore_ary2_cout[72]), .Y(n2616));
AND2X1 mul_U10938(.A(n5624), .B(n5002), .Y(dpath_mulcore_ary2_cout[71]));
INVX1 mul_U10939(.A(dpath_mulcore_ary2_cout[71]), .Y(n2617));
AND2X1 mul_U10940(.A(n5625), .B(n5003), .Y(dpath_mulcore_ary2_cout[70]));
INVX1 mul_U10941(.A(dpath_mulcore_ary2_cout[70]), .Y(n2618));
AND2X1 mul_U10942(.A(n5626), .B(n5004), .Y(dpath_mulcore_ary2_cout[6]));
INVX1 mul_U10943(.A(dpath_mulcore_ary2_cout[6]), .Y(n2619));
AND2X1 mul_U10944(.A(n5627), .B(n5005), .Y(dpath_mulcore_ary2_cout[69]));
INVX1 mul_U10945(.A(dpath_mulcore_ary2_cout[69]), .Y(n2620));
AND2X1 mul_U10946(.A(n5628), .B(n5006), .Y(dpath_mulcore_ary2_cout[68]));
INVX1 mul_U10947(.A(dpath_mulcore_ary2_cout[68]), .Y(n2621));
AND2X1 mul_U10948(.A(n5629), .B(n5007), .Y(dpath_mulcore_ary2_cout[67]));
INVX1 mul_U10949(.A(dpath_mulcore_ary2_cout[67]), .Y(n2622));
AND2X1 mul_U10950(.A(n5630), .B(n5008), .Y(dpath_mulcore_ary2_cout[66]));
INVX1 mul_U10951(.A(dpath_mulcore_ary2_cout[66]), .Y(n2623));
AND2X1 mul_U10952(.A(n5631), .B(n5009), .Y(dpath_mulcore_ary2_cout[65]));
INVX1 mul_U10953(.A(dpath_mulcore_ary2_cout[65]), .Y(n2624));
AND2X1 mul_U10954(.A(n5632), .B(n5010), .Y(dpath_mulcore_ary2_cout[64]));
INVX1 mul_U10955(.A(dpath_mulcore_ary2_cout[64]), .Y(n2625));
AND2X1 mul_U10956(.A(n5633), .B(n5011), .Y(dpath_mulcore_ary2_cout[63]));
INVX1 mul_U10957(.A(dpath_mulcore_ary2_cout[63]), .Y(n2626));
AND2X1 mul_U10958(.A(n5634), .B(n5012), .Y(dpath_mulcore_ary2_cout[62]));
INVX1 mul_U10959(.A(dpath_mulcore_ary2_cout[62]), .Y(n2627));
AND2X1 mul_U10960(.A(n5635), .B(n5013), .Y(dpath_mulcore_ary2_cout[61]));
INVX1 mul_U10961(.A(dpath_mulcore_ary2_cout[61]), .Y(n2628));
AND2X1 mul_U10962(.A(n5636), .B(n5014), .Y(dpath_mulcore_ary2_cout[60]));
INVX1 mul_U10963(.A(dpath_mulcore_ary2_cout[60]), .Y(n2629));
AND2X1 mul_U10964(.A(n5637), .B(n5015), .Y(dpath_mulcore_ary2_cout[5]));
INVX1 mul_U10965(.A(dpath_mulcore_ary2_cout[5]), .Y(n2630));
AND2X1 mul_U10966(.A(n5638), .B(n5016), .Y(dpath_mulcore_ary2_cout[59]));
INVX1 mul_U10967(.A(dpath_mulcore_ary2_cout[59]), .Y(n2631));
AND2X1 mul_U10968(.A(n5639), .B(n5017), .Y(dpath_mulcore_ary2_cout[58]));
INVX1 mul_U10969(.A(dpath_mulcore_ary2_cout[58]), .Y(n2632));
AND2X1 mul_U10970(.A(n5640), .B(n5018), .Y(dpath_mulcore_ary2_cout[57]));
INVX1 mul_U10971(.A(dpath_mulcore_ary2_cout[57]), .Y(n2633));
AND2X1 mul_U10972(.A(n5641), .B(n5019), .Y(dpath_mulcore_ary2_cout[56]));
INVX1 mul_U10973(.A(dpath_mulcore_ary2_cout[56]), .Y(n2634));
AND2X1 mul_U10974(.A(n5642), .B(n5020), .Y(dpath_mulcore_ary2_cout[55]));
INVX1 mul_U10975(.A(dpath_mulcore_ary2_cout[55]), .Y(n2635));
AND2X1 mul_U10976(.A(n5643), .B(n5021), .Y(dpath_mulcore_ary2_cout[54]));
INVX1 mul_U10977(.A(dpath_mulcore_ary2_cout[54]), .Y(n2636));
AND2X1 mul_U10978(.A(n5644), .B(n5022), .Y(dpath_mulcore_ary2_cout[53]));
INVX1 mul_U10979(.A(dpath_mulcore_ary2_cout[53]), .Y(n2637));
AND2X1 mul_U10980(.A(n5645), .B(n5023), .Y(dpath_mulcore_ary2_cout[52]));
INVX1 mul_U10981(.A(dpath_mulcore_ary2_cout[52]), .Y(n2638));
AND2X1 mul_U10982(.A(n5646), .B(n5024), .Y(dpath_mulcore_ary2_cout[51]));
INVX1 mul_U10983(.A(dpath_mulcore_ary2_cout[51]), .Y(n2639));
AND2X1 mul_U10984(.A(n5647), .B(n5025), .Y(dpath_mulcore_ary2_cout[50]));
INVX1 mul_U10985(.A(dpath_mulcore_ary2_cout[50]), .Y(n2640));
AND2X1 mul_U10986(.A(n5648), .B(n5026), .Y(dpath_mulcore_ary2_cout[4]));
INVX1 mul_U10987(.A(dpath_mulcore_ary2_cout[4]), .Y(n2641));
AND2X1 mul_U10988(.A(n5649), .B(n5027), .Y(dpath_mulcore_ary2_cout[49]));
INVX1 mul_U10989(.A(dpath_mulcore_ary2_cout[49]), .Y(n2642));
AND2X1 mul_U10990(.A(n5650), .B(n5028), .Y(dpath_mulcore_ary2_cout[48]));
INVX1 mul_U10991(.A(dpath_mulcore_ary2_cout[48]), .Y(n2643));
AND2X1 mul_U10992(.A(n5651), .B(n5029), .Y(dpath_mulcore_ary2_cout[47]));
INVX1 mul_U10993(.A(dpath_mulcore_ary2_cout[47]), .Y(n2644));
AND2X1 mul_U10994(.A(n5652), .B(n5030), .Y(dpath_mulcore_ary2_cout[46]));
INVX1 mul_U10995(.A(dpath_mulcore_ary2_cout[46]), .Y(n2645));
AND2X1 mul_U10996(.A(n5653), .B(n5031), .Y(dpath_mulcore_ary2_cout[45]));
INVX1 mul_U10997(.A(dpath_mulcore_ary2_cout[45]), .Y(n2646));
AND2X1 mul_U10998(.A(n5654), .B(n5032), .Y(dpath_mulcore_ary2_cout[44]));
INVX1 mul_U10999(.A(dpath_mulcore_ary2_cout[44]), .Y(n2647));
AND2X1 mul_U11000(.A(n5655), .B(n5033), .Y(dpath_mulcore_ary2_cout[43]));
INVX1 mul_U11001(.A(dpath_mulcore_ary2_cout[43]), .Y(n2648));
AND2X1 mul_U11002(.A(n5656), .B(n5034), .Y(dpath_mulcore_ary2_cout[42]));
INVX1 mul_U11003(.A(dpath_mulcore_ary2_cout[42]), .Y(n2649));
AND2X1 mul_U11004(.A(n5657), .B(n5035), .Y(dpath_mulcore_ary2_cout[41]));
INVX1 mul_U11005(.A(dpath_mulcore_ary2_cout[41]), .Y(n2650));
AND2X1 mul_U11006(.A(n5658), .B(n5036), .Y(dpath_mulcore_ary2_cout[40]));
INVX1 mul_U11007(.A(dpath_mulcore_ary2_cout[40]), .Y(n2651));
AND2X1 mul_U11008(.A(n5659), .B(n5037), .Y(dpath_mulcore_ary2_cout[3]));
INVX1 mul_U11009(.A(dpath_mulcore_ary2_cout[3]), .Y(n2652));
AND2X1 mul_U11010(.A(n5660), .B(n5038), .Y(dpath_mulcore_ary2_cout[39]));
INVX1 mul_U11011(.A(dpath_mulcore_ary2_cout[39]), .Y(n2653));
AND2X1 mul_U11012(.A(n5661), .B(n5039), .Y(dpath_mulcore_ary2_cout[38]));
INVX1 mul_U11013(.A(dpath_mulcore_ary2_cout[38]), .Y(n2654));
AND2X1 mul_U11014(.A(n5662), .B(n5040), .Y(dpath_mulcore_ary2_cout[37]));
INVX1 mul_U11015(.A(dpath_mulcore_ary2_cout[37]), .Y(n2655));
AND2X1 mul_U11016(.A(n5663), .B(n5041), .Y(dpath_mulcore_ary2_cout[36]));
INVX1 mul_U11017(.A(dpath_mulcore_ary2_cout[36]), .Y(n2656));
AND2X1 mul_U11018(.A(n5664), .B(n5042), .Y(dpath_mulcore_ary2_cout[35]));
INVX1 mul_U11019(.A(dpath_mulcore_ary2_cout[35]), .Y(n2657));
AND2X1 mul_U11020(.A(n5665), .B(n5043), .Y(dpath_mulcore_ary2_cout[34]));
INVX1 mul_U11021(.A(dpath_mulcore_ary2_cout[34]), .Y(n2658));
AND2X1 mul_U11022(.A(n5666), .B(n5044), .Y(dpath_mulcore_ary2_cout[33]));
INVX1 mul_U11023(.A(dpath_mulcore_ary2_cout[33]), .Y(n2659));
AND2X1 mul_U11024(.A(n5667), .B(n5045), .Y(dpath_mulcore_ary2_cout[32]));
INVX1 mul_U11025(.A(dpath_mulcore_ary2_cout[32]), .Y(n2660));
AND2X1 mul_U11026(.A(n5668), .B(n5046), .Y(dpath_mulcore_ary2_cout[31]));
INVX1 mul_U11027(.A(dpath_mulcore_ary2_cout[31]), .Y(n2661));
AND2X1 mul_U11028(.A(n5669), .B(n5047), .Y(dpath_mulcore_ary2_cout[30]));
INVX1 mul_U11029(.A(dpath_mulcore_ary2_cout[30]), .Y(n2662));
AND2X1 mul_U11030(.A(n5670), .B(n5048), .Y(dpath_mulcore_ary2_cout[2]));
INVX1 mul_U11031(.A(dpath_mulcore_ary2_cout[2]), .Y(n2663));
AND2X1 mul_U11032(.A(n5671), .B(n5049), .Y(dpath_mulcore_ary2_cout[29]));
INVX1 mul_U11033(.A(dpath_mulcore_ary2_cout[29]), .Y(n2664));
AND2X1 mul_U11034(.A(n5672), .B(n5050), .Y(dpath_mulcore_ary2_cout[28]));
INVX1 mul_U11035(.A(dpath_mulcore_ary2_cout[28]), .Y(n2665));
AND2X1 mul_U11036(.A(n5673), .B(n5051), .Y(dpath_mulcore_ary2_cout[27]));
INVX1 mul_U11037(.A(dpath_mulcore_ary2_cout[27]), .Y(n2666));
AND2X1 mul_U11038(.A(n5674), .B(n5052), .Y(dpath_mulcore_ary2_cout[26]));
INVX1 mul_U11039(.A(dpath_mulcore_ary2_cout[26]), .Y(n2667));
AND2X1 mul_U11040(.A(n5675), .B(n5053), .Y(dpath_mulcore_ary2_cout[25]));
INVX1 mul_U11041(.A(dpath_mulcore_ary2_cout[25]), .Y(n2668));
AND2X1 mul_U11042(.A(n5676), .B(n5054), .Y(dpath_mulcore_ary2_cout[24]));
INVX1 mul_U11043(.A(dpath_mulcore_ary2_cout[24]), .Y(n2669));
AND2X1 mul_U11044(.A(n5677), .B(n5055), .Y(dpath_mulcore_ary2_cout[23]));
INVX1 mul_U11045(.A(dpath_mulcore_ary2_cout[23]), .Y(n2670));
AND2X1 mul_U11046(.A(n5678), .B(n5056), .Y(dpath_mulcore_ary2_cout[22]));
INVX1 mul_U11047(.A(dpath_mulcore_ary2_cout[22]), .Y(n2671));
AND2X1 mul_U11048(.A(n5679), .B(n5057), .Y(dpath_mulcore_ary2_cout[21]));
INVX1 mul_U11049(.A(dpath_mulcore_ary2_cout[21]), .Y(n2672));
AND2X1 mul_U11050(.A(n5680), .B(n5058), .Y(dpath_mulcore_ary2_cout[20]));
INVX1 mul_U11051(.A(dpath_mulcore_ary2_cout[20]), .Y(n2673));
AND2X1 mul_U11052(.A(n5681), .B(n5059), .Y(dpath_mulcore_ary2_cout[1]));
INVX1 mul_U11053(.A(dpath_mulcore_ary2_cout[1]), .Y(n2674));
AND2X1 mul_U11054(.A(n5682), .B(n5060), .Y(dpath_mulcore_ary2_cout[19]));
INVX1 mul_U11055(.A(dpath_mulcore_ary2_cout[19]), .Y(n2675));
AND2X1 mul_U11056(.A(n5683), .B(n5061), .Y(dpath_mulcore_ary2_cout[18]));
INVX1 mul_U11057(.A(dpath_mulcore_ary2_cout[18]), .Y(n2676));
AND2X1 mul_U11058(.A(n5684), .B(n5062), .Y(dpath_mulcore_ary2_cout[17]));
INVX1 mul_U11059(.A(dpath_mulcore_ary2_cout[17]), .Y(n2677));
AND2X1 mul_U11060(.A(n5685), .B(n5063), .Y(dpath_mulcore_ary2_cout[16]));
INVX1 mul_U11061(.A(dpath_mulcore_ary2_cout[16]), .Y(n2678));
AND2X1 mul_U11062(.A(n5686), .B(n5064), .Y(dpath_mulcore_ary2_cout[15]));
INVX1 mul_U11063(.A(dpath_mulcore_ary2_cout[15]), .Y(n2679));
AND2X1 mul_U11064(.A(n5687), .B(n5065), .Y(dpath_mulcore_ary2_cout[14]));
INVX1 mul_U11065(.A(dpath_mulcore_ary2_cout[14]), .Y(n2680));
AND2X1 mul_U11066(.A(n5688), .B(n5066), .Y(dpath_mulcore_ary2_cout[13]));
INVX1 mul_U11067(.A(dpath_mulcore_ary2_cout[13]), .Y(n2681));
AND2X1 mul_U11068(.A(n5689), .B(n5067), .Y(dpath_mulcore_ary2_cout[12]));
INVX1 mul_U11069(.A(dpath_mulcore_ary2_cout[12]), .Y(n2682));
AND2X1 mul_U11070(.A(n5690), .B(n5068), .Y(dpath_mulcore_ary2_cout[11]));
INVX1 mul_U11071(.A(dpath_mulcore_ary2_cout[11]), .Y(n2683));
AND2X1 mul_U11072(.A(n5691), .B(n5069), .Y(dpath_mulcore_ary2_cout[10]));
INVX1 mul_U11073(.A(dpath_mulcore_ary2_cout[10]), .Y(n2684));
AND2X1 mul_U11074(.A(n5692), .B(n5070), .Y(dpath_mulcore_ary2_cout[0]));
INVX1 mul_U11075(.A(dpath_mulcore_ary2_cout[0]), .Y(n2685));
OR2X1 mul_U11076(.A(se), .B(n9815), .Y(dpath_mulcore_cyc1_dff_n3));
INVX1 mul_U11077(.A(dpath_mulcore_cyc1_dff_n3), .Y(n2686));
AND2X1 mul_U11078(.A(dpath_n9), .B(dpath_n10), .Y(dpath_mulcore_rs1_l[63]));
INVX1 mul_U11079(.A(dpath_mulcore_rs1_l[63]), .Y(n2687));
AND2X1 mul_U11080(.A(dpath_n11), .B(dpath_n12), .Y(dpath_mulcore_rs1_l[62]));
INVX1 mul_U11081(.A(dpath_mulcore_rs1_l[62]), .Y(n2688));
AND2X1 mul_U11082(.A(dpath_n13), .B(dpath_n14), .Y(dpath_mulcore_rs1_l[61]));
INVX1 mul_U11083(.A(dpath_mulcore_rs1_l[61]), .Y(n2689));
AND2X1 mul_U11084(.A(dpath_n15), .B(dpath_n16), .Y(dpath_mulcore_rs1_l[60]));
INVX1 mul_U11085(.A(dpath_mulcore_rs1_l[60]), .Y(n2690));
AND2X1 mul_U11086(.A(dpath_n17), .B(dpath_n18), .Y(dpath_mulcore_rs1_l[59]));
INVX1 mul_U11087(.A(dpath_mulcore_rs1_l[59]), .Y(n2691));
AND2X1 mul_U11088(.A(dpath_n19), .B(dpath_n20), .Y(dpath_mulcore_rs1_l[58]));
INVX1 mul_U11089(.A(dpath_mulcore_rs1_l[58]), .Y(n2692));
AND2X1 mul_U11090(.A(dpath_n21), .B(dpath_n22), .Y(dpath_mulcore_rs1_l[57]));
INVX1 mul_U11091(.A(dpath_mulcore_rs1_l[57]), .Y(n2693));
AND2X1 mul_U11092(.A(dpath_n23), .B(dpath_n24), .Y(dpath_mulcore_rs1_l[56]));
INVX1 mul_U11093(.A(dpath_mulcore_rs1_l[56]), .Y(n2694));
AND2X1 mul_U11094(.A(dpath_n25), .B(dpath_n26), .Y(dpath_mulcore_rs1_l[55]));
INVX1 mul_U11095(.A(dpath_mulcore_rs1_l[55]), .Y(n2695));
AND2X1 mul_U11096(.A(dpath_n27), .B(dpath_n28), .Y(dpath_mulcore_rs1_l[54]));
INVX1 mul_U11097(.A(dpath_mulcore_rs1_l[54]), .Y(n2696));
AND2X1 mul_U11098(.A(dpath_n29), .B(dpath_n30), .Y(dpath_mulcore_rs1_l[53]));
INVX1 mul_U11099(.A(dpath_mulcore_rs1_l[53]), .Y(n2697));
AND2X1 mul_U11100(.A(dpath_n31), .B(dpath_n32), .Y(dpath_mulcore_rs1_l[52]));
INVX1 mul_U11101(.A(dpath_mulcore_rs1_l[52]), .Y(n2698));
AND2X1 mul_U11102(.A(dpath_n33), .B(dpath_n34), .Y(dpath_mulcore_rs1_l[51]));
INVX1 mul_U11103(.A(dpath_mulcore_rs1_l[51]), .Y(n2699));
AND2X1 mul_U11104(.A(dpath_n35), .B(dpath_n36), .Y(dpath_mulcore_rs1_l[50]));
INVX1 mul_U11105(.A(dpath_mulcore_rs1_l[50]), .Y(n2700));
AND2X1 mul_U11106(.A(dpath_n37), .B(dpath_n38), .Y(dpath_mulcore_rs1_l[49]));
INVX1 mul_U11107(.A(dpath_mulcore_rs1_l[49]), .Y(n2701));
AND2X1 mul_U11108(.A(dpath_n39), .B(dpath_n40), .Y(dpath_mulcore_rs1_l[48]));
INVX1 mul_U11109(.A(dpath_mulcore_rs1_l[48]), .Y(n2702));
AND2X1 mul_U11110(.A(dpath_n41), .B(dpath_n42), .Y(dpath_mulcore_rs1_l[47]));
INVX1 mul_U11111(.A(dpath_mulcore_rs1_l[47]), .Y(n2703));
AND2X1 mul_U11112(.A(dpath_n43), .B(dpath_n44), .Y(dpath_mulcore_rs1_l[46]));
INVX1 mul_U11113(.A(dpath_mulcore_rs1_l[46]), .Y(n2704));
AND2X1 mul_U11114(.A(dpath_n45), .B(dpath_n46), .Y(dpath_mulcore_rs1_l[45]));
INVX1 mul_U11115(.A(dpath_mulcore_rs1_l[45]), .Y(n2705));
AND2X1 mul_U11116(.A(dpath_n47), .B(dpath_n48), .Y(dpath_mulcore_rs1_l[44]));
INVX1 mul_U11117(.A(dpath_mulcore_rs1_l[44]), .Y(n2706));
AND2X1 mul_U11118(.A(dpath_n49), .B(dpath_n50), .Y(dpath_mulcore_rs1_l[43]));
INVX1 mul_U11119(.A(dpath_mulcore_rs1_l[43]), .Y(n2707));
AND2X1 mul_U11120(.A(dpath_n51), .B(dpath_n52), .Y(dpath_mulcore_rs1_l[42]));
INVX1 mul_U11121(.A(dpath_mulcore_rs1_l[42]), .Y(n2708));
AND2X1 mul_U11122(.A(dpath_n53), .B(dpath_n54), .Y(dpath_mulcore_rs1_l[41]));
INVX1 mul_U11123(.A(dpath_mulcore_rs1_l[41]), .Y(n2709));
AND2X1 mul_U11124(.A(dpath_n55), .B(dpath_n56), .Y(dpath_mulcore_rs1_l[40]));
INVX1 mul_U11125(.A(dpath_mulcore_rs1_l[40]), .Y(n2710));
AND2X1 mul_U11126(.A(dpath_n57), .B(dpath_n58), .Y(dpath_mulcore_rs1_l[39]));
INVX1 mul_U11127(.A(dpath_mulcore_rs1_l[39]), .Y(n2711));
AND2X1 mul_U11128(.A(dpath_n59), .B(dpath_n60), .Y(dpath_mulcore_rs1_l[38]));
INVX1 mul_U11129(.A(dpath_mulcore_rs1_l[38]), .Y(n2712));
AND2X1 mul_U11130(.A(dpath_n61), .B(dpath_n62), .Y(dpath_mulcore_rs1_l[37]));
INVX1 mul_U11131(.A(dpath_mulcore_rs1_l[37]), .Y(n2713));
AND2X1 mul_U11132(.A(dpath_n63), .B(dpath_n64), .Y(dpath_mulcore_rs1_l[36]));
INVX1 mul_U11133(.A(dpath_mulcore_rs1_l[36]), .Y(n2714));
AND2X1 mul_U11134(.A(dpath_n65), .B(dpath_n66), .Y(dpath_mulcore_rs1_l[35]));
INVX1 mul_U11135(.A(dpath_mulcore_rs1_l[35]), .Y(n2715));
AND2X1 mul_U11136(.A(dpath_n67), .B(dpath_n68), .Y(dpath_mulcore_rs1_l[34]));
INVX1 mul_U11137(.A(dpath_mulcore_rs1_l[34]), .Y(n2716));
AND2X1 mul_U11138(.A(dpath_n69), .B(dpath_n70), .Y(dpath_mulcore_rs1_l[33]));
INVX1 mul_U11139(.A(dpath_mulcore_rs1_l[33]), .Y(n2717));
AND2X1 mul_U11140(.A(dpath_n71), .B(dpath_n72), .Y(dpath_mulcore_rs1_l[32]));
INVX1 mul_U11141(.A(dpath_mulcore_rs1_l[32]), .Y(n2718));
AND2X1 mul_U11142(.A(dpath_n73), .B(dpath_n74), .Y(dpath_mulcore_rs1_l[31]));
INVX1 mul_U11143(.A(dpath_mulcore_rs1_l[31]), .Y(n2719));
AND2X1 mul_U11144(.A(dpath_n75), .B(dpath_n76), .Y(dpath_mulcore_rs1_l[30]));
INVX1 mul_U11145(.A(dpath_mulcore_rs1_l[30]), .Y(n2720));
AND2X1 mul_U11146(.A(dpath_n77), .B(dpath_n78), .Y(dpath_mulcore_rs1_l[29]));
INVX1 mul_U11147(.A(dpath_mulcore_rs1_l[29]), .Y(n2721));
AND2X1 mul_U11148(.A(dpath_n79), .B(dpath_n80), .Y(dpath_mulcore_rs1_l[28]));
INVX1 mul_U11149(.A(dpath_mulcore_rs1_l[28]), .Y(n2722));
AND2X1 mul_U11150(.A(dpath_n81), .B(dpath_n82), .Y(dpath_mulcore_rs1_l[27]));
INVX1 mul_U11151(.A(dpath_mulcore_rs1_l[27]), .Y(n2723));
AND2X1 mul_U11152(.A(dpath_n83), .B(dpath_n84), .Y(dpath_mulcore_rs1_l[26]));
INVX1 mul_U11153(.A(dpath_mulcore_rs1_l[26]), .Y(n2724));
AND2X1 mul_U11154(.A(dpath_n85), .B(dpath_n86), .Y(dpath_mulcore_rs1_l[25]));
INVX1 mul_U11155(.A(dpath_mulcore_rs1_l[25]), .Y(n2725));
AND2X1 mul_U11156(.A(dpath_n87), .B(dpath_n88), .Y(dpath_mulcore_rs1_l[24]));
INVX1 mul_U11157(.A(dpath_mulcore_rs1_l[24]), .Y(n2726));
AND2X1 mul_U11158(.A(dpath_n89), .B(dpath_n90), .Y(dpath_mulcore_rs1_l[23]));
INVX1 mul_U11159(.A(dpath_mulcore_rs1_l[23]), .Y(n2727));
AND2X1 mul_U11160(.A(dpath_n91), .B(dpath_n92), .Y(dpath_mulcore_rs1_l[22]));
INVX1 mul_U11161(.A(dpath_mulcore_rs1_l[22]), .Y(n2728));
AND2X1 mul_U11162(.A(dpath_n93), .B(dpath_n94), .Y(dpath_mulcore_rs1_l[21]));
INVX1 mul_U11163(.A(dpath_mulcore_rs1_l[21]), .Y(n2729));
AND2X1 mul_U11164(.A(dpath_n95), .B(dpath_n96), .Y(dpath_mulcore_rs1_l[20]));
INVX1 mul_U11165(.A(dpath_mulcore_rs1_l[20]), .Y(n2730));
AND2X1 mul_U11166(.A(dpath_n97), .B(dpath_n98), .Y(dpath_mulcore_rs1_l[19]));
INVX1 mul_U11167(.A(dpath_mulcore_rs1_l[19]), .Y(n2731));
AND2X1 mul_U11168(.A(dpath_n99), .B(dpath_n100), .Y(dpath_mulcore_rs1_l[18]));
INVX1 mul_U11169(.A(dpath_mulcore_rs1_l[18]), .Y(n2732));
AND2X1 mul_U11170(.A(dpath_n101), .B(dpath_n102), .Y(dpath_mulcore_rs1_l[17]));
INVX1 mul_U11171(.A(dpath_mulcore_rs1_l[17]), .Y(n2733));
AND2X1 mul_U11172(.A(dpath_n103), .B(dpath_n104), .Y(dpath_mulcore_rs1_l[16]));
INVX1 mul_U11173(.A(dpath_mulcore_rs1_l[16]), .Y(n2734));
AND2X1 mul_U11174(.A(dpath_n105), .B(dpath_n106), .Y(dpath_mulcore_rs1_l[15]));
INVX1 mul_U11175(.A(dpath_mulcore_rs1_l[15]), .Y(n2735));
AND2X1 mul_U11176(.A(dpath_n107), .B(dpath_n108), .Y(dpath_mulcore_rs1_l[14]));
INVX1 mul_U11177(.A(dpath_mulcore_rs1_l[14]), .Y(n2736));
AND2X1 mul_U11178(.A(dpath_n109), .B(dpath_n110), .Y(dpath_mulcore_rs1_l[13]));
INVX1 mul_U11179(.A(dpath_mulcore_rs1_l[13]), .Y(n2737));
AND2X1 mul_U11180(.A(dpath_n111), .B(dpath_n112), .Y(dpath_mulcore_rs1_l[12]));
INVX1 mul_U11181(.A(dpath_mulcore_rs1_l[12]), .Y(n2738));
AND2X1 mul_U11182(.A(dpath_n113), .B(dpath_n114), .Y(dpath_mulcore_rs1_l[11]));
INVX1 mul_U11183(.A(dpath_mulcore_rs1_l[11]), .Y(n2739));
AND2X1 mul_U11184(.A(dpath_n115), .B(dpath_n116), .Y(dpath_mulcore_rs1_l[10]));
INVX1 mul_U11185(.A(dpath_mulcore_rs1_l[10]), .Y(n2740));
AND2X1 mul_U11186(.A(dpath_n117), .B(dpath_n118), .Y(dpath_mulcore_rs1_l[9]));
INVX1 mul_U11187(.A(dpath_mulcore_rs1_l[9]), .Y(n2741));
AND2X1 mul_U11188(.A(dpath_n119), .B(dpath_n120), .Y(dpath_mulcore_rs1_l[8]));
INVX1 mul_U11189(.A(dpath_mulcore_rs1_l[8]), .Y(n2742));
AND2X1 mul_U11190(.A(dpath_n121), .B(dpath_n122), .Y(dpath_mulcore_rs1_l[7]));
INVX1 mul_U11191(.A(dpath_mulcore_rs1_l[7]), .Y(n2743));
AND2X1 mul_U11192(.A(dpath_n123), .B(dpath_n124), .Y(dpath_mulcore_rs1_l[6]));
INVX1 mul_U11193(.A(dpath_mulcore_rs1_l[6]), .Y(n2744));
AND2X1 mul_U11194(.A(dpath_n125), .B(dpath_n126), .Y(dpath_mulcore_rs1_l[5]));
INVX1 mul_U11195(.A(dpath_mulcore_rs1_l[5]), .Y(n2745));
AND2X1 mul_U11196(.A(dpath_n127), .B(dpath_n128), .Y(dpath_mulcore_rs1_l[4]));
INVX1 mul_U11197(.A(dpath_mulcore_rs1_l[4]), .Y(n2746));
AND2X1 mul_U11198(.A(dpath_n129), .B(dpath_n130), .Y(dpath_mulcore_rs1_l[3]));
INVX1 mul_U11199(.A(dpath_mulcore_rs1_l[3]), .Y(n2747));
AND2X1 mul_U11200(.A(dpath_n131), .B(dpath_n132), .Y(dpath_mulcore_rs1_l[2]));
INVX1 mul_U11201(.A(dpath_mulcore_rs1_l[2]), .Y(n2748));
AND2X1 mul_U11202(.A(dpath_n133), .B(dpath_n134), .Y(dpath_mulcore_rs1_l[1]));
INVX1 mul_U11203(.A(dpath_mulcore_rs1_l[1]), .Y(n2749));
AND2X1 mul_U11204(.A(dpath_n135), .B(dpath_n136), .Y(dpath_mulcore_rs1_l[0]));
INVX1 mul_U11205(.A(dpath_mulcore_rs1_l[0]), .Y(n2750));
AND2X1 mul_U11206(.A(exu_mul_rs2_data[9]), .B(n9772), .Y(dpath_n139));
INVX1 mul_U11207(.A(dpath_n139), .Y(n2751));
AND2X1 mul_U11208(.A(dpath_mout[9]), .B(n9762), .Y(dpath_n142));
INVX1 mul_U11209(.A(dpath_n142), .Y(n2752));
AND2X1 mul_U11210(.A(exu_mul_rs2_data[8]), .B(n9772), .Y(dpath_n148));
INVX1 mul_U11211(.A(dpath_n148), .Y(n2753));
AND2X1 mul_U11212(.A(dpath_mout[8]), .B(n9762), .Y(dpath_n150));
INVX1 mul_U11213(.A(dpath_n150), .Y(n2754));
AND2X1 mul_U11214(.A(exu_mul_rs2_data[7]), .B(n9773), .Y(dpath_n154));
INVX1 mul_U11215(.A(dpath_n154), .Y(n2755));
AND2X1 mul_U11216(.A(dpath_mout[7]), .B(n9762), .Y(dpath_n156));
INVX1 mul_U11217(.A(dpath_n156), .Y(n2756));
AND2X1 mul_U11218(.A(exu_mul_rs2_data[6]), .B(n7198), .Y(dpath_n160));
INVX1 mul_U11219(.A(dpath_n160), .Y(n2757));
AND2X1 mul_U11220(.A(dpath_mout[6]), .B(n9762), .Y(dpath_n162));
INVX1 mul_U11221(.A(dpath_n162), .Y(n2758));
AND2X1 mul_U11222(.A(exu_mul_rs2_data[63]), .B(n9774), .Y(dpath_n166));
INVX1 mul_U11223(.A(dpath_n166), .Y(n2759));
AND2X1 mul_U11224(.A(dpath_mout[63]), .B(n9762), .Y(dpath_n168));
INVX1 mul_U11225(.A(dpath_n168), .Y(n2760));
AND2X1 mul_U11226(.A(exu_mul_rs2_data[62]), .B(n9774), .Y(dpath_n172));
INVX1 mul_U11227(.A(dpath_n172), .Y(n2761));
AND2X1 mul_U11228(.A(dpath_mout[62]), .B(n9762), .Y(dpath_n174));
INVX1 mul_U11229(.A(dpath_n174), .Y(n2762));
AND2X1 mul_U11230(.A(exu_mul_rs2_data[61]), .B(n9773), .Y(dpath_n178));
INVX1 mul_U11231(.A(dpath_n178), .Y(n2763));
AND2X1 mul_U11232(.A(dpath_mout[61]), .B(n9762), .Y(dpath_n180));
INVX1 mul_U11233(.A(dpath_n180), .Y(n2764));
AND2X1 mul_U11234(.A(exu_mul_rs2_data[60]), .B(n9772), .Y(dpath_n184));
INVX1 mul_U11235(.A(dpath_n184), .Y(n2765));
AND2X1 mul_U11236(.A(dpath_mout[60]), .B(n9762), .Y(dpath_n186));
INVX1 mul_U11237(.A(dpath_n186), .Y(n2766));
AND2X1 mul_U11238(.A(exu_mul_rs2_data[5]), .B(n9773), .Y(dpath_n190));
INVX1 mul_U11239(.A(dpath_n190), .Y(n2767));
AND2X1 mul_U11240(.A(dpath_mout[5]), .B(n9762), .Y(dpath_n192));
INVX1 mul_U11241(.A(dpath_n192), .Y(n2768));
AND2X1 mul_U11242(.A(exu_mul_rs2_data[59]), .B(n7198), .Y(dpath_n196));
INVX1 mul_U11243(.A(dpath_n196), .Y(n2769));
AND2X1 mul_U11244(.A(dpath_mout[59]), .B(n9762), .Y(dpath_n198));
INVX1 mul_U11245(.A(dpath_n198), .Y(n2770));
AND2X1 mul_U11246(.A(exu_mul_rs2_data[58]), .B(n9774), .Y(dpath_n202));
INVX1 mul_U11247(.A(dpath_n202), .Y(n2771));
AND2X1 mul_U11248(.A(dpath_mout[58]), .B(n9762), .Y(dpath_n204));
INVX1 mul_U11249(.A(dpath_n204), .Y(n2772));
AND2X1 mul_U11250(.A(exu_mul_rs2_data[57]), .B(n9772), .Y(dpath_n208));
INVX1 mul_U11251(.A(dpath_n208), .Y(n2773));
AND2X1 mul_U11252(.A(dpath_mout[57]), .B(n9762), .Y(dpath_n210));
INVX1 mul_U11253(.A(dpath_n210), .Y(n2774));
AND2X1 mul_U11254(.A(exu_mul_rs2_data[56]), .B(n9772), .Y(dpath_n214));
INVX1 mul_U11255(.A(dpath_n214), .Y(n2775));
AND2X1 mul_U11256(.A(dpath_mout[56]), .B(n9762), .Y(dpath_n216));
INVX1 mul_U11257(.A(dpath_n216), .Y(n2776));
AND2X1 mul_U11258(.A(exu_mul_rs2_data[55]), .B(n9773), .Y(dpath_n220));
INVX1 mul_U11259(.A(dpath_n220), .Y(n2777));
AND2X1 mul_U11260(.A(dpath_mout[55]), .B(dpath_n145), .Y(dpath_n222));
INVX1 mul_U11261(.A(dpath_n222), .Y(n2778));
AND2X1 mul_U11262(.A(exu_mul_rs2_data[54]), .B(n7198), .Y(dpath_n226));
INVX1 mul_U11263(.A(dpath_n226), .Y(n2779));
AND2X1 mul_U11264(.A(dpath_mout[54]), .B(n9762), .Y(dpath_n228));
INVX1 mul_U11265(.A(dpath_n228), .Y(n2780));
AND2X1 mul_U11266(.A(exu_mul_rs2_data[53]), .B(n9774), .Y(dpath_n232));
INVX1 mul_U11267(.A(dpath_n232), .Y(n2781));
AND2X1 mul_U11268(.A(dpath_mout[53]), .B(dpath_n145), .Y(dpath_n234));
INVX1 mul_U11269(.A(dpath_n234), .Y(n2782));
AND2X1 mul_U11270(.A(exu_mul_rs2_data[52]), .B(n9773), .Y(dpath_n238));
INVX1 mul_U11271(.A(dpath_n238), .Y(n2783));
AND2X1 mul_U11272(.A(dpath_mout[52]), .B(n9762), .Y(dpath_n240));
INVX1 mul_U11273(.A(dpath_n240), .Y(n2784));
AND2X1 mul_U11274(.A(exu_mul_rs2_data[51]), .B(n7198), .Y(dpath_n244));
INVX1 mul_U11275(.A(dpath_n244), .Y(n2785));
AND2X1 mul_U11276(.A(dpath_mout[51]), .B(dpath_n145), .Y(dpath_n246));
INVX1 mul_U11277(.A(dpath_n246), .Y(n2786));
AND2X1 mul_U11278(.A(exu_mul_rs2_data[50]), .B(n9774), .Y(dpath_n250));
INVX1 mul_U11279(.A(dpath_n250), .Y(n2787));
AND2X1 mul_U11280(.A(dpath_mout[50]), .B(n9762), .Y(dpath_n252));
INVX1 mul_U11281(.A(dpath_n252), .Y(n2788));
AND2X1 mul_U11282(.A(exu_mul_rs2_data[4]), .B(n9772), .Y(dpath_n256));
INVX1 mul_U11283(.A(dpath_n256), .Y(n2789));
AND2X1 mul_U11284(.A(dpath_mout[4]), .B(dpath_n145), .Y(dpath_n258));
INVX1 mul_U11285(.A(dpath_n258), .Y(n2790));
AND2X1 mul_U11286(.A(exu_mul_rs2_data[49]), .B(n9773), .Y(dpath_n262));
INVX1 mul_U11287(.A(dpath_n262), .Y(n2791));
AND2X1 mul_U11288(.A(dpath_mout[49]), .B(n9762), .Y(dpath_n264));
INVX1 mul_U11289(.A(dpath_n264), .Y(n2792));
AND2X1 mul_U11290(.A(exu_mul_rs2_data[48]), .B(n7198), .Y(dpath_n268));
INVX1 mul_U11291(.A(dpath_n268), .Y(n2793));
AND2X1 mul_U11292(.A(dpath_mout[48]), .B(dpath_n145), .Y(dpath_n270));
INVX1 mul_U11293(.A(dpath_n270), .Y(n2794));
AND2X1 mul_U11294(.A(exu_mul_rs2_data[47]), .B(n9774), .Y(dpath_n274));
INVX1 mul_U11295(.A(dpath_n274), .Y(n2795));
AND2X1 mul_U11296(.A(dpath_mout[47]), .B(n9762), .Y(dpath_n276));
INVX1 mul_U11297(.A(dpath_n276), .Y(n2796));
AND2X1 mul_U11298(.A(exu_mul_rs2_data[46]), .B(n7198), .Y(dpath_n280));
INVX1 mul_U11299(.A(dpath_n280), .Y(n2797));
AND2X1 mul_U11300(.A(dpath_mout[46]), .B(dpath_n145), .Y(dpath_n282));
INVX1 mul_U11301(.A(dpath_n282), .Y(n2798));
AND2X1 mul_U11302(.A(exu_mul_rs2_data[45]), .B(n9774), .Y(dpath_n286));
INVX1 mul_U11303(.A(dpath_n286), .Y(n2799));
AND2X1 mul_U11304(.A(dpath_mout[45]), .B(n9762), .Y(dpath_n288));
INVX1 mul_U11305(.A(dpath_n288), .Y(n2800));
AND2X1 mul_U11306(.A(exu_mul_rs2_data[44]), .B(n9772), .Y(dpath_n292));
INVX1 mul_U11307(.A(dpath_n292), .Y(n2801));
AND2X1 mul_U11308(.A(dpath_mout[44]), .B(dpath_n145), .Y(dpath_n294));
INVX1 mul_U11309(.A(dpath_n294), .Y(n2802));
AND2X1 mul_U11310(.A(exu_mul_rs2_data[43]), .B(n9773), .Y(dpath_n298));
INVX1 mul_U11311(.A(dpath_n298), .Y(n2803));
AND2X1 mul_U11312(.A(dpath_mout[43]), .B(n9762), .Y(dpath_n300));
INVX1 mul_U11313(.A(dpath_n300), .Y(n2804));
AND2X1 mul_U11314(.A(exu_mul_rs2_data[42]), .B(n9774), .Y(dpath_n304));
INVX1 mul_U11315(.A(dpath_n304), .Y(n2805));
AND2X1 mul_U11316(.A(dpath_mout[42]), .B(dpath_n145), .Y(dpath_n306));
INVX1 mul_U11317(.A(dpath_n306), .Y(n2806));
AND2X1 mul_U11318(.A(exu_mul_rs2_data[41]), .B(n9774), .Y(dpath_n310));
INVX1 mul_U11319(.A(dpath_n310), .Y(n2807));
AND2X1 mul_U11320(.A(dpath_mout[41]), .B(dpath_n145), .Y(dpath_n312));
INVX1 mul_U11321(.A(dpath_n312), .Y(n2808));
AND2X1 mul_U11322(.A(exu_mul_rs2_data[40]), .B(n9772), .Y(dpath_n316));
INVX1 mul_U11323(.A(dpath_n316), .Y(n2809));
AND2X1 mul_U11324(.A(dpath_mout[40]), .B(n9762), .Y(dpath_n318));
INVX1 mul_U11325(.A(dpath_n318), .Y(n2810));
AND2X1 mul_U11326(.A(exu_mul_rs2_data[3]), .B(n9773), .Y(dpath_n322));
INVX1 mul_U11327(.A(dpath_n322), .Y(n2811));
AND2X1 mul_U11328(.A(dpath_mout[3]), .B(dpath_n145), .Y(dpath_n324));
INVX1 mul_U11329(.A(dpath_n324), .Y(n2812));
AND2X1 mul_U11330(.A(exu_mul_rs2_data[39]), .B(n7198), .Y(dpath_n328));
INVX1 mul_U11331(.A(dpath_n328), .Y(n2813));
AND2X1 mul_U11332(.A(dpath_mout[39]), .B(n9762), .Y(dpath_n330));
INVX1 mul_U11333(.A(dpath_n330), .Y(n2814));
AND2X1 mul_U11334(.A(exu_mul_rs2_data[38]), .B(n9774), .Y(dpath_n334));
INVX1 mul_U11335(.A(dpath_n334), .Y(n2815));
AND2X1 mul_U11336(.A(dpath_mout[38]), .B(n9762), .Y(dpath_n336));
INVX1 mul_U11337(.A(dpath_n336), .Y(n2816));
AND2X1 mul_U11338(.A(exu_mul_rs2_data[37]), .B(n9772), .Y(dpath_n340));
INVX1 mul_U11339(.A(dpath_n340), .Y(n2817));
AND2X1 mul_U11340(.A(dpath_mout[37]), .B(dpath_n145), .Y(dpath_n342));
INVX1 mul_U11341(.A(dpath_n342), .Y(n2818));
AND2X1 mul_U11342(.A(exu_mul_rs2_data[36]), .B(n7198), .Y(dpath_n346));
INVX1 mul_U11343(.A(dpath_n346), .Y(n2819));
AND2X1 mul_U11344(.A(dpath_mout[36]), .B(dpath_n145), .Y(dpath_n348));
INVX1 mul_U11345(.A(dpath_n348), .Y(n2820));
AND2X1 mul_U11346(.A(exu_mul_rs2_data[35]), .B(n9773), .Y(dpath_n352));
INVX1 mul_U11347(.A(dpath_n352), .Y(n2821));
AND2X1 mul_U11348(.A(dpath_mout[35]), .B(n9762), .Y(dpath_n354));
INVX1 mul_U11349(.A(dpath_n354), .Y(n2822));
AND2X1 mul_U11350(.A(exu_mul_rs2_data[34]), .B(n9774), .Y(dpath_n358));
INVX1 mul_U11351(.A(dpath_n358), .Y(n2823));
AND2X1 mul_U11352(.A(dpath_mout[34]), .B(dpath_n145), .Y(dpath_n360));
INVX1 mul_U11353(.A(dpath_n360), .Y(n2824));
AND2X1 mul_U11354(.A(exu_mul_rs2_data[33]), .B(n9772), .Y(dpath_n364));
INVX1 mul_U11355(.A(dpath_n364), .Y(n2825));
AND2X1 mul_U11356(.A(dpath_mout[33]), .B(n9762), .Y(dpath_n366));
INVX1 mul_U11357(.A(dpath_n366), .Y(n2826));
AND2X1 mul_U11358(.A(exu_mul_rs2_data[32]), .B(n9773), .Y(dpath_n370));
INVX1 mul_U11359(.A(dpath_n370), .Y(n2827));
AND2X1 mul_U11360(.A(dpath_mout[32]), .B(n9762), .Y(dpath_n372));
INVX1 mul_U11361(.A(dpath_n372), .Y(n2828));
AND2X1 mul_U11362(.A(exu_mul_rs2_data[31]), .B(n7198), .Y(dpath_n376));
INVX1 mul_U11363(.A(dpath_n376), .Y(n2829));
AND2X1 mul_U11364(.A(dpath_mout[31]), .B(dpath_n145), .Y(dpath_n378));
INVX1 mul_U11365(.A(dpath_n378), .Y(n2830));
AND2X1 mul_U11366(.A(exu_mul_rs2_data[30]), .B(n9774), .Y(dpath_n382));
INVX1 mul_U11367(.A(dpath_n382), .Y(n2831));
AND2X1 mul_U11368(.A(dpath_mout[30]), .B(dpath_n145), .Y(dpath_n384));
INVX1 mul_U11369(.A(dpath_n384), .Y(n2832));
AND2X1 mul_U11370(.A(exu_mul_rs2_data[2]), .B(n9774), .Y(dpath_n388));
INVX1 mul_U11371(.A(dpath_n388), .Y(n2833));
AND2X1 mul_U11372(.A(dpath_mout[2]), .B(dpath_n145), .Y(dpath_n390));
INVX1 mul_U11373(.A(dpath_n390), .Y(n2834));
AND2X1 mul_U11374(.A(exu_mul_rs2_data[29]), .B(n9774), .Y(dpath_n394));
INVX1 mul_U11375(.A(dpath_n394), .Y(n2835));
AND2X1 mul_U11376(.A(dpath_mout[29]), .B(dpath_n145), .Y(dpath_n396));
INVX1 mul_U11377(.A(dpath_n396), .Y(n2836));
AND2X1 mul_U11378(.A(exu_mul_rs2_data[28]), .B(n9774), .Y(dpath_n400));
INVX1 mul_U11379(.A(dpath_n400), .Y(n2837));
AND2X1 mul_U11380(.A(dpath_mout[28]), .B(dpath_n145), .Y(dpath_n402));
INVX1 mul_U11381(.A(dpath_n402), .Y(n2838));
AND2X1 mul_U11382(.A(exu_mul_rs2_data[27]), .B(n7198), .Y(dpath_n406));
INVX1 mul_U11383(.A(dpath_n406), .Y(n2839));
AND2X1 mul_U11384(.A(dpath_mout[27]), .B(dpath_n145), .Y(dpath_n408));
INVX1 mul_U11385(.A(dpath_n408), .Y(n2840));
AND2X1 mul_U11386(.A(exu_mul_rs2_data[26]), .B(n7198), .Y(dpath_n412));
INVX1 mul_U11387(.A(dpath_n412), .Y(n2841));
AND2X1 mul_U11388(.A(dpath_mout[26]), .B(n9762), .Y(dpath_n414));
INVX1 mul_U11389(.A(dpath_n414), .Y(n2842));
AND2X1 mul_U11390(.A(exu_mul_rs2_data[25]), .B(n9773), .Y(dpath_n418));
INVX1 mul_U11391(.A(dpath_n418), .Y(n2843));
AND2X1 mul_U11392(.A(dpath_mout[25]), .B(n9762), .Y(dpath_n420));
INVX1 mul_U11393(.A(dpath_n420), .Y(n2844));
AND2X1 mul_U11394(.A(exu_mul_rs2_data[24]), .B(n9774), .Y(dpath_n424));
INVX1 mul_U11395(.A(dpath_n424), .Y(n2845));
AND2X1 mul_U11396(.A(dpath_mout[24]), .B(dpath_n145), .Y(dpath_n426));
INVX1 mul_U11397(.A(dpath_n426), .Y(n2846));
AND2X1 mul_U11398(.A(exu_mul_rs2_data[23]), .B(n7198), .Y(dpath_n430));
INVX1 mul_U11399(.A(dpath_n430), .Y(n2847));
AND2X1 mul_U11400(.A(dpath_mout[23]), .B(n9762), .Y(dpath_n432));
INVX1 mul_U11401(.A(dpath_n432), .Y(n2848));
AND2X1 mul_U11402(.A(exu_mul_rs2_data[22]), .B(n9774), .Y(dpath_n436));
INVX1 mul_U11403(.A(dpath_n436), .Y(n2849));
AND2X1 mul_U11404(.A(dpath_mout[22]), .B(n9762), .Y(dpath_n438));
INVX1 mul_U11405(.A(dpath_n438), .Y(n2850));
AND2X1 mul_U11406(.A(exu_mul_rs2_data[21]), .B(n9774), .Y(dpath_n442));
INVX1 mul_U11407(.A(dpath_n442), .Y(n2851));
AND2X1 mul_U11408(.A(dpath_mout[21]), .B(dpath_n145), .Y(dpath_n444));
INVX1 mul_U11409(.A(dpath_n444), .Y(n2852));
AND2X1 mul_U11410(.A(exu_mul_rs2_data[20]), .B(n9772), .Y(dpath_n448));
INVX1 mul_U11411(.A(dpath_n448), .Y(n2853));
AND2X1 mul_U11412(.A(dpath_mout[20]), .B(dpath_n145), .Y(dpath_n450));
INVX1 mul_U11413(.A(dpath_n450), .Y(n2854));
AND2X1 mul_U11414(.A(exu_mul_rs2_data[1]), .B(n9773), .Y(dpath_n454));
INVX1 mul_U11415(.A(dpath_n454), .Y(n2855));
AND2X1 mul_U11416(.A(dpath_mout[1]), .B(dpath_n145), .Y(dpath_n456));
INVX1 mul_U11417(.A(dpath_n456), .Y(n2856));
AND2X1 mul_U11418(.A(exu_mul_rs2_data[19]), .B(n7198), .Y(dpath_n460));
INVX1 mul_U11419(.A(dpath_n460), .Y(n2857));
AND2X1 mul_U11420(.A(dpath_mout[19]), .B(dpath_n145), .Y(dpath_n462));
INVX1 mul_U11421(.A(dpath_n462), .Y(n2858));
AND2X1 mul_U11422(.A(exu_mul_rs2_data[18]), .B(n7198), .Y(dpath_n466));
INVX1 mul_U11423(.A(dpath_n466), .Y(n2859));
AND2X1 mul_U11424(.A(dpath_mout[18]), .B(dpath_n145), .Y(dpath_n468));
INVX1 mul_U11425(.A(dpath_n468), .Y(n2860));
AND2X1 mul_U11426(.A(exu_mul_rs2_data[17]), .B(n7198), .Y(dpath_n472));
INVX1 mul_U11427(.A(dpath_n472), .Y(n2861));
AND2X1 mul_U11428(.A(dpath_mout[17]), .B(dpath_n145), .Y(dpath_n474));
INVX1 mul_U11429(.A(dpath_n474), .Y(n2862));
AND2X1 mul_U11430(.A(exu_mul_rs2_data[16]), .B(n7198), .Y(dpath_n478));
INVX1 mul_U11431(.A(dpath_n478), .Y(n2863));
AND2X1 mul_U11432(.A(dpath_mout[16]), .B(dpath_n145), .Y(dpath_n480));
INVX1 mul_U11433(.A(dpath_n480), .Y(n2864));
AND2X1 mul_U11434(.A(exu_mul_rs2_data[15]), .B(n7198), .Y(dpath_n484));
INVX1 mul_U11435(.A(dpath_n484), .Y(n2865));
AND2X1 mul_U11436(.A(dpath_mout[15]), .B(n9762), .Y(dpath_n486));
INVX1 mul_U11437(.A(dpath_n486), .Y(n2866));
AND2X1 mul_U11438(.A(exu_mul_rs2_data[14]), .B(n7198), .Y(dpath_n490));
INVX1 mul_U11439(.A(dpath_n490), .Y(n2867));
AND2X1 mul_U11440(.A(dpath_mout[14]), .B(dpath_n145), .Y(dpath_n492));
INVX1 mul_U11441(.A(dpath_n492), .Y(n2868));
AND2X1 mul_U11442(.A(exu_mul_rs2_data[13]), .B(n7198), .Y(dpath_n496));
INVX1 mul_U11443(.A(dpath_n496), .Y(n2869));
AND2X1 mul_U11444(.A(dpath_mout[13]), .B(n9762), .Y(dpath_n498));
INVX1 mul_U11445(.A(dpath_n498), .Y(n2870));
AND2X1 mul_U11446(.A(exu_mul_rs2_data[12]), .B(n7198), .Y(dpath_n502));
INVX1 mul_U11447(.A(dpath_n502), .Y(n2871));
AND2X1 mul_U11448(.A(dpath_mout[12]), .B(dpath_n145), .Y(dpath_n504));
INVX1 mul_U11449(.A(dpath_n504), .Y(n2872));
AND2X1 mul_U11450(.A(exu_mul_rs2_data[11]), .B(n7198), .Y(dpath_n508));
INVX1 mul_U11451(.A(dpath_n508), .Y(n2873));
AND2X1 mul_U11452(.A(dpath_mout[11]), .B(dpath_n145), .Y(dpath_n510));
INVX1 mul_U11453(.A(dpath_n510), .Y(n2874));
AND2X1 mul_U11454(.A(exu_mul_rs2_data[10]), .B(n9774), .Y(dpath_n514));
INVX1 mul_U11455(.A(dpath_n514), .Y(n2875));
AND2X1 mul_U11456(.A(dpath_mout[10]), .B(n9762), .Y(dpath_n516));
INVX1 mul_U11457(.A(dpath_n516), .Y(n2876));
AND2X1 mul_U11458(.A(exu_mul_rs2_data[0]), .B(n7198), .Y(dpath_n520));
INVX1 mul_U11459(.A(dpath_n520), .Y(n2877));
AND2X1 mul_U11460(.A(dpath_mout[0]), .B(n9762), .Y(dpath_n523));
INVX1 mul_U11461(.A(dpath_n523), .Y(n2878));
AND2X1 mul_U11462(.A(dpath_n658), .B(dpath_acc_reg[9]), .Y(dpath_n655));
INVX1 mul_U11463(.A(dpath_n655), .Y(n2879));
AND2X1 mul_U11464(.A(n9764), .B(dpath_mout[9]), .Y(dpath_n659));
INVX1 mul_U11465(.A(dpath_n659), .Y(n2880));
AND2X1 mul_U11466(.A(dpath_mout[128]), .B(n9767), .Y(dpath_n663));
INVX1 mul_U11467(.A(dpath_n663), .Y(n2881));
AND2X1 mul_U11468(.A(dpath_mout[127]), .B(n9767), .Y(dpath_n667));
INVX1 mul_U11469(.A(dpath_n667), .Y(n2882));
AND2X1 mul_U11470(.A(dpath_mout[126]), .B(n9767), .Y(dpath_n669));
INVX1 mul_U11471(.A(dpath_n669), .Y(n2883));
AND2X1 mul_U11472(.A(dpath_mout[125]), .B(n9767), .Y(dpath_n671));
INVX1 mul_U11473(.A(dpath_n671), .Y(n2884));
AND2X1 mul_U11474(.A(dpath_mout[124]), .B(n9767), .Y(dpath_n673));
INVX1 mul_U11475(.A(dpath_n673), .Y(n2885));
AND2X1 mul_U11476(.A(dpath_mout[123]), .B(n9767), .Y(dpath_n675));
INVX1 mul_U11477(.A(dpath_n675), .Y(n2886));
AND2X1 mul_U11478(.A(dpath_mout[122]), .B(n9767), .Y(dpath_n677));
INVX1 mul_U11479(.A(dpath_n677), .Y(n2887));
AND2X1 mul_U11480(.A(dpath_n658), .B(dpath_acc_reg[8]), .Y(dpath_n681));
INVX1 mul_U11481(.A(dpath_n681), .Y(n2888));
AND2X1 mul_U11482(.A(n9764), .B(dpath_mout[8]), .Y(dpath_n683));
INVX1 mul_U11483(.A(dpath_n683), .Y(n2889));
AND2X1 mul_U11484(.A(dpath_mout[121]), .B(n9767), .Y(dpath_n685));
INVX1 mul_U11485(.A(dpath_n685), .Y(n2890));
AND2X1 mul_U11486(.A(dpath_mout[120]), .B(n9767), .Y(dpath_n687));
INVX1 mul_U11487(.A(dpath_n687), .Y(n2891));
AND2X1 mul_U11488(.A(dpath_mout[119]), .B(n9767), .Y(dpath_n689));
INVX1 mul_U11489(.A(dpath_n689), .Y(n2892));
AND2X1 mul_U11490(.A(dpath_mout[118]), .B(n9767), .Y(dpath_n691));
INVX1 mul_U11491(.A(dpath_n691), .Y(n2893));
AND2X1 mul_U11492(.A(dpath_mout[117]), .B(n9767), .Y(dpath_n693));
INVX1 mul_U11493(.A(dpath_n693), .Y(n2894));
AND2X1 mul_U11494(.A(dpath_mout[116]), .B(n9767), .Y(dpath_n695));
INVX1 mul_U11495(.A(dpath_n695), .Y(n2895));
AND2X1 mul_U11496(.A(dpath_mout[115]), .B(n9767), .Y(dpath_n697));
INVX1 mul_U11497(.A(dpath_n697), .Y(n2896));
AND2X1 mul_U11498(.A(dpath_mout[114]), .B(dpath_n666), .Y(dpath_n699));
INVX1 mul_U11499(.A(dpath_n699), .Y(n2897));
AND2X1 mul_U11500(.A(dpath_mout[113]), .B(n9767), .Y(dpath_n701));
INVX1 mul_U11501(.A(dpath_n701), .Y(n2898));
AND2X1 mul_U11502(.A(dpath_mout[112]), .B(dpath_n666), .Y(dpath_n703));
INVX1 mul_U11503(.A(dpath_n703), .Y(n2899));
AND2X1 mul_U11504(.A(dpath_n658), .B(dpath_acc_reg[7]), .Y(dpath_n707));
INVX1 mul_U11505(.A(dpath_n707), .Y(n2900));
AND2X1 mul_U11506(.A(n9764), .B(dpath_mout[7]), .Y(dpath_n709));
INVX1 mul_U11507(.A(dpath_n709), .Y(n2901));
AND2X1 mul_U11508(.A(dpath_mout[111]), .B(n9767), .Y(dpath_n711));
INVX1 mul_U11509(.A(dpath_n711), .Y(n2902));
AND2X1 mul_U11510(.A(dpath_mout[110]), .B(dpath_n666), .Y(dpath_n713));
INVX1 mul_U11511(.A(dpath_n713), .Y(n2903));
AND2X1 mul_U11512(.A(dpath_mout[109]), .B(n9767), .Y(dpath_n715));
INVX1 mul_U11513(.A(dpath_n715), .Y(n2904));
AND2X1 mul_U11514(.A(dpath_mout[108]), .B(dpath_n666), .Y(dpath_n717));
INVX1 mul_U11515(.A(dpath_n717), .Y(n2905));
AND2X1 mul_U11516(.A(dpath_mout[107]), .B(n9767), .Y(dpath_n719));
INVX1 mul_U11517(.A(dpath_n719), .Y(n2906));
AND2X1 mul_U11518(.A(dpath_mout[106]), .B(dpath_n666), .Y(dpath_n721));
INVX1 mul_U11519(.A(dpath_n721), .Y(n2907));
AND2X1 mul_U11520(.A(dpath_mout[105]), .B(n9767), .Y(dpath_n723));
INVX1 mul_U11521(.A(dpath_n723), .Y(n2908));
AND2X1 mul_U11522(.A(dpath_mout[104]), .B(dpath_n666), .Y(dpath_n725));
INVX1 mul_U11523(.A(dpath_n725), .Y(n2909));
AND2X1 mul_U11524(.A(dpath_mout[103]), .B(n9767), .Y(dpath_n727));
INVX1 mul_U11525(.A(dpath_n727), .Y(n2910));
AND2X1 mul_U11526(.A(dpath_mout[102]), .B(n9767), .Y(dpath_n729));
INVX1 mul_U11527(.A(dpath_n729), .Y(n2911));
AND2X1 mul_U11528(.A(dpath_n658), .B(dpath_acc_reg[6]), .Y(dpath_n733));
INVX1 mul_U11529(.A(dpath_n733), .Y(n2912));
AND2X1 mul_U11530(.A(n9764), .B(dpath_mout[6]), .Y(dpath_n735));
INVX1 mul_U11531(.A(dpath_n735), .Y(n2913));
AND2X1 mul_U11532(.A(dpath_mout[101]), .B(dpath_n666), .Y(dpath_n737));
INVX1 mul_U11533(.A(dpath_n737), .Y(n2914));
AND2X1 mul_U11534(.A(dpath_mout[100]), .B(dpath_n666), .Y(dpath_n739));
INVX1 mul_U11535(.A(dpath_n739), .Y(n2915));
AND2X1 mul_U11536(.A(dpath_mout[99]), .B(n9767), .Y(dpath_n741));
INVX1 mul_U11537(.A(dpath_n741), .Y(n2916));
AND2X1 mul_U11538(.A(dpath_mout[98]), .B(dpath_n666), .Y(dpath_n743));
INVX1 mul_U11539(.A(dpath_n743), .Y(n2917));
AND2X1 mul_U11540(.A(dpath_mout[97]), .B(n9767), .Y(dpath_n745));
INVX1 mul_U11541(.A(dpath_n745), .Y(n2918));
AND2X1 mul_U11542(.A(dpath_mout[96]), .B(n9767), .Y(dpath_n747));
INVX1 mul_U11543(.A(dpath_n747), .Y(n2919));
AND2X1 mul_U11544(.A(dpath_mout[95]), .B(dpath_n666), .Y(dpath_n749));
INVX1 mul_U11545(.A(dpath_n749), .Y(n2920));
AND2X1 mul_U11546(.A(dpath_mout[94]), .B(dpath_n666), .Y(dpath_n751));
INVX1 mul_U11547(.A(dpath_n751), .Y(n2921));
AND2X1 mul_U11548(.A(dpath_mout[93]), .B(n9767), .Y(dpath_n753));
INVX1 mul_U11549(.A(dpath_n753), .Y(n2922));
AND2X1 mul_U11550(.A(dpath_mout[92]), .B(dpath_n666), .Y(dpath_n755));
INVX1 mul_U11551(.A(dpath_n755), .Y(n2923));
AND2X1 mul_U11552(.A(dpath_n658), .B(dpath_acc_reg[5]), .Y(dpath_n759));
INVX1 mul_U11553(.A(dpath_n759), .Y(n2924));
AND2X1 mul_U11554(.A(n9764), .B(dpath_mout[5]), .Y(dpath_n761));
INVX1 mul_U11555(.A(dpath_n761), .Y(n2925));
AND2X1 mul_U11556(.A(dpath_mout[91]), .B(n9767), .Y(dpath_n763));
INVX1 mul_U11557(.A(dpath_n763), .Y(n2926));
AND2X1 mul_U11558(.A(dpath_mout[90]), .B(n9767), .Y(dpath_n765));
INVX1 mul_U11559(.A(dpath_n765), .Y(n2927));
AND2X1 mul_U11560(.A(dpath_mout[89]), .B(n9767), .Y(dpath_n767));
INVX1 mul_U11561(.A(dpath_n767), .Y(n2928));
AND2X1 mul_U11562(.A(dpath_mout[88]), .B(dpath_n666), .Y(dpath_n769));
INVX1 mul_U11563(.A(dpath_n769), .Y(n2929));
AND2X1 mul_U11564(.A(dpath_mout[87]), .B(dpath_n666), .Y(dpath_n771));
INVX1 mul_U11565(.A(dpath_n771), .Y(n2930));
AND2X1 mul_U11566(.A(dpath_mout[86]), .B(dpath_n666), .Y(dpath_n773));
INVX1 mul_U11567(.A(dpath_n773), .Y(n2931));
AND2X1 mul_U11568(.A(dpath_mout[85]), .B(n9767), .Y(dpath_n775));
INVX1 mul_U11569(.A(dpath_n775), .Y(n2932));
AND2X1 mul_U11570(.A(dpath_mout[84]), .B(n9767), .Y(dpath_n777));
INVX1 mul_U11571(.A(dpath_n777), .Y(n2933));
AND2X1 mul_U11572(.A(dpath_mout[83]), .B(dpath_n666), .Y(dpath_n779));
INVX1 mul_U11573(.A(dpath_n779), .Y(n2934));
AND2X1 mul_U11574(.A(dpath_mout[82]), .B(dpath_n666), .Y(dpath_n781));
INVX1 mul_U11575(.A(dpath_n781), .Y(n2935));
AND2X1 mul_U11576(.A(dpath_n658), .B(dpath_acc_reg[4]), .Y(dpath_n785));
INVX1 mul_U11577(.A(dpath_n785), .Y(n2936));
AND2X1 mul_U11578(.A(n9764), .B(dpath_mout[4]), .Y(dpath_n787));
INVX1 mul_U11579(.A(dpath_n787), .Y(n2937));
AND2X1 mul_U11580(.A(dpath_mout[81]), .B(n9767), .Y(dpath_n789));
INVX1 mul_U11581(.A(dpath_n789), .Y(n2938));
AND2X1 mul_U11582(.A(dpath_mout[80]), .B(dpath_n666), .Y(dpath_n791));
INVX1 mul_U11583(.A(dpath_n791), .Y(n2939));
AND2X1 mul_U11584(.A(dpath_mout[79]), .B(n9767), .Y(dpath_n793));
INVX1 mul_U11585(.A(dpath_n793), .Y(n2940));
AND2X1 mul_U11586(.A(dpath_mout[78]), .B(dpath_n666), .Y(dpath_n795));
INVX1 mul_U11587(.A(dpath_n795), .Y(n2941));
AND2X1 mul_U11588(.A(dpath_mout[77]), .B(n9767), .Y(dpath_n797));
INVX1 mul_U11589(.A(dpath_n797), .Y(n2942));
AND2X1 mul_U11590(.A(dpath_mout[76]), .B(dpath_n666), .Y(dpath_n799));
INVX1 mul_U11591(.A(dpath_n799), .Y(n2943));
AND2X1 mul_U11592(.A(dpath_mout[75]), .B(dpath_n666), .Y(dpath_n801));
INVX1 mul_U11593(.A(dpath_n801), .Y(n2944));
AND2X1 mul_U11594(.A(dpath_mout[74]), .B(dpath_n666), .Y(dpath_n803));
INVX1 mul_U11595(.A(dpath_n803), .Y(n2945));
AND2X1 mul_U11596(.A(dpath_mout[73]), .B(dpath_n666), .Y(dpath_n805));
INVX1 mul_U11597(.A(dpath_n805), .Y(n2946));
AND2X1 mul_U11598(.A(dpath_mout[72]), .B(dpath_n666), .Y(dpath_n807));
INVX1 mul_U11599(.A(dpath_n807), .Y(n2947));
AND2X1 mul_U11600(.A(dpath_n658), .B(dpath_acc_reg[3]), .Y(dpath_n811));
INVX1 mul_U11601(.A(dpath_n811), .Y(n2948));
AND2X1 mul_U11602(.A(n9764), .B(dpath_mout[3]), .Y(dpath_n813));
INVX1 mul_U11603(.A(dpath_n813), .Y(n2949));
AND2X1 mul_U11604(.A(dpath_mout[71]), .B(dpath_n666), .Y(dpath_n815));
INVX1 mul_U11605(.A(dpath_n815), .Y(n2950));
AND2X1 mul_U11606(.A(dpath_mout[70]), .B(dpath_n666), .Y(dpath_n817));
INVX1 mul_U11607(.A(dpath_n817), .Y(n2951));
AND2X1 mul_U11608(.A(dpath_mout[69]), .B(dpath_n666), .Y(dpath_n819));
INVX1 mul_U11609(.A(dpath_n819), .Y(n2952));
AND2X1 mul_U11610(.A(dpath_mout[68]), .B(dpath_n666), .Y(dpath_n821));
INVX1 mul_U11611(.A(dpath_n821), .Y(n2953));
AND2X1 mul_U11612(.A(dpath_mout[67]), .B(dpath_n666), .Y(dpath_n823));
INVX1 mul_U11613(.A(dpath_n823), .Y(n2954));
AND2X1 mul_U11614(.A(dpath_mout[66]), .B(dpath_n666), .Y(dpath_n825));
INVX1 mul_U11615(.A(dpath_n825), .Y(n2955));
AND2X1 mul_U11616(.A(dpath_mout[65]), .B(dpath_n666), .Y(dpath_n827));
INVX1 mul_U11617(.A(dpath_n827), .Y(n2956));
AND2X1 mul_U11618(.A(dpath_mout[64]), .B(dpath_n666), .Y(dpath_n829));
INVX1 mul_U11619(.A(dpath_n829), .Y(n2957));
AND2X1 mul_U11620(.A(dpath_n658), .B(dpath_acc_reg[31]), .Y(dpath_n833));
INVX1 mul_U11621(.A(dpath_n833), .Y(n2958));
AND2X1 mul_U11622(.A(n9764), .B(dpath_mout[31]), .Y(dpath_n835));
INVX1 mul_U11623(.A(dpath_n835), .Y(n2959));
AND2X1 mul_U11624(.A(dpath_n658), .B(dpath_acc_reg[30]), .Y(dpath_n839));
INVX1 mul_U11625(.A(dpath_n839), .Y(n2960));
AND2X1 mul_U11626(.A(n9764), .B(dpath_mout[30]), .Y(dpath_n841));
INVX1 mul_U11627(.A(dpath_n841), .Y(n2961));
AND2X1 mul_U11628(.A(dpath_n658), .B(dpath_acc_reg[2]), .Y(dpath_n845));
INVX1 mul_U11629(.A(dpath_n845), .Y(n2962));
AND2X1 mul_U11630(.A(n9764), .B(dpath_mout[2]), .Y(dpath_n847));
INVX1 mul_U11631(.A(dpath_n847), .Y(n2963));
AND2X1 mul_U11632(.A(dpath_n658), .B(dpath_acc_reg[29]), .Y(dpath_n851));
INVX1 mul_U11633(.A(dpath_n851), .Y(n2964));
AND2X1 mul_U11634(.A(n9764), .B(dpath_mout[29]), .Y(dpath_n853));
INVX1 mul_U11635(.A(dpath_n853), .Y(n2965));
AND2X1 mul_U11636(.A(dpath_n658), .B(dpath_acc_reg[28]), .Y(dpath_n857));
INVX1 mul_U11637(.A(dpath_n857), .Y(n2966));
AND2X1 mul_U11638(.A(n9764), .B(dpath_mout[28]), .Y(dpath_n859));
INVX1 mul_U11639(.A(dpath_n859), .Y(n2967));
AND2X1 mul_U11640(.A(dpath_n658), .B(dpath_acc_reg[27]), .Y(dpath_n863));
INVX1 mul_U11641(.A(dpath_n863), .Y(n2968));
AND2X1 mul_U11642(.A(n9764), .B(dpath_mout[27]), .Y(dpath_n865));
INVX1 mul_U11643(.A(dpath_n865), .Y(n2969));
AND2X1 mul_U11644(.A(dpath_n658), .B(dpath_acc_reg[26]), .Y(dpath_n869));
INVX1 mul_U11645(.A(dpath_n869), .Y(n2970));
AND2X1 mul_U11646(.A(n9764), .B(dpath_mout[26]), .Y(dpath_n871));
INVX1 mul_U11647(.A(dpath_n871), .Y(n2971));
AND2X1 mul_U11648(.A(dpath_n658), .B(dpath_acc_reg[25]), .Y(dpath_n875));
INVX1 mul_U11649(.A(dpath_n875), .Y(n2972));
AND2X1 mul_U11650(.A(n9764), .B(dpath_mout[25]), .Y(dpath_n877));
INVX1 mul_U11651(.A(dpath_n877), .Y(n2973));
AND2X1 mul_U11652(.A(dpath_n658), .B(dpath_acc_reg[24]), .Y(dpath_n881));
INVX1 mul_U11653(.A(dpath_n881), .Y(n2974));
AND2X1 mul_U11654(.A(n9764), .B(dpath_mout[24]), .Y(dpath_n883));
INVX1 mul_U11655(.A(dpath_n883), .Y(n2975));
AND2X1 mul_U11656(.A(dpath_n658), .B(dpath_acc_reg[23]), .Y(dpath_n887));
INVX1 mul_U11657(.A(dpath_n887), .Y(n2976));
AND2X1 mul_U11658(.A(n9764), .B(dpath_mout[23]), .Y(dpath_n889));
INVX1 mul_U11659(.A(dpath_n889), .Y(n2977));
AND2X1 mul_U11660(.A(dpath_n658), .B(dpath_acc_reg[22]), .Y(dpath_n893));
INVX1 mul_U11661(.A(dpath_n893), .Y(n2978));
AND2X1 mul_U11662(.A(n9764), .B(dpath_mout[22]), .Y(dpath_n895));
INVX1 mul_U11663(.A(dpath_n895), .Y(n2979));
AND2X1 mul_U11664(.A(dpath_n658), .B(dpath_acc_reg[21]), .Y(dpath_n899));
INVX1 mul_U11665(.A(dpath_n899), .Y(n2980));
AND2X1 mul_U11666(.A(n9764), .B(dpath_mout[21]), .Y(dpath_n901));
INVX1 mul_U11667(.A(dpath_n901), .Y(n2981));
AND2X1 mul_U11668(.A(dpath_n658), .B(dpath_acc_reg[20]), .Y(dpath_n905));
INVX1 mul_U11669(.A(dpath_n905), .Y(n2982));
AND2X1 mul_U11670(.A(n9764), .B(dpath_mout[20]), .Y(dpath_n907));
INVX1 mul_U11671(.A(dpath_n907), .Y(n2983));
AND2X1 mul_U11672(.A(dpath_n658), .B(dpath_acc_reg[1]), .Y(dpath_n911));
INVX1 mul_U11673(.A(dpath_n911), .Y(n2984));
AND2X1 mul_U11674(.A(n9764), .B(dpath_mout[1]), .Y(dpath_n913));
INVX1 mul_U11675(.A(dpath_n913), .Y(n2985));
AND2X1 mul_U11676(.A(dpath_n658), .B(dpath_acc_reg[19]), .Y(dpath_n917));
INVX1 mul_U11677(.A(dpath_n917), .Y(n2986));
AND2X1 mul_U11678(.A(n9764), .B(dpath_mout[19]), .Y(dpath_n919));
INVX1 mul_U11679(.A(dpath_n919), .Y(n2987));
AND2X1 mul_U11680(.A(dpath_n658), .B(dpath_acc_reg[18]), .Y(dpath_n923));
INVX1 mul_U11681(.A(dpath_n923), .Y(n2988));
AND2X1 mul_U11682(.A(n9764), .B(dpath_mout[18]), .Y(dpath_n925));
INVX1 mul_U11683(.A(dpath_n925), .Y(n2989));
AND2X1 mul_U11684(.A(dpath_n658), .B(dpath_acc_reg[17]), .Y(dpath_n929));
INVX1 mul_U11685(.A(dpath_n929), .Y(n2990));
AND2X1 mul_U11686(.A(n9764), .B(dpath_mout[17]), .Y(dpath_n931));
INVX1 mul_U11687(.A(dpath_n931), .Y(n2991));
AND2X1 mul_U11688(.A(dpath_n658), .B(dpath_acc_reg[16]), .Y(dpath_n935));
INVX1 mul_U11689(.A(dpath_n935), .Y(n2992));
AND2X1 mul_U11690(.A(n9764), .B(dpath_mout[16]), .Y(dpath_n937));
INVX1 mul_U11691(.A(dpath_n937), .Y(n2993));
AND2X1 mul_U11692(.A(dpath_n658), .B(dpath_acc_reg[15]), .Y(dpath_n941));
INVX1 mul_U11693(.A(dpath_n941), .Y(n2994));
AND2X1 mul_U11694(.A(n9764), .B(dpath_mout[15]), .Y(dpath_n943));
INVX1 mul_U11695(.A(dpath_n943), .Y(n2995));
AND2X1 mul_U11696(.A(dpath_n658), .B(dpath_acc_reg[14]), .Y(dpath_n947));
INVX1 mul_U11697(.A(dpath_n947), .Y(n2996));
AND2X1 mul_U11698(.A(n9764), .B(dpath_mout[14]), .Y(dpath_n949));
INVX1 mul_U11699(.A(dpath_n949), .Y(n2997));
AND2X1 mul_U11700(.A(dpath_n658), .B(dpath_acc_reg[13]), .Y(dpath_n953));
INVX1 mul_U11701(.A(dpath_n953), .Y(n2998));
AND2X1 mul_U11702(.A(n9764), .B(dpath_mout[13]), .Y(dpath_n955));
INVX1 mul_U11703(.A(dpath_n955), .Y(n2999));
AND2X1 mul_U11704(.A(dpath_n658), .B(dpath_acc_reg[12]), .Y(dpath_n959));
INVX1 mul_U11705(.A(dpath_n959), .Y(n3000));
AND2X1 mul_U11706(.A(n9764), .B(dpath_mout[12]), .Y(dpath_n961));
INVX1 mul_U11707(.A(dpath_n961), .Y(n3001));
AND2X1 mul_U11708(.A(dpath_n658), .B(dpath_acc_reg[11]), .Y(dpath_n965));
INVX1 mul_U11709(.A(dpath_n965), .Y(n3002));
AND2X1 mul_U11710(.A(n9764), .B(dpath_mout[11]), .Y(dpath_n967));
INVX1 mul_U11711(.A(dpath_n967), .Y(n3003));
AND2X1 mul_U11712(.A(dpath_n658), .B(dpath_acc_reg[10]), .Y(dpath_n971));
INVX1 mul_U11713(.A(dpath_n971), .Y(n3004));
AND2X1 mul_U11714(.A(n9764), .B(dpath_mout[10]), .Y(dpath_n973));
INVX1 mul_U11715(.A(dpath_n973), .Y(n3005));
AND2X1 mul_U11716(.A(dpath_n658), .B(dpath_acc_reg[0]), .Y(dpath_n977));
INVX1 mul_U11717(.A(dpath_n977), .Y(n3006));
AND2X1 mul_U11718(.A(n9764), .B(dpath_mout[0]), .Y(dpath_n981));
INVX1 mul_U11719(.A(dpath_n981), .Y(n3007));
AND2X1 mul_U11720(.A(n5757), .B(n5136), .Y(dpath_acc_reg_in[9]));
INVX1 mul_U11721(.A(dpath_acc_reg_in[9]), .Y(n3008));
AND2X1 mul_U11722(.A(n5758), .B(n5137), .Y(dpath_acc_reg_in[8]));
INVX1 mul_U11723(.A(dpath_acc_reg_in[8]), .Y(n3009));
AND2X1 mul_U11724(.A(n5759), .B(n5138), .Y(dpath_acc_reg_in[7]));
INVX1 mul_U11725(.A(dpath_acc_reg_in[7]), .Y(n3010));
AND2X1 mul_U11726(.A(n5760), .B(n5139), .Y(dpath_acc_reg_in[71]));
INVX1 mul_U11727(.A(dpath_acc_reg_in[71]), .Y(n3011));
AND2X1 mul_U11728(.A(n5761), .B(n5140), .Y(dpath_acc_reg_in[70]));
INVX1 mul_U11729(.A(dpath_acc_reg_in[70]), .Y(n3012));
AND2X1 mul_U11730(.A(n5762), .B(n5141), .Y(dpath_acc_reg_in[6]));
INVX1 mul_U11731(.A(dpath_acc_reg_in[6]), .Y(n3013));
AND2X1 mul_U11732(.A(n5763), .B(n5142), .Y(dpath_acc_reg_in[69]));
INVX1 mul_U11733(.A(dpath_acc_reg_in[69]), .Y(n3014));
AND2X1 mul_U11734(.A(n5764), .B(n5143), .Y(dpath_acc_reg_in[68]));
INVX1 mul_U11735(.A(dpath_acc_reg_in[68]), .Y(n3015));
AND2X1 mul_U11736(.A(n5765), .B(n5144), .Y(dpath_acc_reg_in[67]));
INVX1 mul_U11737(.A(dpath_acc_reg_in[67]), .Y(n3016));
AND2X1 mul_U11738(.A(n5766), .B(n5145), .Y(dpath_acc_reg_in[66]));
INVX1 mul_U11739(.A(dpath_acc_reg_in[66]), .Y(n3017));
AND2X1 mul_U11740(.A(n5767), .B(n5146), .Y(dpath_acc_reg_in[65]));
INVX1 mul_U11741(.A(dpath_acc_reg_in[65]), .Y(n3018));
AND2X1 mul_U11742(.A(n5768), .B(n5147), .Y(dpath_acc_reg_in[64]));
INVX1 mul_U11743(.A(dpath_acc_reg_in[64]), .Y(n3019));
AND2X1 mul_U11744(.A(n5769), .B(n5148), .Y(dpath_acc_reg_in[63]));
INVX1 mul_U11745(.A(dpath_acc_reg_in[63]), .Y(n3020));
AND2X1 mul_U11746(.A(n5770), .B(n5149), .Y(dpath_acc_reg_in[62]));
INVX1 mul_U11747(.A(dpath_acc_reg_in[62]), .Y(n3021));
AND2X1 mul_U11748(.A(n5771), .B(n5150), .Y(dpath_acc_reg_in[61]));
INVX1 mul_U11749(.A(dpath_acc_reg_in[61]), .Y(n3022));
AND2X1 mul_U11750(.A(n5772), .B(n5151), .Y(dpath_acc_reg_in[60]));
INVX1 mul_U11751(.A(dpath_acc_reg_in[60]), .Y(n3023));
AND2X1 mul_U11752(.A(n5773), .B(n5152), .Y(dpath_acc_reg_in[5]));
INVX1 mul_U11753(.A(dpath_acc_reg_in[5]), .Y(n3024));
AND2X1 mul_U11754(.A(n5774), .B(n5153), .Y(dpath_acc_reg_in[59]));
INVX1 mul_U11755(.A(dpath_acc_reg_in[59]), .Y(n3025));
AND2X1 mul_U11756(.A(n5775), .B(n5154), .Y(dpath_acc_reg_in[58]));
INVX1 mul_U11757(.A(dpath_acc_reg_in[58]), .Y(n3026));
AND2X1 mul_U11758(.A(n5776), .B(n5155), .Y(dpath_acc_reg_in[57]));
INVX1 mul_U11759(.A(dpath_acc_reg_in[57]), .Y(n3027));
AND2X1 mul_U11760(.A(n5777), .B(n5156), .Y(dpath_acc_reg_in[56]));
INVX1 mul_U11761(.A(dpath_acc_reg_in[56]), .Y(n3028));
AND2X1 mul_U11762(.A(n5778), .B(n5157), .Y(dpath_acc_reg_in[55]));
INVX1 mul_U11763(.A(dpath_acc_reg_in[55]), .Y(n3029));
AND2X1 mul_U11764(.A(n5779), .B(n5158), .Y(dpath_acc_reg_in[54]));
INVX1 mul_U11765(.A(dpath_acc_reg_in[54]), .Y(n3030));
AND2X1 mul_U11766(.A(n5780), .B(n5159), .Y(dpath_acc_reg_in[53]));
INVX1 mul_U11767(.A(dpath_acc_reg_in[53]), .Y(n3031));
AND2X1 mul_U11768(.A(n5781), .B(n5160), .Y(dpath_acc_reg_in[52]));
INVX1 mul_U11769(.A(dpath_acc_reg_in[52]), .Y(n3032));
AND2X1 mul_U11770(.A(n5782), .B(n5161), .Y(dpath_acc_reg_in[51]));
INVX1 mul_U11771(.A(dpath_acc_reg_in[51]), .Y(n3033));
AND2X1 mul_U11772(.A(n5783), .B(n5162), .Y(dpath_acc_reg_in[50]));
INVX1 mul_U11773(.A(dpath_acc_reg_in[50]), .Y(n3034));
AND2X1 mul_U11774(.A(n5784), .B(n5163), .Y(dpath_acc_reg_in[4]));
INVX1 mul_U11775(.A(dpath_acc_reg_in[4]), .Y(n3035));
AND2X1 mul_U11776(.A(n5785), .B(n5164), .Y(dpath_acc_reg_in[49]));
INVX1 mul_U11777(.A(dpath_acc_reg_in[49]), .Y(n3036));
AND2X1 mul_U11778(.A(n5786), .B(n5165), .Y(dpath_acc_reg_in[48]));
INVX1 mul_U11779(.A(dpath_acc_reg_in[48]), .Y(n3037));
AND2X1 mul_U11780(.A(n5787), .B(n5166), .Y(dpath_acc_reg_in[47]));
INVX1 mul_U11781(.A(dpath_acc_reg_in[47]), .Y(n3038));
AND2X1 mul_U11782(.A(n5788), .B(n5167), .Y(dpath_acc_reg_in[46]));
INVX1 mul_U11783(.A(dpath_acc_reg_in[46]), .Y(n3039));
AND2X1 mul_U11784(.A(n5789), .B(n5168), .Y(dpath_acc_reg_in[45]));
INVX1 mul_U11785(.A(dpath_acc_reg_in[45]), .Y(n3040));
AND2X1 mul_U11786(.A(n5790), .B(n5169), .Y(dpath_acc_reg_in[44]));
INVX1 mul_U11787(.A(dpath_acc_reg_in[44]), .Y(n3041));
AND2X1 mul_U11788(.A(n5791), .B(n5170), .Y(dpath_acc_reg_in[43]));
INVX1 mul_U11789(.A(dpath_acc_reg_in[43]), .Y(n3042));
AND2X1 mul_U11790(.A(n5792), .B(n5171), .Y(dpath_acc_reg_in[42]));
INVX1 mul_U11791(.A(dpath_acc_reg_in[42]), .Y(n3043));
AND2X1 mul_U11792(.A(n5793), .B(n5172), .Y(dpath_acc_reg_in[41]));
INVX1 mul_U11793(.A(dpath_acc_reg_in[41]), .Y(n3044));
AND2X1 mul_U11794(.A(n5794), .B(n5173), .Y(dpath_acc_reg_in[40]));
INVX1 mul_U11795(.A(dpath_acc_reg_in[40]), .Y(n3045));
AND2X1 mul_U11796(.A(n5795), .B(n5174), .Y(dpath_acc_reg_in[3]));
INVX1 mul_U11797(.A(dpath_acc_reg_in[3]), .Y(n3046));
AND2X1 mul_U11798(.A(n5796), .B(n5175), .Y(dpath_acc_reg_in[39]));
INVX1 mul_U11799(.A(dpath_acc_reg_in[39]), .Y(n3047));
AND2X1 mul_U11800(.A(n5797), .B(n5176), .Y(dpath_acc_reg_in[38]));
INVX1 mul_U11801(.A(dpath_acc_reg_in[38]), .Y(n3048));
AND2X1 mul_U11802(.A(n5798), .B(n5177), .Y(dpath_acc_reg_in[37]));
INVX1 mul_U11803(.A(dpath_acc_reg_in[37]), .Y(n3049));
AND2X1 mul_U11804(.A(n5799), .B(n5178), .Y(dpath_acc_reg_in[36]));
INVX1 mul_U11805(.A(dpath_acc_reg_in[36]), .Y(n3050));
AND2X1 mul_U11806(.A(n5800), .B(n5179), .Y(dpath_acc_reg_in[35]));
INVX1 mul_U11807(.A(dpath_acc_reg_in[35]), .Y(n3051));
AND2X1 mul_U11808(.A(n5801), .B(n5180), .Y(dpath_acc_reg_in[34]));
INVX1 mul_U11809(.A(dpath_acc_reg_in[34]), .Y(n3052));
AND2X1 mul_U11810(.A(n5802), .B(n5181), .Y(dpath_acc_reg_in[33]));
INVX1 mul_U11811(.A(dpath_acc_reg_in[33]), .Y(n3053));
AND2X1 mul_U11812(.A(n5803), .B(n5182), .Y(dpath_acc_reg_in[32]));
INVX1 mul_U11813(.A(dpath_acc_reg_in[32]), .Y(n3054));
AND2X1 mul_U11814(.A(n5804), .B(n5183), .Y(dpath_acc_reg_in[31]));
INVX1 mul_U11815(.A(dpath_acc_reg_in[31]), .Y(n3055));
AND2X1 mul_U11816(.A(n5805), .B(n5184), .Y(dpath_acc_reg_in[30]));
INVX1 mul_U11817(.A(dpath_acc_reg_in[30]), .Y(n3056));
AND2X1 mul_U11818(.A(n5806), .B(n5185), .Y(dpath_acc_reg_in[2]));
INVX1 mul_U11819(.A(dpath_acc_reg_in[2]), .Y(n3057));
AND2X1 mul_U11820(.A(n5807), .B(n5186), .Y(dpath_acc_reg_in[29]));
INVX1 mul_U11821(.A(dpath_acc_reg_in[29]), .Y(n3058));
AND2X1 mul_U11822(.A(n5808), .B(n5187), .Y(dpath_acc_reg_in[28]));
INVX1 mul_U11823(.A(dpath_acc_reg_in[28]), .Y(n3059));
AND2X1 mul_U11824(.A(n5809), .B(n5188), .Y(dpath_acc_reg_in[27]));
INVX1 mul_U11825(.A(dpath_acc_reg_in[27]), .Y(n3060));
AND2X1 mul_U11826(.A(n5810), .B(n5189), .Y(dpath_acc_reg_in[26]));
INVX1 mul_U11827(.A(dpath_acc_reg_in[26]), .Y(n3061));
AND2X1 mul_U11828(.A(n5811), .B(n5190), .Y(dpath_acc_reg_in[25]));
INVX1 mul_U11829(.A(dpath_acc_reg_in[25]), .Y(n3062));
AND2X1 mul_U11830(.A(n5812), .B(n5191), .Y(dpath_acc_reg_in[24]));
INVX1 mul_U11831(.A(dpath_acc_reg_in[24]), .Y(n3063));
AND2X1 mul_U11832(.A(n5813), .B(n5192), .Y(dpath_acc_reg_in[23]));
INVX1 mul_U11833(.A(dpath_acc_reg_in[23]), .Y(n3064));
AND2X1 mul_U11834(.A(n5814), .B(n5193), .Y(dpath_acc_reg_in[22]));
INVX1 mul_U11835(.A(dpath_acc_reg_in[22]), .Y(n3065));
AND2X1 mul_U11836(.A(n5815), .B(n5194), .Y(dpath_acc_reg_in[21]));
INVX1 mul_U11837(.A(dpath_acc_reg_in[21]), .Y(n3066));
AND2X1 mul_U11838(.A(n5816), .B(n5195), .Y(dpath_acc_reg_in[20]));
INVX1 mul_U11839(.A(dpath_acc_reg_in[20]), .Y(n3067));
AND2X1 mul_U11840(.A(n5817), .B(n5196), .Y(dpath_acc_reg_in[1]));
INVX1 mul_U11841(.A(dpath_acc_reg_in[1]), .Y(n3068));
AND2X1 mul_U11842(.A(n5818), .B(n5197), .Y(dpath_acc_reg_in[19]));
INVX1 mul_U11843(.A(dpath_acc_reg_in[19]), .Y(n3069));
AND2X1 mul_U11844(.A(n5819), .B(n5198), .Y(dpath_acc_reg_in[18]));
INVX1 mul_U11845(.A(dpath_acc_reg_in[18]), .Y(n3070));
AND2X1 mul_U11846(.A(n5820), .B(n5199), .Y(dpath_acc_reg_in[17]));
INVX1 mul_U11847(.A(dpath_acc_reg_in[17]), .Y(n3071));
AND2X1 mul_U11848(.A(n5821), .B(n5200), .Y(dpath_acc_reg_in[16]));
INVX1 mul_U11849(.A(dpath_acc_reg_in[16]), .Y(n3072));
AND2X1 mul_U11850(.A(n5822), .B(n5201), .Y(dpath_acc_reg_in[15]));
INVX1 mul_U11851(.A(dpath_acc_reg_in[15]), .Y(n3073));
AND2X1 mul_U11852(.A(n5823), .B(n5202), .Y(dpath_acc_reg_in[14]));
INVX1 mul_U11853(.A(dpath_acc_reg_in[14]), .Y(n3074));
AND2X1 mul_U11854(.A(n5824), .B(n5203), .Y(dpath_acc_reg_in[13]));
INVX1 mul_U11855(.A(dpath_acc_reg_in[13]), .Y(n3075));
AND2X1 mul_U11856(.A(n5825), .B(n5204), .Y(dpath_acc_reg_in[12]));
INVX1 mul_U11857(.A(dpath_acc_reg_in[12]), .Y(n3076));
AND2X1 mul_U11858(.A(n5826), .B(n5205), .Y(dpath_acc_reg_in[11]));
INVX1 mul_U11859(.A(dpath_acc_reg_in[11]), .Y(n3077));
AND2X1 mul_U11860(.A(n5827), .B(n5206), .Y(dpath_acc_reg_in[10]));
INVX1 mul_U11861(.A(dpath_acc_reg_in[10]), .Y(n3078));
AND2X1 mul_U11862(.A(n5828), .B(n5207), .Y(dpath_acc_reg_in[0]));
INVX1 mul_U11863(.A(dpath_acc_reg_in[0]), .Y(n3079));
OR2X1 mul_U11864(.A(spu_mul_acc), .B(n9774), .Y(byp_sel));
INVX1 mul_U11865(.A(byp_sel), .Y(n3080));
AND2X1 mul_U11866(.A(control_acc_actc4), .B(acc_actc2), .Y(control_n8));
INVX1 mul_U11867(.A(control_n8), .Y(n3081));
OR2X1 mul_U11868(.A(control_mul_ecl_ack_d), .B(n9815), .Y(control_n11));
INVX1 mul_U11869(.A(control_n11), .Y(n3082));
OR2X1 mul_U11870(.A(n9815), .B(control_acc_actc1), .Y(control_n15));
INVX1 mul_U11871(.A(control_n15), .Y(n3083));
OR2X1 mul_U11872(.A(control_acc_actc4), .B(acc_actc2), .Y(control_n16));
INVX1 mul_U11873(.A(control_n16), .Y(n3084));
AND2X1 mul_U11874(.A(control_n18), .B(n9817), .Y(control_n21));
INVX1 mul_U11875(.A(control_n21), .Y(n3085));
AND2X1 mul_U11876(.A(n9814), .B(n5208), .Y(control_n23));
INVX1 mul_U11877(.A(control_n23), .Y(n3086));
OR2X1 mul_U11878(.A(n5831), .B(n6063), .Y(control_N10));
INVX1 mul_U11879(.A(control_N10), .Y(n3087));
AND2X1 mul_U11880(.A(dpath_mulcore_addin_cout[0]), .B(n10110), .Y(n10111));
INVX1 mul_U11881(.A(n10111), .Y(n3088));
AND2X1 mul_U11882(.A(dpath_mulcore_addin_cout[1]), .B(n10113), .Y(n10114));
INVX1 mul_U11883(.A(n10114), .Y(n3089));
AND2X1 mul_U11884(.A(dpath_mulcore_addin_cout[2]), .B(n10116), .Y(n10117));
INVX1 mul_U11885(.A(n10117), .Y(n3090));
AND2X1 mul_U11886(.A(dpath_mulcore_addin_cout[3]), .B(n10119), .Y(n10120));
INVX1 mul_U11887(.A(n10120), .Y(n3091));
AND2X1 mul_U11888(.A(dpath_mulcore_addin_cout[4]), .B(n10122), .Y(n10123));
INVX1 mul_U11889(.A(n10123), .Y(n3092));
AND2X1 mul_U11890(.A(dpath_mulcore_addin_cout[5]), .B(n10125), .Y(n10126));
INVX1 mul_U11891(.A(n10126), .Y(n3093));
AND2X1 mul_U11892(.A(dpath_mulcore_addin_cout[6]), .B(n10128), .Y(n10129));
INVX1 mul_U11893(.A(n10129), .Y(n3094));
AND2X1 mul_U11894(.A(dpath_mulcore_addin_cout[7]), .B(n10131), .Y(n10132));
INVX1 mul_U11895(.A(n10132), .Y(n3095));
AND2X1 mul_U11896(.A(dpath_mulcore_addin_cout[8]), .B(n10134), .Y(n10135));
INVX1 mul_U11897(.A(n10135), .Y(n3096));
AND2X1 mul_U11898(.A(dpath_mulcore_addin_cout[9]), .B(n10139), .Y(n10140));
INVX1 mul_U11899(.A(n10140), .Y(n3097));
AND2X1 mul_U11900(.A(dpath_mulcore_addin_cout[10]), .B(n10144), .Y(n10145));
INVX1 mul_U11901(.A(n10145), .Y(n3098));
AND2X1 mul_U11902(.A(dpath_mulcore_addin_cout[11]), .B(n10149), .Y(n10150));
INVX1 mul_U11903(.A(n10150), .Y(n3099));
AND2X1 mul_U11904(.A(dpath_mulcore_addin_cout[12]), .B(n10154), .Y(n10155));
INVX1 mul_U11905(.A(n10155), .Y(n3100));
AND2X1 mul_U11906(.A(dpath_mulcore_addin_cout[13]), .B(n10159), .Y(n10160));
INVX1 mul_U11907(.A(n10160), .Y(n3101));
AND2X1 mul_U11908(.A(dpath_mulcore_addin_cout[14]), .B(n10164), .Y(n10165));
INVX1 mul_U11909(.A(n10165), .Y(n3102));
AND2X1 mul_U11910(.A(dpath_mulcore_addin_cout[15]), .B(n10169), .Y(n10170));
INVX1 mul_U11911(.A(n10170), .Y(n3103));
AND2X1 mul_U11912(.A(dpath_mulcore_addin_cout[16]), .B(n10174), .Y(n10175));
INVX1 mul_U11913(.A(n10175), .Y(n3104));
AND2X1 mul_U11914(.A(dpath_mulcore_addin_cout[17]), .B(n10179), .Y(n10180));
INVX1 mul_U11915(.A(n10180), .Y(n3105));
AND2X1 mul_U11916(.A(dpath_mulcore_addin_cout[18]), .B(n10186), .Y(n10187));
INVX1 mul_U11917(.A(n10187), .Y(n3106));
AND2X1 mul_U11918(.A(dpath_mulcore_addin_cout[19]), .B(n10191), .Y(n10192));
INVX1 mul_U11919(.A(n10192), .Y(n3107));
AND2X1 mul_U11920(.A(dpath_mulcore_addin_cout[20]), .B(n10196), .Y(n10197));
INVX1 mul_U11921(.A(n10197), .Y(n3108));
AND2X1 mul_U11922(.A(dpath_mulcore_addin_cout[21]), .B(n10201), .Y(n10202));
INVX1 mul_U11923(.A(n10202), .Y(n3109));
AND2X1 mul_U11924(.A(dpath_mulcore_addin_cout[22]), .B(n10206), .Y(n10207));
INVX1 mul_U11925(.A(n10207), .Y(n3110));
AND2X1 mul_U11926(.A(dpath_mulcore_addin_cout[23]), .B(n10211), .Y(n10212));
INVX1 mul_U11927(.A(n10212), .Y(n3111));
AND2X1 mul_U11928(.A(dpath_mulcore_addin_cout[24]), .B(n10216), .Y(n10217));
INVX1 mul_U11929(.A(n10217), .Y(n3112));
AND2X1 mul_U11930(.A(dpath_mulcore_addin_cout[25]), .B(n10221), .Y(n10222));
INVX1 mul_U11931(.A(n10222), .Y(n3113));
AND2X1 mul_U11932(.A(dpath_mulcore_addin_cout[26]), .B(n10226), .Y(n10227));
INVX1 mul_U11933(.A(n10227), .Y(n3114));
AND2X1 mul_U11934(.A(dpath_mulcore_addin_cout[27]), .B(n10231), .Y(n10232));
INVX1 mul_U11935(.A(n10232), .Y(n3115));
AND2X1 mul_U11936(.A(dpath_mulcore_addin_cout[28]), .B(n10238), .Y(n10239));
INVX1 mul_U11937(.A(n10239), .Y(n3116));
AND2X1 mul_U11938(.A(dpath_mulcore_addin_cout[29]), .B(n10243), .Y(n10244));
INVX1 mul_U11939(.A(n10244), .Y(n3117));
AND2X1 mul_U11940(.A(dpath_mulcore_addin_cout[30]), .B(n10248), .Y(n10249));
INVX1 mul_U11941(.A(n10249), .Y(n3118));
AND2X1 mul_U11942(.A(n9216), .B(n10266), .Y(n10267));
INVX1 mul_U11943(.A(n10267), .Y(n3119));
AND2X1 mul_U11944(.A(dpath_mulcore_addin_cout[32]), .B(n10269), .Y(n10270));
INVX1 mul_U11945(.A(n10270), .Y(n3120));
AND2X1 mul_U11946(.A(dpath_mulcore_addin_cout[33]), .B(n10272), .Y(n10273));
INVX1 mul_U11947(.A(n10273), .Y(n3121));
AND2X1 mul_U11948(.A(dpath_mulcore_addin_cout[34]), .B(n10275), .Y(n10276));
INVX1 mul_U11949(.A(n10276), .Y(n3122));
AND2X1 mul_U11950(.A(dpath_mulcore_addin_cout[35]), .B(n10278), .Y(n10279));
INVX1 mul_U11951(.A(n10279), .Y(n3123));
AND2X1 mul_U11952(.A(dpath_mulcore_addin_cout[36]), .B(n10281), .Y(n10282));
INVX1 mul_U11953(.A(n10282), .Y(n3124));
AND2X1 mul_U11954(.A(dpath_mulcore_addin_cout[37]), .B(n10284), .Y(n10285));
INVX1 mul_U11955(.A(n10285), .Y(n3125));
AND2X1 mul_U11956(.A(dpath_mulcore_addin_cout[38]), .B(n10287), .Y(n10288));
INVX1 mul_U11957(.A(n10288), .Y(n3126));
AND2X1 mul_U11958(.A(dpath_mulcore_addin_cout[39]), .B(n10290), .Y(n10291));
INVX1 mul_U11959(.A(n10291), .Y(n3127));
AND2X1 mul_U11960(.A(dpath_mulcore_addin_cout[40]), .B(n10293), .Y(n10294));
INVX1 mul_U11961(.A(n10294), .Y(n3128));
AND2X1 mul_U11962(.A(dpath_mulcore_addin_cout[41]), .B(n10298), .Y(n10299));
INVX1 mul_U11963(.A(n10299), .Y(n3129));
AND2X1 mul_U11964(.A(dpath_mulcore_addin_cout[42]), .B(n10303), .Y(n10304));
INVX1 mul_U11965(.A(n10304), .Y(n3130));
AND2X1 mul_U11966(.A(dpath_mulcore_addin_cout[43]), .B(n10308), .Y(n10309));
INVX1 mul_U11967(.A(n10309), .Y(n3131));
AND2X1 mul_U11968(.A(dpath_mulcore_addin_cout[44]), .B(n10313), .Y(n10314));
INVX1 mul_U11969(.A(n10314), .Y(n3132));
AND2X1 mul_U11970(.A(dpath_mulcore_addin_cout[45]), .B(n10318), .Y(n10319));
INVX1 mul_U11971(.A(n10319), .Y(n3133));
AND2X1 mul_U11972(.A(dpath_mulcore_addin_cout[46]), .B(n10323), .Y(n10324));
INVX1 mul_U11973(.A(n10324), .Y(n3134));
AND2X1 mul_U11974(.A(dpath_mulcore_addin_cout[47]), .B(n10328), .Y(n10329));
INVX1 mul_U11975(.A(n10329), .Y(n3135));
AND2X1 mul_U11976(.A(dpath_mulcore_addin_cout[48]), .B(n10333), .Y(n10334));
INVX1 mul_U11977(.A(n10334), .Y(n3136));
AND2X1 mul_U11978(.A(dpath_mulcore_addin_cout[49]), .B(n10338), .Y(n10339));
INVX1 mul_U11979(.A(n10339), .Y(n3137));
AND2X1 mul_U11980(.A(dpath_mulcore_addin_cout[50]), .B(n10345), .Y(n10346));
INVX1 mul_U11981(.A(n10346), .Y(n3138));
AND2X1 mul_U11982(.A(dpath_mulcore_addin_cout[51]), .B(n10350), .Y(n10351));
INVX1 mul_U11983(.A(n10351), .Y(n3139));
AND2X1 mul_U11984(.A(dpath_mulcore_addin_cout[52]), .B(n10355), .Y(n10356));
INVX1 mul_U11985(.A(n10356), .Y(n3140));
AND2X1 mul_U11986(.A(dpath_mulcore_addin_cout[53]), .B(n10360), .Y(n10361));
INVX1 mul_U11987(.A(n10361), .Y(n3141));
AND2X1 mul_U11988(.A(dpath_mulcore_addin_cout[54]), .B(n10365), .Y(n10366));
INVX1 mul_U11989(.A(n10366), .Y(n3142));
AND2X1 mul_U11990(.A(dpath_mulcore_addin_cout[55]), .B(n10370), .Y(n10371));
INVX1 mul_U11991(.A(n10371), .Y(n3143));
AND2X1 mul_U11992(.A(dpath_mulcore_addin_cout[56]), .B(n10375), .Y(n10376));
INVX1 mul_U11993(.A(n10376), .Y(n3144));
AND2X1 mul_U11994(.A(dpath_mulcore_addin_cout[57]), .B(n10380), .Y(n10381));
INVX1 mul_U11995(.A(n10381), .Y(n3145));
AND2X1 mul_U11996(.A(dpath_mulcore_addin_cout[58]), .B(n10385), .Y(n10386));
INVX1 mul_U11997(.A(n10386), .Y(n3146));
AND2X1 mul_U11998(.A(dpath_mulcore_addin_cout[59]), .B(n10390), .Y(n10391));
INVX1 mul_U11999(.A(n10391), .Y(n3147));
AND2X1 mul_U12000(.A(dpath_mulcore_addin_cout[60]), .B(n10397), .Y(n10398));
INVX1 mul_U12001(.A(n10398), .Y(n3148));
AND2X1 mul_U12002(.A(dpath_mulcore_addin_cout[61]), .B(n10402), .Y(n10403));
INVX1 mul_U12003(.A(n10403), .Y(n3149));
AND2X1 mul_U12004(.A(dpath_mulcore_addin_cout[62]), .B(n10407), .Y(n10408));
INVX1 mul_U12005(.A(n10408), .Y(n3150));
AND2X1 mul_U12006(.A(dpath_mulcore_addin_cout[63]), .B(n10412), .Y(n10413));
INVX1 mul_U12007(.A(n10413), .Y(n3151));
AND2X1 mul_U12008(.A(dpath_mulcore_addin_cout[64]), .B(n10417), .Y(n10418));
INVX1 mul_U12009(.A(n10418), .Y(n3152));
AND2X1 mul_U12010(.A(dpath_mulcore_addin_cout[65]), .B(n10422), .Y(n10423));
INVX1 mul_U12011(.A(n10423), .Y(n3153));
AND2X1 mul_U12012(.A(dpath_mulcore_addin_cout[66]), .B(n10427), .Y(n10428));
INVX1 mul_U12013(.A(n10428), .Y(n3154));
AND2X1 mul_U12014(.A(dpath_mulcore_addin_cout[67]), .B(n10432), .Y(n10433));
INVX1 mul_U12015(.A(n10433), .Y(n3155));
AND2X1 mul_U12016(.A(dpath_mulcore_addin_cout[68]), .B(n10437), .Y(n10438));
INVX1 mul_U12017(.A(n10438), .Y(n3156));
AND2X1 mul_U12018(.A(dpath_mulcore_addin_cout[69]), .B(n10442), .Y(n10443));
INVX1 mul_U12019(.A(n10443), .Y(n3157));
AND2X1 mul_U12020(.A(dpath_mulcore_addin_cout[70]), .B(n10449), .Y(n10450));
INVX1 mul_U12021(.A(n10450), .Y(n3158));
AND2X1 mul_U12022(.A(dpath_mulcore_addin_cout[71]), .B(n10454), .Y(n10455));
INVX1 mul_U12023(.A(n10455), .Y(n3159));
AND2X1 mul_U12024(.A(dpath_mulcore_addin_cout[72]), .B(n10459), .Y(n10460));
INVX1 mul_U12025(.A(n10460), .Y(n3160));
AND2X1 mul_U12026(.A(dpath_mulcore_addin_cout[73]), .B(n10464), .Y(n10465));
INVX1 mul_U12027(.A(n10465), .Y(n3161));
AND2X1 mul_U12028(.A(dpath_mulcore_addin_cout[74]), .B(n10469), .Y(n10470));
INVX1 mul_U12029(.A(n10470), .Y(n3162));
AND2X1 mul_U12030(.A(dpath_mulcore_addin_cout[75]), .B(n10474), .Y(n10475));
INVX1 mul_U12031(.A(n10475), .Y(n3163));
AND2X1 mul_U12032(.A(dpath_mulcore_addin_cout[76]), .B(n10479), .Y(n10480));
INVX1 mul_U12033(.A(n10480), .Y(n3164));
AND2X1 mul_U12034(.A(dpath_mulcore_addin_cout[77]), .B(n10484), .Y(n10485));
INVX1 mul_U12035(.A(n10485), .Y(n3165));
AND2X1 mul_U12036(.A(dpath_mulcore_addin_cout[78]), .B(n10489), .Y(n10490));
INVX1 mul_U12037(.A(n10490), .Y(n3166));
AND2X1 mul_U12038(.A(dpath_mulcore_addin_cout[79]), .B(n10494), .Y(n10495));
INVX1 mul_U12039(.A(n10495), .Y(n3167));
AND2X1 mul_U12040(.A(dpath_mulcore_addin_cout[80]), .B(n10501), .Y(n10502));
INVX1 mul_U12041(.A(n10502), .Y(n3168));
AND2X1 mul_U12042(.A(dpath_mulcore_addin_cout[81]), .B(n10506), .Y(n10507));
INVX1 mul_U12043(.A(n10507), .Y(n3169));
AND2X1 mul_U12044(.A(dpath_mulcore_addin_cout[82]), .B(n10511), .Y(n10512));
INVX1 mul_U12045(.A(n10512), .Y(n3170));
AND2X1 mul_U12046(.A(dpath_mulcore_addin_cout[83]), .B(n10516), .Y(n10517));
INVX1 mul_U12047(.A(n10517), .Y(n3171));
AND2X1 mul_U12048(.A(dpath_mulcore_addin_cout[84]), .B(n10521), .Y(n10522));
INVX1 mul_U12049(.A(n10522), .Y(n3172));
AND2X1 mul_U12050(.A(dpath_mulcore_addin_cout[85]), .B(n10526), .Y(n10527));
INVX1 mul_U12051(.A(n10527), .Y(n3173));
AND2X1 mul_U12052(.A(dpath_mulcore_addin_cout[86]), .B(n10531), .Y(n10532));
INVX1 mul_U12053(.A(n10532), .Y(n3174));
AND2X1 mul_U12054(.A(dpath_mulcore_addin_cout[87]), .B(n10536), .Y(n10537));
INVX1 mul_U12055(.A(n10537), .Y(n3175));
AND2X1 mul_U12056(.A(dpath_mulcore_addin_cout[88]), .B(n10541), .Y(n10542));
INVX1 mul_U12057(.A(n10542), .Y(n3176));
AND2X1 mul_U12058(.A(dpath_mulcore_addin_cout[89]), .B(n10546), .Y(n10547));
INVX1 mul_U12059(.A(n10547), .Y(n3177));
AND2X1 mul_U12060(.A(dpath_mulcore_addin_cout[90]), .B(n10553), .Y(n10554));
INVX1 mul_U12061(.A(n10554), .Y(n3178));
AND2X1 mul_U12062(.A(dpath_mulcore_addin_cout[91]), .B(n10558), .Y(n10559));
INVX1 mul_U12063(.A(n10559), .Y(n3179));
AND2X1 mul_U12064(.A(dpath_mulcore_addin_cout[92]), .B(n10563), .Y(n10564));
INVX1 mul_U12065(.A(n10564), .Y(n3180));
AND2X1 mul_U12066(.A(dpath_mulcore_addin_cout[93]), .B(n10568), .Y(n10569));
INVX1 mul_U12067(.A(n10569), .Y(n3181));
AND2X1 mul_U12068(.A(dpath_mulcore_addin_cout[94]), .B(n10573), .Y(n10574));
INVX1 mul_U12069(.A(n10574), .Y(n3182));
AND2X1 mul_U12070(.A(dpath_mulcore_addin_cout[95]), .B(n10578), .Y(n10579));
INVX1 mul_U12071(.A(n10579), .Y(n3183));
OR2X1 mul_U12072(.A(n5830), .B(n6056), .Y(n10601));
INVX1 mul_U12073(.A(n10601), .Y(n3184));
AND2X1 mul_U12074(.A(n8055), .B(n13697), .Y(n13695));
INVX1 mul_U12075(.A(n13695), .Y(n3185));
AND2X1 mul_U12076(.A(n8054), .B(n13700), .Y(n13698));
INVX1 mul_U12077(.A(n13698), .Y(n3186));
AND2X1 mul_U12078(.A(n8059), .B(n13708), .Y(n13706));
INVX1 mul_U12079(.A(n13706), .Y(n3187));
AND2X1 mul_U12080(.A(n8058), .B(n13711), .Y(n13709));
INVX1 mul_U12081(.A(n13709), .Y(n3188));
AND2X1 mul_U12082(.A(n8061), .B(n13719), .Y(n13717));
INVX1 mul_U12083(.A(n13717), .Y(n3189));
AND2X1 mul_U12084(.A(n8060), .B(n13722), .Y(n13720));
INVX1 mul_U12085(.A(n13720), .Y(n3190));
AND2X1 mul_U12086(.A(n8063), .B(n13730), .Y(n13728));
INVX1 mul_U12087(.A(n13728), .Y(n3191));
AND2X1 mul_U12088(.A(n8062), .B(n13733), .Y(n13731));
INVX1 mul_U12089(.A(n13731), .Y(n3192));
AND2X1 mul_U12090(.A(n8067), .B(n13741), .Y(n13739));
INVX1 mul_U12091(.A(n13739), .Y(n3193));
AND2X1 mul_U12092(.A(n8066), .B(n13744), .Y(n13742));
INVX1 mul_U12093(.A(n13742), .Y(n3194));
AND2X1 mul_U12094(.A(n7487), .B(n13865), .Y(n13863));
INVX1 mul_U12095(.A(n13863), .Y(n3195));
AND2X1 mul_U12096(.A(n7489), .B(n13868), .Y(n13866));
INVX1 mul_U12097(.A(n13866), .Y(n3196));
AND2X1 mul_U12098(.A(n7491), .B(n13871), .Y(n13869));
INVX1 mul_U12099(.A(n13869), .Y(n3197));
AND2X1 mul_U12100(.A(n7493), .B(n13874), .Y(n13872));
INVX1 mul_U12101(.A(n13872), .Y(n3198));
AND2X1 mul_U12102(.A(n7495), .B(n13877), .Y(n13875));
INVX1 mul_U12103(.A(n13875), .Y(n3199));
AND2X1 mul_U12104(.A(n7497), .B(n13880), .Y(n13878));
INVX1 mul_U12105(.A(n13878), .Y(n3200));
AND2X1 mul_U12106(.A(n7499), .B(n13883), .Y(n13881));
INVX1 mul_U12107(.A(n13881), .Y(n3201));
AND2X1 mul_U12108(.A(n7501), .B(n13886), .Y(n13884));
INVX1 mul_U12109(.A(n13884), .Y(n3202));
AND2X1 mul_U12110(.A(n7503), .B(n13889), .Y(n13887));
INVX1 mul_U12111(.A(n13887), .Y(n3203));
AND2X1 mul_U12112(.A(n7505), .B(n13892), .Y(n13890));
INVX1 mul_U12113(.A(n13890), .Y(n3204));
AND2X1 mul_U12114(.A(n7507), .B(n13895), .Y(n13893));
INVX1 mul_U12115(.A(n13893), .Y(n3205));
AND2X1 mul_U12116(.A(n7509), .B(n13898), .Y(n13896));
INVX1 mul_U12117(.A(n13896), .Y(n3206));
AND2X1 mul_U12118(.A(n7511), .B(n13901), .Y(n13899));
INVX1 mul_U12119(.A(n13899), .Y(n3207));
AND2X1 mul_U12120(.A(n7513), .B(n13904), .Y(n13902));
INVX1 mul_U12121(.A(n13902), .Y(n3208));
AND2X1 mul_U12122(.A(n7515), .B(n13907), .Y(n13905));
INVX1 mul_U12123(.A(n13905), .Y(n3209));
AND2X1 mul_U12124(.A(n7517), .B(n13910), .Y(n13908));
INVX1 mul_U12125(.A(n13908), .Y(n3210));
AND2X1 mul_U12126(.A(n7519), .B(n13913), .Y(n13911));
INVX1 mul_U12127(.A(n13911), .Y(n3211));
AND2X1 mul_U12128(.A(n7521), .B(n13916), .Y(n13914));
INVX1 mul_U12129(.A(n13914), .Y(n3212));
AND2X1 mul_U12130(.A(n7523), .B(n13919), .Y(n13917));
INVX1 mul_U12131(.A(n13917), .Y(n3213));
AND2X1 mul_U12132(.A(n7525), .B(n13922), .Y(n13920));
INVX1 mul_U12133(.A(n13920), .Y(n3214));
AND2X1 mul_U12134(.A(n7527), .B(n13925), .Y(n13923));
INVX1 mul_U12135(.A(n13923), .Y(n3215));
AND2X1 mul_U12136(.A(n7529), .B(n13928), .Y(n13926));
INVX1 mul_U12137(.A(n13926), .Y(n3216));
AND2X1 mul_U12138(.A(n7531), .B(n13931), .Y(n13929));
INVX1 mul_U12139(.A(n13929), .Y(n3217));
AND2X1 mul_U12140(.A(n7533), .B(n13934), .Y(n13932));
INVX1 mul_U12141(.A(n13932), .Y(n3218));
AND2X1 mul_U12142(.A(n7535), .B(n13937), .Y(n13935));
INVX1 mul_U12143(.A(n13935), .Y(n3219));
AND2X1 mul_U12144(.A(n7537), .B(n13940), .Y(n13938));
INVX1 mul_U12145(.A(n13938), .Y(n3220));
AND2X1 mul_U12146(.A(n7539), .B(n13943), .Y(n13941));
INVX1 mul_U12147(.A(n13941), .Y(n3221));
AND2X1 mul_U12148(.A(n7541), .B(n13946), .Y(n13944));
INVX1 mul_U12149(.A(n13944), .Y(n3222));
AND2X1 mul_U12150(.A(n7543), .B(n13949), .Y(n13947));
INVX1 mul_U12151(.A(n13947), .Y(n3223));
AND2X1 mul_U12152(.A(n7545), .B(n13952), .Y(n13950));
INVX1 mul_U12153(.A(n13950), .Y(n3224));
AND2X1 mul_U12154(.A(n7547), .B(n13955), .Y(n13953));
INVX1 mul_U12155(.A(n13953), .Y(n3225));
AND2X1 mul_U12156(.A(n7549), .B(n13958), .Y(n13956));
INVX1 mul_U12157(.A(n13956), .Y(n3226));
AND2X1 mul_U12158(.A(n7551), .B(n13961), .Y(n13959));
INVX1 mul_U12159(.A(n13959), .Y(n3227));
AND2X1 mul_U12160(.A(n7553), .B(n13964), .Y(n13962));
INVX1 mul_U12161(.A(n13962), .Y(n3228));
AND2X1 mul_U12162(.A(n7555), .B(n13967), .Y(n13965));
INVX1 mul_U12163(.A(n13965), .Y(n3229));
AND2X1 mul_U12164(.A(n7557), .B(n13970), .Y(n13968));
INVX1 mul_U12165(.A(n13968), .Y(n3230));
AND2X1 mul_U12166(.A(n7559), .B(n13973), .Y(n13971));
INVX1 mul_U12167(.A(n13971), .Y(n3231));
AND2X1 mul_U12168(.A(n7561), .B(n13976), .Y(n13974));
INVX1 mul_U12169(.A(n13974), .Y(n3232));
AND2X1 mul_U12170(.A(n7563), .B(n13979), .Y(n13977));
INVX1 mul_U12171(.A(n13977), .Y(n3233));
AND2X1 mul_U12172(.A(n7565), .B(n13982), .Y(n13980));
INVX1 mul_U12173(.A(n13980), .Y(n3234));
AND2X1 mul_U12174(.A(n7567), .B(n13985), .Y(n13983));
INVX1 mul_U12175(.A(n13983), .Y(n3235));
AND2X1 mul_U12176(.A(n7569), .B(n13988), .Y(n13986));
INVX1 mul_U12177(.A(n13986), .Y(n3236));
AND2X1 mul_U12178(.A(n7571), .B(n13991), .Y(n13989));
INVX1 mul_U12179(.A(n13989), .Y(n3237));
AND2X1 mul_U12180(.A(n7573), .B(n13994), .Y(n13992));
INVX1 mul_U12181(.A(n13992), .Y(n3238));
AND2X1 mul_U12182(.A(n7575), .B(n13997), .Y(n13995));
INVX1 mul_U12183(.A(n13995), .Y(n3239));
AND2X1 mul_U12184(.A(n7577), .B(n14000), .Y(n13998));
INVX1 mul_U12185(.A(n13998), .Y(n3240));
AND2X1 mul_U12186(.A(n7579), .B(n14003), .Y(n14001));
INVX1 mul_U12187(.A(n14001), .Y(n3241));
AND2X1 mul_U12188(.A(n7581), .B(n14006), .Y(n14004));
INVX1 mul_U12189(.A(n14004), .Y(n3242));
AND2X1 mul_U12190(.A(n7583), .B(n14009), .Y(n14007));
INVX1 mul_U12191(.A(n14007), .Y(n3243));
AND2X1 mul_U12192(.A(n7585), .B(n14012), .Y(n14010));
INVX1 mul_U12193(.A(n14010), .Y(n3244));
AND2X1 mul_U12194(.A(n7587), .B(n14015), .Y(n14013));
INVX1 mul_U12195(.A(n14013), .Y(n3245));
AND2X1 mul_U12196(.A(n7589), .B(n14018), .Y(n14016));
INVX1 mul_U12197(.A(n14016), .Y(n3246));
AND2X1 mul_U12198(.A(n7591), .B(n14021), .Y(n14019));
INVX1 mul_U12199(.A(n14019), .Y(n3247));
AND2X1 mul_U12200(.A(n7593), .B(n14024), .Y(n14022));
INVX1 mul_U12201(.A(n14022), .Y(n3248));
AND2X1 mul_U12202(.A(n7595), .B(n14027), .Y(n14025));
INVX1 mul_U12203(.A(n14025), .Y(n3249));
AND2X1 mul_U12204(.A(n7597), .B(n14030), .Y(n14028));
INVX1 mul_U12205(.A(n14028), .Y(n3250));
AND2X1 mul_U12206(.A(n7599), .B(n14033), .Y(n14031));
INVX1 mul_U12207(.A(n14031), .Y(n3251));
AND2X1 mul_U12208(.A(n7601), .B(n14036), .Y(n14034));
INVX1 mul_U12209(.A(n14034), .Y(n3252));
AND2X1 mul_U12210(.A(n7603), .B(n14039), .Y(n14037));
INVX1 mul_U12211(.A(n14037), .Y(n3253));
AND2X1 mul_U12212(.A(n9848), .B(n14042), .Y(n14040));
INVX1 mul_U12213(.A(n14040), .Y(n3254));
AND2X1 mul_U12214(.A(n7614), .B(n14045), .Y(n14043));
INVX1 mul_U12215(.A(n14043), .Y(n3255));
AND2X1 mul_U12216(.A(n7616), .B(n14048), .Y(n14046));
INVX1 mul_U12217(.A(n14046), .Y(n3256));
AND2X1 mul_U12218(.A(n7618), .B(n14051), .Y(n14049));
INVX1 mul_U12219(.A(n14049), .Y(n3257));
AND2X1 mul_U12220(.A(n7620), .B(n14054), .Y(n14052));
INVX1 mul_U12221(.A(n14052), .Y(n3258));
AND2X1 mul_U12222(.A(n7622), .B(n14057), .Y(n14055));
INVX1 mul_U12223(.A(n14055), .Y(n3259));
AND2X1 mul_U12224(.A(n7624), .B(n14060), .Y(n14058));
INVX1 mul_U12225(.A(n14058), .Y(n3260));
AND2X1 mul_U12226(.A(n7626), .B(n14063), .Y(n14061));
INVX1 mul_U12227(.A(n14061), .Y(n3261));
AND2X1 mul_U12228(.A(n7628), .B(n14066), .Y(n14064));
INVX1 mul_U12229(.A(n14064), .Y(n3262));
AND2X1 mul_U12230(.A(n7630), .B(n14069), .Y(n14067));
INVX1 mul_U12231(.A(n14067), .Y(n3263));
AND2X1 mul_U12232(.A(n7632), .B(n14072), .Y(n14070));
INVX1 mul_U12233(.A(n14070), .Y(n3264));
AND2X1 mul_U12234(.A(n7634), .B(n14075), .Y(n14073));
INVX1 mul_U12235(.A(n14073), .Y(n3265));
AND2X1 mul_U12236(.A(n7636), .B(n14078), .Y(n14076));
INVX1 mul_U12237(.A(n14076), .Y(n3266));
AND2X1 mul_U12238(.A(n7638), .B(n14081), .Y(n14079));
INVX1 mul_U12239(.A(n14079), .Y(n3267));
AND2X1 mul_U12240(.A(n7640), .B(n14084), .Y(n14082));
INVX1 mul_U12241(.A(n14082), .Y(n3268));
AND2X1 mul_U12242(.A(n7642), .B(n14087), .Y(n14085));
INVX1 mul_U12243(.A(n14085), .Y(n3269));
AND2X1 mul_U12244(.A(n7644), .B(n14090), .Y(n14088));
INVX1 mul_U12245(.A(n14088), .Y(n3270));
AND2X1 mul_U12246(.A(n7646), .B(n14093), .Y(n14091));
INVX1 mul_U12247(.A(n14091), .Y(n3271));
AND2X1 mul_U12248(.A(n7648), .B(n14096), .Y(n14094));
INVX1 mul_U12249(.A(n14094), .Y(n3272));
AND2X1 mul_U12250(.A(n7650), .B(n14099), .Y(n14097));
INVX1 mul_U12251(.A(n14097), .Y(n3273));
AND2X1 mul_U12252(.A(n7652), .B(n14102), .Y(n14100));
INVX1 mul_U12253(.A(n14100), .Y(n3274));
AND2X1 mul_U12254(.A(n7654), .B(n14105), .Y(n14103));
INVX1 mul_U12255(.A(n14103), .Y(n3275));
AND2X1 mul_U12256(.A(n7656), .B(n14108), .Y(n14106));
INVX1 mul_U12257(.A(n14106), .Y(n3276));
AND2X1 mul_U12258(.A(n7658), .B(n14111), .Y(n14109));
INVX1 mul_U12259(.A(n14109), .Y(n3277));
AND2X1 mul_U12260(.A(n7660), .B(n14114), .Y(n14112));
INVX1 mul_U12261(.A(n14112), .Y(n3278));
AND2X1 mul_U12262(.A(n7662), .B(n14117), .Y(n14115));
INVX1 mul_U12263(.A(n14115), .Y(n3279));
AND2X1 mul_U12264(.A(n7664), .B(n14120), .Y(n14118));
INVX1 mul_U12265(.A(n14118), .Y(n3280));
AND2X1 mul_U12266(.A(n7666), .B(n14123), .Y(n14121));
INVX1 mul_U12267(.A(n14121), .Y(n3281));
AND2X1 mul_U12268(.A(n7668), .B(n14126), .Y(n14124));
INVX1 mul_U12269(.A(n14124), .Y(n3282));
AND2X1 mul_U12270(.A(n7670), .B(n14129), .Y(n14127));
INVX1 mul_U12271(.A(n14127), .Y(n3283));
AND2X1 mul_U12272(.A(n7672), .B(n14132), .Y(n14130));
INVX1 mul_U12273(.A(n14130), .Y(n3284));
AND2X1 mul_U12274(.A(n7674), .B(n14135), .Y(n14133));
INVX1 mul_U12275(.A(n14133), .Y(n3285));
AND2X1 mul_U12276(.A(n7676), .B(n14138), .Y(n14136));
INVX1 mul_U12277(.A(n14136), .Y(n3286));
AND2X1 mul_U12278(.A(n7678), .B(n14141), .Y(n14139));
INVX1 mul_U12279(.A(n14139), .Y(n3287));
AND2X1 mul_U12280(.A(n7680), .B(n14144), .Y(n14142));
INVX1 mul_U12281(.A(n14142), .Y(n3288));
AND2X1 mul_U12282(.A(n7682), .B(n14147), .Y(n14145));
INVX1 mul_U12283(.A(n14145), .Y(n3289));
AND2X1 mul_U12284(.A(n7684), .B(n14150), .Y(n14148));
INVX1 mul_U12285(.A(n14148), .Y(n3290));
AND2X1 mul_U12286(.A(n7686), .B(n14153), .Y(n14151));
INVX1 mul_U12287(.A(n14151), .Y(n3291));
AND2X1 mul_U12288(.A(n7688), .B(n14156), .Y(n14154));
INVX1 mul_U12289(.A(n14154), .Y(n3292));
AND2X1 mul_U12290(.A(n7690), .B(n14159), .Y(n14157));
INVX1 mul_U12291(.A(n14157), .Y(n3293));
AND2X1 mul_U12292(.A(n7692), .B(n14162), .Y(n14160));
INVX1 mul_U12293(.A(n14160), .Y(n3294));
AND2X1 mul_U12294(.A(n7694), .B(n14165), .Y(n14163));
INVX1 mul_U12295(.A(n14163), .Y(n3295));
AND2X1 mul_U12296(.A(n7696), .B(n14168), .Y(n14166));
INVX1 mul_U12297(.A(n14166), .Y(n3296));
AND2X1 mul_U12298(.A(n7698), .B(n14171), .Y(n14169));
INVX1 mul_U12299(.A(n14169), .Y(n3297));
AND2X1 mul_U12300(.A(n7700), .B(n14174), .Y(n14172));
INVX1 mul_U12301(.A(n14172), .Y(n3298));
AND2X1 mul_U12302(.A(n7702), .B(n14177), .Y(n14175));
INVX1 mul_U12303(.A(n14175), .Y(n3299));
AND2X1 mul_U12304(.A(n7704), .B(n14180), .Y(n14178));
INVX1 mul_U12305(.A(n14178), .Y(n3300));
AND2X1 mul_U12306(.A(n7706), .B(n14183), .Y(n14181));
INVX1 mul_U12307(.A(n14181), .Y(n3301));
AND2X1 mul_U12308(.A(n7708), .B(n14186), .Y(n14184));
INVX1 mul_U12309(.A(n14184), .Y(n3302));
AND2X1 mul_U12310(.A(n7710), .B(n14189), .Y(n14187));
INVX1 mul_U12311(.A(n14187), .Y(n3303));
AND2X1 mul_U12312(.A(n7712), .B(n14192), .Y(n14190));
INVX1 mul_U12313(.A(n14190), .Y(n3304));
AND2X1 mul_U12314(.A(n7714), .B(n14195), .Y(n14193));
INVX1 mul_U12315(.A(n14193), .Y(n3305));
AND2X1 mul_U12316(.A(n7716), .B(n14198), .Y(n14196));
INVX1 mul_U12317(.A(n14196), .Y(n3306));
AND2X1 mul_U12318(.A(n7718), .B(n14201), .Y(n14199));
INVX1 mul_U12319(.A(n14199), .Y(n3307));
AND2X1 mul_U12320(.A(n7720), .B(n14204), .Y(n14202));
INVX1 mul_U12321(.A(n14202), .Y(n3308));
AND2X1 mul_U12322(.A(n7722), .B(n14207), .Y(n14205));
INVX1 mul_U12323(.A(n14205), .Y(n3309));
AND2X1 mul_U12324(.A(n7724), .B(n14210), .Y(n14208));
INVX1 mul_U12325(.A(n14208), .Y(n3310));
AND2X1 mul_U12326(.A(n7726), .B(n14213), .Y(n14211));
INVX1 mul_U12327(.A(n14211), .Y(n3311));
AND2X1 mul_U12328(.A(n7728), .B(n14216), .Y(n14214));
INVX1 mul_U12329(.A(n14214), .Y(n3312));
AND2X1 mul_U12330(.A(n7730), .B(n14219), .Y(n14217));
INVX1 mul_U12331(.A(n14217), .Y(n3313));
AND2X1 mul_U12332(.A(n9842), .B(n14222), .Y(n14220));
INVX1 mul_U12333(.A(n14220), .Y(n3314));
AND2X1 mul_U12334(.A(dpath_mulcore_ary1_a1_I2_p2_l[63]), .B(n14225), .Y(n14223));
INVX1 mul_U12335(.A(n14223), .Y(n3315));
AND2X1 mul_U12336(.A(dpath_mulcore_ary1_a1_I2_p2_l[62]), .B(n14228), .Y(n14226));
INVX1 mul_U12337(.A(n14226), .Y(n3316));
AND2X1 mul_U12338(.A(dpath_mulcore_ary1_a1_I2_p2_l[61]), .B(n14231), .Y(n14229));
INVX1 mul_U12339(.A(n14229), .Y(n3317));
AND2X1 mul_U12340(.A(dpath_mulcore_ary1_a1_I2_p2_l[60]), .B(n14234), .Y(n14232));
INVX1 mul_U12341(.A(n14232), .Y(n3318));
AND2X1 mul_U12342(.A(dpath_mulcore_ary1_a1_I2_p2_l[59]), .B(n14237), .Y(n14235));
INVX1 mul_U12343(.A(n14235), .Y(n3319));
AND2X1 mul_U12344(.A(dpath_mulcore_ary1_a1_I2_p2_l[58]), .B(n14240), .Y(n14238));
INVX1 mul_U12345(.A(n14238), .Y(n3320));
AND2X1 mul_U12346(.A(dpath_mulcore_ary1_a1_I2_p2_l[57]), .B(n14243), .Y(n14241));
INVX1 mul_U12347(.A(n14241), .Y(n3321));
AND2X1 mul_U12348(.A(dpath_mulcore_ary1_a1_I2_p2_l[56]), .B(n14246), .Y(n14244));
INVX1 mul_U12349(.A(n14244), .Y(n3322));
AND2X1 mul_U12350(.A(dpath_mulcore_ary1_a1_I2_p2_l[55]), .B(n14249), .Y(n14247));
INVX1 mul_U12351(.A(n14247), .Y(n3323));
AND2X1 mul_U12352(.A(dpath_mulcore_ary1_a1_I2_p2_l[54]), .B(n14252), .Y(n14250));
INVX1 mul_U12353(.A(n14250), .Y(n3324));
AND2X1 mul_U12354(.A(dpath_mulcore_ary1_a1_I2_p2_l[53]), .B(n14255), .Y(n14253));
INVX1 mul_U12355(.A(n14253), .Y(n3325));
AND2X1 mul_U12356(.A(dpath_mulcore_ary1_a1_I2_p2_l[52]), .B(n14258), .Y(n14256));
INVX1 mul_U12357(.A(n14256), .Y(n3326));
AND2X1 mul_U12358(.A(dpath_mulcore_ary1_a1_I2_p2_l[51]), .B(n14261), .Y(n14259));
INVX1 mul_U12359(.A(n14259), .Y(n3327));
AND2X1 mul_U12360(.A(dpath_mulcore_ary1_a1_I2_p2_l[50]), .B(n14264), .Y(n14262));
INVX1 mul_U12361(.A(n14262), .Y(n3328));
AND2X1 mul_U12362(.A(dpath_mulcore_ary1_a1_I2_p2_l[49]), .B(n14267), .Y(n14265));
INVX1 mul_U12363(.A(n14265), .Y(n3329));
AND2X1 mul_U12364(.A(dpath_mulcore_ary1_a1_I2_p2_l[48]), .B(n14270), .Y(n14268));
INVX1 mul_U12365(.A(n14268), .Y(n3330));
AND2X1 mul_U12366(.A(dpath_mulcore_ary1_a1_I2_p2_l[47]), .B(n14273), .Y(n14271));
INVX1 mul_U12367(.A(n14271), .Y(n3331));
AND2X1 mul_U12368(.A(dpath_mulcore_ary1_a1_I2_p2_l[46]), .B(n14276), .Y(n14274));
INVX1 mul_U12369(.A(n14274), .Y(n3332));
AND2X1 mul_U12370(.A(dpath_mulcore_ary1_a1_I2_p2_l[45]), .B(n14279), .Y(n14277));
INVX1 mul_U12371(.A(n14277), .Y(n3333));
AND2X1 mul_U12372(.A(dpath_mulcore_ary1_a1_I2_p2_l[44]), .B(n14282), .Y(n14280));
INVX1 mul_U12373(.A(n14280), .Y(n3334));
AND2X1 mul_U12374(.A(dpath_mulcore_ary1_a1_I2_p2_l[43]), .B(n14285), .Y(n14283));
INVX1 mul_U12375(.A(n14283), .Y(n3335));
AND2X1 mul_U12376(.A(dpath_mulcore_ary1_a1_I2_p2_l[42]), .B(n14288), .Y(n14286));
INVX1 mul_U12377(.A(n14286), .Y(n3336));
AND2X1 mul_U12378(.A(dpath_mulcore_ary1_a1_I2_p2_l[41]), .B(n14291), .Y(n14289));
INVX1 mul_U12379(.A(n14289), .Y(n3337));
AND2X1 mul_U12380(.A(dpath_mulcore_ary1_a1_I2_p2_l[40]), .B(n14294), .Y(n14292));
INVX1 mul_U12381(.A(n14292), .Y(n3338));
AND2X1 mul_U12382(.A(dpath_mulcore_ary1_a1_I2_p2_l[39]), .B(n14297), .Y(n14295));
INVX1 mul_U12383(.A(n14295), .Y(n3339));
AND2X1 mul_U12384(.A(dpath_mulcore_ary1_a1_I2_p2_l[38]), .B(n14300), .Y(n14298));
INVX1 mul_U12385(.A(n14298), .Y(n3340));
AND2X1 mul_U12386(.A(dpath_mulcore_ary1_a1_I2_p2_l[37]), .B(n14303), .Y(n14301));
INVX1 mul_U12387(.A(n14301), .Y(n3341));
AND2X1 mul_U12388(.A(dpath_mulcore_ary1_a1_I2_p2_l[36]), .B(n14306), .Y(n14304));
INVX1 mul_U12389(.A(n14304), .Y(n3342));
AND2X1 mul_U12390(.A(dpath_mulcore_ary1_a1_I2_p2_l[35]), .B(n14309), .Y(n14307));
INVX1 mul_U12391(.A(n14307), .Y(n3343));
AND2X1 mul_U12392(.A(dpath_mulcore_ary1_a1_I2_p2_l[34]), .B(n14312), .Y(n14310));
INVX1 mul_U12393(.A(n14310), .Y(n3344));
AND2X1 mul_U12394(.A(dpath_mulcore_ary1_a1_I2_p2_l[33]), .B(n14315), .Y(n14313));
INVX1 mul_U12395(.A(n14313), .Y(n3345));
AND2X1 mul_U12396(.A(dpath_mulcore_ary1_a1_I2_p2_l[32]), .B(n14318), .Y(n14316));
INVX1 mul_U12397(.A(n14316), .Y(n3346));
AND2X1 mul_U12398(.A(dpath_mulcore_ary1_a1_I2_p2_l[31]), .B(n14321), .Y(n14319));
INVX1 mul_U12399(.A(n14319), .Y(n3347));
AND2X1 mul_U12400(.A(dpath_mulcore_ary1_a1_I2_p2_l[30]), .B(n14324), .Y(n14322));
INVX1 mul_U12401(.A(n14322), .Y(n3348));
AND2X1 mul_U12402(.A(dpath_mulcore_ary1_a1_I2_p2_l[29]), .B(n14327), .Y(n14325));
INVX1 mul_U12403(.A(n14325), .Y(n3349));
AND2X1 mul_U12404(.A(dpath_mulcore_ary1_a1_I2_p2_l[28]), .B(n14330), .Y(n14328));
INVX1 mul_U12405(.A(n14328), .Y(n3350));
AND2X1 mul_U12406(.A(dpath_mulcore_ary1_a1_I2_p2_l[27]), .B(n14333), .Y(n14331));
INVX1 mul_U12407(.A(n14331), .Y(n3351));
AND2X1 mul_U12408(.A(dpath_mulcore_ary1_a1_I2_p2_l[26]), .B(n14336), .Y(n14334));
INVX1 mul_U12409(.A(n14334), .Y(n3352));
AND2X1 mul_U12410(.A(dpath_mulcore_ary1_a1_I2_p2_l[25]), .B(n14339), .Y(n14337));
INVX1 mul_U12411(.A(n14337), .Y(n3353));
AND2X1 mul_U12412(.A(dpath_mulcore_ary1_a1_I2_p2_l[24]), .B(n14342), .Y(n14340));
INVX1 mul_U12413(.A(n14340), .Y(n3354));
AND2X1 mul_U12414(.A(dpath_mulcore_ary1_a1_I2_p2_l[23]), .B(n14345), .Y(n14343));
INVX1 mul_U12415(.A(n14343), .Y(n3355));
AND2X1 mul_U12416(.A(dpath_mulcore_ary1_a1_I2_p2_l[22]), .B(n14348), .Y(n14346));
INVX1 mul_U12417(.A(n14346), .Y(n3356));
AND2X1 mul_U12418(.A(dpath_mulcore_ary1_a1_I2_p2_l[21]), .B(n14351), .Y(n14349));
INVX1 mul_U12419(.A(n14349), .Y(n3357));
AND2X1 mul_U12420(.A(dpath_mulcore_ary1_a1_I2_p2_l[20]), .B(n14354), .Y(n14352));
INVX1 mul_U12421(.A(n14352), .Y(n3358));
AND2X1 mul_U12422(.A(dpath_mulcore_ary1_a1_I2_p2_l[19]), .B(n14357), .Y(n14355));
INVX1 mul_U12423(.A(n14355), .Y(n3359));
AND2X1 mul_U12424(.A(dpath_mulcore_ary1_a1_I2_p2_l[18]), .B(n14360), .Y(n14358));
INVX1 mul_U12425(.A(n14358), .Y(n3360));
AND2X1 mul_U12426(.A(dpath_mulcore_ary1_a1_I2_p2_l[17]), .B(n14363), .Y(n14361));
INVX1 mul_U12427(.A(n14361), .Y(n3361));
AND2X1 mul_U12428(.A(dpath_mulcore_ary1_a1_I2_p2_l[16]), .B(n14366), .Y(n14364));
INVX1 mul_U12429(.A(n14364), .Y(n3362));
AND2X1 mul_U12430(.A(dpath_mulcore_ary1_a1_I2_p2_l[15]), .B(n14369), .Y(n14367));
INVX1 mul_U12431(.A(n14367), .Y(n3363));
AND2X1 mul_U12432(.A(dpath_mulcore_ary1_a1_I2_p2_l[14]), .B(n14372), .Y(n14370));
INVX1 mul_U12433(.A(n14370), .Y(n3364));
AND2X1 mul_U12434(.A(dpath_mulcore_ary1_a1_I2_p2_l[13]), .B(n14375), .Y(n14373));
INVX1 mul_U12435(.A(n14373), .Y(n3365));
AND2X1 mul_U12436(.A(dpath_mulcore_ary1_a1_I2_p2_l[12]), .B(n14378), .Y(n14376));
INVX1 mul_U12437(.A(n14376), .Y(n3366));
AND2X1 mul_U12438(.A(dpath_mulcore_ary1_a1_I2_p2_l[11]), .B(n14381), .Y(n14379));
INVX1 mul_U12439(.A(n14379), .Y(n3367));
AND2X1 mul_U12440(.A(dpath_mulcore_ary1_a1_I2_p2_l[10]), .B(n14384), .Y(n14382));
INVX1 mul_U12441(.A(n14382), .Y(n3368));
AND2X1 mul_U12442(.A(dpath_mulcore_ary1_a1_I2_p2_l[9]), .B(n14387), .Y(n14385));
INVX1 mul_U12443(.A(n14385), .Y(n3369));
AND2X1 mul_U12444(.A(dpath_mulcore_ary1_a1_I2_p2_l[8]), .B(n14390), .Y(n14388));
INVX1 mul_U12445(.A(n14388), .Y(n3370));
AND2X1 mul_U12446(.A(dpath_mulcore_ary1_a1_I2_p2_l[7]), .B(n14393), .Y(n14391));
INVX1 mul_U12447(.A(n14391), .Y(n3371));
AND2X1 mul_U12448(.A(dpath_mulcore_ary1_a1_I2_p2_l[6]), .B(n14396), .Y(n14394));
INVX1 mul_U12449(.A(n14394), .Y(n3372));
AND2X1 mul_U12450(.A(dpath_mulcore_ary1_a1_I2_p2_l[5]), .B(n14399), .Y(n14397));
INVX1 mul_U12451(.A(n14397), .Y(n3373));
AND2X1 mul_U12452(.A(dpath_mulcore_ary1_a1_I2_p2_l[4]), .B(n14402), .Y(n14400));
INVX1 mul_U12453(.A(n14400), .Y(n3374));
AND2X1 mul_U12454(.A(n7805), .B(n14405), .Y(n14403));
INVX1 mul_U12455(.A(n14403), .Y(n3375));
AND2X1 mul_U12456(.A(n7807), .B(n14408), .Y(n14406));
INVX1 mul_U12457(.A(n14406), .Y(n3376));
AND2X1 mul_U12458(.A(n7809), .B(n14411), .Y(n14409));
INVX1 mul_U12459(.A(n14409), .Y(n3377));
AND2X1 mul_U12460(.A(n7811), .B(n14414), .Y(n14412));
INVX1 mul_U12461(.A(n14412), .Y(n3378));
AND2X1 mul_U12462(.A(n7813), .B(n14417), .Y(n14415));
INVX1 mul_U12463(.A(n14415), .Y(n3379));
AND2X1 mul_U12464(.A(n7815), .B(n14420), .Y(n14418));
INVX1 mul_U12465(.A(n14418), .Y(n3380));
AND2X1 mul_U12466(.A(n7817), .B(n14423), .Y(n14421));
INVX1 mul_U12467(.A(n14421), .Y(n3381));
AND2X1 mul_U12468(.A(n7819), .B(n14426), .Y(n14424));
INVX1 mul_U12469(.A(n14424), .Y(n3382));
AND2X1 mul_U12470(.A(n7821), .B(n14429), .Y(n14427));
INVX1 mul_U12471(.A(n14427), .Y(n3383));
AND2X1 mul_U12472(.A(n7823), .B(n14432), .Y(n14430));
INVX1 mul_U12473(.A(n14430), .Y(n3384));
AND2X1 mul_U12474(.A(n7825), .B(n14435), .Y(n14433));
INVX1 mul_U12475(.A(n14433), .Y(n3385));
AND2X1 mul_U12476(.A(n7827), .B(n14438), .Y(n14436));
INVX1 mul_U12477(.A(n14436), .Y(n3386));
AND2X1 mul_U12478(.A(n7829), .B(n14441), .Y(n14439));
INVX1 mul_U12479(.A(n14439), .Y(n3387));
AND2X1 mul_U12480(.A(n7831), .B(n14444), .Y(n14442));
INVX1 mul_U12481(.A(n14442), .Y(n3388));
AND2X1 mul_U12482(.A(n7833), .B(n14447), .Y(n14445));
INVX1 mul_U12483(.A(n14445), .Y(n3389));
AND2X1 mul_U12484(.A(n7835), .B(n14450), .Y(n14448));
INVX1 mul_U12485(.A(n14448), .Y(n3390));
AND2X1 mul_U12486(.A(n7837), .B(n14453), .Y(n14451));
INVX1 mul_U12487(.A(n14451), .Y(n3391));
AND2X1 mul_U12488(.A(n7839), .B(n14456), .Y(n14454));
INVX1 mul_U12489(.A(n14454), .Y(n3392));
AND2X1 mul_U12490(.A(n7841), .B(n14459), .Y(n14457));
INVX1 mul_U12491(.A(n14457), .Y(n3393));
AND2X1 mul_U12492(.A(n7843), .B(n14462), .Y(n14460));
INVX1 mul_U12493(.A(n14460), .Y(n3394));
AND2X1 mul_U12494(.A(n7845), .B(n14465), .Y(n14463));
INVX1 mul_U12495(.A(n14463), .Y(n3395));
AND2X1 mul_U12496(.A(n7847), .B(n14468), .Y(n14466));
INVX1 mul_U12497(.A(n14466), .Y(n3396));
AND2X1 mul_U12498(.A(n7849), .B(n14471), .Y(n14469));
INVX1 mul_U12499(.A(n14469), .Y(n3397));
AND2X1 mul_U12500(.A(n7851), .B(n14474), .Y(n14472));
INVX1 mul_U12501(.A(n14472), .Y(n3398));
AND2X1 mul_U12502(.A(n7853), .B(n14477), .Y(n14475));
INVX1 mul_U12503(.A(n14475), .Y(n3399));
AND2X1 mul_U12504(.A(n7855), .B(n14480), .Y(n14478));
INVX1 mul_U12505(.A(n14478), .Y(n3400));
AND2X1 mul_U12506(.A(n7857), .B(n14483), .Y(n14481));
INVX1 mul_U12507(.A(n14481), .Y(n3401));
AND2X1 mul_U12508(.A(n7859), .B(n14486), .Y(n14484));
INVX1 mul_U12509(.A(n14484), .Y(n3402));
AND2X1 mul_U12510(.A(n7861), .B(n14489), .Y(n14487));
INVX1 mul_U12511(.A(n14487), .Y(n3403));
AND2X1 mul_U12512(.A(n7863), .B(n14492), .Y(n14490));
INVX1 mul_U12513(.A(n14490), .Y(n3404));
AND2X1 mul_U12514(.A(n7865), .B(n14495), .Y(n14493));
INVX1 mul_U12515(.A(n14493), .Y(n3405));
AND2X1 mul_U12516(.A(n7867), .B(n14498), .Y(n14496));
INVX1 mul_U12517(.A(n14496), .Y(n3406));
AND2X1 mul_U12518(.A(n7869), .B(n14501), .Y(n14499));
INVX1 mul_U12519(.A(n14499), .Y(n3407));
AND2X1 mul_U12520(.A(n7871), .B(n14504), .Y(n14502));
INVX1 mul_U12521(.A(n14502), .Y(n3408));
AND2X1 mul_U12522(.A(n7873), .B(n14507), .Y(n14505));
INVX1 mul_U12523(.A(n14505), .Y(n3409));
AND2X1 mul_U12524(.A(n7875), .B(n14510), .Y(n14508));
INVX1 mul_U12525(.A(n14508), .Y(n3410));
AND2X1 mul_U12526(.A(n7877), .B(n14513), .Y(n14511));
INVX1 mul_U12527(.A(n14511), .Y(n3411));
AND2X1 mul_U12528(.A(n7879), .B(n14516), .Y(n14514));
INVX1 mul_U12529(.A(n14514), .Y(n3412));
AND2X1 mul_U12530(.A(n7881), .B(n14519), .Y(n14517));
INVX1 mul_U12531(.A(n14517), .Y(n3413));
AND2X1 mul_U12532(.A(n7883), .B(n14522), .Y(n14520));
INVX1 mul_U12533(.A(n14520), .Y(n3414));
AND2X1 mul_U12534(.A(n7885), .B(n14525), .Y(n14523));
INVX1 mul_U12535(.A(n14523), .Y(n3415));
AND2X1 mul_U12536(.A(n7887), .B(n14528), .Y(n14526));
INVX1 mul_U12537(.A(n14526), .Y(n3416));
AND2X1 mul_U12538(.A(n7889), .B(n14531), .Y(n14529));
INVX1 mul_U12539(.A(n14529), .Y(n3417));
AND2X1 mul_U12540(.A(n7891), .B(n14534), .Y(n14532));
INVX1 mul_U12541(.A(n14532), .Y(n3418));
AND2X1 mul_U12542(.A(n7893), .B(n14537), .Y(n14535));
INVX1 mul_U12543(.A(n14535), .Y(n3419));
AND2X1 mul_U12544(.A(n7895), .B(n14540), .Y(n14538));
INVX1 mul_U12545(.A(n14538), .Y(n3420));
AND2X1 mul_U12546(.A(n7897), .B(n14543), .Y(n14541));
INVX1 mul_U12547(.A(n14541), .Y(n3421));
AND2X1 mul_U12548(.A(n7899), .B(n14546), .Y(n14544));
INVX1 mul_U12549(.A(n14544), .Y(n3422));
AND2X1 mul_U12550(.A(n7901), .B(n14549), .Y(n14547));
INVX1 mul_U12551(.A(n14547), .Y(n3423));
AND2X1 mul_U12552(.A(n7903), .B(n14552), .Y(n14550));
INVX1 mul_U12553(.A(n14550), .Y(n3424));
AND2X1 mul_U12554(.A(n7905), .B(n14555), .Y(n14553));
INVX1 mul_U12555(.A(n14553), .Y(n3425));
AND2X1 mul_U12556(.A(n7907), .B(n14558), .Y(n14556));
INVX1 mul_U12557(.A(n14556), .Y(n3426));
AND2X1 mul_U12558(.A(n7909), .B(n14561), .Y(n14559));
INVX1 mul_U12559(.A(n14559), .Y(n3427));
AND2X1 mul_U12560(.A(n7911), .B(n14564), .Y(n14562));
INVX1 mul_U12561(.A(n14562), .Y(n3428));
AND2X1 mul_U12562(.A(n7913), .B(n14567), .Y(n14565));
INVX1 mul_U12563(.A(n14565), .Y(n3429));
AND2X1 mul_U12564(.A(n7915), .B(n14570), .Y(n14568));
INVX1 mul_U12565(.A(n14568), .Y(n3430));
AND2X1 mul_U12566(.A(n7917), .B(n14573), .Y(n14571));
INVX1 mul_U12567(.A(n14571), .Y(n3431));
AND2X1 mul_U12568(.A(n7919), .B(n14576), .Y(n14574));
INVX1 mul_U12569(.A(n14574), .Y(n3432));
AND2X1 mul_U12570(.A(n7921), .B(n14579), .Y(n14577));
INVX1 mul_U12571(.A(n14577), .Y(n3433));
AND2X1 mul_U12572(.A(n9835), .B(n14582), .Y(n14580));
INVX1 mul_U12573(.A(n14580), .Y(n3434));
AND2X1 mul_U12574(.A(n7932), .B(n14585), .Y(n14583));
INVX1 mul_U12575(.A(n14583), .Y(n3435));
AND2X1 mul_U12576(.A(n7934), .B(n14588), .Y(n14586));
INVX1 mul_U12577(.A(n14586), .Y(n3436));
AND2X1 mul_U12578(.A(n7936), .B(n14591), .Y(n14589));
INVX1 mul_U12579(.A(n14589), .Y(n3437));
AND2X1 mul_U12580(.A(n7938), .B(n14594), .Y(n14592));
INVX1 mul_U12581(.A(n14592), .Y(n3438));
AND2X1 mul_U12582(.A(n7940), .B(n14597), .Y(n14595));
INVX1 mul_U12583(.A(n14595), .Y(n3439));
AND2X1 mul_U12584(.A(n7942), .B(n14600), .Y(n14598));
INVX1 mul_U12585(.A(n14598), .Y(n3440));
AND2X1 mul_U12586(.A(n7944), .B(n14603), .Y(n14601));
INVX1 mul_U12587(.A(n14601), .Y(n3441));
AND2X1 mul_U12588(.A(n7946), .B(n14606), .Y(n14604));
INVX1 mul_U12589(.A(n14604), .Y(n3442));
AND2X1 mul_U12590(.A(n7948), .B(n14609), .Y(n14607));
INVX1 mul_U12591(.A(n14607), .Y(n3443));
AND2X1 mul_U12592(.A(n7950), .B(n14612), .Y(n14610));
INVX1 mul_U12593(.A(n14610), .Y(n3444));
AND2X1 mul_U12594(.A(n7952), .B(n14615), .Y(n14613));
INVX1 mul_U12595(.A(n14613), .Y(n3445));
AND2X1 mul_U12596(.A(n7954), .B(n14618), .Y(n14616));
INVX1 mul_U12597(.A(n14616), .Y(n3446));
AND2X1 mul_U12598(.A(n7956), .B(n14621), .Y(n14619));
INVX1 mul_U12599(.A(n14619), .Y(n3447));
AND2X1 mul_U12600(.A(n7958), .B(n14624), .Y(n14622));
INVX1 mul_U12601(.A(n14622), .Y(n3448));
AND2X1 mul_U12602(.A(n7960), .B(n14627), .Y(n14625));
INVX1 mul_U12603(.A(n14625), .Y(n3449));
AND2X1 mul_U12604(.A(n7962), .B(n14630), .Y(n14628));
INVX1 mul_U12605(.A(n14628), .Y(n3450));
AND2X1 mul_U12606(.A(n7964), .B(n14633), .Y(n14631));
INVX1 mul_U12607(.A(n14631), .Y(n3451));
AND2X1 mul_U12608(.A(n7966), .B(n14636), .Y(n14634));
INVX1 mul_U12609(.A(n14634), .Y(n3452));
AND2X1 mul_U12610(.A(n7968), .B(n14639), .Y(n14637));
INVX1 mul_U12611(.A(n14637), .Y(n3453));
AND2X1 mul_U12612(.A(n7970), .B(n14642), .Y(n14640));
INVX1 mul_U12613(.A(n14640), .Y(n3454));
AND2X1 mul_U12614(.A(n7972), .B(n14645), .Y(n14643));
INVX1 mul_U12615(.A(n14643), .Y(n3455));
AND2X1 mul_U12616(.A(n7974), .B(n14648), .Y(n14646));
INVX1 mul_U12617(.A(n14646), .Y(n3456));
AND2X1 mul_U12618(.A(n7976), .B(n14651), .Y(n14649));
INVX1 mul_U12619(.A(n14649), .Y(n3457));
AND2X1 mul_U12620(.A(n7978), .B(n14654), .Y(n14652));
INVX1 mul_U12621(.A(n14652), .Y(n3458));
AND2X1 mul_U12622(.A(n7980), .B(n14657), .Y(n14655));
INVX1 mul_U12623(.A(n14655), .Y(n3459));
AND2X1 mul_U12624(.A(n7982), .B(n14660), .Y(n14658));
INVX1 mul_U12625(.A(n14658), .Y(n3460));
AND2X1 mul_U12626(.A(n7984), .B(n14663), .Y(n14661));
INVX1 mul_U12627(.A(n14661), .Y(n3461));
AND2X1 mul_U12628(.A(n7986), .B(n14666), .Y(n14664));
INVX1 mul_U12629(.A(n14664), .Y(n3462));
AND2X1 mul_U12630(.A(n7988), .B(n14669), .Y(n14667));
INVX1 mul_U12631(.A(n14667), .Y(n3463));
AND2X1 mul_U12632(.A(n7990), .B(n14672), .Y(n14670));
INVX1 mul_U12633(.A(n14670), .Y(n3464));
AND2X1 mul_U12634(.A(n7992), .B(n14675), .Y(n14673));
INVX1 mul_U12635(.A(n14673), .Y(n3465));
AND2X1 mul_U12636(.A(n7994), .B(n14678), .Y(n14676));
INVX1 mul_U12637(.A(n14676), .Y(n3466));
AND2X1 mul_U12638(.A(n7996), .B(n14681), .Y(n14679));
INVX1 mul_U12639(.A(n14679), .Y(n3467));
AND2X1 mul_U12640(.A(n7998), .B(n14684), .Y(n14682));
INVX1 mul_U12641(.A(n14682), .Y(n3468));
AND2X1 mul_U12642(.A(n8000), .B(n14687), .Y(n14685));
INVX1 mul_U12643(.A(n14685), .Y(n3469));
AND2X1 mul_U12644(.A(n8002), .B(n14690), .Y(n14688));
INVX1 mul_U12645(.A(n14688), .Y(n3470));
AND2X1 mul_U12646(.A(n8004), .B(n14693), .Y(n14691));
INVX1 mul_U12647(.A(n14691), .Y(n3471));
AND2X1 mul_U12648(.A(n8006), .B(n14696), .Y(n14694));
INVX1 mul_U12649(.A(n14694), .Y(n3472));
AND2X1 mul_U12650(.A(n8008), .B(n14699), .Y(n14697));
INVX1 mul_U12651(.A(n14697), .Y(n3473));
AND2X1 mul_U12652(.A(n8010), .B(n14702), .Y(n14700));
INVX1 mul_U12653(.A(n14700), .Y(n3474));
AND2X1 mul_U12654(.A(n8012), .B(n14705), .Y(n14703));
INVX1 mul_U12655(.A(n14703), .Y(n3475));
AND2X1 mul_U12656(.A(n8014), .B(n14708), .Y(n14706));
INVX1 mul_U12657(.A(n14706), .Y(n3476));
AND2X1 mul_U12658(.A(n8016), .B(n14711), .Y(n14709));
INVX1 mul_U12659(.A(n14709), .Y(n3477));
AND2X1 mul_U12660(.A(n8018), .B(n14714), .Y(n14712));
INVX1 mul_U12661(.A(n14712), .Y(n3478));
AND2X1 mul_U12662(.A(n8020), .B(n14717), .Y(n14715));
INVX1 mul_U12663(.A(n14715), .Y(n3479));
AND2X1 mul_U12664(.A(n8022), .B(n14720), .Y(n14718));
INVX1 mul_U12665(.A(n14718), .Y(n3480));
AND2X1 mul_U12666(.A(n8024), .B(n14723), .Y(n14721));
INVX1 mul_U12667(.A(n14721), .Y(n3481));
AND2X1 mul_U12668(.A(n8026), .B(n14726), .Y(n14724));
INVX1 mul_U12669(.A(n14724), .Y(n3482));
AND2X1 mul_U12670(.A(n8028), .B(n14729), .Y(n14727));
INVX1 mul_U12671(.A(n14727), .Y(n3483));
AND2X1 mul_U12672(.A(n8030), .B(n14732), .Y(n14730));
INVX1 mul_U12673(.A(n14730), .Y(n3484));
AND2X1 mul_U12674(.A(n8032), .B(n14735), .Y(n14733));
INVX1 mul_U12675(.A(n14733), .Y(n3485));
AND2X1 mul_U12676(.A(n8034), .B(n14738), .Y(n14736));
INVX1 mul_U12677(.A(n14736), .Y(n3486));
AND2X1 mul_U12678(.A(n8036), .B(n14741), .Y(n14739));
INVX1 mul_U12679(.A(n14739), .Y(n3487));
AND2X1 mul_U12680(.A(n8038), .B(n14744), .Y(n14742));
INVX1 mul_U12681(.A(n14742), .Y(n3488));
AND2X1 mul_U12682(.A(n8040), .B(n14747), .Y(n14745));
INVX1 mul_U12683(.A(n14745), .Y(n3489));
AND2X1 mul_U12684(.A(n8042), .B(n14750), .Y(n14748));
INVX1 mul_U12685(.A(n14748), .Y(n3490));
AND2X1 mul_U12686(.A(n8044), .B(n14753), .Y(n14751));
INVX1 mul_U12687(.A(n14751), .Y(n3491));
AND2X1 mul_U12688(.A(n8046), .B(n14756), .Y(n14754));
INVX1 mul_U12689(.A(n14754), .Y(n3492));
AND2X1 mul_U12690(.A(n8048), .B(n14759), .Y(n14757));
INVX1 mul_U12691(.A(n14757), .Y(n3493));
AND2X1 mul_U12692(.A(n9829), .B(n14762), .Y(n14760));
INVX1 mul_U12693(.A(n14760), .Y(n3494));
AND2X1 mul_U12694(.A(n7613), .B(n14765), .Y(n14763));
INVX1 mul_U12695(.A(n14763), .Y(n3495));
AND2X1 mul_U12696(.A(n7610), .B(n14768), .Y(n14766));
INVX1 mul_U12697(.A(n14766), .Y(n3496));
AND2X1 mul_U12698(.A(n7609), .B(n14771), .Y(n14769));
INVX1 mul_U12699(.A(n14769), .Y(n3497));
AND2X1 mul_U12700(.A(n7608), .B(n14774), .Y(n14772));
INVX1 mul_U12701(.A(n14772), .Y(n3498));
AND2X1 mul_U12702(.A(dpath_mulcore_ary1_a1_I2_I2_p2_l_64), .B(n14777), .Y(n14775));
INVX1 mul_U12703(.A(n14775), .Y(n3499));
AND2X1 mul_U12704(.A(dpath_mulcore_ary1_a1_I2_I2_p2_l_65), .B(n14780), .Y(n14778));
INVX1 mul_U12705(.A(n14778), .Y(n3500));
AND2X1 mul_U12706(.A(dpath_mulcore_ary1_a1_I2_I2_p2_l_66), .B(dpath_mulcore_ary1_a1_I2_I2_net38), .Y(n14781));
INVX1 mul_U12707(.A(n14781), .Y(n3501));
AND2X1 mul_U12708(.A(n7804), .B(n14785), .Y(n14783));
INVX1 mul_U12709(.A(n14783), .Y(n3502));
AND2X1 mul_U12710(.A(n7801), .B(n14788), .Y(n14786));
INVX1 mul_U12711(.A(n14786), .Y(n3503));
AND2X1 mul_U12712(.A(n7800), .B(dpath_mulcore_ary1_a1_I1_I2_net38), .Y(n14789));
INVX1 mul_U12713(.A(n14789), .Y(n3504));
AND2X1 mul_U12714(.A(n7931), .B(n14793), .Y(n14791));
INVX1 mul_U12715(.A(n14791), .Y(n3505));
AND2X1 mul_U12716(.A(n7928), .B(n14796), .Y(n14794));
INVX1 mul_U12717(.A(n14794), .Y(n3506));
AND2X1 mul_U12718(.A(n7927), .B(dpath_mulcore_ary1_a1_I0_I2_net38), .Y(n14797));
INVX1 mul_U12719(.A(n14797), .Y(n3507));
AND2X1 mul_U12720(.A(n6103), .B(n9682), .Y(n14800));
INVX1 mul_U12721(.A(n14800), .Y(n3508));
AND2X1 mul_U12722(.A(n6104), .B(n9682), .Y(n14802));
INVX1 mul_U12723(.A(n14802), .Y(n3509));
AND2X1 mul_U12724(.A(n6105), .B(n9681), .Y(n14804));
INVX1 mul_U12725(.A(n14804), .Y(n3510));
AND2X1 mul_U12726(.A(n6106), .B(n9682), .Y(n14806));
INVX1 mul_U12727(.A(n14806), .Y(n3511));
AND2X1 mul_U12728(.A(n6107), .B(n9701), .Y(n14808));
INVX1 mul_U12729(.A(n14808), .Y(n3512));
AND2X1 mul_U12730(.A(n6108), .B(n9698), .Y(n14810));
INVX1 mul_U12731(.A(n14810), .Y(n3513));
AND2X1 mul_U12732(.A(n6109), .B(n9681), .Y(n14812));
INVX1 mul_U12733(.A(n14812), .Y(n3514));
AND2X1 mul_U12734(.A(n6110), .B(n9682), .Y(n14814));
INVX1 mul_U12735(.A(n14814), .Y(n3515));
AND2X1 mul_U12736(.A(n6111), .B(n9701), .Y(n14816));
INVX1 mul_U12737(.A(n14816), .Y(n3516));
AND2X1 mul_U12738(.A(n6112), .B(n9698), .Y(n14818));
INVX1 mul_U12739(.A(n14818), .Y(n3517));
AND2X1 mul_U12740(.A(n6113), .B(n9681), .Y(n14820));
INVX1 mul_U12741(.A(n14820), .Y(n3518));
AND2X1 mul_U12742(.A(n6114), .B(n9682), .Y(n14822));
INVX1 mul_U12743(.A(n14822), .Y(n3519));
AND2X1 mul_U12744(.A(n6115), .B(n9701), .Y(n14824));
INVX1 mul_U12745(.A(n14824), .Y(n3520));
AND2X1 mul_U12746(.A(n6116), .B(n9698), .Y(n14826));
INVX1 mul_U12747(.A(n14826), .Y(n3521));
AND2X1 mul_U12748(.A(n6117), .B(n9717), .Y(n14828));
INVX1 mul_U12749(.A(n14828), .Y(n3522));
AND2X1 mul_U12750(.A(n6118), .B(n9717), .Y(n14830));
INVX1 mul_U12751(.A(n14830), .Y(n3523));
AND2X1 mul_U12752(.A(n6119), .B(n9717), .Y(n14832));
INVX1 mul_U12753(.A(n14832), .Y(n3524));
AND2X1 mul_U12754(.A(n6120), .B(n9717), .Y(n14834));
INVX1 mul_U12755(.A(n14834), .Y(n3525));
AND2X1 mul_U12756(.A(n6121), .B(n9717), .Y(n14836));
INVX1 mul_U12757(.A(n14836), .Y(n3526));
AND2X1 mul_U12758(.A(n6122), .B(n9717), .Y(n14838));
INVX1 mul_U12759(.A(n14838), .Y(n3527));
AND2X1 mul_U12760(.A(n6123), .B(n9717), .Y(n14840));
INVX1 mul_U12761(.A(n14840), .Y(n3528));
AND2X1 mul_U12762(.A(n6124), .B(n9717), .Y(n14842));
INVX1 mul_U12763(.A(n14842), .Y(n3529));
AND2X1 mul_U12764(.A(n6125), .B(n9717), .Y(n14844));
INVX1 mul_U12765(.A(n14844), .Y(n3530));
AND2X1 mul_U12766(.A(n6126), .B(n9717), .Y(n14846));
INVX1 mul_U12767(.A(n14846), .Y(n3531));
AND2X1 mul_U12768(.A(n6127), .B(n9717), .Y(n14848));
INVX1 mul_U12769(.A(n14848), .Y(n3532));
AND2X1 mul_U12770(.A(n6128), .B(n9717), .Y(n14850));
INVX1 mul_U12771(.A(n14850), .Y(n3533));
AND2X1 mul_U12772(.A(n6129), .B(n9717), .Y(n14852));
INVX1 mul_U12773(.A(n14852), .Y(n3534));
AND2X1 mul_U12774(.A(n6130), .B(n9717), .Y(n14854));
INVX1 mul_U12775(.A(n14854), .Y(n3535));
AND2X1 mul_U12776(.A(n6131), .B(n9717), .Y(n14856));
INVX1 mul_U12777(.A(n14856), .Y(n3536));
AND2X1 mul_U12778(.A(n6132), .B(n9716), .Y(n14858));
INVX1 mul_U12779(.A(n14858), .Y(n3537));
AND2X1 mul_U12780(.A(n6133), .B(n9716), .Y(n14860));
INVX1 mul_U12781(.A(n14860), .Y(n3538));
AND2X1 mul_U12782(.A(n6134), .B(n9716), .Y(n14862));
INVX1 mul_U12783(.A(n14862), .Y(n3539));
AND2X1 mul_U12784(.A(n6135), .B(n9716), .Y(n14864));
INVX1 mul_U12785(.A(n14864), .Y(n3540));
AND2X1 mul_U12786(.A(n6136), .B(n9716), .Y(n14866));
INVX1 mul_U12787(.A(n14866), .Y(n3541));
AND2X1 mul_U12788(.A(n6137), .B(n9716), .Y(n14868));
INVX1 mul_U12789(.A(n14868), .Y(n3542));
AND2X1 mul_U12790(.A(n6138), .B(n9716), .Y(n14870));
INVX1 mul_U12791(.A(n14870), .Y(n3543));
AND2X1 mul_U12792(.A(n6139), .B(n9716), .Y(n14872));
INVX1 mul_U12793(.A(n14872), .Y(n3544));
AND2X1 mul_U12794(.A(dpath_areg[31]), .B(n9716), .Y(n14874));
INVX1 mul_U12795(.A(n14874), .Y(n3545));
AND2X1 mul_U12796(.A(dpath_areg[30]), .B(n9716), .Y(n14876));
INVX1 mul_U12797(.A(n14876), .Y(n3546));
AND2X1 mul_U12798(.A(dpath_areg[29]), .B(n9716), .Y(n14878));
INVX1 mul_U12799(.A(n14878), .Y(n3547));
AND2X1 mul_U12800(.A(dpath_areg[28]), .B(n9716), .Y(n14880));
INVX1 mul_U12801(.A(n14880), .Y(n3548));
AND2X1 mul_U12802(.A(dpath_areg[27]), .B(n9716), .Y(n14882));
INVX1 mul_U12803(.A(n14882), .Y(n3549));
AND2X1 mul_U12804(.A(dpath_areg[26]), .B(n9716), .Y(n14884));
INVX1 mul_U12805(.A(n14884), .Y(n3550));
AND2X1 mul_U12806(.A(dpath_areg[25]), .B(n9716), .Y(n14886));
INVX1 mul_U12807(.A(n14886), .Y(n3551));
AND2X1 mul_U12808(.A(dpath_areg[24]), .B(n9680), .Y(n14888));
INVX1 mul_U12809(.A(n14888), .Y(n3552));
AND2X1 mul_U12810(.A(dpath_areg[23]), .B(n9680), .Y(n14890));
INVX1 mul_U12811(.A(n14890), .Y(n3553));
AND2X1 mul_U12812(.A(dpath_areg[22]), .B(n9680), .Y(n14892));
INVX1 mul_U12813(.A(n14892), .Y(n3554));
AND2X1 mul_U12814(.A(dpath_areg[21]), .B(n9680), .Y(n14894));
INVX1 mul_U12815(.A(n14894), .Y(n3555));
AND2X1 mul_U12816(.A(dpath_areg[20]), .B(n9681), .Y(n14896));
INVX1 mul_U12817(.A(n14896), .Y(n3556));
AND2X1 mul_U12818(.A(n6076), .B(n9682), .Y(n14899));
INVX1 mul_U12819(.A(n14899), .Y(n3557));
AND2X1 mul_U12820(.A(n6077), .B(n9699), .Y(n14901));
INVX1 mul_U12821(.A(n14901), .Y(n3558));
AND2X1 mul_U12822(.A(n6078), .B(n9700), .Y(n14903));
INVX1 mul_U12823(.A(n14903), .Y(n3559));
AND2X1 mul_U12824(.A(n6079), .B(n9696), .Y(n14905));
INVX1 mul_U12825(.A(n14905), .Y(n3560));
AND2X1 mul_U12826(.A(n6080), .B(n9680), .Y(n14907));
INVX1 mul_U12827(.A(n14907), .Y(n3561));
AND2X1 mul_U12828(.A(n6081), .B(n9701), .Y(n14909));
INVX1 mul_U12829(.A(n14909), .Y(n3562));
AND2X1 mul_U12830(.A(n6082), .B(n9698), .Y(n14911));
INVX1 mul_U12831(.A(n14911), .Y(n3563));
AND2X1 mul_U12832(.A(n6083), .B(n9681), .Y(n14913));
INVX1 mul_U12833(.A(n14913), .Y(n3564));
AND2X1 mul_U12834(.A(n6084), .B(n9682), .Y(n14915));
INVX1 mul_U12835(.A(n14915), .Y(n3565));
AND2X1 mul_U12836(.A(n6085), .B(n9715), .Y(n14917));
INVX1 mul_U12837(.A(n14917), .Y(n3566));
AND2X1 mul_U12838(.A(n6086), .B(n9715), .Y(n14919));
INVX1 mul_U12839(.A(n14919), .Y(n3567));
AND2X1 mul_U12840(.A(n6087), .B(n9715), .Y(n14921));
INVX1 mul_U12841(.A(n14921), .Y(n3568));
AND2X1 mul_U12842(.A(dpath_areg[0]), .B(n9715), .Y(n14923));
INVX1 mul_U12843(.A(n14923), .Y(n3569));
AND2X1 mul_U12844(.A(n6090), .B(n9715), .Y(n14925));
INVX1 mul_U12845(.A(n14925), .Y(n3570));
AND2X1 mul_U12846(.A(n6091), .B(n9715), .Y(n14927));
INVX1 mul_U12847(.A(n14927), .Y(n3571));
AND2X1 mul_U12848(.A(n6092), .B(n9715), .Y(n14929));
INVX1 mul_U12849(.A(n14929), .Y(n3572));
AND2X1 mul_U12850(.A(n6093), .B(n9715), .Y(n14931));
INVX1 mul_U12851(.A(n14931), .Y(n3573));
AND2X1 mul_U12852(.A(n6094), .B(n9715), .Y(n14933));
INVX1 mul_U12853(.A(n14933), .Y(n3574));
AND2X1 mul_U12854(.A(n6095), .B(n9715), .Y(n14935));
INVX1 mul_U12855(.A(n14935), .Y(n3575));
AND2X1 mul_U12856(.A(n6096), .B(n9715), .Y(n14937));
INVX1 mul_U12857(.A(n14937), .Y(n3576));
AND2X1 mul_U12858(.A(n6097), .B(n9715), .Y(n14939));
INVX1 mul_U12859(.A(n14939), .Y(n3577));
AND2X1 mul_U12860(.A(n6098), .B(n9715), .Y(n14941));
INVX1 mul_U12861(.A(n14941), .Y(n3578));
AND2X1 mul_U12862(.A(n6099), .B(n9715), .Y(n14943));
INVX1 mul_U12863(.A(n14943), .Y(n3579));
AND2X1 mul_U12864(.A(n6100), .B(n9715), .Y(n14945));
INVX1 mul_U12865(.A(n14945), .Y(n3580));
AND2X1 mul_U12866(.A(n6101), .B(n9714), .Y(n14947));
INVX1 mul_U12867(.A(n14947), .Y(n3581));
AND2X1 mul_U12868(.A(n6102), .B(n9714), .Y(n14949));
INVX1 mul_U12869(.A(n14949), .Y(n3582));
AND2X1 mul_U12870(.A(dpath_areg[19]), .B(n9714), .Y(n14951));
INVX1 mul_U12871(.A(n14951), .Y(n3583));
AND2X1 mul_U12872(.A(dpath_areg[18]), .B(n9714), .Y(n14953));
INVX1 mul_U12873(.A(n14953), .Y(n3584));
AND2X1 mul_U12874(.A(dpath_areg[17]), .B(n9714), .Y(n14955));
INVX1 mul_U12875(.A(n14955), .Y(n3585));
AND2X1 mul_U12876(.A(dpath_areg[16]), .B(n9714), .Y(n14957));
INVX1 mul_U12877(.A(n14957), .Y(n3586));
AND2X1 mul_U12878(.A(dpath_areg[15]), .B(n9714), .Y(n14959));
INVX1 mul_U12879(.A(n14959), .Y(n3587));
AND2X1 mul_U12880(.A(dpath_areg[4]), .B(n9714), .Y(n14961));
INVX1 mul_U12881(.A(n14961), .Y(n3588));
AND2X1 mul_U12882(.A(dpath_areg[3]), .B(n9714), .Y(n14963));
INVX1 mul_U12883(.A(n14963), .Y(n3589));
AND2X1 mul_U12884(.A(dpath_areg[2]), .B(n9714), .Y(n14965));
INVX1 mul_U12885(.A(n14965), .Y(n3590));
AND2X1 mul_U12886(.A(dpath_areg[1]), .B(n9714), .Y(n14967));
INVX1 mul_U12887(.A(n14967), .Y(n3591));
AND2X1 mul_U12888(.A(n6088), .B(n9714), .Y(n14970));
INVX1 mul_U12889(.A(n14970), .Y(n3592));
AND2X1 mul_U12890(.A(dpath_areg[14]), .B(n9714), .Y(n14972));
INVX1 mul_U12891(.A(n14972), .Y(n3593));
AND2X1 mul_U12892(.A(dpath_areg[13]), .B(n9714), .Y(n14974));
INVX1 mul_U12893(.A(n14974), .Y(n3594));
AND2X1 mul_U12894(.A(dpath_areg[12]), .B(n9714), .Y(n14976));
INVX1 mul_U12895(.A(n14976), .Y(n3595));
AND2X1 mul_U12896(.A(dpath_areg[11]), .B(n9713), .Y(n14978));
INVX1 mul_U12897(.A(n14978), .Y(n3596));
AND2X1 mul_U12898(.A(dpath_areg[10]), .B(n9713), .Y(n14980));
INVX1 mul_U12899(.A(n14980), .Y(n3597));
AND2X1 mul_U12900(.A(dpath_areg[9]), .B(n9713), .Y(n14982));
INVX1 mul_U12901(.A(n14982), .Y(n3598));
AND2X1 mul_U12902(.A(dpath_areg[8]), .B(n9713), .Y(n14984));
INVX1 mul_U12903(.A(n14984), .Y(n3599));
AND2X1 mul_U12904(.A(dpath_areg[7]), .B(n9713), .Y(n14986));
INVX1 mul_U12905(.A(n14986), .Y(n3600));
AND2X1 mul_U12906(.A(dpath_areg[6]), .B(n9713), .Y(n14988));
INVX1 mul_U12907(.A(n14988), .Y(n3601));
AND2X1 mul_U12908(.A(dpath_areg[5]), .B(n9713), .Y(n14990));
INVX1 mul_U12909(.A(n14990), .Y(n3602));
AND2X1 mul_U12910(.A(n8069), .B(n14991), .Y(n14993));
INVX1 mul_U12911(.A(n14993), .Y(n3603));
AND2X1 mul_U12912(.A(n8070), .B(n14994), .Y(n14996));
INVX1 mul_U12913(.A(n14996), .Y(n3604));
AND2X1 mul_U12914(.A(n8071), .B(n14997), .Y(n14999));
INVX1 mul_U12915(.A(n14999), .Y(n3605));
AND2X1 mul_U12916(.A(n8072), .B(n15000), .Y(n15002));
INVX1 mul_U12917(.A(n15002), .Y(n3606));
AND2X1 mul_U12918(.A(n8073), .B(n15003), .Y(n15005));
INVX1 mul_U12919(.A(n15005), .Y(n3607));
AND2X1 mul_U12920(.A(n8074), .B(n15006), .Y(n15008));
INVX1 mul_U12921(.A(n15008), .Y(n3608));
AND2X1 mul_U12922(.A(n8075), .B(n15009), .Y(n15011));
INVX1 mul_U12923(.A(n15011), .Y(n3609));
AND2X1 mul_U12924(.A(n8076), .B(n15012), .Y(n15014));
INVX1 mul_U12925(.A(n15014), .Y(n3610));
AND2X1 mul_U12926(.A(n8077), .B(n15015), .Y(n15017));
INVX1 mul_U12927(.A(n15017), .Y(n3611));
AND2X1 mul_U12928(.A(n8078), .B(n15018), .Y(n15020));
INVX1 mul_U12929(.A(n15020), .Y(n3612));
AND2X1 mul_U12930(.A(n8079), .B(n15021), .Y(n15023));
INVX1 mul_U12931(.A(n15023), .Y(n3613));
AND2X1 mul_U12932(.A(n8080), .B(n15024), .Y(n15026));
INVX1 mul_U12933(.A(n15026), .Y(n3614));
AND2X1 mul_U12934(.A(n8081), .B(n15027), .Y(n15029));
INVX1 mul_U12935(.A(n15029), .Y(n3615));
AND2X1 mul_U12936(.A(n8082), .B(n15030), .Y(n15032));
INVX1 mul_U12937(.A(n15032), .Y(n3616));
AND2X1 mul_U12938(.A(n8083), .B(n15033), .Y(n15035));
INVX1 mul_U12939(.A(n15035), .Y(n3617));
AND2X1 mul_U12940(.A(n8084), .B(n15036), .Y(n15038));
INVX1 mul_U12941(.A(n15038), .Y(n3618));
AND2X1 mul_U12942(.A(n8085), .B(n15039), .Y(n15041));
INVX1 mul_U12943(.A(n15041), .Y(n3619));
AND2X1 mul_U12944(.A(n8086), .B(n15042), .Y(n15044));
INVX1 mul_U12945(.A(n15044), .Y(n3620));
AND2X1 mul_U12946(.A(n8087), .B(n15045), .Y(n15047));
INVX1 mul_U12947(.A(n15047), .Y(n3621));
AND2X1 mul_U12948(.A(n8088), .B(n15048), .Y(n15050));
INVX1 mul_U12949(.A(n15050), .Y(n3622));
AND2X1 mul_U12950(.A(n8089), .B(n15051), .Y(n15053));
INVX1 mul_U12951(.A(n15053), .Y(n3623));
AND2X1 mul_U12952(.A(n8090), .B(n15054), .Y(n15056));
INVX1 mul_U12953(.A(n15056), .Y(n3624));
AND2X1 mul_U12954(.A(n8091), .B(n15057), .Y(n15059));
INVX1 mul_U12955(.A(n15059), .Y(n3625));
AND2X1 mul_U12956(.A(n8092), .B(n15060), .Y(n15062));
INVX1 mul_U12957(.A(n15062), .Y(n3626));
AND2X1 mul_U12958(.A(n8093), .B(n15063), .Y(n15065));
INVX1 mul_U12959(.A(n15065), .Y(n3627));
AND2X1 mul_U12960(.A(n8094), .B(n15066), .Y(n15068));
INVX1 mul_U12961(.A(n15068), .Y(n3628));
AND2X1 mul_U12962(.A(n8095), .B(n15069), .Y(n15071));
INVX1 mul_U12963(.A(n15071), .Y(n3629));
AND2X1 mul_U12964(.A(n8096), .B(n15072), .Y(n15074));
INVX1 mul_U12965(.A(n15074), .Y(n3630));
AND2X1 mul_U12966(.A(n8097), .B(n15075), .Y(n15077));
INVX1 mul_U12967(.A(n15077), .Y(n3631));
AND2X1 mul_U12968(.A(n8098), .B(n15078), .Y(n15080));
INVX1 mul_U12969(.A(n15080), .Y(n3632));
AND2X1 mul_U12970(.A(n8099), .B(n15081), .Y(n15083));
INVX1 mul_U12971(.A(n15083), .Y(n3633));
AND2X1 mul_U12972(.A(n8100), .B(n15084), .Y(n15086));
INVX1 mul_U12973(.A(n15086), .Y(n3634));
AND2X1 mul_U12974(.A(n8101), .B(n15087), .Y(n15089));
INVX1 mul_U12975(.A(n15089), .Y(n3635));
AND2X1 mul_U12976(.A(n8102), .B(n15090), .Y(n15092));
INVX1 mul_U12977(.A(n15092), .Y(n3636));
AND2X1 mul_U12978(.A(n8103), .B(n15093), .Y(n15095));
INVX1 mul_U12979(.A(n15095), .Y(n3637));
AND2X1 mul_U12980(.A(n8104), .B(n15096), .Y(n15098));
INVX1 mul_U12981(.A(n15098), .Y(n3638));
AND2X1 mul_U12982(.A(n8105), .B(n15099), .Y(n15101));
INVX1 mul_U12983(.A(n15101), .Y(n3639));
AND2X1 mul_U12984(.A(n8106), .B(n15102), .Y(n15104));
INVX1 mul_U12985(.A(n15104), .Y(n3640));
AND2X1 mul_U12986(.A(n8107), .B(n15105), .Y(n15107));
INVX1 mul_U12987(.A(n15107), .Y(n3641));
AND2X1 mul_U12988(.A(n8108), .B(n15108), .Y(n15110));
INVX1 mul_U12989(.A(n15110), .Y(n3642));
AND2X1 mul_U12990(.A(n8109), .B(n15111), .Y(n15113));
INVX1 mul_U12991(.A(n15113), .Y(n3643));
AND2X1 mul_U12992(.A(n8110), .B(n15114), .Y(n15116));
INVX1 mul_U12993(.A(n15116), .Y(n3644));
AND2X1 mul_U12994(.A(n8111), .B(n15117), .Y(n15119));
INVX1 mul_U12995(.A(n15119), .Y(n3645));
AND2X1 mul_U12996(.A(n8112), .B(n15120), .Y(n15122));
INVX1 mul_U12997(.A(n15122), .Y(n3646));
AND2X1 mul_U12998(.A(n8113), .B(n15123), .Y(n15125));
INVX1 mul_U12999(.A(n15125), .Y(n3647));
AND2X1 mul_U13000(.A(n8114), .B(n15126), .Y(n15128));
INVX1 mul_U13001(.A(n15128), .Y(n3648));
AND2X1 mul_U13002(.A(n8115), .B(n15129), .Y(n15131));
INVX1 mul_U13003(.A(n15131), .Y(n3649));
AND2X1 mul_U13004(.A(n8116), .B(n15132), .Y(n15134));
INVX1 mul_U13005(.A(n15134), .Y(n3650));
AND2X1 mul_U13006(.A(n8117), .B(n15135), .Y(n15137));
INVX1 mul_U13007(.A(n15137), .Y(n3651));
AND2X1 mul_U13008(.A(n8118), .B(n15138), .Y(n15140));
INVX1 mul_U13009(.A(n15140), .Y(n3652));
AND2X1 mul_U13010(.A(n8119), .B(n15141), .Y(n15143));
INVX1 mul_U13011(.A(n15143), .Y(n3653));
AND2X1 mul_U13012(.A(n8120), .B(n15144), .Y(n15146));
INVX1 mul_U13013(.A(n15146), .Y(n3654));
AND2X1 mul_U13014(.A(n8121), .B(n15147), .Y(n15149));
INVX1 mul_U13015(.A(n15149), .Y(n3655));
AND2X1 mul_U13016(.A(n8122), .B(n15150), .Y(n15152));
INVX1 mul_U13017(.A(n15152), .Y(n3656));
AND2X1 mul_U13018(.A(n8123), .B(n15153), .Y(n15155));
INVX1 mul_U13019(.A(n15155), .Y(n3657));
AND2X1 mul_U13020(.A(n8124), .B(n15156), .Y(n15158));
INVX1 mul_U13021(.A(n15158), .Y(n3658));
AND2X1 mul_U13022(.A(n8125), .B(n15159), .Y(n15161));
INVX1 mul_U13023(.A(n15161), .Y(n3659));
AND2X1 mul_U13024(.A(n8126), .B(n15162), .Y(n15164));
INVX1 mul_U13025(.A(n15164), .Y(n3660));
AND2X1 mul_U13026(.A(n8127), .B(n15165), .Y(n15167));
INVX1 mul_U13027(.A(n15167), .Y(n3661));
AND2X1 mul_U13028(.A(n8056), .B(n15168), .Y(n15170));
INVX1 mul_U13029(.A(n15170), .Y(n3662));
AND2X1 mul_U13030(.A(dpath_mulcore_ary1_a0_s1[3]), .B(n15175), .Y(n15177));
INVX1 mul_U13031(.A(n15177), .Y(n3663));
AND2X1 mul_U13032(.A(dpath_mulcore_ary1_a0_s1[2]), .B(n15178), .Y(n15180));
INVX1 mul_U13033(.A(n15180), .Y(n3664));
AND2X1 mul_U13034(.A(dpath_mulcore_ary1_a0_c_1[2]), .B(n15181), .Y(n15183));
INVX1 mul_U13035(.A(n15183), .Y(n3665));
AND2X1 mul_U13036(.A(n8328), .B(n15193), .Y(n15195));
INVX1 mul_U13037(.A(n15195), .Y(n3666));
AND2X1 mul_U13038(.A(n9486), .B(n15196), .Y(n15198));
INVX1 mul_U13039(.A(n15198), .Y(n3667));
AND2X1 mul_U13040(.A(n16580), .B(n15199), .Y(n15201));
INVX1 mul_U13041(.A(n15201), .Y(n3668));
AND2X1 mul_U13042(.A(n8326), .B(n15202), .Y(n15204));
INVX1 mul_U13043(.A(n15204), .Y(n3669));
AND2X1 mul_U13044(.A(n8327), .B(n15205), .Y(n15207));
INVX1 mul_U13045(.A(n15207), .Y(n3670));
AND2X1 mul_U13046(.A(dpath_mulcore_ary1_a0_s1[63]), .B(n15208), .Y(n15210));
INVX1 mul_U13047(.A(n15210), .Y(n3671));
AND2X1 mul_U13048(.A(dpath_mulcore_ary1_a0_s1[62]), .B(n15211), .Y(n15213));
INVX1 mul_U13049(.A(n15213), .Y(n3672));
AND2X1 mul_U13050(.A(dpath_mulcore_ary1_a0_s1[61]), .B(n15214), .Y(n15216));
INVX1 mul_U13051(.A(n15216), .Y(n3673));
AND2X1 mul_U13052(.A(dpath_mulcore_ary1_a0_s1[60]), .B(n15217), .Y(n15219));
INVX1 mul_U13053(.A(n15219), .Y(n3674));
AND2X1 mul_U13054(.A(dpath_mulcore_ary1_a0_s1[59]), .B(n15220), .Y(n15222));
INVX1 mul_U13055(.A(n15222), .Y(n3675));
AND2X1 mul_U13056(.A(dpath_mulcore_ary1_a0_s1[58]), .B(n15223), .Y(n15225));
INVX1 mul_U13057(.A(n15225), .Y(n3676));
AND2X1 mul_U13058(.A(dpath_mulcore_ary1_a0_s1[57]), .B(n15226), .Y(n15228));
INVX1 mul_U13059(.A(n15228), .Y(n3677));
AND2X1 mul_U13060(.A(dpath_mulcore_ary1_a0_s1[56]), .B(n15229), .Y(n15231));
INVX1 mul_U13061(.A(n15231), .Y(n3678));
AND2X1 mul_U13062(.A(dpath_mulcore_ary1_a0_s1[55]), .B(n15232), .Y(n15234));
INVX1 mul_U13063(.A(n15234), .Y(n3679));
AND2X1 mul_U13064(.A(dpath_mulcore_ary1_a0_s1[54]), .B(n15235), .Y(n15237));
INVX1 mul_U13065(.A(n15237), .Y(n3680));
AND2X1 mul_U13066(.A(dpath_mulcore_ary1_a0_s1[53]), .B(n15238), .Y(n15240));
INVX1 mul_U13067(.A(n15240), .Y(n3681));
AND2X1 mul_U13068(.A(dpath_mulcore_ary1_a0_s1[52]), .B(n15241), .Y(n15243));
INVX1 mul_U13069(.A(n15243), .Y(n3682));
AND2X1 mul_U13070(.A(dpath_mulcore_ary1_a0_s1[51]), .B(n15244), .Y(n15246));
INVX1 mul_U13071(.A(n15246), .Y(n3683));
AND2X1 mul_U13072(.A(dpath_mulcore_ary1_a0_s1[50]), .B(n15247), .Y(n15249));
INVX1 mul_U13073(.A(n15249), .Y(n3684));
AND2X1 mul_U13074(.A(dpath_mulcore_ary1_a0_s1[49]), .B(n15250), .Y(n15252));
INVX1 mul_U13075(.A(n15252), .Y(n3685));
AND2X1 mul_U13076(.A(dpath_mulcore_ary1_a0_s1[48]), .B(n15253), .Y(n15255));
INVX1 mul_U13077(.A(n15255), .Y(n3686));
AND2X1 mul_U13078(.A(dpath_mulcore_ary1_a0_s1[47]), .B(n15256), .Y(n15258));
INVX1 mul_U13079(.A(n15258), .Y(n3687));
AND2X1 mul_U13080(.A(dpath_mulcore_ary1_a0_s1[46]), .B(n15259), .Y(n15261));
INVX1 mul_U13081(.A(n15261), .Y(n3688));
AND2X1 mul_U13082(.A(dpath_mulcore_ary1_a0_s1[45]), .B(n15262), .Y(n15264));
INVX1 mul_U13083(.A(n15264), .Y(n3689));
AND2X1 mul_U13084(.A(dpath_mulcore_ary1_a0_s1[44]), .B(n15265), .Y(n15267));
INVX1 mul_U13085(.A(n15267), .Y(n3690));
AND2X1 mul_U13086(.A(dpath_mulcore_ary1_a0_s1[43]), .B(n15268), .Y(n15270));
INVX1 mul_U13087(.A(n15270), .Y(n3691));
AND2X1 mul_U13088(.A(dpath_mulcore_ary1_a0_s1[42]), .B(n15271), .Y(n15273));
INVX1 mul_U13089(.A(n15273), .Y(n3692));
AND2X1 mul_U13090(.A(dpath_mulcore_ary1_a0_s1[41]), .B(n15274), .Y(n15276));
INVX1 mul_U13091(.A(n15276), .Y(n3693));
AND2X1 mul_U13092(.A(dpath_mulcore_ary1_a0_s1[40]), .B(n15277), .Y(n15279));
INVX1 mul_U13093(.A(n15279), .Y(n3694));
AND2X1 mul_U13094(.A(dpath_mulcore_ary1_a0_s1[39]), .B(n15280), .Y(n15282));
INVX1 mul_U13095(.A(n15282), .Y(n3695));
AND2X1 mul_U13096(.A(dpath_mulcore_ary1_a0_s1[38]), .B(n15283), .Y(n15285));
INVX1 mul_U13097(.A(n15285), .Y(n3696));
AND2X1 mul_U13098(.A(dpath_mulcore_ary1_a0_s1[37]), .B(n15286), .Y(n15288));
INVX1 mul_U13099(.A(n15288), .Y(n3697));
AND2X1 mul_U13100(.A(dpath_mulcore_ary1_a0_s1[36]), .B(n15289), .Y(n15291));
INVX1 mul_U13101(.A(n15291), .Y(n3698));
AND2X1 mul_U13102(.A(dpath_mulcore_ary1_a0_s1[35]), .B(n15292), .Y(n15294));
INVX1 mul_U13103(.A(n15294), .Y(n3699));
AND2X1 mul_U13104(.A(dpath_mulcore_ary1_a0_s1[34]), .B(n15295), .Y(n15297));
INVX1 mul_U13105(.A(n15297), .Y(n3700));
AND2X1 mul_U13106(.A(dpath_mulcore_ary1_a0_s1[33]), .B(n15298), .Y(n15300));
INVX1 mul_U13107(.A(n15300), .Y(n3701));
AND2X1 mul_U13108(.A(dpath_mulcore_ary1_a0_s1[32]), .B(n15301), .Y(n15303));
INVX1 mul_U13109(.A(n15303), .Y(n3702));
AND2X1 mul_U13110(.A(dpath_mulcore_ary1_a0_s1[31]), .B(n15304), .Y(n15306));
INVX1 mul_U13111(.A(n15306), .Y(n3703));
AND2X1 mul_U13112(.A(dpath_mulcore_ary1_a0_s1[30]), .B(n15307), .Y(n15309));
INVX1 mul_U13113(.A(n15309), .Y(n3704));
AND2X1 mul_U13114(.A(dpath_mulcore_ary1_a0_s1[29]), .B(n15310), .Y(n15312));
INVX1 mul_U13115(.A(n15312), .Y(n3705));
AND2X1 mul_U13116(.A(dpath_mulcore_ary1_a0_s1[28]), .B(n15313), .Y(n15315));
INVX1 mul_U13117(.A(n15315), .Y(n3706));
AND2X1 mul_U13118(.A(dpath_mulcore_ary1_a0_s1[27]), .B(n15316), .Y(n15318));
INVX1 mul_U13119(.A(n15318), .Y(n3707));
AND2X1 mul_U13120(.A(dpath_mulcore_ary1_a0_s1[26]), .B(n15319), .Y(n15321));
INVX1 mul_U13121(.A(n15321), .Y(n3708));
AND2X1 mul_U13122(.A(dpath_mulcore_ary1_a0_s1[25]), .B(n15322), .Y(n15324));
INVX1 mul_U13123(.A(n15324), .Y(n3709));
AND2X1 mul_U13124(.A(dpath_mulcore_ary1_a0_s1[24]), .B(n15325), .Y(n15327));
INVX1 mul_U13125(.A(n15327), .Y(n3710));
AND2X1 mul_U13126(.A(dpath_mulcore_ary1_a0_s1[23]), .B(n15328), .Y(n15330));
INVX1 mul_U13127(.A(n15330), .Y(n3711));
AND2X1 mul_U13128(.A(dpath_mulcore_ary1_a0_s1[22]), .B(n15331), .Y(n15333));
INVX1 mul_U13129(.A(n15333), .Y(n3712));
AND2X1 mul_U13130(.A(dpath_mulcore_ary1_a0_s1[21]), .B(n15334), .Y(n15336));
INVX1 mul_U13131(.A(n15336), .Y(n3713));
AND2X1 mul_U13132(.A(dpath_mulcore_ary1_a0_s1[20]), .B(n15337), .Y(n15339));
INVX1 mul_U13133(.A(n15339), .Y(n3714));
AND2X1 mul_U13134(.A(dpath_mulcore_ary1_a0_s1[19]), .B(n15340), .Y(n15342));
INVX1 mul_U13135(.A(n15342), .Y(n3715));
AND2X1 mul_U13136(.A(dpath_mulcore_ary1_a0_s1[18]), .B(n15343), .Y(n15345));
INVX1 mul_U13137(.A(n15345), .Y(n3716));
AND2X1 mul_U13138(.A(dpath_mulcore_ary1_a0_s1[17]), .B(n15346), .Y(n15348));
INVX1 mul_U13139(.A(n15348), .Y(n3717));
AND2X1 mul_U13140(.A(dpath_mulcore_ary1_a0_s1[16]), .B(n15349), .Y(n15351));
INVX1 mul_U13141(.A(n15351), .Y(n3718));
AND2X1 mul_U13142(.A(dpath_mulcore_ary1_a0_s1[15]), .B(n15352), .Y(n15354));
INVX1 mul_U13143(.A(n15354), .Y(n3719));
AND2X1 mul_U13144(.A(dpath_mulcore_ary1_a0_s1[14]), .B(n15355), .Y(n15357));
INVX1 mul_U13145(.A(n15357), .Y(n3720));
AND2X1 mul_U13146(.A(dpath_mulcore_ary1_a0_s1[13]), .B(n15358), .Y(n15360));
INVX1 mul_U13147(.A(n15360), .Y(n3721));
AND2X1 mul_U13148(.A(dpath_mulcore_ary1_a0_s1[12]), .B(n15361), .Y(n15363));
INVX1 mul_U13149(.A(n15363), .Y(n3722));
AND2X1 mul_U13150(.A(dpath_mulcore_ary1_a0_s1[11]), .B(n15364), .Y(n15366));
INVX1 mul_U13151(.A(n15366), .Y(n3723));
AND2X1 mul_U13152(.A(dpath_mulcore_ary1_a0_s1[10]), .B(n15367), .Y(n15369));
INVX1 mul_U13153(.A(n15369), .Y(n3724));
AND2X1 mul_U13154(.A(dpath_mulcore_ary1_a0_s1[9]), .B(n15370), .Y(n15372));
INVX1 mul_U13155(.A(n15372), .Y(n3725));
AND2X1 mul_U13156(.A(dpath_mulcore_ary1_a0_s1[8]), .B(n15373), .Y(n15375));
INVX1 mul_U13157(.A(n15375), .Y(n3726));
AND2X1 mul_U13158(.A(dpath_mulcore_ary1_a0_s1[1]), .B(n15376), .Y(n15378));
INVX1 mul_U13159(.A(n15378), .Y(n3727));
AND2X1 mul_U13160(.A(dpath_mulcore_ary1_a0_s1[0]), .B(n15379), .Y(n15381));
INVX1 mul_U13161(.A(n15381), .Y(n3728));
AND2X1 mul_U13162(.A(n8377), .B(n15382), .Y(n15384));
INVX1 mul_U13163(.A(n15384), .Y(n3729));
AND2X1 mul_U13164(.A(n8378), .B(n15385), .Y(n15387));
INVX1 mul_U13165(.A(n15387), .Y(n3730));
AND2X1 mul_U13166(.A(n8128), .B(n15388), .Y(n15390));
INVX1 mul_U13167(.A(n15390), .Y(n3731));
AND2X1 mul_U13168(.A(n8129), .B(n15391), .Y(n15393));
INVX1 mul_U13169(.A(n15393), .Y(n3732));
AND2X1 mul_U13170(.A(n8130), .B(n15394), .Y(n15396));
INVX1 mul_U13171(.A(n15396), .Y(n3733));
AND2X1 mul_U13172(.A(n8131), .B(n15397), .Y(n15399));
INVX1 mul_U13173(.A(n15399), .Y(n3734));
AND2X1 mul_U13174(.A(n8132), .B(n15400), .Y(n15402));
INVX1 mul_U13175(.A(n15402), .Y(n3735));
AND2X1 mul_U13176(.A(n8133), .B(n15403), .Y(n15405));
INVX1 mul_U13177(.A(n15405), .Y(n3736));
AND2X1 mul_U13178(.A(n8134), .B(n15406), .Y(n15408));
INVX1 mul_U13179(.A(n15408), .Y(n3737));
AND2X1 mul_U13180(.A(n8135), .B(n15409), .Y(n15411));
INVX1 mul_U13181(.A(n15411), .Y(n3738));
AND2X1 mul_U13182(.A(n8136), .B(n15412), .Y(n15414));
INVX1 mul_U13183(.A(n15414), .Y(n3739));
AND2X1 mul_U13184(.A(n8137), .B(n15415), .Y(n15417));
INVX1 mul_U13185(.A(n15417), .Y(n3740));
AND2X1 mul_U13186(.A(n8138), .B(n15418), .Y(n15420));
INVX1 mul_U13187(.A(n15420), .Y(n3741));
AND2X1 mul_U13188(.A(n8139), .B(n15421), .Y(n15423));
INVX1 mul_U13189(.A(n15423), .Y(n3742));
AND2X1 mul_U13190(.A(n8140), .B(n15424), .Y(n15426));
INVX1 mul_U13191(.A(n15426), .Y(n3743));
AND2X1 mul_U13192(.A(n8141), .B(n15427), .Y(n15429));
INVX1 mul_U13193(.A(n15429), .Y(n3744));
AND2X1 mul_U13194(.A(n8142), .B(n15430), .Y(n15432));
INVX1 mul_U13195(.A(n15432), .Y(n3745));
AND2X1 mul_U13196(.A(n8143), .B(n15433), .Y(n15435));
INVX1 mul_U13197(.A(n15435), .Y(n3746));
AND2X1 mul_U13198(.A(n8144), .B(n15436), .Y(n15438));
INVX1 mul_U13199(.A(n15438), .Y(n3747));
AND2X1 mul_U13200(.A(n8145), .B(n15439), .Y(n15441));
INVX1 mul_U13201(.A(n15441), .Y(n3748));
AND2X1 mul_U13202(.A(n8146), .B(n15442), .Y(n15444));
INVX1 mul_U13203(.A(n15444), .Y(n3749));
AND2X1 mul_U13204(.A(n8147), .B(n15445), .Y(n15447));
INVX1 mul_U13205(.A(n15447), .Y(n3750));
AND2X1 mul_U13206(.A(n8148), .B(n15448), .Y(n15450));
INVX1 mul_U13207(.A(n15450), .Y(n3751));
AND2X1 mul_U13208(.A(n8149), .B(n15451), .Y(n15453));
INVX1 mul_U13209(.A(n15453), .Y(n3752));
AND2X1 mul_U13210(.A(n8150), .B(n15454), .Y(n15456));
INVX1 mul_U13211(.A(n15456), .Y(n3753));
AND2X1 mul_U13212(.A(n8151), .B(n15457), .Y(n15459));
INVX1 mul_U13213(.A(n15459), .Y(n3754));
AND2X1 mul_U13214(.A(n8152), .B(n15460), .Y(n15462));
INVX1 mul_U13215(.A(n15462), .Y(n3755));
AND2X1 mul_U13216(.A(n8153), .B(n15463), .Y(n15465));
INVX1 mul_U13217(.A(n15465), .Y(n3756));
AND2X1 mul_U13218(.A(n8154), .B(n15466), .Y(n15468));
INVX1 mul_U13219(.A(n15468), .Y(n3757));
AND2X1 mul_U13220(.A(n8155), .B(n15469), .Y(n15471));
INVX1 mul_U13221(.A(n15471), .Y(n3758));
AND2X1 mul_U13222(.A(n8156), .B(n15472), .Y(n15474));
INVX1 mul_U13223(.A(n15474), .Y(n3759));
AND2X1 mul_U13224(.A(n8157), .B(n15475), .Y(n15477));
INVX1 mul_U13225(.A(n15477), .Y(n3760));
AND2X1 mul_U13226(.A(n8158), .B(n15478), .Y(n15480));
INVX1 mul_U13227(.A(n15480), .Y(n3761));
AND2X1 mul_U13228(.A(n8159), .B(n15481), .Y(n15483));
INVX1 mul_U13229(.A(n15483), .Y(n3762));
AND2X1 mul_U13230(.A(n8160), .B(n15484), .Y(n15486));
INVX1 mul_U13231(.A(n15486), .Y(n3763));
AND2X1 mul_U13232(.A(n8161), .B(n15487), .Y(n15489));
INVX1 mul_U13233(.A(n15489), .Y(n3764));
AND2X1 mul_U13234(.A(n8162), .B(n15490), .Y(n15492));
INVX1 mul_U13235(.A(n15492), .Y(n3765));
AND2X1 mul_U13236(.A(n8163), .B(n15493), .Y(n15495));
INVX1 mul_U13237(.A(n15495), .Y(n3766));
AND2X1 mul_U13238(.A(n8164), .B(n15496), .Y(n15498));
INVX1 mul_U13239(.A(n15498), .Y(n3767));
AND2X1 mul_U13240(.A(n8165), .B(n15499), .Y(n15501));
INVX1 mul_U13241(.A(n15501), .Y(n3768));
AND2X1 mul_U13242(.A(n8166), .B(n15502), .Y(n15504));
INVX1 mul_U13243(.A(n15504), .Y(n3769));
AND2X1 mul_U13244(.A(n8167), .B(n15505), .Y(n15507));
INVX1 mul_U13245(.A(n15507), .Y(n3770));
AND2X1 mul_U13246(.A(n8168), .B(n15508), .Y(n15510));
INVX1 mul_U13247(.A(n15510), .Y(n3771));
AND2X1 mul_U13248(.A(n8169), .B(n15511), .Y(n15513));
INVX1 mul_U13249(.A(n15513), .Y(n3772));
AND2X1 mul_U13250(.A(n8170), .B(n15514), .Y(n15516));
INVX1 mul_U13251(.A(n15516), .Y(n3773));
AND2X1 mul_U13252(.A(n8171), .B(n15517), .Y(n15519));
INVX1 mul_U13253(.A(n15519), .Y(n3774));
AND2X1 mul_U13254(.A(n8172), .B(n15520), .Y(n15522));
INVX1 mul_U13255(.A(n15522), .Y(n3775));
AND2X1 mul_U13256(.A(n8173), .B(n15523), .Y(n15525));
INVX1 mul_U13257(.A(n15525), .Y(n3776));
AND2X1 mul_U13258(.A(n8174), .B(n15526), .Y(n15528));
INVX1 mul_U13259(.A(n15528), .Y(n3777));
AND2X1 mul_U13260(.A(n8175), .B(n15529), .Y(n15531));
INVX1 mul_U13261(.A(n15531), .Y(n3778));
AND2X1 mul_U13262(.A(n8176), .B(n15532), .Y(n15534));
INVX1 mul_U13263(.A(n15534), .Y(n3779));
AND2X1 mul_U13264(.A(n8177), .B(n15535), .Y(n15537));
INVX1 mul_U13265(.A(n15537), .Y(n3780));
AND2X1 mul_U13266(.A(n8178), .B(n15538), .Y(n15540));
INVX1 mul_U13267(.A(n15540), .Y(n3781));
AND2X1 mul_U13268(.A(n8179), .B(n15541), .Y(n15543));
INVX1 mul_U13269(.A(n15543), .Y(n3782));
AND2X1 mul_U13270(.A(n8180), .B(n15544), .Y(n15546));
INVX1 mul_U13271(.A(n15546), .Y(n3783));
AND2X1 mul_U13272(.A(n8181), .B(n15547), .Y(n15549));
INVX1 mul_U13273(.A(n15549), .Y(n3784));
AND2X1 mul_U13274(.A(n8182), .B(n15550), .Y(n15552));
INVX1 mul_U13275(.A(n15552), .Y(n3785));
AND2X1 mul_U13276(.A(n8183), .B(n15553), .Y(n15555));
INVX1 mul_U13277(.A(n15555), .Y(n3786));
AND2X1 mul_U13278(.A(n8184), .B(n15556), .Y(n15558));
INVX1 mul_U13279(.A(n15558), .Y(n3787));
AND2X1 mul_U13280(.A(n8185), .B(n15559), .Y(n15561));
INVX1 mul_U13281(.A(n15561), .Y(n3788));
AND2X1 mul_U13282(.A(n8186), .B(n15562), .Y(n15564));
INVX1 mul_U13283(.A(n15564), .Y(n3789));
AND2X1 mul_U13284(.A(n8187), .B(n15565), .Y(n15567));
INVX1 mul_U13285(.A(n15567), .Y(n3790));
AND2X1 mul_U13286(.A(n8064), .B(n15568), .Y(n15570));
INVX1 mul_U13287(.A(n15570), .Y(n3791));
AND2X1 mul_U13288(.A(dpath_mulcore_ary1_a1_s1[3]), .B(n15575), .Y(n15577));
INVX1 mul_U13289(.A(n15577), .Y(n3792));
AND2X1 mul_U13290(.A(dpath_mulcore_ary1_a1_s1[2]), .B(n15578), .Y(n15580));
INVX1 mul_U13291(.A(n15580), .Y(n3793));
AND2X1 mul_U13292(.A(dpath_mulcore_ary1_a1_c_1[2]), .B(n15581), .Y(n15583));
INVX1 mul_U13293(.A(n15583), .Y(n3794));
AND2X1 mul_U13294(.A(n8188), .B(n15593), .Y(n15595));
INVX1 mul_U13295(.A(n15595), .Y(n3795));
AND2X1 mul_U13296(.A(n9487), .B(n15596), .Y(n15598));
INVX1 mul_U13297(.A(n15598), .Y(n3796));
AND2X1 mul_U13298(.A(n14790), .B(n15599), .Y(n15601));
INVX1 mul_U13299(.A(n15601), .Y(n3797));
AND2X1 mul_U13300(.A(n8190), .B(n15602), .Y(n15604));
INVX1 mul_U13301(.A(n15604), .Y(n3798));
AND2X1 mul_U13302(.A(n8189), .B(n15605), .Y(n15607));
INVX1 mul_U13303(.A(n15607), .Y(n3799));
AND2X1 mul_U13304(.A(dpath_mulcore_ary1_a1_s1[63]), .B(n15608), .Y(n15610));
INVX1 mul_U13305(.A(n15610), .Y(n3800));
AND2X1 mul_U13306(.A(dpath_mulcore_ary1_a1_s1[62]), .B(n15611), .Y(n15613));
INVX1 mul_U13307(.A(n15613), .Y(n3801));
AND2X1 mul_U13308(.A(dpath_mulcore_ary1_a1_s1[61]), .B(n15614), .Y(n15616));
INVX1 mul_U13309(.A(n15616), .Y(n3802));
AND2X1 mul_U13310(.A(dpath_mulcore_ary1_a1_s1[60]), .B(n15617), .Y(n15619));
INVX1 mul_U13311(.A(n15619), .Y(n3803));
AND2X1 mul_U13312(.A(dpath_mulcore_ary1_a1_s1[59]), .B(n15620), .Y(n15622));
INVX1 mul_U13313(.A(n15622), .Y(n3804));
AND2X1 mul_U13314(.A(dpath_mulcore_ary1_a1_s1[58]), .B(n15623), .Y(n15625));
INVX1 mul_U13315(.A(n15625), .Y(n3805));
AND2X1 mul_U13316(.A(dpath_mulcore_ary1_a1_s1[57]), .B(n15626), .Y(n15628));
INVX1 mul_U13317(.A(n15628), .Y(n3806));
AND2X1 mul_U13318(.A(dpath_mulcore_ary1_a1_s1[56]), .B(n15629), .Y(n15631));
INVX1 mul_U13319(.A(n15631), .Y(n3807));
AND2X1 mul_U13320(.A(dpath_mulcore_ary1_a1_s1[55]), .B(n15632), .Y(n15634));
INVX1 mul_U13321(.A(n15634), .Y(n3808));
AND2X1 mul_U13322(.A(dpath_mulcore_ary1_a1_s1[54]), .B(n15635), .Y(n15637));
INVX1 mul_U13323(.A(n15637), .Y(n3809));
AND2X1 mul_U13324(.A(dpath_mulcore_ary1_a1_s1[53]), .B(n15638), .Y(n15640));
INVX1 mul_U13325(.A(n15640), .Y(n3810));
AND2X1 mul_U13326(.A(dpath_mulcore_ary1_a1_s1[52]), .B(n15641), .Y(n15643));
INVX1 mul_U13327(.A(n15643), .Y(n3811));
AND2X1 mul_U13328(.A(dpath_mulcore_ary1_a1_s1[51]), .B(n15644), .Y(n15646));
INVX1 mul_U13329(.A(n15646), .Y(n3812));
AND2X1 mul_U13330(.A(dpath_mulcore_ary1_a1_s1[50]), .B(n15647), .Y(n15649));
INVX1 mul_U13331(.A(n15649), .Y(n3813));
AND2X1 mul_U13332(.A(dpath_mulcore_ary1_a1_s1[49]), .B(n15650), .Y(n15652));
INVX1 mul_U13333(.A(n15652), .Y(n3814));
AND2X1 mul_U13334(.A(dpath_mulcore_ary1_a1_s1[48]), .B(n15653), .Y(n15655));
INVX1 mul_U13335(.A(n15655), .Y(n3815));
AND2X1 mul_U13336(.A(dpath_mulcore_ary1_a1_s1[47]), .B(n15656), .Y(n15658));
INVX1 mul_U13337(.A(n15658), .Y(n3816));
AND2X1 mul_U13338(.A(dpath_mulcore_ary1_a1_s1[46]), .B(n15659), .Y(n15661));
INVX1 mul_U13339(.A(n15661), .Y(n3817));
AND2X1 mul_U13340(.A(dpath_mulcore_ary1_a1_s1[45]), .B(n15662), .Y(n15664));
INVX1 mul_U13341(.A(n15664), .Y(n3818));
AND2X1 mul_U13342(.A(dpath_mulcore_ary1_a1_s1[44]), .B(n15665), .Y(n15667));
INVX1 mul_U13343(.A(n15667), .Y(n3819));
AND2X1 mul_U13344(.A(dpath_mulcore_ary1_a1_s1[43]), .B(n15668), .Y(n15670));
INVX1 mul_U13345(.A(n15670), .Y(n3820));
AND2X1 mul_U13346(.A(dpath_mulcore_ary1_a1_s1[42]), .B(n15671), .Y(n15673));
INVX1 mul_U13347(.A(n15673), .Y(n3821));
AND2X1 mul_U13348(.A(dpath_mulcore_ary1_a1_s1[41]), .B(n15674), .Y(n15676));
INVX1 mul_U13349(.A(n15676), .Y(n3822));
AND2X1 mul_U13350(.A(dpath_mulcore_ary1_a1_s1[40]), .B(n15677), .Y(n15679));
INVX1 mul_U13351(.A(n15679), .Y(n3823));
AND2X1 mul_U13352(.A(dpath_mulcore_ary1_a1_s1[39]), .B(n15680), .Y(n15682));
INVX1 mul_U13353(.A(n15682), .Y(n3824));
AND2X1 mul_U13354(.A(dpath_mulcore_ary1_a1_s1[38]), .B(n15683), .Y(n15685));
INVX1 mul_U13355(.A(n15685), .Y(n3825));
AND2X1 mul_U13356(.A(dpath_mulcore_ary1_a1_s1[37]), .B(n15686), .Y(n15688));
INVX1 mul_U13357(.A(n15688), .Y(n3826));
AND2X1 mul_U13358(.A(dpath_mulcore_ary1_a1_s1[36]), .B(n15689), .Y(n15691));
INVX1 mul_U13359(.A(n15691), .Y(n3827));
AND2X1 mul_U13360(.A(dpath_mulcore_ary1_a1_s1[35]), .B(n15692), .Y(n15694));
INVX1 mul_U13361(.A(n15694), .Y(n3828));
AND2X1 mul_U13362(.A(dpath_mulcore_ary1_a1_s1[34]), .B(n15695), .Y(n15697));
INVX1 mul_U13363(.A(n15697), .Y(n3829));
AND2X1 mul_U13364(.A(dpath_mulcore_ary1_a1_s1[33]), .B(n15698), .Y(n15700));
INVX1 mul_U13365(.A(n15700), .Y(n3830));
AND2X1 mul_U13366(.A(dpath_mulcore_ary1_a1_s1[32]), .B(n15701), .Y(n15703));
INVX1 mul_U13367(.A(n15703), .Y(n3831));
AND2X1 mul_U13368(.A(dpath_mulcore_ary1_a1_s1[31]), .B(n15704), .Y(n15706));
INVX1 mul_U13369(.A(n15706), .Y(n3832));
AND2X1 mul_U13370(.A(dpath_mulcore_ary1_a1_s1[30]), .B(n15707), .Y(n15709));
INVX1 mul_U13371(.A(n15709), .Y(n3833));
AND2X1 mul_U13372(.A(dpath_mulcore_ary1_a1_s1[29]), .B(n15710), .Y(n15712));
INVX1 mul_U13373(.A(n15712), .Y(n3834));
AND2X1 mul_U13374(.A(dpath_mulcore_ary1_a1_s1[28]), .B(n15713), .Y(n15715));
INVX1 mul_U13375(.A(n15715), .Y(n3835));
AND2X1 mul_U13376(.A(dpath_mulcore_ary1_a1_s1[27]), .B(n15716), .Y(n15718));
INVX1 mul_U13377(.A(n15718), .Y(n3836));
AND2X1 mul_U13378(.A(dpath_mulcore_ary1_a1_s1[26]), .B(n15719), .Y(n15721));
INVX1 mul_U13379(.A(n15721), .Y(n3837));
AND2X1 mul_U13380(.A(dpath_mulcore_ary1_a1_s1[25]), .B(n15722), .Y(n15724));
INVX1 mul_U13381(.A(n15724), .Y(n3838));
AND2X1 mul_U13382(.A(dpath_mulcore_ary1_a1_s1[24]), .B(n15725), .Y(n15727));
INVX1 mul_U13383(.A(n15727), .Y(n3839));
AND2X1 mul_U13384(.A(dpath_mulcore_ary1_a1_s1[23]), .B(n15728), .Y(n15730));
INVX1 mul_U13385(.A(n15730), .Y(n3840));
AND2X1 mul_U13386(.A(dpath_mulcore_ary1_a1_s1[22]), .B(n15731), .Y(n15733));
INVX1 mul_U13387(.A(n15733), .Y(n3841));
AND2X1 mul_U13388(.A(dpath_mulcore_ary1_a1_s1[21]), .B(n15734), .Y(n15736));
INVX1 mul_U13389(.A(n15736), .Y(n3842));
AND2X1 mul_U13390(.A(dpath_mulcore_ary1_a1_s1[20]), .B(n15737), .Y(n15739));
INVX1 mul_U13391(.A(n15739), .Y(n3843));
AND2X1 mul_U13392(.A(dpath_mulcore_ary1_a1_s1[19]), .B(n15740), .Y(n15742));
INVX1 mul_U13393(.A(n15742), .Y(n3844));
AND2X1 mul_U13394(.A(dpath_mulcore_ary1_a1_s1[18]), .B(n15743), .Y(n15745));
INVX1 mul_U13395(.A(n15745), .Y(n3845));
AND2X1 mul_U13396(.A(dpath_mulcore_ary1_a1_s1[17]), .B(n15746), .Y(n15748));
INVX1 mul_U13397(.A(n15748), .Y(n3846));
AND2X1 mul_U13398(.A(dpath_mulcore_ary1_a1_s1[16]), .B(n15749), .Y(n15751));
INVX1 mul_U13399(.A(n15751), .Y(n3847));
AND2X1 mul_U13400(.A(dpath_mulcore_ary1_a1_s1[15]), .B(n15752), .Y(n15754));
INVX1 mul_U13401(.A(n15754), .Y(n3848));
AND2X1 mul_U13402(.A(dpath_mulcore_ary1_a1_s1[14]), .B(n15755), .Y(n15757));
INVX1 mul_U13403(.A(n15757), .Y(n3849));
AND2X1 mul_U13404(.A(dpath_mulcore_ary1_a1_s1[13]), .B(n15758), .Y(n15760));
INVX1 mul_U13405(.A(n15760), .Y(n3850));
AND2X1 mul_U13406(.A(dpath_mulcore_ary1_a1_s1[12]), .B(n15761), .Y(n15763));
INVX1 mul_U13407(.A(n15763), .Y(n3851));
AND2X1 mul_U13408(.A(dpath_mulcore_ary1_a1_s1[11]), .B(n15764), .Y(n15766));
INVX1 mul_U13409(.A(n15766), .Y(n3852));
AND2X1 mul_U13410(.A(dpath_mulcore_ary1_a1_s1[10]), .B(n15767), .Y(n15769));
INVX1 mul_U13411(.A(n15769), .Y(n3853));
AND2X1 mul_U13412(.A(dpath_mulcore_ary1_a1_s1[9]), .B(n15770), .Y(n15772));
INVX1 mul_U13413(.A(n15772), .Y(n3854));
AND2X1 mul_U13414(.A(dpath_mulcore_ary1_a1_s1[8]), .B(n15773), .Y(n15775));
INVX1 mul_U13415(.A(n15775), .Y(n3855));
AND2X1 mul_U13416(.A(dpath_mulcore_ary1_a1_s1[1]), .B(n15776), .Y(n15778));
INVX1 mul_U13417(.A(n15778), .Y(n3856));
AND2X1 mul_U13418(.A(dpath_mulcore_ary1_a1_s1[0]), .B(n15779), .Y(n15781));
INVX1 mul_U13419(.A(n15781), .Y(n3857));
AND2X1 mul_U13420(.A(n8381), .B(n15782), .Y(n15784));
INVX1 mul_U13421(.A(n15784), .Y(n3858));
AND2X1 mul_U13422(.A(n8382), .B(n15785), .Y(n15787));
INVX1 mul_U13423(.A(n15787), .Y(n3859));
AND2X1 mul_U13424(.A(dpath_mulcore_array2_c3[81]), .B(n15788), .Y(n15790));
INVX1 mul_U13425(.A(n15790), .Y(n3860));
AND2X1 mul_U13426(.A(n8330), .B(n15791), .Y(n15793));
INVX1 mul_U13427(.A(n15793), .Y(n3861));
AND2X1 mul_U13428(.A(n8331), .B(n15794), .Y(n15796));
INVX1 mul_U13429(.A(n15796), .Y(n3862));
AND2X1 mul_U13430(.A(n8332), .B(n15797), .Y(n15799));
INVX1 mul_U13431(.A(n15799), .Y(n3863));
AND2X1 mul_U13432(.A(n8333), .B(n15800), .Y(n15802));
INVX1 mul_U13433(.A(n15802), .Y(n3864));
AND2X1 mul_U13434(.A(n8334), .B(n15803), .Y(n15805));
INVX1 mul_U13435(.A(n15805), .Y(n3865));
AND2X1 mul_U13436(.A(n8335), .B(n15806), .Y(n15808));
INVX1 mul_U13437(.A(n15808), .Y(n3866));
AND2X1 mul_U13438(.A(n8336), .B(n15809), .Y(n15811));
INVX1 mul_U13439(.A(n15811), .Y(n3867));
AND2X1 mul_U13440(.A(n8337), .B(n15812), .Y(n15814));
INVX1 mul_U13441(.A(n15814), .Y(n3868));
AND2X1 mul_U13442(.A(n8338), .B(n15815), .Y(n15817));
INVX1 mul_U13443(.A(n15817), .Y(n3869));
AND2X1 mul_U13444(.A(n8339), .B(n15818), .Y(n15820));
INVX1 mul_U13445(.A(n15820), .Y(n3870));
AND2X1 mul_U13446(.A(n8340), .B(n15821), .Y(n15823));
INVX1 mul_U13447(.A(n15823), .Y(n3871));
AND2X1 mul_U13448(.A(n8341), .B(n15824), .Y(n15826));
INVX1 mul_U13449(.A(n15826), .Y(n3872));
AND2X1 mul_U13450(.A(n8342), .B(n15827), .Y(n15829));
INVX1 mul_U13451(.A(n15829), .Y(n3873));
AND2X1 mul_U13452(.A(n8343), .B(n15830), .Y(n15832));
INVX1 mul_U13453(.A(n15832), .Y(n3874));
AND2X1 mul_U13454(.A(n8344), .B(n15833), .Y(n15835));
INVX1 mul_U13455(.A(n15835), .Y(n3875));
AND2X1 mul_U13456(.A(n8345), .B(n15836), .Y(n15838));
INVX1 mul_U13457(.A(n15838), .Y(n3876));
AND2X1 mul_U13458(.A(n8346), .B(n15839), .Y(n15841));
INVX1 mul_U13459(.A(n15841), .Y(n3877));
AND2X1 mul_U13460(.A(n8347), .B(n15842), .Y(n15844));
INVX1 mul_U13461(.A(n15844), .Y(n3878));
AND2X1 mul_U13462(.A(n8348), .B(n15845), .Y(n15847));
INVX1 mul_U13463(.A(n15847), .Y(n3879));
AND2X1 mul_U13464(.A(n8349), .B(n15848), .Y(n15850));
INVX1 mul_U13465(.A(n15850), .Y(n3880));
AND2X1 mul_U13466(.A(n8350), .B(n15851), .Y(n15853));
INVX1 mul_U13467(.A(n15853), .Y(n3881));
AND2X1 mul_U13468(.A(n8351), .B(n15854), .Y(n15856));
INVX1 mul_U13469(.A(n15856), .Y(n3882));
AND2X1 mul_U13470(.A(n8352), .B(n15857), .Y(n15859));
INVX1 mul_U13471(.A(n15859), .Y(n3883));
AND2X1 mul_U13472(.A(n8353), .B(n15860), .Y(n15862));
INVX1 mul_U13473(.A(n15862), .Y(n3884));
AND2X1 mul_U13474(.A(n8354), .B(n15863), .Y(n15865));
INVX1 mul_U13475(.A(n15865), .Y(n3885));
AND2X1 mul_U13476(.A(n8355), .B(n15866), .Y(n15868));
INVX1 mul_U13477(.A(n15868), .Y(n3886));
AND2X1 mul_U13478(.A(n8356), .B(n15869), .Y(n15871));
INVX1 mul_U13479(.A(n15871), .Y(n3887));
AND2X1 mul_U13480(.A(n8357), .B(n15872), .Y(n15874));
INVX1 mul_U13481(.A(n15874), .Y(n3888));
AND2X1 mul_U13482(.A(n8358), .B(n15875), .Y(n15877));
INVX1 mul_U13483(.A(n15877), .Y(n3889));
AND2X1 mul_U13484(.A(n8359), .B(n15878), .Y(n15880));
INVX1 mul_U13485(.A(n15880), .Y(n3890));
AND2X1 mul_U13486(.A(n8360), .B(n15881), .Y(n15883));
INVX1 mul_U13487(.A(n15883), .Y(n3891));
AND2X1 mul_U13488(.A(n8361), .B(n15884), .Y(n15886));
INVX1 mul_U13489(.A(n15886), .Y(n3892));
AND2X1 mul_U13490(.A(n8362), .B(n15887), .Y(n15889));
INVX1 mul_U13491(.A(n15889), .Y(n3893));
AND2X1 mul_U13492(.A(n8363), .B(n15890), .Y(n15892));
INVX1 mul_U13493(.A(n15892), .Y(n3894));
AND2X1 mul_U13494(.A(n8364), .B(n15893), .Y(n15895));
INVX1 mul_U13495(.A(n15895), .Y(n3895));
AND2X1 mul_U13496(.A(n8365), .B(n15896), .Y(n15898));
INVX1 mul_U13497(.A(n15898), .Y(n3896));
AND2X1 mul_U13498(.A(n8366), .B(n15899), .Y(n15901));
INVX1 mul_U13499(.A(n15901), .Y(n3897));
AND2X1 mul_U13500(.A(n8367), .B(n15902), .Y(n15904));
INVX1 mul_U13501(.A(n15904), .Y(n3898));
AND2X1 mul_U13502(.A(n8368), .B(n15905), .Y(n15907));
INVX1 mul_U13503(.A(n15907), .Y(n3899));
AND2X1 mul_U13504(.A(n8369), .B(n15908), .Y(n15910));
INVX1 mul_U13505(.A(n15910), .Y(n3900));
AND2X1 mul_U13506(.A(n8370), .B(n15911), .Y(n15913));
INVX1 mul_U13507(.A(n15913), .Y(n3901));
AND2X1 mul_U13508(.A(n8371), .B(n15914), .Y(n15916));
INVX1 mul_U13509(.A(n15916), .Y(n3902));
AND2X1 mul_U13510(.A(n8372), .B(n15917), .Y(n15919));
INVX1 mul_U13511(.A(n15919), .Y(n3903));
AND2X1 mul_U13512(.A(n8373), .B(n15920), .Y(n15922));
INVX1 mul_U13513(.A(n15922), .Y(n3904));
AND2X1 mul_U13514(.A(n8374), .B(n15923), .Y(n15925));
INVX1 mul_U13515(.A(n15925), .Y(n3905));
AND2X1 mul_U13516(.A(n8375), .B(n15926), .Y(n15928));
INVX1 mul_U13517(.A(n15928), .Y(n3906));
AND2X1 mul_U13518(.A(n8376), .B(n15929), .Y(n15931));
INVX1 mul_U13519(.A(n15931), .Y(n3907));
AND2X1 mul_U13520(.A(n17800), .B(n15932), .Y(n15934));
INVX1 mul_U13521(.A(n15934), .Y(n3908));
AND2X1 mul_U13522(.A(n8308), .B(n15935), .Y(n15937));
INVX1 mul_U13523(.A(n15937), .Y(n3909));
AND2X1 mul_U13524(.A(dpath_mulcore_array2_c2[95]), .B(n15938), .Y(n15940));
INVX1 mul_U13525(.A(n15940), .Y(n3910));
AND2X1 mul_U13526(.A(dpath_mulcore_array2_c2[94]), .B(n15941), .Y(n15943));
INVX1 mul_U13527(.A(n15943), .Y(n3911));
AND2X1 mul_U13528(.A(dpath_mulcore_array2_c2[93]), .B(n15944), .Y(n15946));
INVX1 mul_U13529(.A(n15946), .Y(n3912));
AND2X1 mul_U13530(.A(dpath_mulcore_array2_c2[92]), .B(n15947), .Y(n15949));
INVX1 mul_U13531(.A(n15949), .Y(n3913));
AND2X1 mul_U13532(.A(dpath_mulcore_array2_c2[91]), .B(n15950), .Y(n15952));
INVX1 mul_U13533(.A(n15952), .Y(n3914));
AND2X1 mul_U13534(.A(dpath_mulcore_array2_c2[90]), .B(n15953), .Y(n15955));
INVX1 mul_U13535(.A(n15955), .Y(n3915));
AND2X1 mul_U13536(.A(dpath_mulcore_array2_c2[89]), .B(n15956), .Y(n15958));
INVX1 mul_U13537(.A(n15958), .Y(n3916));
AND2X1 mul_U13538(.A(dpath_mulcore_array2_c2[88]), .B(n15959), .Y(n15961));
INVX1 mul_U13539(.A(n15961), .Y(n3917));
AND2X1 mul_U13540(.A(dpath_mulcore_array2_c2[87]), .B(n15962), .Y(n15964));
INVX1 mul_U13541(.A(n15964), .Y(n3918));
AND2X1 mul_U13542(.A(dpath_mulcore_array2_c2[86]), .B(n15965), .Y(n15967));
INVX1 mul_U13543(.A(n15967), .Y(n3919));
AND2X1 mul_U13544(.A(dpath_mulcore_array2_c2[85]), .B(n15968), .Y(n15970));
INVX1 mul_U13545(.A(n15970), .Y(n3920));
AND2X1 mul_U13546(.A(dpath_mulcore_array2_c2[84]), .B(n15971), .Y(n15973));
INVX1 mul_U13547(.A(n15973), .Y(n3921));
AND2X1 mul_U13548(.A(n8303), .B(n15974), .Y(n15976));
INVX1 mul_U13549(.A(n15976), .Y(n3922));
AND2X1 mul_U13550(.A(dpath_mulcore_array2_c3[80]), .B(n15977), .Y(n15979));
INVX1 mul_U13551(.A(n15979), .Y(n3923));
AND2X1 mul_U13552(.A(dpath_mulcore_array2_c3[79]), .B(n15980), .Y(n15982));
INVX1 mul_U13553(.A(n15982), .Y(n3924));
AND2X1 mul_U13554(.A(dpath_mulcore_array2_c3[78]), .B(n15983), .Y(n15985));
INVX1 mul_U13555(.A(n15985), .Y(n3925));
AND2X1 mul_U13556(.A(dpath_mulcore_array2_c3[77]), .B(n15986), .Y(n15988));
INVX1 mul_U13557(.A(n15988), .Y(n3926));
AND2X1 mul_U13558(.A(dpath_mulcore_array2_c3[76]), .B(n15989), .Y(n15991));
INVX1 mul_U13559(.A(n15991), .Y(n3927));
AND2X1 mul_U13560(.A(dpath_mulcore_array2_c3[75]), .B(n15992), .Y(n15994));
INVX1 mul_U13561(.A(n15994), .Y(n3928));
AND2X1 mul_U13562(.A(dpath_mulcore_array2_c3[74]), .B(n15995), .Y(n15997));
INVX1 mul_U13563(.A(n15997), .Y(n3929));
AND2X1 mul_U13564(.A(dpath_mulcore_array2_c3[73]), .B(n15998), .Y(n16000));
INVX1 mul_U13565(.A(n16000), .Y(n3930));
AND2X1 mul_U13566(.A(dpath_mulcore_array2_c3[72]), .B(n16001), .Y(n16003));
INVX1 mul_U13567(.A(n16003), .Y(n3931));
AND2X1 mul_U13568(.A(dpath_mulcore_array2_c3[71]), .B(n16004), .Y(n16006));
INVX1 mul_U13569(.A(n16006), .Y(n3932));
AND2X1 mul_U13570(.A(dpath_mulcore_array2_c3[70]), .B(n16007), .Y(n16009));
INVX1 mul_U13571(.A(n16009), .Y(n3933));
AND2X1 mul_U13572(.A(dpath_mulcore_array2_c3[69]), .B(n16010), .Y(n16012));
INVX1 mul_U13573(.A(n16012), .Y(n3934));
AND2X1 mul_U13574(.A(n8329), .B(n16013), .Y(n16015));
INVX1 mul_U13575(.A(n16015), .Y(n3935));
AND2X1 mul_U13576(.A(dpath_mulcore_array2_c2[3]), .B(n16016), .Y(n16018));
INVX1 mul_U13577(.A(n16018), .Y(n3936));
AND2X1 mul_U13578(.A(dpath_mulcore_array2_c2[2]), .B(n16019), .Y(n16021));
INVX1 mul_U13579(.A(n16021), .Y(n3937));
AND2X1 mul_U13580(.A(dpath_mulcore_array2_c2[1]), .B(n16022), .Y(n16024));
INVX1 mul_U13581(.A(n16024), .Y(n3938));
AND2X1 mul_U13582(.A(dpath_mulcore_array2_c2[0]), .B(n16025), .Y(n16027));
INVX1 mul_U13583(.A(n16027), .Y(n3939));
AND2X1 mul_U13584(.A(dpath_mulcore_a1s[3]), .B(n16031), .Y(n16033));
INVX1 mul_U13585(.A(n16033), .Y(n3940));
AND2X1 mul_U13586(.A(dpath_mulcore_a1s[2]), .B(n16034), .Y(n16036));
INVX1 mul_U13587(.A(n16036), .Y(n3941));
AND2X1 mul_U13588(.A(dpath_mulcore_a1s[1]), .B(n16037), .Y(n16039));
INVX1 mul_U13589(.A(n16039), .Y(n3942));
AND2X1 mul_U13590(.A(dpath_mulcore_a1s[0]), .B(n16040), .Y(n16042));
INVX1 mul_U13591(.A(n16042), .Y(n3943));
AND2X1 mul_U13592(.A(n8324), .B(n16045), .Y(n16047));
INVX1 mul_U13593(.A(n16047), .Y(n3944));
AND2X1 mul_U13594(.A(n8313), .B(n16048), .Y(n16050));
INVX1 mul_U13595(.A(n16050), .Y(n3945));
AND2X1 mul_U13596(.A(dpath_mulcore_a0c[18]), .B(n16051), .Y(n16053));
INVX1 mul_U13597(.A(n16053), .Y(n3946));
AND2X1 mul_U13598(.A(dpath_mulcore_a0c[17]), .B(n16054), .Y(n16056));
INVX1 mul_U13599(.A(n16056), .Y(n3947));
AND2X1 mul_U13600(.A(dpath_mulcore_a0c[16]), .B(n16057), .Y(n16059));
INVX1 mul_U13601(.A(n16059), .Y(n3948));
AND2X1 mul_U13602(.A(dpath_mulcore_a0c[15]), .B(n16060), .Y(n16062));
INVX1 mul_U13603(.A(n16062), .Y(n3949));
AND2X1 mul_U13604(.A(dpath_mulcore_a0c[14]), .B(n16063), .Y(n16065));
INVX1 mul_U13605(.A(n16065), .Y(n3950));
AND2X1 mul_U13606(.A(dpath_mulcore_a0s[80]), .B(n16067), .Y(n16069));
INVX1 mul_U13607(.A(n16069), .Y(n3951));
AND2X1 mul_U13608(.A(dpath_mulcore_a0s[79]), .B(n16070), .Y(n16072));
INVX1 mul_U13609(.A(n16072), .Y(n3952));
AND2X1 mul_U13610(.A(dpath_mulcore_a0s[78]), .B(n16073), .Y(n16075));
INVX1 mul_U13611(.A(n16075), .Y(n3953));
AND2X1 mul_U13612(.A(dpath_mulcore_a0s[77]), .B(n16076), .Y(n16078));
INVX1 mul_U13613(.A(n16078), .Y(n3954));
AND2X1 mul_U13614(.A(dpath_mulcore_a0s[76]), .B(n16079), .Y(n16081));
INVX1 mul_U13615(.A(n16081), .Y(n3955));
AND2X1 mul_U13616(.A(dpath_mulcore_a0s[75]), .B(n16082), .Y(n16084));
INVX1 mul_U13617(.A(n16084), .Y(n3956));
AND2X1 mul_U13618(.A(dpath_mulcore_a0s[74]), .B(n16085), .Y(n16087));
INVX1 mul_U13619(.A(n16087), .Y(n3957));
AND2X1 mul_U13620(.A(dpath_mulcore_a0s[73]), .B(n16088), .Y(n16090));
INVX1 mul_U13621(.A(n16090), .Y(n3958));
AND2X1 mul_U13622(.A(dpath_mulcore_a0s[72]), .B(n16091), .Y(n16093));
INVX1 mul_U13623(.A(n16093), .Y(n3959));
AND2X1 mul_U13624(.A(dpath_mulcore_a0s[71]), .B(n16094), .Y(n16096));
INVX1 mul_U13625(.A(n16096), .Y(n3960));
AND2X1 mul_U13626(.A(dpath_mulcore_a0s[70]), .B(n16097), .Y(n16099));
INVX1 mul_U13627(.A(n16099), .Y(n3961));
AND2X1 mul_U13628(.A(dpath_mulcore_a0s[69]), .B(n16100), .Y(n16102));
INVX1 mul_U13629(.A(n16102), .Y(n3962));
AND2X1 mul_U13630(.A(dpath_mulcore_a0s[68]), .B(n16103), .Y(n16105));
INVX1 mul_U13631(.A(n16105), .Y(n3963));
AND2X1 mul_U13632(.A(n8304), .B(n16106), .Y(n16108));
INVX1 mul_U13633(.A(n16108), .Y(n3964));
AND2X1 mul_U13634(.A(n8305), .B(n16109), .Y(n16111));
INVX1 mul_U13635(.A(n16111), .Y(n3965));
AND2X1 mul_U13636(.A(n8306), .B(n16112), .Y(n16114));
INVX1 mul_U13637(.A(n16114), .Y(n3966));
AND2X1 mul_U13638(.A(n8307), .B(n16115), .Y(n16117));
INVX1 mul_U13639(.A(n16117), .Y(n3967));
AND2X1 mul_U13640(.A(n8314), .B(n16118), .Y(n16120));
INVX1 mul_U13641(.A(n16120), .Y(n3968));
AND2X1 mul_U13642(.A(n8315), .B(n16122), .Y(n16124));
INVX1 mul_U13643(.A(n16124), .Y(n3969));
AND2X1 mul_U13644(.A(n8316), .B(n16125), .Y(n16127));
INVX1 mul_U13645(.A(n16127), .Y(n3970));
AND2X1 mul_U13646(.A(n8317), .B(n16128), .Y(n16130));
INVX1 mul_U13647(.A(n16130), .Y(n3971));
AND2X1 mul_U13648(.A(n8318), .B(n16131), .Y(n16133));
INVX1 mul_U13649(.A(n16133), .Y(n3972));
AND2X1 mul_U13650(.A(n8319), .B(n16134), .Y(n16136));
INVX1 mul_U13651(.A(n16136), .Y(n3973));
AND2X1 mul_U13652(.A(n8320), .B(n16137), .Y(n16139));
INVX1 mul_U13653(.A(n16139), .Y(n3974));
AND2X1 mul_U13654(.A(n8321), .B(n16140), .Y(n16142));
INVX1 mul_U13655(.A(n16142), .Y(n3975));
AND2X1 mul_U13656(.A(n8322), .B(n16143), .Y(n16145));
INVX1 mul_U13657(.A(n16145), .Y(n3976));
AND2X1 mul_U13658(.A(n8323), .B(n16146), .Y(n16148));
INVX1 mul_U13659(.A(n16148), .Y(n3977));
AND2X1 mul_U13660(.A(dpath_mulcore_array2_c2[4]), .B(n16149), .Y(n16151));
INVX1 mul_U13661(.A(n16151), .Y(n3978));
AND2X1 mul_U13662(.A(dpath_mulcore_a0c[66]), .B(n16152), .Y(n16154));
INVX1 mul_U13663(.A(n16154), .Y(n3979));
AND2X1 mul_U13664(.A(dpath_mulcore_a0s[14]), .B(n16155), .Y(n16157));
INVX1 mul_U13665(.A(n16157), .Y(n3980));
AND2X1 mul_U13666(.A(dpath_mulcore_a0s[13]), .B(n16158), .Y(n16160));
INVX1 mul_U13667(.A(n16160), .Y(n3981));
AND2X1 mul_U13668(.A(dpath_mulcore_a0s[12]), .B(n16161), .Y(n16163));
INVX1 mul_U13669(.A(n16163), .Y(n3982));
AND2X1 mul_U13670(.A(dpath_mulcore_a0s[11]), .B(n16164), .Y(n16166));
INVX1 mul_U13671(.A(n16166), .Y(n3983));
AND2X1 mul_U13672(.A(dpath_mulcore_a0s[10]), .B(n16167), .Y(n16169));
INVX1 mul_U13673(.A(n16169), .Y(n3984));
AND2X1 mul_U13674(.A(dpath_mulcore_a0s[9]), .B(n16170), .Y(n16172));
INVX1 mul_U13675(.A(n16172), .Y(n3985));
AND2X1 mul_U13676(.A(dpath_mulcore_a0s[8]), .B(n16173), .Y(n16175));
INVX1 mul_U13677(.A(n16175), .Y(n3986));
AND2X1 mul_U13678(.A(dpath_mulcore_a0s[7]), .B(n16176), .Y(n16178));
INVX1 mul_U13679(.A(n16178), .Y(n3987));
AND2X1 mul_U13680(.A(dpath_mulcore_a0s[6]), .B(n16179), .Y(n16181));
INVX1 mul_U13681(.A(n16181), .Y(n3988));
AND2X1 mul_U13682(.A(dpath_mulcore_a0s[5]), .B(n16182), .Y(n16184));
INVX1 mul_U13683(.A(n16184), .Y(n3989));
AND2X1 mul_U13684(.A(dpath_mulcore_a0c[13]), .B(n16185), .Y(n16187));
INVX1 mul_U13685(.A(n16187), .Y(n3990));
AND2X1 mul_U13686(.A(dpath_mulcore_a0c[12]), .B(n16188), .Y(n16190));
INVX1 mul_U13687(.A(n16190), .Y(n3991));
AND2X1 mul_U13688(.A(dpath_mulcore_a0c[11]), .B(n16191), .Y(n16193));
INVX1 mul_U13689(.A(n16193), .Y(n3992));
AND2X1 mul_U13690(.A(dpath_mulcore_a0c[10]), .B(n16194), .Y(n16196));
INVX1 mul_U13691(.A(n16196), .Y(n3993));
AND2X1 mul_U13692(.A(dpath_mulcore_a0c[9]), .B(n16197), .Y(n16199));
INVX1 mul_U13693(.A(n16199), .Y(n3994));
AND2X1 mul_U13694(.A(dpath_mulcore_a0c[8]), .B(n16200), .Y(n16202));
INVX1 mul_U13695(.A(n16202), .Y(n3995));
AND2X1 mul_U13696(.A(dpath_mulcore_a0c[7]), .B(n16203), .Y(n16205));
INVX1 mul_U13697(.A(n16205), .Y(n3996));
AND2X1 mul_U13698(.A(dpath_mulcore_a0c[6]), .B(n16206), .Y(n16208));
INVX1 mul_U13699(.A(n16208), .Y(n3997));
AND2X1 mul_U13700(.A(dpath_mulcore_a0c[5]), .B(n16209), .Y(n16211));
INVX1 mul_U13701(.A(n16211), .Y(n3998));
AND2X1 mul_U13702(.A(dpath_mulcore_a0c[4]), .B(n16212), .Y(n16214));
INVX1 mul_U13703(.A(n16214), .Y(n3999));
AND2X1 mul_U13704(.A(n8325), .B(n16215), .Y(n16217));
INVX1 mul_U13705(.A(n16217), .Y(n4000));
AND2X1 mul_U13706(.A(dpath_mulcore_a0s[4]), .B(n16218), .Y(n16220));
INVX1 mul_U13707(.A(n16220), .Y(n4001));
AND2X1 mul_U13708(.A(dpath_mulcore_a0s[3]), .B(n16221), .Y(n16223));
INVX1 mul_U13709(.A(n16223), .Y(n4002));
AND2X1 mul_U13710(.A(dpath_mulcore_a0s[2]), .B(n16224), .Y(n16226));
INVX1 mul_U13711(.A(n16226), .Y(n4003));
AND2X1 mul_U13712(.A(dpath_mulcore_a0s[1]), .B(n16227), .Y(n16229));
INVX1 mul_U13713(.A(n16229), .Y(n4004));
AND2X1 mul_U13714(.A(dpath_mulcore_a0c[65]), .B(n16230), .Y(n16232));
INVX1 mul_U13715(.A(n16232), .Y(n4005));
AND2X1 mul_U13716(.A(dpath_mulcore_a0c[64]), .B(n16233), .Y(n16235));
INVX1 mul_U13717(.A(n16235), .Y(n4006));
AND2X1 mul_U13718(.A(dpath_mulcore_a0c[63]), .B(n16236), .Y(n16238));
INVX1 mul_U13719(.A(n16238), .Y(n4007));
AND2X1 mul_U13720(.A(dpath_mulcore_a0c[62]), .B(n16239), .Y(n16241));
INVX1 mul_U13721(.A(n16241), .Y(n4008));
AND2X1 mul_U13722(.A(dpath_mulcore_a0c[61]), .B(n16242), .Y(n16244));
INVX1 mul_U13723(.A(n16244), .Y(n4009));
AND2X1 mul_U13724(.A(dpath_mulcore_a0c[60]), .B(n16245), .Y(n16247));
INVX1 mul_U13725(.A(n16247), .Y(n4010));
AND2X1 mul_U13726(.A(dpath_mulcore_a0c[59]), .B(n16248), .Y(n16250));
INVX1 mul_U13727(.A(n16250), .Y(n4011));
AND2X1 mul_U13728(.A(dpath_mulcore_a0c[58]), .B(n16251), .Y(n16253));
INVX1 mul_U13729(.A(n16253), .Y(n4012));
AND2X1 mul_U13730(.A(dpath_mulcore_a0c[57]), .B(n16254), .Y(n16256));
INVX1 mul_U13731(.A(n16256), .Y(n4013));
AND2X1 mul_U13732(.A(dpath_mulcore_a0c[56]), .B(n16257), .Y(n16259));
INVX1 mul_U13733(.A(n16259), .Y(n4014));
AND2X1 mul_U13734(.A(dpath_mulcore_a0c[55]), .B(n16260), .Y(n16262));
INVX1 mul_U13735(.A(n16262), .Y(n4015));
AND2X1 mul_U13736(.A(dpath_mulcore_a0c[54]), .B(n16263), .Y(n16265));
INVX1 mul_U13737(.A(n16265), .Y(n4016));
AND2X1 mul_U13738(.A(dpath_mulcore_a0c[53]), .B(n16266), .Y(n16268));
INVX1 mul_U13739(.A(n16268), .Y(n4017));
AND2X1 mul_U13740(.A(dpath_mulcore_a0c[52]), .B(n16269), .Y(n16271));
INVX1 mul_U13741(.A(n16271), .Y(n4018));
AND2X1 mul_U13742(.A(dpath_mulcore_a0c[51]), .B(n16272), .Y(n16274));
INVX1 mul_U13743(.A(n16274), .Y(n4019));
AND2X1 mul_U13744(.A(dpath_mulcore_a0c[50]), .B(n16275), .Y(n16277));
INVX1 mul_U13745(.A(n16277), .Y(n4020));
AND2X1 mul_U13746(.A(dpath_mulcore_a0c[49]), .B(n16278), .Y(n16280));
INVX1 mul_U13747(.A(n16280), .Y(n4021));
AND2X1 mul_U13748(.A(dpath_mulcore_a0c[48]), .B(n16281), .Y(n16283));
INVX1 mul_U13749(.A(n16283), .Y(n4022));
AND2X1 mul_U13750(.A(dpath_mulcore_a0c[47]), .B(n16284), .Y(n16286));
INVX1 mul_U13751(.A(n16286), .Y(n4023));
AND2X1 mul_U13752(.A(dpath_mulcore_a0c[46]), .B(n16287), .Y(n16289));
INVX1 mul_U13753(.A(n16289), .Y(n4024));
AND2X1 mul_U13754(.A(dpath_mulcore_a0c[45]), .B(n16290), .Y(n16292));
INVX1 mul_U13755(.A(n16292), .Y(n4025));
AND2X1 mul_U13756(.A(dpath_mulcore_a0c[44]), .B(n16293), .Y(n16295));
INVX1 mul_U13757(.A(n16295), .Y(n4026));
AND2X1 mul_U13758(.A(dpath_mulcore_a0c[43]), .B(n16296), .Y(n16298));
INVX1 mul_U13759(.A(n16298), .Y(n4027));
AND2X1 mul_U13760(.A(dpath_mulcore_a0c[42]), .B(n16299), .Y(n16301));
INVX1 mul_U13761(.A(n16301), .Y(n4028));
AND2X1 mul_U13762(.A(dpath_mulcore_a0c[41]), .B(n16302), .Y(n16304));
INVX1 mul_U13763(.A(n16304), .Y(n4029));
AND2X1 mul_U13764(.A(dpath_mulcore_a0c[40]), .B(n16305), .Y(n16307));
INVX1 mul_U13765(.A(n16307), .Y(n4030));
AND2X1 mul_U13766(.A(dpath_mulcore_a0c[39]), .B(n16308), .Y(n16310));
INVX1 mul_U13767(.A(n16310), .Y(n4031));
AND2X1 mul_U13768(.A(dpath_mulcore_a0c[38]), .B(n16311), .Y(n16313));
INVX1 mul_U13769(.A(n16313), .Y(n4032));
AND2X1 mul_U13770(.A(dpath_mulcore_a0c[37]), .B(n16314), .Y(n16316));
INVX1 mul_U13771(.A(n16316), .Y(n4033));
AND2X1 mul_U13772(.A(dpath_mulcore_a0c[36]), .B(n16317), .Y(n16319));
INVX1 mul_U13773(.A(n16319), .Y(n4034));
AND2X1 mul_U13774(.A(dpath_mulcore_a0c[35]), .B(n16320), .Y(n16322));
INVX1 mul_U13775(.A(n16322), .Y(n4035));
AND2X1 mul_U13776(.A(dpath_mulcore_a0c[34]), .B(n16323), .Y(n16325));
INVX1 mul_U13777(.A(n16325), .Y(n4036));
AND2X1 mul_U13778(.A(dpath_mulcore_a0c[33]), .B(n16326), .Y(n16328));
INVX1 mul_U13779(.A(n16328), .Y(n4037));
AND2X1 mul_U13780(.A(dpath_mulcore_a0c[32]), .B(n16329), .Y(n16331));
INVX1 mul_U13781(.A(n16331), .Y(n4038));
AND2X1 mul_U13782(.A(dpath_mulcore_a0c[31]), .B(n16332), .Y(n16334));
INVX1 mul_U13783(.A(n16334), .Y(n4039));
AND2X1 mul_U13784(.A(dpath_mulcore_a0c[30]), .B(n16335), .Y(n16337));
INVX1 mul_U13785(.A(n16337), .Y(n4040));
AND2X1 mul_U13786(.A(dpath_mulcore_a0c[29]), .B(n16338), .Y(n16340));
INVX1 mul_U13787(.A(n16340), .Y(n4041));
AND2X1 mul_U13788(.A(dpath_mulcore_a0c[28]), .B(n16341), .Y(n16343));
INVX1 mul_U13789(.A(n16343), .Y(n4042));
AND2X1 mul_U13790(.A(dpath_mulcore_a0c[27]), .B(n16344), .Y(n16346));
INVX1 mul_U13791(.A(n16346), .Y(n4043));
AND2X1 mul_U13792(.A(dpath_mulcore_a0c[26]), .B(n16347), .Y(n16349));
INVX1 mul_U13793(.A(n16349), .Y(n4044));
AND2X1 mul_U13794(.A(dpath_mulcore_a0c[25]), .B(n16350), .Y(n16352));
INVX1 mul_U13795(.A(n16352), .Y(n4045));
AND2X1 mul_U13796(.A(dpath_mulcore_a0c[24]), .B(n16353), .Y(n16355));
INVX1 mul_U13797(.A(n16355), .Y(n4046));
AND2X1 mul_U13798(.A(dpath_mulcore_a0c[23]), .B(n16356), .Y(n16358));
INVX1 mul_U13799(.A(n16358), .Y(n4047));
AND2X1 mul_U13800(.A(dpath_mulcore_a0c[22]), .B(n16359), .Y(n16361));
INVX1 mul_U13801(.A(n16361), .Y(n4048));
AND2X1 mul_U13802(.A(dpath_mulcore_a0c[21]), .B(n16362), .Y(n16364));
INVX1 mul_U13803(.A(n16364), .Y(n4049));
AND2X1 mul_U13804(.A(dpath_mulcore_a0c[20]), .B(n16365), .Y(n16367));
INVX1 mul_U13805(.A(n16367), .Y(n4050));
AND2X1 mul_U13806(.A(dpath_mulcore_a1s[50]), .B(n16369), .Y(n16371));
INVX1 mul_U13807(.A(n16371), .Y(n4051));
AND2X1 mul_U13808(.A(dpath_mulcore_a1s[49]), .B(n16372), .Y(n16374));
INVX1 mul_U13809(.A(n16374), .Y(n4052));
AND2X1 mul_U13810(.A(dpath_mulcore_a1s[48]), .B(n16375), .Y(n16377));
INVX1 mul_U13811(.A(n16377), .Y(n4053));
AND2X1 mul_U13812(.A(dpath_mulcore_a1s[47]), .B(n16378), .Y(n16380));
INVX1 mul_U13813(.A(n16380), .Y(n4054));
AND2X1 mul_U13814(.A(dpath_mulcore_a1s[46]), .B(n16381), .Y(n16383));
INVX1 mul_U13815(.A(n16383), .Y(n4055));
AND2X1 mul_U13816(.A(dpath_mulcore_a1s[45]), .B(n16384), .Y(n16386));
INVX1 mul_U13817(.A(n16386), .Y(n4056));
AND2X1 mul_U13818(.A(dpath_mulcore_a1s[44]), .B(n16387), .Y(n16389));
INVX1 mul_U13819(.A(n16389), .Y(n4057));
AND2X1 mul_U13820(.A(dpath_mulcore_a1s[43]), .B(n16390), .Y(n16392));
INVX1 mul_U13821(.A(n16392), .Y(n4058));
AND2X1 mul_U13822(.A(dpath_mulcore_a1s[42]), .B(n16393), .Y(n16395));
INVX1 mul_U13823(.A(n16395), .Y(n4059));
AND2X1 mul_U13824(.A(dpath_mulcore_a1s[41]), .B(n16396), .Y(n16398));
INVX1 mul_U13825(.A(n16398), .Y(n4060));
AND2X1 mul_U13826(.A(dpath_mulcore_a1s[40]), .B(n16399), .Y(n16401));
INVX1 mul_U13827(.A(n16401), .Y(n4061));
AND2X1 mul_U13828(.A(dpath_mulcore_a1s[39]), .B(n16402), .Y(n16404));
INVX1 mul_U13829(.A(n16404), .Y(n4062));
AND2X1 mul_U13830(.A(dpath_mulcore_a1s[38]), .B(n16405), .Y(n16407));
INVX1 mul_U13831(.A(n16407), .Y(n4063));
AND2X1 mul_U13832(.A(dpath_mulcore_a1s[37]), .B(n16408), .Y(n16410));
INVX1 mul_U13833(.A(n16410), .Y(n4064));
AND2X1 mul_U13834(.A(dpath_mulcore_a1s[36]), .B(n16411), .Y(n16413));
INVX1 mul_U13835(.A(n16413), .Y(n4065));
AND2X1 mul_U13836(.A(dpath_mulcore_a1s[35]), .B(n16414), .Y(n16416));
INVX1 mul_U13837(.A(n16416), .Y(n4066));
AND2X1 mul_U13838(.A(dpath_mulcore_a1s[34]), .B(n16417), .Y(n16419));
INVX1 mul_U13839(.A(n16419), .Y(n4067));
AND2X1 mul_U13840(.A(dpath_mulcore_a1s[33]), .B(n16420), .Y(n16422));
INVX1 mul_U13841(.A(n16422), .Y(n4068));
AND2X1 mul_U13842(.A(dpath_mulcore_a1s[32]), .B(n16423), .Y(n16425));
INVX1 mul_U13843(.A(n16425), .Y(n4069));
AND2X1 mul_U13844(.A(dpath_mulcore_a1s[31]), .B(n16426), .Y(n16428));
INVX1 mul_U13845(.A(n16428), .Y(n4070));
AND2X1 mul_U13846(.A(dpath_mulcore_a1s[30]), .B(n16429), .Y(n16431));
INVX1 mul_U13847(.A(n16431), .Y(n4071));
AND2X1 mul_U13848(.A(dpath_mulcore_a1s[29]), .B(n16432), .Y(n16434));
INVX1 mul_U13849(.A(n16434), .Y(n4072));
AND2X1 mul_U13850(.A(dpath_mulcore_a1s[28]), .B(n16435), .Y(n16437));
INVX1 mul_U13851(.A(n16437), .Y(n4073));
AND2X1 mul_U13852(.A(dpath_mulcore_a1s[27]), .B(n16438), .Y(n16440));
INVX1 mul_U13853(.A(n16440), .Y(n4074));
AND2X1 mul_U13854(.A(dpath_mulcore_a1s[26]), .B(n16441), .Y(n16443));
INVX1 mul_U13855(.A(n16443), .Y(n4075));
AND2X1 mul_U13856(.A(dpath_mulcore_a1s[25]), .B(n16444), .Y(n16446));
INVX1 mul_U13857(.A(n16446), .Y(n4076));
AND2X1 mul_U13858(.A(dpath_mulcore_a1s[24]), .B(n16447), .Y(n16449));
INVX1 mul_U13859(.A(n16449), .Y(n4077));
AND2X1 mul_U13860(.A(dpath_mulcore_a1s[23]), .B(n16450), .Y(n16452));
INVX1 mul_U13861(.A(n16452), .Y(n4078));
AND2X1 mul_U13862(.A(dpath_mulcore_a1s[22]), .B(n16453), .Y(n16455));
INVX1 mul_U13863(.A(n16455), .Y(n4079));
AND2X1 mul_U13864(.A(dpath_mulcore_a1s[21]), .B(n16456), .Y(n16458));
INVX1 mul_U13865(.A(n16458), .Y(n4080));
AND2X1 mul_U13866(.A(dpath_mulcore_a1s[20]), .B(n16459), .Y(n16461));
INVX1 mul_U13867(.A(n16461), .Y(n4081));
AND2X1 mul_U13868(.A(dpath_mulcore_a1s[19]), .B(n16462), .Y(n16464));
INVX1 mul_U13869(.A(n16464), .Y(n4082));
AND2X1 mul_U13870(.A(dpath_mulcore_a1s[18]), .B(n16465), .Y(n16467));
INVX1 mul_U13871(.A(n16467), .Y(n4083));
AND2X1 mul_U13872(.A(dpath_mulcore_a1s[17]), .B(n16468), .Y(n16470));
INVX1 mul_U13873(.A(n16470), .Y(n4084));
AND2X1 mul_U13874(.A(dpath_mulcore_a1s[16]), .B(n16471), .Y(n16473));
INVX1 mul_U13875(.A(n16473), .Y(n4085));
AND2X1 mul_U13876(.A(dpath_mulcore_a1s[15]), .B(n16474), .Y(n16476));
INVX1 mul_U13877(.A(n16476), .Y(n4086));
AND2X1 mul_U13878(.A(dpath_mulcore_a1s[14]), .B(n16477), .Y(n16479));
INVX1 mul_U13879(.A(n16479), .Y(n4087));
AND2X1 mul_U13880(.A(dpath_mulcore_a1s[13]), .B(n16480), .Y(n16482));
INVX1 mul_U13881(.A(n16482), .Y(n4088));
AND2X1 mul_U13882(.A(dpath_mulcore_a1s[12]), .B(n16483), .Y(n16485));
INVX1 mul_U13883(.A(n16485), .Y(n4089));
AND2X1 mul_U13884(.A(dpath_mulcore_a1s[11]), .B(n16486), .Y(n16488));
INVX1 mul_U13885(.A(n16488), .Y(n4090));
AND2X1 mul_U13886(.A(dpath_mulcore_a1s[10]), .B(n16489), .Y(n16491));
INVX1 mul_U13887(.A(n16491), .Y(n4091));
AND2X1 mul_U13888(.A(dpath_mulcore_a1s[9]), .B(n16492), .Y(n16494));
INVX1 mul_U13889(.A(n16494), .Y(n4092));
AND2X1 mul_U13890(.A(dpath_mulcore_a1s[8]), .B(n16495), .Y(n16497));
INVX1 mul_U13891(.A(n16497), .Y(n4093));
AND2X1 mul_U13892(.A(dpath_mulcore_a1s[7]), .B(n16498), .Y(n16500));
INVX1 mul_U13893(.A(n16500), .Y(n4094));
AND2X1 mul_U13894(.A(dpath_mulcore_a1s[6]), .B(n16501), .Y(n16503));
INVX1 mul_U13895(.A(n16503), .Y(n4095));
AND2X1 mul_U13896(.A(dpath_mulcore_a1s[5]), .B(n16504), .Y(n16506));
INVX1 mul_U13897(.A(n16506), .Y(n4096));
AND2X1 mul_U13898(.A(dpath_mulcore_a1s[4]), .B(n16507), .Y(n16509));
INVX1 mul_U13899(.A(n16509), .Y(n4097));
AND2X1 mul_U13900(.A(dpath_mulcore_a0c[79]), .B(n16511), .Y(n16513));
INVX1 mul_U13901(.A(n16513), .Y(n4098));
AND2X1 mul_U13902(.A(dpath_mulcore_a0c[78]), .B(n16514), .Y(n16516));
INVX1 mul_U13903(.A(n16516), .Y(n4099));
AND2X1 mul_U13904(.A(dpath_mulcore_a0c[77]), .B(n16517), .Y(n16519));
INVX1 mul_U13905(.A(n16519), .Y(n4100));
AND2X1 mul_U13906(.A(dpath_mulcore_a0c[76]), .B(n16520), .Y(n16522));
INVX1 mul_U13907(.A(n16522), .Y(n4101));
AND2X1 mul_U13908(.A(dpath_mulcore_a0c[75]), .B(n16523), .Y(n16525));
INVX1 mul_U13909(.A(n16525), .Y(n4102));
AND2X1 mul_U13910(.A(dpath_mulcore_a0c[74]), .B(n16526), .Y(n16528));
INVX1 mul_U13911(.A(n16528), .Y(n4103));
AND2X1 mul_U13912(.A(dpath_mulcore_a0c[73]), .B(n16529), .Y(n16531));
INVX1 mul_U13913(.A(n16531), .Y(n4104));
AND2X1 mul_U13914(.A(dpath_mulcore_a0c[72]), .B(n16532), .Y(n16534));
INVX1 mul_U13915(.A(n16534), .Y(n4105));
AND2X1 mul_U13916(.A(dpath_mulcore_a0c[71]), .B(n16535), .Y(n16537));
INVX1 mul_U13917(.A(n16537), .Y(n4106));
AND2X1 mul_U13918(.A(dpath_mulcore_a0c[70]), .B(n16538), .Y(n16540));
INVX1 mul_U13919(.A(n16540), .Y(n4107));
AND2X1 mul_U13920(.A(dpath_mulcore_a0c[69]), .B(n16541), .Y(n16543));
INVX1 mul_U13921(.A(n16543), .Y(n4108));
AND2X1 mul_U13922(.A(dpath_mulcore_a0c[68]), .B(n16544), .Y(n16546));
INVX1 mul_U13923(.A(n16546), .Y(n4109));
AND2X1 mul_U13924(.A(dpath_mulcore_a0c[67]), .B(n16547), .Y(n16549));
INVX1 mul_U13925(.A(n16549), .Y(n4110));
AND2X1 mul_U13926(.A(n8309), .B(n16550), .Y(n16552));
INVX1 mul_U13927(.A(n16552), .Y(n4111));
AND2X1 mul_U13928(.A(n8310), .B(n16553), .Y(n16555));
INVX1 mul_U13929(.A(n16555), .Y(n4112));
AND2X1 mul_U13930(.A(n8311), .B(n16556), .Y(n16558));
INVX1 mul_U13931(.A(n16558), .Y(n4113));
AND2X1 mul_U13932(.A(n8312), .B(n16559), .Y(n16561));
INVX1 mul_U13933(.A(n16561), .Y(n4114));
AND2X1 mul_U13934(.A(dpath_mulcore_a0s[0]), .B(n16564), .Y(n16566));
INVX1 mul_U13935(.A(n16566), .Y(n4115));
AND2X1 mul_U13936(.A(dpath_mulcore_a1c[50]), .B(dpath_mulcore_a1s[51]), .Y(n16567));
INVX1 mul_U13937(.A(n16567), .Y(dpath_mulcore_array2_c1[67]));
AND2X1 mul_U13938(.A(n8384), .B(n16574), .Y(n16576));
INVX1 mul_U13939(.A(n16576), .Y(n4116));
AND2X1 mul_U13940(.A(n8383), .B(n16577), .Y(n16579));
INVX1 mul_U13941(.A(n16579), .Y(n4117));
AND2X1 mul_U13942(.A(n7482), .B(dpath_mulcore_ary1_a0_I1_I2_net38), .Y(n16581));
INVX1 mul_U13943(.A(n16581), .Y(n4118));
AND2X1 mul_U13944(.A(n7483), .B(n16582), .Y(n16584));
INVX1 mul_U13945(.A(n16584), .Y(n4119));
AND2X1 mul_U13946(.A(n7486), .B(n16585), .Y(n16587));
INVX1 mul_U13947(.A(n16587), .Y(n4120));
AND2X1 mul_U13948(.A(n10026), .B(n16608), .Y(n16607));
INVX1 mul_U13949(.A(n16607), .Y(n4121));
AND2X1 mul_U13950(.A(dpath_mulcore_ary1_a0_s_1[69]), .B(n16615), .Y(n16614));
INVX1 mul_U13951(.A(n16614), .Y(n4122));
AND2X1 mul_U13952(.A(dpath_mulcore_ary1_a0_s_1[68]), .B(n16622), .Y(n16621));
INVX1 mul_U13953(.A(n16621), .Y(n4123));
AND2X1 mul_U13954(.A(dpath_mulcore_ary1_a0_s_1[67]), .B(n16629), .Y(n16628));
INVX1 mul_U13955(.A(n16628), .Y(n4124));
AND2X1 mul_U13956(.A(dpath_mulcore_ary1_a0_s_1[66]), .B(n16636), .Y(n16635));
INVX1 mul_U13957(.A(n16635), .Y(n4125));
AND2X1 mul_U13958(.A(dpath_mulcore_ary1_a0_s_1[65]), .B(n16643), .Y(n16642));
INVX1 mul_U13959(.A(n16642), .Y(n4126));
AND2X1 mul_U13960(.A(dpath_mulcore_ary1_a0_s_1[64]), .B(n16650), .Y(n16649));
INVX1 mul_U13961(.A(n16649), .Y(n4127));
AND2X1 mul_U13962(.A(dpath_mulcore_ary1_a0_s_1[63]), .B(n16657), .Y(n16656));
INVX1 mul_U13963(.A(n16656), .Y(n4128));
AND2X1 mul_U13964(.A(dpath_mulcore_ary1_a0_s_1[62]), .B(n16664), .Y(n16663));
INVX1 mul_U13965(.A(n16663), .Y(n4129));
AND2X1 mul_U13966(.A(dpath_mulcore_ary1_a0_s_1[61]), .B(n16671), .Y(n16670));
INVX1 mul_U13967(.A(n16670), .Y(n4130));
AND2X1 mul_U13968(.A(dpath_mulcore_ary1_a0_s_1[60]), .B(n16678), .Y(n16677));
INVX1 mul_U13969(.A(n16677), .Y(n4131));
AND2X1 mul_U13970(.A(dpath_mulcore_ary1_a0_s_1[59]), .B(n16685), .Y(n16684));
INVX1 mul_U13971(.A(n16684), .Y(n4132));
AND2X1 mul_U13972(.A(dpath_mulcore_ary1_a0_s_1[58]), .B(n16692), .Y(n16691));
INVX1 mul_U13973(.A(n16691), .Y(n4133));
AND2X1 mul_U13974(.A(dpath_mulcore_ary1_a0_s_1[57]), .B(n16699), .Y(n16698));
INVX1 mul_U13975(.A(n16698), .Y(n4134));
AND2X1 mul_U13976(.A(dpath_mulcore_ary1_a0_s_1[56]), .B(n16706), .Y(n16705));
INVX1 mul_U13977(.A(n16705), .Y(n4135));
AND2X1 mul_U13978(.A(dpath_mulcore_ary1_a0_s_1[55]), .B(n16713), .Y(n16712));
INVX1 mul_U13979(.A(n16712), .Y(n4136));
AND2X1 mul_U13980(.A(dpath_mulcore_ary1_a0_s_1[54]), .B(n16720), .Y(n16719));
INVX1 mul_U13981(.A(n16719), .Y(n4137));
AND2X1 mul_U13982(.A(dpath_mulcore_ary1_a0_s_1[53]), .B(n16727), .Y(n16726));
INVX1 mul_U13983(.A(n16726), .Y(n4138));
AND2X1 mul_U13984(.A(dpath_mulcore_ary1_a0_s_1[52]), .B(n16734), .Y(n16733));
INVX1 mul_U13985(.A(n16733), .Y(n4139));
AND2X1 mul_U13986(.A(dpath_mulcore_ary1_a0_s_1[51]), .B(n16741), .Y(n16740));
INVX1 mul_U13987(.A(n16740), .Y(n4140));
AND2X1 mul_U13988(.A(dpath_mulcore_ary1_a0_s_1[50]), .B(n16748), .Y(n16747));
INVX1 mul_U13989(.A(n16747), .Y(n4141));
AND2X1 mul_U13990(.A(dpath_mulcore_ary1_a0_s_1[49]), .B(n16755), .Y(n16754));
INVX1 mul_U13991(.A(n16754), .Y(n4142));
AND2X1 mul_U13992(.A(dpath_mulcore_ary1_a0_s_1[48]), .B(n16762), .Y(n16761));
INVX1 mul_U13993(.A(n16761), .Y(n4143));
AND2X1 mul_U13994(.A(dpath_mulcore_ary1_a0_s_1[47]), .B(n16769), .Y(n16768));
INVX1 mul_U13995(.A(n16768), .Y(n4144));
AND2X1 mul_U13996(.A(dpath_mulcore_ary1_a0_s_1[46]), .B(n16776), .Y(n16775));
INVX1 mul_U13997(.A(n16775), .Y(n4145));
AND2X1 mul_U13998(.A(dpath_mulcore_ary1_a0_s_1[45]), .B(n16783), .Y(n16782));
INVX1 mul_U13999(.A(n16782), .Y(n4146));
AND2X1 mul_U14000(.A(dpath_mulcore_ary1_a0_s_1[44]), .B(n16790), .Y(n16789));
INVX1 mul_U14001(.A(n16789), .Y(n4147));
AND2X1 mul_U14002(.A(dpath_mulcore_ary1_a0_s_1[43]), .B(n16797), .Y(n16796));
INVX1 mul_U14003(.A(n16796), .Y(n4148));
AND2X1 mul_U14004(.A(dpath_mulcore_ary1_a0_s_1[42]), .B(n16804), .Y(n16803));
INVX1 mul_U14005(.A(n16803), .Y(n4149));
AND2X1 mul_U14006(.A(dpath_mulcore_ary1_a0_s_1[41]), .B(n16811), .Y(n16810));
INVX1 mul_U14007(.A(n16810), .Y(n4150));
AND2X1 mul_U14008(.A(dpath_mulcore_ary1_a0_s_1[40]), .B(n16818), .Y(n16817));
INVX1 mul_U14009(.A(n16817), .Y(n4151));
AND2X1 mul_U14010(.A(dpath_mulcore_ary1_a0_s_1[39]), .B(n16825), .Y(n16824));
INVX1 mul_U14011(.A(n16824), .Y(n4152));
AND2X1 mul_U14012(.A(dpath_mulcore_ary1_a0_s_1[38]), .B(n16832), .Y(n16831));
INVX1 mul_U14013(.A(n16831), .Y(n4153));
AND2X1 mul_U14014(.A(dpath_mulcore_ary1_a0_s_1[37]), .B(n16839), .Y(n16838));
INVX1 mul_U14015(.A(n16838), .Y(n4154));
AND2X1 mul_U14016(.A(dpath_mulcore_ary1_a0_s_1[36]), .B(n16846), .Y(n16845));
INVX1 mul_U14017(.A(n16845), .Y(n4155));
AND2X1 mul_U14018(.A(dpath_mulcore_ary1_a0_s_1[35]), .B(n16853), .Y(n16852));
INVX1 mul_U14019(.A(n16852), .Y(n4156));
AND2X1 mul_U14020(.A(dpath_mulcore_ary1_a0_s_1[34]), .B(n16860), .Y(n16859));
INVX1 mul_U14021(.A(n16859), .Y(n4157));
AND2X1 mul_U14022(.A(dpath_mulcore_ary1_a0_s_1[33]), .B(n16867), .Y(n16866));
INVX1 mul_U14023(.A(n16866), .Y(n4158));
AND2X1 mul_U14024(.A(dpath_mulcore_ary1_a0_s_1[32]), .B(n16874), .Y(n16873));
INVX1 mul_U14025(.A(n16873), .Y(n4159));
AND2X1 mul_U14026(.A(dpath_mulcore_ary1_a0_s_1[31]), .B(n16881), .Y(n16880));
INVX1 mul_U14027(.A(n16880), .Y(n4160));
AND2X1 mul_U14028(.A(dpath_mulcore_ary1_a0_s_1[30]), .B(n16888), .Y(n16887));
INVX1 mul_U14029(.A(n16887), .Y(n4161));
AND2X1 mul_U14030(.A(dpath_mulcore_ary1_a0_s_1[29]), .B(n16895), .Y(n16894));
INVX1 mul_U14031(.A(n16894), .Y(n4162));
AND2X1 mul_U14032(.A(dpath_mulcore_ary1_a0_s_1[28]), .B(n16902), .Y(n16901));
INVX1 mul_U14033(.A(n16901), .Y(n4163));
AND2X1 mul_U14034(.A(dpath_mulcore_ary1_a0_s_1[27]), .B(n16909), .Y(n16908));
INVX1 mul_U14035(.A(n16908), .Y(n4164));
AND2X1 mul_U14036(.A(dpath_mulcore_ary1_a0_s_1[26]), .B(n16916), .Y(n16915));
INVX1 mul_U14037(.A(n16915), .Y(n4165));
AND2X1 mul_U14038(.A(dpath_mulcore_ary1_a0_s_1[25]), .B(n16923), .Y(n16922));
INVX1 mul_U14039(.A(n16922), .Y(n4166));
AND2X1 mul_U14040(.A(dpath_mulcore_ary1_a0_s_1[24]), .B(n16930), .Y(n16929));
INVX1 mul_U14041(.A(n16929), .Y(n4167));
AND2X1 mul_U14042(.A(dpath_mulcore_ary1_a0_s_1[23]), .B(n16937), .Y(n16936));
INVX1 mul_U14043(.A(n16936), .Y(n4168));
AND2X1 mul_U14044(.A(dpath_mulcore_ary1_a0_s_1[22]), .B(n16944), .Y(n16943));
INVX1 mul_U14045(.A(n16943), .Y(n4169));
AND2X1 mul_U14046(.A(dpath_mulcore_ary1_a0_s_1[21]), .B(n16951), .Y(n16950));
INVX1 mul_U14047(.A(n16950), .Y(n4170));
AND2X1 mul_U14048(.A(dpath_mulcore_ary1_a0_s_1[20]), .B(n16958), .Y(n16957));
INVX1 mul_U14049(.A(n16957), .Y(n4171));
AND2X1 mul_U14050(.A(dpath_mulcore_ary1_a0_s_1[19]), .B(n16965), .Y(n16964));
INVX1 mul_U14051(.A(n16964), .Y(n4172));
AND2X1 mul_U14052(.A(dpath_mulcore_ary1_a0_s_1[18]), .B(n16972), .Y(n16971));
INVX1 mul_U14053(.A(n16971), .Y(n4173));
AND2X1 mul_U14054(.A(dpath_mulcore_ary1_a0_s_1[17]), .B(n16979), .Y(n16978));
INVX1 mul_U14055(.A(n16978), .Y(n4174));
AND2X1 mul_U14056(.A(dpath_mulcore_ary1_a0_s_1[16]), .B(n16986), .Y(n16985));
INVX1 mul_U14057(.A(n16985), .Y(n4175));
AND2X1 mul_U14058(.A(dpath_mulcore_ary1_a0_s_1[15]), .B(n16993), .Y(n16992));
INVX1 mul_U14059(.A(n16992), .Y(n4176));
AND2X1 mul_U14060(.A(dpath_mulcore_ary1_a0_s_1[14]), .B(n17000), .Y(n16999));
INVX1 mul_U14061(.A(n16999), .Y(n4177));
AND2X1 mul_U14062(.A(dpath_mulcore_ary1_a0_s_1[13]), .B(n17007), .Y(n17006));
INVX1 mul_U14063(.A(n17006), .Y(n4178));
AND2X1 mul_U14064(.A(dpath_mulcore_ary1_a0_s_1[12]), .B(n17014), .Y(n17013));
INVX1 mul_U14065(.A(n17013), .Y(n4179));
AND2X1 mul_U14066(.A(dpath_mulcore_ary1_a0_s_1[11]), .B(n17021), .Y(n17020));
INVX1 mul_U14067(.A(n17020), .Y(n4180));
AND2X1 mul_U14068(.A(dpath_mulcore_ary1_a1_s1[65]), .B(n17027), .Y(n17026));
INVX1 mul_U14069(.A(n17026), .Y(n4181));
AND2X1 mul_U14070(.A(n10025), .B(n17052), .Y(n17051));
INVX1 mul_U14071(.A(n17051), .Y(n4182));
AND2X1 mul_U14072(.A(dpath_mulcore_ary1_a1_s_1[69]), .B(n17059), .Y(n17058));
INVX1 mul_U14073(.A(n17058), .Y(n4183));
AND2X1 mul_U14074(.A(dpath_mulcore_ary1_a1_s_1[68]), .B(n17066), .Y(n17065));
INVX1 mul_U14075(.A(n17065), .Y(n4184));
AND2X1 mul_U14076(.A(dpath_mulcore_ary1_a1_s_1[67]), .B(n17073), .Y(n17072));
INVX1 mul_U14077(.A(n17072), .Y(n4185));
AND2X1 mul_U14078(.A(dpath_mulcore_ary1_a1_s_1[66]), .B(n17080), .Y(n17079));
INVX1 mul_U14079(.A(n17079), .Y(n4186));
AND2X1 mul_U14080(.A(dpath_mulcore_ary1_a1_s_1[65]), .B(n17087), .Y(n17086));
INVX1 mul_U14081(.A(n17086), .Y(n4187));
AND2X1 mul_U14082(.A(dpath_mulcore_ary1_a1_s_1[64]), .B(n17094), .Y(n17093));
INVX1 mul_U14083(.A(n17093), .Y(n4188));
AND2X1 mul_U14084(.A(dpath_mulcore_ary1_a1_s_1[63]), .B(n17101), .Y(n17100));
INVX1 mul_U14085(.A(n17100), .Y(n4189));
AND2X1 mul_U14086(.A(dpath_mulcore_ary1_a1_s_1[62]), .B(n17108), .Y(n17107));
INVX1 mul_U14087(.A(n17107), .Y(n4190));
AND2X1 mul_U14088(.A(dpath_mulcore_ary1_a1_s_1[61]), .B(n17115), .Y(n17114));
INVX1 mul_U14089(.A(n17114), .Y(n4191));
AND2X1 mul_U14090(.A(dpath_mulcore_ary1_a1_s_1[60]), .B(n17122), .Y(n17121));
INVX1 mul_U14091(.A(n17121), .Y(n4192));
AND2X1 mul_U14092(.A(dpath_mulcore_ary1_a1_s_1[59]), .B(n17129), .Y(n17128));
INVX1 mul_U14093(.A(n17128), .Y(n4193));
AND2X1 mul_U14094(.A(dpath_mulcore_ary1_a1_s_1[58]), .B(n17136), .Y(n17135));
INVX1 mul_U14095(.A(n17135), .Y(n4194));
AND2X1 mul_U14096(.A(dpath_mulcore_ary1_a1_s_1[57]), .B(n17143), .Y(n17142));
INVX1 mul_U14097(.A(n17142), .Y(n4195));
AND2X1 mul_U14098(.A(dpath_mulcore_ary1_a1_s_1[56]), .B(n17150), .Y(n17149));
INVX1 mul_U14099(.A(n17149), .Y(n4196));
AND2X1 mul_U14100(.A(dpath_mulcore_ary1_a1_s_1[55]), .B(n17157), .Y(n17156));
INVX1 mul_U14101(.A(n17156), .Y(n4197));
AND2X1 mul_U14102(.A(dpath_mulcore_ary1_a1_s_1[54]), .B(n17164), .Y(n17163));
INVX1 mul_U14103(.A(n17163), .Y(n4198));
AND2X1 mul_U14104(.A(dpath_mulcore_ary1_a1_s_1[53]), .B(n17171), .Y(n17170));
INVX1 mul_U14105(.A(n17170), .Y(n4199));
AND2X1 mul_U14106(.A(dpath_mulcore_ary1_a1_s_1[52]), .B(n17178), .Y(n17177));
INVX1 mul_U14107(.A(n17177), .Y(n4200));
AND2X1 mul_U14108(.A(dpath_mulcore_ary1_a1_s_1[51]), .B(n17185), .Y(n17184));
INVX1 mul_U14109(.A(n17184), .Y(n4201));
AND2X1 mul_U14110(.A(dpath_mulcore_ary1_a1_s_1[50]), .B(n17192), .Y(n17191));
INVX1 mul_U14111(.A(n17191), .Y(n4202));
AND2X1 mul_U14112(.A(dpath_mulcore_ary1_a1_s_1[49]), .B(n17199), .Y(n17198));
INVX1 mul_U14113(.A(n17198), .Y(n4203));
AND2X1 mul_U14114(.A(dpath_mulcore_ary1_a1_s_1[48]), .B(n17206), .Y(n17205));
INVX1 mul_U14115(.A(n17205), .Y(n4204));
AND2X1 mul_U14116(.A(dpath_mulcore_ary1_a1_s_1[47]), .B(n17213), .Y(n17212));
INVX1 mul_U14117(.A(n17212), .Y(n4205));
AND2X1 mul_U14118(.A(dpath_mulcore_ary1_a1_s_1[46]), .B(n17220), .Y(n17219));
INVX1 mul_U14119(.A(n17219), .Y(n4206));
AND2X1 mul_U14120(.A(dpath_mulcore_ary1_a1_s_1[45]), .B(n17227), .Y(n17226));
INVX1 mul_U14121(.A(n17226), .Y(n4207));
AND2X1 mul_U14122(.A(dpath_mulcore_ary1_a1_s_1[44]), .B(n17234), .Y(n17233));
INVX1 mul_U14123(.A(n17233), .Y(n4208));
AND2X1 mul_U14124(.A(dpath_mulcore_ary1_a1_s_1[43]), .B(n17241), .Y(n17240));
INVX1 mul_U14125(.A(n17240), .Y(n4209));
AND2X1 mul_U14126(.A(dpath_mulcore_ary1_a1_s_1[42]), .B(n17248), .Y(n17247));
INVX1 mul_U14127(.A(n17247), .Y(n4210));
AND2X1 mul_U14128(.A(dpath_mulcore_ary1_a1_s_1[41]), .B(n17255), .Y(n17254));
INVX1 mul_U14129(.A(n17254), .Y(n4211));
AND2X1 mul_U14130(.A(dpath_mulcore_ary1_a1_s_1[40]), .B(n17262), .Y(n17261));
INVX1 mul_U14131(.A(n17261), .Y(n4212));
AND2X1 mul_U14132(.A(dpath_mulcore_ary1_a1_s_1[39]), .B(n17269), .Y(n17268));
INVX1 mul_U14133(.A(n17268), .Y(n4213));
AND2X1 mul_U14134(.A(dpath_mulcore_ary1_a1_s_1[38]), .B(n17276), .Y(n17275));
INVX1 mul_U14135(.A(n17275), .Y(n4214));
AND2X1 mul_U14136(.A(dpath_mulcore_ary1_a1_s_1[37]), .B(n17283), .Y(n17282));
INVX1 mul_U14137(.A(n17282), .Y(n4215));
AND2X1 mul_U14138(.A(dpath_mulcore_ary1_a1_s_1[36]), .B(n17290), .Y(n17289));
INVX1 mul_U14139(.A(n17289), .Y(n4216));
AND2X1 mul_U14140(.A(dpath_mulcore_ary1_a1_s_1[35]), .B(n17297), .Y(n17296));
INVX1 mul_U14141(.A(n17296), .Y(n4217));
AND2X1 mul_U14142(.A(dpath_mulcore_ary1_a1_s_1[34]), .B(n17304), .Y(n17303));
INVX1 mul_U14143(.A(n17303), .Y(n4218));
AND2X1 mul_U14144(.A(dpath_mulcore_ary1_a1_s_1[33]), .B(n17311), .Y(n17310));
INVX1 mul_U14145(.A(n17310), .Y(n4219));
AND2X1 mul_U14146(.A(dpath_mulcore_ary1_a1_s_1[32]), .B(n17318), .Y(n17317));
INVX1 mul_U14147(.A(n17317), .Y(n4220));
AND2X1 mul_U14148(.A(dpath_mulcore_ary1_a1_s_1[31]), .B(n17325), .Y(n17324));
INVX1 mul_U14149(.A(n17324), .Y(n4221));
AND2X1 mul_U14150(.A(dpath_mulcore_ary1_a1_s_1[30]), .B(n17332), .Y(n17331));
INVX1 mul_U14151(.A(n17331), .Y(n4222));
AND2X1 mul_U14152(.A(dpath_mulcore_ary1_a1_s_1[29]), .B(n17339), .Y(n17338));
INVX1 mul_U14153(.A(n17338), .Y(n4223));
AND2X1 mul_U14154(.A(dpath_mulcore_ary1_a1_s_1[28]), .B(n17346), .Y(n17345));
INVX1 mul_U14155(.A(n17345), .Y(n4224));
AND2X1 mul_U14156(.A(dpath_mulcore_ary1_a1_s_1[27]), .B(n17353), .Y(n17352));
INVX1 mul_U14157(.A(n17352), .Y(n4225));
AND2X1 mul_U14158(.A(dpath_mulcore_ary1_a1_s_1[26]), .B(n17360), .Y(n17359));
INVX1 mul_U14159(.A(n17359), .Y(n4226));
AND2X1 mul_U14160(.A(dpath_mulcore_ary1_a1_s_1[25]), .B(n17367), .Y(n17366));
INVX1 mul_U14161(.A(n17366), .Y(n4227));
AND2X1 mul_U14162(.A(dpath_mulcore_ary1_a1_s_1[24]), .B(n17374), .Y(n17373));
INVX1 mul_U14163(.A(n17373), .Y(n4228));
AND2X1 mul_U14164(.A(dpath_mulcore_ary1_a1_s_1[23]), .B(n17381), .Y(n17380));
INVX1 mul_U14165(.A(n17380), .Y(n4229));
AND2X1 mul_U14166(.A(dpath_mulcore_ary1_a1_s_1[22]), .B(n17388), .Y(n17387));
INVX1 mul_U14167(.A(n17387), .Y(n4230));
AND2X1 mul_U14168(.A(dpath_mulcore_ary1_a1_s_1[21]), .B(n17395), .Y(n17394));
INVX1 mul_U14169(.A(n17394), .Y(n4231));
AND2X1 mul_U14170(.A(dpath_mulcore_ary1_a1_s_1[20]), .B(n17402), .Y(n17401));
INVX1 mul_U14171(.A(n17401), .Y(n4232));
AND2X1 mul_U14172(.A(dpath_mulcore_ary1_a1_s_1[19]), .B(n17409), .Y(n17408));
INVX1 mul_U14173(.A(n17408), .Y(n4233));
AND2X1 mul_U14174(.A(dpath_mulcore_ary1_a1_s_1[18]), .B(n17416), .Y(n17415));
INVX1 mul_U14175(.A(n17415), .Y(n4234));
AND2X1 mul_U14176(.A(dpath_mulcore_ary1_a1_s_1[17]), .B(n17423), .Y(n17422));
INVX1 mul_U14177(.A(n17422), .Y(n4235));
AND2X1 mul_U14178(.A(dpath_mulcore_ary1_a1_s_1[16]), .B(n17430), .Y(n17429));
INVX1 mul_U14179(.A(n17429), .Y(n4236));
AND2X1 mul_U14180(.A(dpath_mulcore_ary1_a1_s_1[15]), .B(n17437), .Y(n17436));
INVX1 mul_U14181(.A(n17436), .Y(n4237));
AND2X1 mul_U14182(.A(dpath_mulcore_ary1_a1_s_1[14]), .B(n17444), .Y(n17443));
INVX1 mul_U14183(.A(n17443), .Y(n4238));
AND2X1 mul_U14184(.A(dpath_mulcore_ary1_a1_s_1[13]), .B(n17451), .Y(n17450));
INVX1 mul_U14185(.A(n17450), .Y(n4239));
AND2X1 mul_U14186(.A(dpath_mulcore_ary1_a1_s_1[12]), .B(n17458), .Y(n17457));
INVX1 mul_U14187(.A(n17457), .Y(n4240));
AND2X1 mul_U14188(.A(dpath_mulcore_ary1_a1_s_1[11]), .B(n17465), .Y(n17464));
INVX1 mul_U14189(.A(n17464), .Y(n4241));
AND2X1 mul_U14190(.A(dpath_mulcore_array2_s2[68]), .B(n10081), .Y(n17470));
INVX1 mul_U14191(.A(n17470), .Y(n4242));
AND2X1 mul_U14192(.A(dpath_mulcore_array2_s2[67]), .B(n10080), .Y(n17473));
INVX1 mul_U14193(.A(n17473), .Y(n4243));
AND2X1 mul_U14194(.A(n9101), .B(n17477), .Y(n17476));
INVX1 mul_U14195(.A(n17476), .Y(n4244));
AND2X1 mul_U14196(.A(dpath_mulcore_array2_s2[66]), .B(n10079), .Y(n17479));
INVX1 mul_U14197(.A(n17479), .Y(n4245));
AND2X1 mul_U14198(.A(n9102), .B(n17484), .Y(n17483));
INVX1 mul_U14199(.A(n17483), .Y(n4246));
AND2X1 mul_U14200(.A(dpath_mulcore_array2_s2[65]), .B(n10078), .Y(n17486));
INVX1 mul_U14201(.A(n17486), .Y(n4247));
AND2X1 mul_U14202(.A(n9103), .B(n17491), .Y(n17490));
INVX1 mul_U14203(.A(n17490), .Y(n4248));
AND2X1 mul_U14204(.A(dpath_mulcore_array2_s2[64]), .B(n10077), .Y(n17493));
INVX1 mul_U14205(.A(n17493), .Y(n4249));
AND2X1 mul_U14206(.A(n9104), .B(n17498), .Y(n17497));
INVX1 mul_U14207(.A(n17497), .Y(n4250));
AND2X1 mul_U14208(.A(dpath_mulcore_array2_s2[63]), .B(n10076), .Y(n17500));
INVX1 mul_U14209(.A(n17500), .Y(n4251));
AND2X1 mul_U14210(.A(n9105), .B(n17505), .Y(n17504));
INVX1 mul_U14211(.A(n17504), .Y(n4252));
AND2X1 mul_U14212(.A(dpath_mulcore_array2_s2[62]), .B(n10075), .Y(n17507));
INVX1 mul_U14213(.A(n17507), .Y(n4253));
AND2X1 mul_U14214(.A(n9106), .B(n17512), .Y(n17511));
INVX1 mul_U14215(.A(n17511), .Y(n4254));
AND2X1 mul_U14216(.A(dpath_mulcore_array2_s2[61]), .B(n10074), .Y(n17514));
INVX1 mul_U14217(.A(n17514), .Y(n4255));
AND2X1 mul_U14218(.A(n9107), .B(n17519), .Y(n17518));
INVX1 mul_U14219(.A(n17518), .Y(n4256));
AND2X1 mul_U14220(.A(dpath_mulcore_array2_s2[60]), .B(n10073), .Y(n17521));
INVX1 mul_U14221(.A(n17521), .Y(n4257));
AND2X1 mul_U14222(.A(n9108), .B(n17526), .Y(n17525));
INVX1 mul_U14223(.A(n17525), .Y(n4258));
AND2X1 mul_U14224(.A(dpath_mulcore_array2_s2[59]), .B(n10072), .Y(n17528));
INVX1 mul_U14225(.A(n17528), .Y(n4259));
AND2X1 mul_U14226(.A(n9109), .B(n17533), .Y(n17532));
INVX1 mul_U14227(.A(n17532), .Y(n4260));
AND2X1 mul_U14228(.A(dpath_mulcore_array2_s2[58]), .B(n10071), .Y(n17535));
INVX1 mul_U14229(.A(n17535), .Y(n4261));
AND2X1 mul_U14230(.A(n9110), .B(n17540), .Y(n17539));
INVX1 mul_U14231(.A(n17539), .Y(n4262));
AND2X1 mul_U14232(.A(dpath_mulcore_array2_s2[57]), .B(n10070), .Y(n17542));
INVX1 mul_U14233(.A(n17542), .Y(n4263));
AND2X1 mul_U14234(.A(n9111), .B(n17547), .Y(n17546));
INVX1 mul_U14235(.A(n17546), .Y(n4264));
AND2X1 mul_U14236(.A(dpath_mulcore_array2_s2[56]), .B(n10069), .Y(n17549));
INVX1 mul_U14237(.A(n17549), .Y(n4265));
AND2X1 mul_U14238(.A(n9112), .B(n17554), .Y(n17553));
INVX1 mul_U14239(.A(n17553), .Y(n4266));
AND2X1 mul_U14240(.A(dpath_mulcore_array2_s2[55]), .B(n10068), .Y(n17556));
INVX1 mul_U14241(.A(n17556), .Y(n4267));
AND2X1 mul_U14242(.A(n9113), .B(n17561), .Y(n17560));
INVX1 mul_U14243(.A(n17560), .Y(n4268));
AND2X1 mul_U14244(.A(dpath_mulcore_array2_s2[54]), .B(n10067), .Y(n17563));
INVX1 mul_U14245(.A(n17563), .Y(n4269));
AND2X1 mul_U14246(.A(n9114), .B(n17568), .Y(n17567));
INVX1 mul_U14247(.A(n17567), .Y(n4270));
AND2X1 mul_U14248(.A(dpath_mulcore_array2_s2[53]), .B(n10066), .Y(n17570));
INVX1 mul_U14249(.A(n17570), .Y(n4271));
AND2X1 mul_U14250(.A(n9115), .B(n17575), .Y(n17574));
INVX1 mul_U14251(.A(n17574), .Y(n4272));
AND2X1 mul_U14252(.A(dpath_mulcore_array2_s2[52]), .B(n10065), .Y(n17577));
INVX1 mul_U14253(.A(n17577), .Y(n4273));
AND2X1 mul_U14254(.A(n9116), .B(n17582), .Y(n17581));
INVX1 mul_U14255(.A(n17581), .Y(n4274));
AND2X1 mul_U14256(.A(dpath_mulcore_array2_s2[51]), .B(n10064), .Y(n17584));
INVX1 mul_U14257(.A(n17584), .Y(n4275));
AND2X1 mul_U14258(.A(n9117), .B(n17589), .Y(n17588));
INVX1 mul_U14259(.A(n17588), .Y(n4276));
AND2X1 mul_U14260(.A(dpath_mulcore_array2_s2[50]), .B(n10063), .Y(n17591));
INVX1 mul_U14261(.A(n17591), .Y(n4277));
AND2X1 mul_U14262(.A(n9118), .B(n17596), .Y(n17595));
INVX1 mul_U14263(.A(n17595), .Y(n4278));
AND2X1 mul_U14264(.A(dpath_mulcore_array2_s2[49]), .B(n10062), .Y(n17598));
INVX1 mul_U14265(.A(n17598), .Y(n4279));
AND2X1 mul_U14266(.A(n9119), .B(n17603), .Y(n17602));
INVX1 mul_U14267(.A(n17602), .Y(n4280));
AND2X1 mul_U14268(.A(dpath_mulcore_array2_s2[48]), .B(n10061), .Y(n17605));
INVX1 mul_U14269(.A(n17605), .Y(n4281));
AND2X1 mul_U14270(.A(n9120), .B(n17610), .Y(n17609));
INVX1 mul_U14271(.A(n17609), .Y(n4282));
AND2X1 mul_U14272(.A(dpath_mulcore_array2_s2[47]), .B(n10060), .Y(n17612));
INVX1 mul_U14273(.A(n17612), .Y(n4283));
AND2X1 mul_U14274(.A(n9121), .B(n17617), .Y(n17616));
INVX1 mul_U14275(.A(n17616), .Y(n4284));
AND2X1 mul_U14276(.A(dpath_mulcore_array2_s2[46]), .B(n10059), .Y(n17619));
INVX1 mul_U14277(.A(n17619), .Y(n4285));
AND2X1 mul_U14278(.A(n9122), .B(n17624), .Y(n17623));
INVX1 mul_U14279(.A(n17623), .Y(n4286));
AND2X1 mul_U14280(.A(dpath_mulcore_array2_s2[45]), .B(n10058), .Y(n17626));
INVX1 mul_U14281(.A(n17626), .Y(n4287));
AND2X1 mul_U14282(.A(n9123), .B(n17631), .Y(n17630));
INVX1 mul_U14283(.A(n17630), .Y(n4288));
AND2X1 mul_U14284(.A(dpath_mulcore_array2_s2[44]), .B(n10057), .Y(n17633));
INVX1 mul_U14285(.A(n17633), .Y(n4289));
AND2X1 mul_U14286(.A(n9124), .B(n17638), .Y(n17637));
INVX1 mul_U14287(.A(n17637), .Y(n4290));
AND2X1 mul_U14288(.A(dpath_mulcore_array2_s2[43]), .B(n10056), .Y(n17640));
INVX1 mul_U14289(.A(n17640), .Y(n4291));
AND2X1 mul_U14290(.A(n9125), .B(n17645), .Y(n17644));
INVX1 mul_U14291(.A(n17644), .Y(n4292));
AND2X1 mul_U14292(.A(dpath_mulcore_array2_s2[42]), .B(n10055), .Y(n17647));
INVX1 mul_U14293(.A(n17647), .Y(n4293));
AND2X1 mul_U14294(.A(n9126), .B(n17652), .Y(n17651));
INVX1 mul_U14295(.A(n17651), .Y(n4294));
AND2X1 mul_U14296(.A(dpath_mulcore_array2_s2[41]), .B(n10054), .Y(n17654));
INVX1 mul_U14297(.A(n17654), .Y(n4295));
AND2X1 mul_U14298(.A(n9127), .B(n17659), .Y(n17658));
INVX1 mul_U14299(.A(n17658), .Y(n4296));
AND2X1 mul_U14300(.A(dpath_mulcore_array2_s2[40]), .B(n10053), .Y(n17661));
INVX1 mul_U14301(.A(n17661), .Y(n4297));
AND2X1 mul_U14302(.A(n9128), .B(n17666), .Y(n17665));
INVX1 mul_U14303(.A(n17665), .Y(n4298));
AND2X1 mul_U14304(.A(dpath_mulcore_array2_s2[39]), .B(n10052), .Y(n17668));
INVX1 mul_U14305(.A(n17668), .Y(n4299));
AND2X1 mul_U14306(.A(n9129), .B(n17673), .Y(n17672));
INVX1 mul_U14307(.A(n17672), .Y(n4300));
AND2X1 mul_U14308(.A(dpath_mulcore_array2_s2[38]), .B(n10051), .Y(n17675));
INVX1 mul_U14309(.A(n17675), .Y(n4301));
AND2X1 mul_U14310(.A(n9130), .B(n17680), .Y(n17679));
INVX1 mul_U14311(.A(n17679), .Y(n4302));
AND2X1 mul_U14312(.A(dpath_mulcore_array2_s2[37]), .B(n10050), .Y(n17682));
INVX1 mul_U14313(.A(n17682), .Y(n4303));
AND2X1 mul_U14314(.A(n9131), .B(n17687), .Y(n17686));
INVX1 mul_U14315(.A(n17686), .Y(n4304));
AND2X1 mul_U14316(.A(dpath_mulcore_array2_s2[36]), .B(n10049), .Y(n17689));
INVX1 mul_U14317(.A(n17689), .Y(n4305));
AND2X1 mul_U14318(.A(n9132), .B(n17694), .Y(n17693));
INVX1 mul_U14319(.A(n17693), .Y(n4306));
AND2X1 mul_U14320(.A(dpath_mulcore_array2_s2[35]), .B(n10048), .Y(n17696));
INVX1 mul_U14321(.A(n17696), .Y(n4307));
AND2X1 mul_U14322(.A(n9133), .B(n17701), .Y(n17700));
INVX1 mul_U14323(.A(n17700), .Y(n4308));
AND2X1 mul_U14324(.A(dpath_mulcore_array2_s2[34]), .B(n10047), .Y(n17703));
INVX1 mul_U14325(.A(n17703), .Y(n4309));
AND2X1 mul_U14326(.A(n9134), .B(n17708), .Y(n17707));
INVX1 mul_U14327(.A(n17707), .Y(n4310));
AND2X1 mul_U14328(.A(dpath_mulcore_array2_s2[33]), .B(n10046), .Y(n17710));
INVX1 mul_U14329(.A(n17710), .Y(n4311));
AND2X1 mul_U14330(.A(n9135), .B(n17715), .Y(n17714));
INVX1 mul_U14331(.A(n17714), .Y(n4312));
AND2X1 mul_U14332(.A(dpath_mulcore_array2_s2[32]), .B(n10045), .Y(n17717));
INVX1 mul_U14333(.A(n17717), .Y(n4313));
AND2X1 mul_U14334(.A(n9136), .B(n17722), .Y(n17721));
INVX1 mul_U14335(.A(n17721), .Y(n4314));
AND2X1 mul_U14336(.A(dpath_mulcore_array2_s2[31]), .B(n10044), .Y(n17724));
INVX1 mul_U14337(.A(n17724), .Y(n4315));
AND2X1 mul_U14338(.A(n9137), .B(n17729), .Y(n17728));
INVX1 mul_U14339(.A(n17728), .Y(n4316));
AND2X1 mul_U14340(.A(dpath_mulcore_array2_s2[30]), .B(n10043), .Y(n17731));
INVX1 mul_U14341(.A(n17731), .Y(n4317));
AND2X1 mul_U14342(.A(n9138), .B(n17736), .Y(n17735));
INVX1 mul_U14343(.A(n17735), .Y(n4318));
AND2X1 mul_U14344(.A(dpath_mulcore_array2_s2[29]), .B(n10042), .Y(n17738));
INVX1 mul_U14345(.A(n17738), .Y(n4319));
AND2X1 mul_U14346(.A(n9139), .B(n17743), .Y(n17742));
INVX1 mul_U14347(.A(n17742), .Y(n4320));
AND2X1 mul_U14348(.A(dpath_mulcore_array2_s2[28]), .B(n10041), .Y(n17745));
INVX1 mul_U14349(.A(n17745), .Y(n4321));
AND2X1 mul_U14350(.A(n9140), .B(n17750), .Y(n17749));
INVX1 mul_U14351(.A(n17749), .Y(n4322));
AND2X1 mul_U14352(.A(dpath_mulcore_array2_s2[27]), .B(n10040), .Y(n17752));
INVX1 mul_U14353(.A(n17752), .Y(n4323));
AND2X1 mul_U14354(.A(n9141), .B(n17757), .Y(n17756));
INVX1 mul_U14355(.A(n17756), .Y(n4324));
AND2X1 mul_U14356(.A(dpath_mulcore_array2_s2[26]), .B(n10039), .Y(n17759));
INVX1 mul_U14357(.A(n17759), .Y(n4325));
AND2X1 mul_U14358(.A(n9142), .B(n17764), .Y(n17763));
INVX1 mul_U14359(.A(n17763), .Y(n4326));
AND2X1 mul_U14360(.A(dpath_mulcore_array2_s2[25]), .B(n10038), .Y(n17766));
INVX1 mul_U14361(.A(n17766), .Y(n4327));
AND2X1 mul_U14362(.A(n9143), .B(n17771), .Y(n17770));
INVX1 mul_U14363(.A(n17770), .Y(n4328));
AND2X1 mul_U14364(.A(dpath_mulcore_array2_s2[24]), .B(n10037), .Y(n17773));
INVX1 mul_U14365(.A(n17773), .Y(n4329));
AND2X1 mul_U14366(.A(n9144), .B(n17778), .Y(n17777));
INVX1 mul_U14367(.A(n17777), .Y(n4330));
AND2X1 mul_U14368(.A(dpath_mulcore_array2_s2[23]), .B(n10036), .Y(n17780));
INVX1 mul_U14369(.A(n17780), .Y(n4331));
AND2X1 mul_U14370(.A(n9145), .B(n17785), .Y(n17784));
INVX1 mul_U14371(.A(n17784), .Y(n4332));
AND2X1 mul_U14372(.A(dpath_mulcore_array2_s2[22]), .B(n10035), .Y(n17787));
INVX1 mul_U14373(.A(n17787), .Y(n4333));
AND2X1 mul_U14374(.A(n9146), .B(n17792), .Y(n17791));
INVX1 mul_U14375(.A(n17791), .Y(n4334));
AND2X1 mul_U14376(.A(dpath_mulcore_array2_s2[21]), .B(n10034), .Y(n17794));
INVX1 mul_U14377(.A(n17794), .Y(n4335));
AND2X1 mul_U14378(.A(n9099), .B(n17799), .Y(n17798));
INVX1 mul_U14379(.A(n17798), .Y(n4336));
AND2X1 mul_U14380(.A(dpath_mul_op2_d[16]), .B(n9792), .Y(n17948));
INVX1 mul_U14381(.A(n17948), .Y(n4337));
AND2X1 mul_U14382(.A(dpath_mulcore_booth_b7_in0[2]), .B(n9793), .Y(n17950));
INVX1 mul_U14383(.A(n17950), .Y(n4338));
AND2X1 mul_U14384(.A(dpath_mulcore_booth_b15_in0[2]), .B(n9806), .Y(n17952));
INVX1 mul_U14385(.A(n17952), .Y(n4339));
AND2X1 mul_U14386(.A(dpath_mul_op2_d[30]), .B(n9805), .Y(n17954));
INVX1 mul_U14387(.A(n17954), .Y(n4340));
AND2X1 mul_U14388(.A(dpath_mulcore_booth_b14_in0[2]), .B(n9804), .Y(n17956));
INVX1 mul_U14389(.A(n17956), .Y(n4341));
AND2X1 mul_U14390(.A(dpath_mul_op2_d[28]), .B(n9803), .Y(n17958));
INVX1 mul_U14391(.A(n17958), .Y(n4342));
AND2X1 mul_U14392(.A(dpath_mulcore_booth_b13_in0[2]), .B(n9802), .Y(n17960));
INVX1 mul_U14393(.A(n17960), .Y(n4343));
AND2X1 mul_U14394(.A(dpath_mul_op2_d[26]), .B(n9801), .Y(n17962));
INVX1 mul_U14395(.A(n17962), .Y(n4344));
AND2X1 mul_U14396(.A(dpath_mulcore_booth_b12_in0[2]), .B(n9800), .Y(n17964));
INVX1 mul_U14397(.A(n17964), .Y(n4345));
AND2X1 mul_U14398(.A(dpath_mul_op2_d[24]), .B(n9799), .Y(n17966));
INVX1 mul_U14399(.A(n17966), .Y(n4346));
AND2X1 mul_U14400(.A(dpath_mulcore_booth_b11_in0[2]), .B(n9798), .Y(n17968));
INVX1 mul_U14401(.A(n17968), .Y(n4347));
AND2X1 mul_U14402(.A(dpath_mul_op2_d[22]), .B(n9797), .Y(n17970));
INVX1 mul_U14403(.A(n17970), .Y(n4348));
AND2X1 mul_U14404(.A(dpath_mulcore_booth_b10_in0[2]), .B(n9796), .Y(n17972));
INVX1 mul_U14405(.A(n17972), .Y(n4349));
AND2X1 mul_U14406(.A(dpath_mul_op2_d[20]), .B(n9794), .Y(n17974));
INVX1 mul_U14407(.A(n17974), .Y(n4350));
AND2X1 mul_U14408(.A(dpath_mul_op2_d[18]), .B(n9793), .Y(n17978));
INVX1 mul_U14409(.A(n17978), .Y(n4351));
AND2X1 mul_U14410(.A(n17981), .B(dpath_mulcore_booth_b15_in0[2]), .Y(n17980));
INVX1 mul_U14411(.A(n17980), .Y(n4352));
AND2X1 mul_U14412(.A(n17985), .B(dpath_mulcore_booth_b14_in0[2]), .Y(n17984));
INVX1 mul_U14413(.A(n17984), .Y(n4353));
AND2X1 mul_U14414(.A(n17989), .B(dpath_mulcore_booth_b13_in0[2]), .Y(n17988));
INVX1 mul_U14415(.A(n17988), .Y(n4354));
AND2X1 mul_U14416(.A(n17993), .B(dpath_mulcore_booth_b12_in0[2]), .Y(n17992));
INVX1 mul_U14417(.A(n17992), .Y(n4355));
AND2X1 mul_U14418(.A(n17997), .B(dpath_mulcore_booth_b11_in0[2]), .Y(n17996));
INVX1 mul_U14419(.A(n17996), .Y(n4356));
AND2X1 mul_U14420(.A(n18001), .B(dpath_mulcore_booth_b10_in0[2]), .Y(n18000));
INVX1 mul_U14421(.A(n18000), .Y(n4357));
AND2X1 mul_U14422(.A(n5413), .B(dpath_mulcore_booth_b9_in0[2]), .Y(n18004));
INVX1 mul_U14423(.A(n18004), .Y(n4358));
AND2X1 mul_U14424(.A(n18009), .B(dpath_mul_op2_d[16]), .Y(n18008));
INVX1 mul_U14425(.A(n18008), .Y(n4359));
AND2X1 mul_U14426(.A(dpath_mulcore_booth_b[31]), .B(n10083), .Y(n18014));
INVX1 mul_U14427(.A(n18014), .Y(n4360));
AND2X1 mul_U14428(.A(dpath_mulcore_booth_b7_in1[2]), .B(n10095), .Y(n18016));
INVX1 mul_U14429(.A(n18016), .Y(n4361));
AND2X1 mul_U14430(.A(dpath_mulcore_booth_b[46]), .B(n10094), .Y(n18018));
INVX1 mul_U14431(.A(n18018), .Y(n4362));
AND2X1 mul_U14432(.A(dpath_mulcore_booth_b6_in1[2]), .B(n10093), .Y(n18020));
INVX1 mul_U14433(.A(n18020), .Y(n4363));
AND2X1 mul_U14434(.A(dpath_mulcore_booth_b[44]), .B(n10092), .Y(n18022));
INVX1 mul_U14435(.A(n18022), .Y(n4364));
AND2X1 mul_U14436(.A(dpath_mulcore_booth_b5_in1[2]), .B(n10091), .Y(n18024));
INVX1 mul_U14437(.A(n18024), .Y(n4365));
AND2X1 mul_U14438(.A(dpath_mulcore_booth_b[42]), .B(n10090), .Y(n18026));
INVX1 mul_U14439(.A(n18026), .Y(n4366));
AND2X1 mul_U14440(.A(dpath_mulcore_booth_b4_in1[2]), .B(n10089), .Y(n18028));
INVX1 mul_U14441(.A(n18028), .Y(n4367));
AND2X1 mul_U14442(.A(dpath_mulcore_booth_b[40]), .B(n10088), .Y(n18030));
INVX1 mul_U14443(.A(n18030), .Y(n4368));
AND2X1 mul_U14444(.A(dpath_mulcore_booth_b3_in1[2]), .B(n10087), .Y(n18032));
INVX1 mul_U14445(.A(n18032), .Y(n4369));
AND2X1 mul_U14446(.A(dpath_mulcore_booth_b[38]), .B(n10086), .Y(n18034));
INVX1 mul_U14447(.A(n18034), .Y(n4370));
AND2X1 mul_U14448(.A(dpath_mulcore_booth_b2_in1[2]), .B(n10085), .Y(n18036));
INVX1 mul_U14449(.A(n18036), .Y(n4371));
AND2X1 mul_U14450(.A(dpath_mulcore_booth_b[36]), .B(n10084), .Y(n18038));
INVX1 mul_U14451(.A(n18038), .Y(n4372));
AND2X1 mul_U14452(.A(dpath_mulcore_booth_b[34]), .B(n10083), .Y(n18042));
INVX1 mul_U14453(.A(n18042), .Y(n4373));
AND2X1 mul_U14454(.A(n18045), .B(dpath_mulcore_booth_b7_in1[2]), .Y(n18044));
INVX1 mul_U14455(.A(n18044), .Y(n4374));
AND2X1 mul_U14456(.A(n18049), .B(dpath_mulcore_booth_b6_in1[2]), .Y(n18048));
INVX1 mul_U14457(.A(n18048), .Y(n4375));
AND2X1 mul_U14458(.A(n18053), .B(dpath_mulcore_booth_b5_in1[2]), .Y(n18052));
INVX1 mul_U14459(.A(n18052), .Y(n4376));
AND2X1 mul_U14460(.A(n18057), .B(dpath_mulcore_booth_b4_in1[2]), .Y(n18056));
INVX1 mul_U14461(.A(n18056), .Y(n4377));
AND2X1 mul_U14462(.A(n18061), .B(dpath_mulcore_booth_b3_in1[2]), .Y(n18060));
INVX1 mul_U14463(.A(n18060), .Y(n4378));
AND2X1 mul_U14464(.A(n18065), .B(dpath_mulcore_booth_b2_in1[2]), .Y(n18064));
INVX1 mul_U14465(.A(n18064), .Y(n4379));
AND2X1 mul_U14466(.A(n5439), .B(dpath_mulcore_booth_b1_in1[2]), .Y(n18068));
INVX1 mul_U14467(.A(n18068), .Y(n4380));
AND2X1 mul_U14468(.A(dpath_mulcore_booth_b[48]), .B(n10096), .Y(n18076));
INVX1 mul_U14469(.A(n18076), .Y(n4381));
AND2X1 mul_U14470(.A(dpath_mulcore_booth_b7_in1[2]), .B(n10097), .Y(n18078));
INVX1 mul_U14471(.A(n18078), .Y(n4382));
AND2X1 mul_U14472(.A(dpath_mulcore_booth_b15_in1[2]), .B(n10109), .Y(n18080));
INVX1 mul_U14473(.A(n18080), .Y(n4383));
AND2X1 mul_U14474(.A(dpath_mulcore_booth_b[62]), .B(n10108), .Y(n18082));
INVX1 mul_U14475(.A(n18082), .Y(n4384));
AND2X1 mul_U14476(.A(dpath_mulcore_booth_b14_in1[2]), .B(n10107), .Y(n18084));
INVX1 mul_U14477(.A(n18084), .Y(n4385));
AND2X1 mul_U14478(.A(dpath_mulcore_booth_b[60]), .B(n10106), .Y(n18086));
INVX1 mul_U14479(.A(n18086), .Y(n4386));
AND2X1 mul_U14480(.A(dpath_mulcore_booth_b13_in1[2]), .B(n10105), .Y(n18088));
INVX1 mul_U14481(.A(n18088), .Y(n4387));
AND2X1 mul_U14482(.A(dpath_mulcore_booth_b[58]), .B(n10104), .Y(n18090));
INVX1 mul_U14483(.A(n18090), .Y(n4388));
AND2X1 mul_U14484(.A(dpath_mulcore_booth_b12_in1[2]), .B(n10103), .Y(n18092));
INVX1 mul_U14485(.A(n18092), .Y(n4389));
AND2X1 mul_U14486(.A(dpath_mulcore_booth_b[56]), .B(n10102), .Y(n18094));
INVX1 mul_U14487(.A(n18094), .Y(n4390));
AND2X1 mul_U14488(.A(dpath_mulcore_booth_b11_in1[2]), .B(n10101), .Y(n18096));
INVX1 mul_U14489(.A(n18096), .Y(n4391));
AND2X1 mul_U14490(.A(dpath_mulcore_booth_b[54]), .B(n10100), .Y(n18098));
INVX1 mul_U14491(.A(n18098), .Y(n4392));
AND2X1 mul_U14492(.A(dpath_mulcore_booth_b10_in1[2]), .B(n10099), .Y(n18100));
INVX1 mul_U14493(.A(n18100), .Y(n4393));
AND2X1 mul_U14494(.A(dpath_mulcore_booth_b[52]), .B(n10098), .Y(n18102));
INVX1 mul_U14495(.A(n18102), .Y(n4394));
AND2X1 mul_U14496(.A(dpath_mulcore_booth_b[50]), .B(n10097), .Y(n18106));
INVX1 mul_U14497(.A(n18106), .Y(n4395));
AND2X1 mul_U14498(.A(n18109), .B(dpath_mulcore_booth_b15_in1[2]), .Y(n18108));
INVX1 mul_U14499(.A(n18108), .Y(n4396));
AND2X1 mul_U14500(.A(n18113), .B(dpath_mulcore_booth_b14_in1[2]), .Y(n18112));
INVX1 mul_U14501(.A(n18112), .Y(n4397));
AND2X1 mul_U14502(.A(n18117), .B(dpath_mulcore_booth_b13_in1[2]), .Y(n18116));
INVX1 mul_U14503(.A(n18116), .Y(n4398));
AND2X1 mul_U14504(.A(n18121), .B(dpath_mulcore_booth_b12_in1[2]), .Y(n18120));
INVX1 mul_U14505(.A(n18120), .Y(n4399));
AND2X1 mul_U14506(.A(n18125), .B(dpath_mulcore_booth_b11_in1[2]), .Y(n18124));
INVX1 mul_U14507(.A(n18124), .Y(n4400));
AND2X1 mul_U14508(.A(n18129), .B(dpath_mulcore_booth_b10_in1[2]), .Y(n18128));
INVX1 mul_U14509(.A(n18128), .Y(n4401));
AND2X1 mul_U14510(.A(n5465), .B(dpath_mulcore_booth_b9_in1[2]), .Y(n18132));
INVX1 mul_U14511(.A(n18132), .Y(n4402));
AND2X1 mul_U14512(.A(n18137), .B(dpath_mulcore_booth_b[48]), .Y(n18136));
INVX1 mul_U14513(.A(n18136), .Y(n4403));
AND2X1 mul_U14514(.A(n6089), .B(n9713), .Y(dpath_mulcore_array2_sh_82__n3));
INVX1 mul_U14515(.A(dpath_mulcore_array2_sh_82__n3), .Y(n4404));
AND2X1 mul_U14516(.A(n8068), .B(dpath_mulcore_ary1_a0_sc2_2_70__n1), .Y(dpath_mulcore_ary1_a0_sc2_2_70__n3));
INVX1 mul_U14517(.A(dpath_mulcore_ary1_a0_sc2_2_70__n3), .Y(n4405));
AND2X1 mul_U14518(.A(dpath_mulcore_ary1_a0_s1[65]), .B(dpath_mulcore_ary1_a0_sc3_71__n4), .Y(dpath_mulcore_ary1_a0_sc3_71__n3));
INVX1 mul_U14519(.A(dpath_mulcore_ary1_a0_sc3_71__n3), .Y(n4406));
AND2X1 mul_U14520(.A(dpath_mulcore_booth_b7_in0[2]), .B(n9791), .Y(dpath_mulcore_booth_encode0_a_n20));
INVX1 mul_U14521(.A(dpath_mulcore_booth_encode0_a_n20), .Y(n4407));
AND2X1 mul_U14522(.A(dpath_mul_op2_d[14]), .B(n9790), .Y(dpath_mulcore_booth_encode0_a_n22));
INVX1 mul_U14523(.A(dpath_mulcore_booth_encode0_a_n22), .Y(n4408));
AND2X1 mul_U14524(.A(dpath_mulcore_booth_b6_in0[2]), .B(n9789), .Y(dpath_mulcore_booth_encode0_a_n24));
INVX1 mul_U14525(.A(dpath_mulcore_booth_encode0_a_n24), .Y(n4409));
AND2X1 mul_U14526(.A(dpath_mul_op2_d[12]), .B(n9788), .Y(dpath_mulcore_booth_encode0_a_n26));
INVX1 mul_U14527(.A(dpath_mulcore_booth_encode0_a_n26), .Y(n4410));
AND2X1 mul_U14528(.A(dpath_mulcore_booth_b5_in0[2]), .B(n9787), .Y(dpath_mulcore_booth_encode0_a_n28));
INVX1 mul_U14529(.A(dpath_mulcore_booth_encode0_a_n28), .Y(n4411));
AND2X1 mul_U14530(.A(dpath_mul_op2_d[10]), .B(n9813), .Y(dpath_mulcore_booth_encode0_a_n30));
INVX1 mul_U14531(.A(dpath_mulcore_booth_encode0_a_n30), .Y(n4412));
AND2X1 mul_U14532(.A(dpath_mulcore_booth_b4_in0[2]), .B(n9812), .Y(dpath_mulcore_booth_encode0_a_n32));
INVX1 mul_U14533(.A(dpath_mulcore_booth_encode0_a_n32), .Y(n4413));
AND2X1 mul_U14534(.A(dpath_mul_op2_d[8]), .B(n9811), .Y(dpath_mulcore_booth_encode0_a_n34));
INVX1 mul_U14535(.A(dpath_mulcore_booth_encode0_a_n34), .Y(n4414));
AND2X1 mul_U14536(.A(dpath_mulcore_booth_b3_in0[2]), .B(n9810), .Y(dpath_mulcore_booth_encode0_a_n36));
INVX1 mul_U14537(.A(dpath_mulcore_booth_encode0_a_n36), .Y(n4415));
AND2X1 mul_U14538(.A(dpath_mul_op2_d[6]), .B(n9809), .Y(dpath_mulcore_booth_encode0_a_n38));
INVX1 mul_U14539(.A(dpath_mulcore_booth_encode0_a_n38), .Y(n4416));
AND2X1 mul_U14540(.A(dpath_mulcore_booth_b2_in0[2]), .B(n9808), .Y(dpath_mulcore_booth_encode0_a_n40));
INVX1 mul_U14541(.A(dpath_mulcore_booth_encode0_a_n40), .Y(n4417));
AND2X1 mul_U14542(.A(dpath_mul_op2_d[4]), .B(n9807), .Y(dpath_mulcore_booth_encode0_a_n42));
INVX1 mul_U14543(.A(dpath_mulcore_booth_encode0_a_n42), .Y(n4418));
AND2X1 mul_U14544(.A(dpath_mul_op2_d[2]), .B(n9795), .Y(dpath_mulcore_booth_encode0_a_n46));
INVX1 mul_U14545(.A(dpath_mulcore_booth_encode0_a_n46), .Y(n4419));
AND2X1 mul_U14546(.A(dpath_mulcore_booth_encode0_a_n49), .B(dpath_mulcore_booth_b7_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n48));
INVX1 mul_U14547(.A(dpath_mulcore_booth_encode0_a_n48), .Y(n4420));
AND2X1 mul_U14548(.A(dpath_mulcore_booth_encode0_a_n53), .B(dpath_mulcore_booth_b6_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n52));
INVX1 mul_U14549(.A(dpath_mulcore_booth_encode0_a_n52), .Y(n4421));
AND2X1 mul_U14550(.A(dpath_mulcore_booth_encode0_a_n57), .B(dpath_mulcore_booth_b5_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n56));
INVX1 mul_U14551(.A(dpath_mulcore_booth_encode0_a_n56), .Y(n4422));
AND2X1 mul_U14552(.A(dpath_mulcore_booth_encode0_a_n61), .B(dpath_mulcore_booth_b4_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n60));
INVX1 mul_U14553(.A(dpath_mulcore_booth_encode0_a_n60), .Y(n4423));
AND2X1 mul_U14554(.A(dpath_mulcore_booth_encode0_a_n65), .B(dpath_mulcore_booth_b3_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n64));
INVX1 mul_U14555(.A(dpath_mulcore_booth_encode0_a_n64), .Y(n4424));
AND2X1 mul_U14556(.A(dpath_mulcore_booth_encode0_a_n69), .B(dpath_mulcore_booth_b2_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n68));
INVX1 mul_U14557(.A(dpath_mulcore_booth_encode0_a_n68), .Y(n4425));
AND2X1 mul_U14558(.A(n5496), .B(dpath_mulcore_booth_b1_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n72));
INVX1 mul_U14559(.A(dpath_mulcore_booth_encode0_a_n72), .Y(n4426));
AND2X1 mul_U14560(.A(spu_mul_op2_data[9]), .B(dpath_n141), .Y(dpath_n140));
INVX1 mul_U14561(.A(dpath_n140), .Y(n4427));
AND2X1 mul_U14562(.A(dpath_acc_reg[9]), .B(n7196), .Y(dpath_n143));
INVX1 mul_U14563(.A(dpath_n143), .Y(n4428));
AND2X1 mul_U14564(.A(spu_mul_op2_data[8]), .B(n9760), .Y(dpath_n149));
INVX1 mul_U14565(.A(dpath_n149), .Y(n4429));
AND2X1 mul_U14566(.A(dpath_acc_reg[8]), .B(n7196), .Y(dpath_n151));
INVX1 mul_U14567(.A(dpath_n151), .Y(n4430));
AND2X1 mul_U14568(.A(spu_mul_op2_data[7]), .B(dpath_n141), .Y(dpath_n155));
INVX1 mul_U14569(.A(dpath_n155), .Y(n4431));
AND2X1 mul_U14570(.A(dpath_acc_reg[7]), .B(n7196), .Y(dpath_n157));
INVX1 mul_U14571(.A(dpath_n157), .Y(n4432));
AND2X1 mul_U14572(.A(spu_mul_op2_data[6]), .B(n9760), .Y(dpath_n161));
INVX1 mul_U14573(.A(dpath_n161), .Y(n4433));
AND2X1 mul_U14574(.A(dpath_acc_reg[6]), .B(n7196), .Y(dpath_n163));
INVX1 mul_U14575(.A(dpath_n163), .Y(n4434));
AND2X1 mul_U14576(.A(spu_mul_op2_data[63]), .B(dpath_n141), .Y(dpath_n167));
INVX1 mul_U14577(.A(dpath_n167), .Y(n4435));
AND2X1 mul_U14578(.A(dpath_acc_reg[63]), .B(n7196), .Y(dpath_n169));
INVX1 mul_U14579(.A(dpath_n169), .Y(n4436));
AND2X1 mul_U14580(.A(spu_mul_op2_data[62]), .B(n9760), .Y(dpath_n173));
INVX1 mul_U14581(.A(dpath_n173), .Y(n4437));
AND2X1 mul_U14582(.A(dpath_acc_reg[62]), .B(n7196), .Y(dpath_n175));
INVX1 mul_U14583(.A(dpath_n175), .Y(n4438));
AND2X1 mul_U14584(.A(spu_mul_op2_data[61]), .B(dpath_n141), .Y(dpath_n179));
INVX1 mul_U14585(.A(dpath_n179), .Y(n4439));
AND2X1 mul_U14586(.A(dpath_acc_reg[61]), .B(n7196), .Y(dpath_n181));
INVX1 mul_U14587(.A(dpath_n181), .Y(n4440));
AND2X1 mul_U14588(.A(spu_mul_op2_data[60]), .B(n9760), .Y(dpath_n185));
INVX1 mul_U14589(.A(dpath_n185), .Y(n4441));
AND2X1 mul_U14590(.A(dpath_acc_reg[60]), .B(n7196), .Y(dpath_n187));
INVX1 mul_U14591(.A(dpath_n187), .Y(n4442));
AND2X1 mul_U14592(.A(spu_mul_op2_data[5]), .B(dpath_n141), .Y(dpath_n191));
INVX1 mul_U14593(.A(dpath_n191), .Y(n4443));
AND2X1 mul_U14594(.A(dpath_acc_reg[5]), .B(n7196), .Y(dpath_n193));
INVX1 mul_U14595(.A(dpath_n193), .Y(n4444));
AND2X1 mul_U14596(.A(spu_mul_op2_data[59]), .B(n9760), .Y(dpath_n197));
INVX1 mul_U14597(.A(dpath_n197), .Y(n4445));
AND2X1 mul_U14598(.A(dpath_acc_reg[59]), .B(n7196), .Y(dpath_n199));
INVX1 mul_U14599(.A(dpath_n199), .Y(n4446));
AND2X1 mul_U14600(.A(spu_mul_op2_data[58]), .B(dpath_n141), .Y(dpath_n203));
INVX1 mul_U14601(.A(dpath_n203), .Y(n4447));
AND2X1 mul_U14602(.A(dpath_acc_reg[58]), .B(n7196), .Y(dpath_n205));
INVX1 mul_U14603(.A(dpath_n205), .Y(n4448));
AND2X1 mul_U14604(.A(spu_mul_op2_data[57]), .B(n9760), .Y(dpath_n209));
INVX1 mul_U14605(.A(dpath_n209), .Y(n4449));
AND2X1 mul_U14606(.A(dpath_acc_reg[57]), .B(n7196), .Y(dpath_n211));
INVX1 mul_U14607(.A(dpath_n211), .Y(n4450));
AND2X1 mul_U14608(.A(spu_mul_op2_data[56]), .B(dpath_n141), .Y(dpath_n215));
INVX1 mul_U14609(.A(dpath_n215), .Y(n4451));
AND2X1 mul_U14610(.A(dpath_acc_reg[56]), .B(n7196), .Y(dpath_n217));
INVX1 mul_U14611(.A(dpath_n217), .Y(n4452));
AND2X1 mul_U14612(.A(spu_mul_op2_data[55]), .B(n9760), .Y(dpath_n221));
INVX1 mul_U14613(.A(dpath_n221), .Y(n4453));
AND2X1 mul_U14614(.A(dpath_acc_reg[55]), .B(n7196), .Y(dpath_n223));
INVX1 mul_U14615(.A(dpath_n223), .Y(n4454));
AND2X1 mul_U14616(.A(spu_mul_op2_data[54]), .B(n9760), .Y(dpath_n227));
INVX1 mul_U14617(.A(dpath_n227), .Y(n4455));
AND2X1 mul_U14618(.A(dpath_acc_reg[54]), .B(n7196), .Y(dpath_n229));
INVX1 mul_U14619(.A(dpath_n229), .Y(n4456));
AND2X1 mul_U14620(.A(spu_mul_op2_data[53]), .B(n9760), .Y(dpath_n233));
INVX1 mul_U14621(.A(dpath_n233), .Y(n4457));
AND2X1 mul_U14622(.A(dpath_acc_reg[53]), .B(n7196), .Y(dpath_n235));
INVX1 mul_U14623(.A(dpath_n235), .Y(n4458));
AND2X1 mul_U14624(.A(spu_mul_op2_data[52]), .B(n9760), .Y(dpath_n239));
INVX1 mul_U14625(.A(dpath_n239), .Y(n4459));
AND2X1 mul_U14626(.A(dpath_acc_reg[52]), .B(n7196), .Y(dpath_n241));
INVX1 mul_U14627(.A(dpath_n241), .Y(n4460));
AND2X1 mul_U14628(.A(spu_mul_op2_data[51]), .B(n9760), .Y(dpath_n245));
INVX1 mul_U14629(.A(dpath_n245), .Y(n4461));
AND2X1 mul_U14630(.A(dpath_acc_reg[51]), .B(n7196), .Y(dpath_n247));
INVX1 mul_U14631(.A(dpath_n247), .Y(n4462));
AND2X1 mul_U14632(.A(spu_mul_op2_data[50]), .B(n9760), .Y(dpath_n251));
INVX1 mul_U14633(.A(dpath_n251), .Y(n4463));
AND2X1 mul_U14634(.A(dpath_acc_reg[50]), .B(n7196), .Y(dpath_n253));
INVX1 mul_U14635(.A(dpath_n253), .Y(n4464));
AND2X1 mul_U14636(.A(spu_mul_op2_data[4]), .B(n9760), .Y(dpath_n257));
INVX1 mul_U14637(.A(dpath_n257), .Y(n4465));
AND2X1 mul_U14638(.A(dpath_acc_reg[4]), .B(n7196), .Y(dpath_n259));
INVX1 mul_U14639(.A(dpath_n259), .Y(n4466));
AND2X1 mul_U14640(.A(spu_mul_op2_data[49]), .B(n9760), .Y(dpath_n263));
INVX1 mul_U14641(.A(dpath_n263), .Y(n4467));
AND2X1 mul_U14642(.A(dpath_acc_reg[49]), .B(n7196), .Y(dpath_n265));
INVX1 mul_U14643(.A(dpath_n265), .Y(n4468));
AND2X1 mul_U14644(.A(spu_mul_op2_data[48]), .B(n9760), .Y(dpath_n269));
INVX1 mul_U14645(.A(dpath_n269), .Y(n4469));
AND2X1 mul_U14646(.A(dpath_acc_reg[48]), .B(n7196), .Y(dpath_n271));
INVX1 mul_U14647(.A(dpath_n271), .Y(n4470));
AND2X1 mul_U14648(.A(spu_mul_op2_data[47]), .B(n9760), .Y(dpath_n275));
INVX1 mul_U14649(.A(dpath_n275), .Y(n4471));
AND2X1 mul_U14650(.A(dpath_acc_reg[47]), .B(n7196), .Y(dpath_n277));
INVX1 mul_U14651(.A(dpath_n277), .Y(n4472));
AND2X1 mul_U14652(.A(spu_mul_op2_data[46]), .B(n9760), .Y(dpath_n281));
INVX1 mul_U14653(.A(dpath_n281), .Y(n4473));
AND2X1 mul_U14654(.A(dpath_acc_reg[46]), .B(n7196), .Y(dpath_n283));
INVX1 mul_U14655(.A(dpath_n283), .Y(n4474));
AND2X1 mul_U14656(.A(spu_mul_op2_data[45]), .B(n9760), .Y(dpath_n287));
INVX1 mul_U14657(.A(dpath_n287), .Y(n4475));
AND2X1 mul_U14658(.A(dpath_acc_reg[45]), .B(n7196), .Y(dpath_n289));
INVX1 mul_U14659(.A(dpath_n289), .Y(n4476));
AND2X1 mul_U14660(.A(spu_mul_op2_data[44]), .B(n9760), .Y(dpath_n293));
INVX1 mul_U14661(.A(dpath_n293), .Y(n4477));
AND2X1 mul_U14662(.A(dpath_acc_reg[44]), .B(n7196), .Y(dpath_n295));
INVX1 mul_U14663(.A(dpath_n295), .Y(n4478));
AND2X1 mul_U14664(.A(spu_mul_op2_data[43]), .B(n9760), .Y(dpath_n299));
INVX1 mul_U14665(.A(dpath_n299), .Y(n4479));
AND2X1 mul_U14666(.A(dpath_acc_reg[43]), .B(n7196), .Y(dpath_n301));
INVX1 mul_U14667(.A(dpath_n301), .Y(n4480));
AND2X1 mul_U14668(.A(spu_mul_op2_data[42]), .B(n9760), .Y(dpath_n305));
INVX1 mul_U14669(.A(dpath_n305), .Y(n4481));
AND2X1 mul_U14670(.A(dpath_acc_reg[42]), .B(n7196), .Y(dpath_n307));
INVX1 mul_U14671(.A(dpath_n307), .Y(n4482));
AND2X1 mul_U14672(.A(spu_mul_op2_data[41]), .B(dpath_n141), .Y(dpath_n311));
INVX1 mul_U14673(.A(dpath_n311), .Y(n4483));
AND2X1 mul_U14674(.A(dpath_acc_reg[41]), .B(n7196), .Y(dpath_n313));
INVX1 mul_U14675(.A(dpath_n313), .Y(n4484));
AND2X1 mul_U14676(.A(spu_mul_op2_data[40]), .B(n9760), .Y(dpath_n317));
INVX1 mul_U14677(.A(dpath_n317), .Y(n4485));
AND2X1 mul_U14678(.A(dpath_acc_reg[40]), .B(n7196), .Y(dpath_n319));
INVX1 mul_U14679(.A(dpath_n319), .Y(n4486));
AND2X1 mul_U14680(.A(spu_mul_op2_data[3]), .B(dpath_n141), .Y(dpath_n323));
INVX1 mul_U14681(.A(dpath_n323), .Y(n4487));
AND2X1 mul_U14682(.A(dpath_acc_reg[3]), .B(n7196), .Y(dpath_n325));
INVX1 mul_U14683(.A(dpath_n325), .Y(n4488));
AND2X1 mul_U14684(.A(spu_mul_op2_data[39]), .B(dpath_n141), .Y(dpath_n329));
INVX1 mul_U14685(.A(dpath_n329), .Y(n4489));
AND2X1 mul_U14686(.A(dpath_acc_reg[39]), .B(n7196), .Y(dpath_n331));
INVX1 mul_U14687(.A(dpath_n331), .Y(n4490));
AND2X1 mul_U14688(.A(spu_mul_op2_data[38]), .B(n9760), .Y(dpath_n335));
INVX1 mul_U14689(.A(dpath_n335), .Y(n4491));
AND2X1 mul_U14690(.A(dpath_acc_reg[38]), .B(n7196), .Y(dpath_n337));
INVX1 mul_U14691(.A(dpath_n337), .Y(n4492));
AND2X1 mul_U14692(.A(spu_mul_op2_data[37]), .B(n9760), .Y(dpath_n341));
INVX1 mul_U14693(.A(dpath_n341), .Y(n4493));
AND2X1 mul_U14694(.A(dpath_acc_reg[37]), .B(n7196), .Y(dpath_n343));
INVX1 mul_U14695(.A(dpath_n343), .Y(n4494));
AND2X1 mul_U14696(.A(spu_mul_op2_data[36]), .B(dpath_n141), .Y(dpath_n347));
INVX1 mul_U14697(.A(dpath_n347), .Y(n4495));
AND2X1 mul_U14698(.A(dpath_acc_reg[36]), .B(n7196), .Y(dpath_n349));
INVX1 mul_U14699(.A(dpath_n349), .Y(n4496));
AND2X1 mul_U14700(.A(spu_mul_op2_data[35]), .B(n9760), .Y(dpath_n353));
INVX1 mul_U14701(.A(dpath_n353), .Y(n4497));
AND2X1 mul_U14702(.A(dpath_acc_reg[35]), .B(n7196), .Y(dpath_n355));
INVX1 mul_U14703(.A(dpath_n355), .Y(n4498));
AND2X1 mul_U14704(.A(spu_mul_op2_data[34]), .B(dpath_n141), .Y(dpath_n359));
INVX1 mul_U14705(.A(dpath_n359), .Y(n4499));
AND2X1 mul_U14706(.A(dpath_acc_reg[34]), .B(n7196), .Y(dpath_n361));
INVX1 mul_U14707(.A(dpath_n361), .Y(n4500));
AND2X1 mul_U14708(.A(spu_mul_op2_data[33]), .B(dpath_n141), .Y(dpath_n365));
INVX1 mul_U14709(.A(dpath_n365), .Y(n4501));
AND2X1 mul_U14710(.A(dpath_acc_reg[33]), .B(n7196), .Y(dpath_n367));
INVX1 mul_U14711(.A(dpath_n367), .Y(n4502));
AND2X1 mul_U14712(.A(spu_mul_op2_data[32]), .B(n9760), .Y(dpath_n371));
INVX1 mul_U14713(.A(dpath_n371), .Y(n4503));
AND2X1 mul_U14714(.A(dpath_acc_reg[32]), .B(n7196), .Y(dpath_n373));
INVX1 mul_U14715(.A(dpath_n373), .Y(n4504));
AND2X1 mul_U14716(.A(spu_mul_op2_data[31]), .B(dpath_n141), .Y(dpath_n377));
INVX1 mul_U14717(.A(dpath_n377), .Y(n4505));
AND2X1 mul_U14718(.A(dpath_acc_reg[31]), .B(n7196), .Y(dpath_n379));
INVX1 mul_U14719(.A(dpath_n379), .Y(n4506));
AND2X1 mul_U14720(.A(spu_mul_op2_data[30]), .B(dpath_n141), .Y(dpath_n383));
INVX1 mul_U14721(.A(dpath_n383), .Y(n4507));
AND2X1 mul_U14722(.A(dpath_acc_reg[30]), .B(n7196), .Y(dpath_n385));
INVX1 mul_U14723(.A(dpath_n385), .Y(n4508));
AND2X1 mul_U14724(.A(spu_mul_op2_data[2]), .B(dpath_n141), .Y(dpath_n389));
INVX1 mul_U14725(.A(dpath_n389), .Y(n4509));
AND2X1 mul_U14726(.A(dpath_acc_reg[2]), .B(n7196), .Y(dpath_n391));
INVX1 mul_U14727(.A(dpath_n391), .Y(n4510));
AND2X1 mul_U14728(.A(spu_mul_op2_data[29]), .B(dpath_n141), .Y(dpath_n395));
INVX1 mul_U14729(.A(dpath_n395), .Y(n4511));
AND2X1 mul_U14730(.A(dpath_acc_reg[29]), .B(n7196), .Y(dpath_n397));
INVX1 mul_U14731(.A(dpath_n397), .Y(n4512));
AND2X1 mul_U14732(.A(spu_mul_op2_data[28]), .B(dpath_n141), .Y(dpath_n401));
INVX1 mul_U14733(.A(dpath_n401), .Y(n4513));
AND2X1 mul_U14734(.A(dpath_acc_reg[28]), .B(n7196), .Y(dpath_n403));
INVX1 mul_U14735(.A(dpath_n403), .Y(n4514));
AND2X1 mul_U14736(.A(spu_mul_op2_data[27]), .B(dpath_n141), .Y(dpath_n407));
INVX1 mul_U14737(.A(dpath_n407), .Y(n4515));
AND2X1 mul_U14738(.A(dpath_acc_reg[27]), .B(n7196), .Y(dpath_n409));
INVX1 mul_U14739(.A(dpath_n409), .Y(n4516));
AND2X1 mul_U14740(.A(spu_mul_op2_data[26]), .B(dpath_n141), .Y(dpath_n413));
INVX1 mul_U14741(.A(dpath_n413), .Y(n4517));
AND2X1 mul_U14742(.A(dpath_acc_reg[26]), .B(n7196), .Y(dpath_n415));
INVX1 mul_U14743(.A(dpath_n415), .Y(n4518));
AND2X1 mul_U14744(.A(spu_mul_op2_data[25]), .B(n9760), .Y(dpath_n419));
INVX1 mul_U14745(.A(dpath_n419), .Y(n4519));
AND2X1 mul_U14746(.A(dpath_acc_reg[25]), .B(n7196), .Y(dpath_n421));
INVX1 mul_U14747(.A(dpath_n421), .Y(n4520));
AND2X1 mul_U14748(.A(spu_mul_op2_data[24]), .B(dpath_n141), .Y(dpath_n425));
INVX1 mul_U14749(.A(dpath_n425), .Y(n4521));
AND2X1 mul_U14750(.A(dpath_acc_reg[24]), .B(n7196), .Y(dpath_n427));
INVX1 mul_U14751(.A(dpath_n427), .Y(n4522));
AND2X1 mul_U14752(.A(spu_mul_op2_data[23]), .B(n9760), .Y(dpath_n431));
INVX1 mul_U14753(.A(dpath_n431), .Y(n4523));
AND2X1 mul_U14754(.A(dpath_acc_reg[23]), .B(n7196), .Y(dpath_n433));
INVX1 mul_U14755(.A(dpath_n433), .Y(n4524));
AND2X1 mul_U14756(.A(spu_mul_op2_data[22]), .B(n9760), .Y(dpath_n437));
INVX1 mul_U14757(.A(dpath_n437), .Y(n4525));
AND2X1 mul_U14758(.A(dpath_acc_reg[22]), .B(n7196), .Y(dpath_n439));
INVX1 mul_U14759(.A(dpath_n439), .Y(n4526));
AND2X1 mul_U14760(.A(spu_mul_op2_data[21]), .B(dpath_n141), .Y(dpath_n443));
INVX1 mul_U14761(.A(dpath_n443), .Y(n4527));
AND2X1 mul_U14762(.A(dpath_acc_reg[21]), .B(n7196), .Y(dpath_n445));
INVX1 mul_U14763(.A(dpath_n445), .Y(n4528));
AND2X1 mul_U14764(.A(spu_mul_op2_data[20]), .B(dpath_n141), .Y(dpath_n449));
INVX1 mul_U14765(.A(dpath_n449), .Y(n4529));
AND2X1 mul_U14766(.A(dpath_acc_reg[20]), .B(n7196), .Y(dpath_n451));
INVX1 mul_U14767(.A(dpath_n451), .Y(n4530));
AND2X1 mul_U14768(.A(spu_mul_op2_data[1]), .B(dpath_n141), .Y(dpath_n455));
INVX1 mul_U14769(.A(dpath_n455), .Y(n4531));
AND2X1 mul_U14770(.A(dpath_acc_reg[1]), .B(n7196), .Y(dpath_n457));
INVX1 mul_U14771(.A(dpath_n457), .Y(n4532));
AND2X1 mul_U14772(.A(spu_mul_op2_data[19]), .B(dpath_n141), .Y(dpath_n461));
INVX1 mul_U14773(.A(dpath_n461), .Y(n4533));
AND2X1 mul_U14774(.A(dpath_acc_reg[19]), .B(n7196), .Y(dpath_n463));
INVX1 mul_U14775(.A(dpath_n463), .Y(n4534));
AND2X1 mul_U14776(.A(spu_mul_op2_data[18]), .B(dpath_n141), .Y(dpath_n467));
INVX1 mul_U14777(.A(dpath_n467), .Y(n4535));
AND2X1 mul_U14778(.A(dpath_acc_reg[18]), .B(n7196), .Y(dpath_n469));
INVX1 mul_U14779(.A(dpath_n469), .Y(n4536));
AND2X1 mul_U14780(.A(spu_mul_op2_data[17]), .B(dpath_n141), .Y(dpath_n473));
INVX1 mul_U14781(.A(dpath_n473), .Y(n4537));
AND2X1 mul_U14782(.A(dpath_acc_reg[17]), .B(n7196), .Y(dpath_n475));
INVX1 mul_U14783(.A(dpath_n475), .Y(n4538));
AND2X1 mul_U14784(.A(spu_mul_op2_data[16]), .B(dpath_n141), .Y(dpath_n479));
INVX1 mul_U14785(.A(dpath_n479), .Y(n4539));
AND2X1 mul_U14786(.A(dpath_acc_reg[16]), .B(n7196), .Y(dpath_n481));
INVX1 mul_U14787(.A(dpath_n481), .Y(n4540));
AND2X1 mul_U14788(.A(spu_mul_op2_data[15]), .B(dpath_n141), .Y(dpath_n485));
INVX1 mul_U14789(.A(dpath_n485), .Y(n4541));
AND2X1 mul_U14790(.A(dpath_acc_reg[15]), .B(n7196), .Y(dpath_n487));
INVX1 mul_U14791(.A(dpath_n487), .Y(n4542));
AND2X1 mul_U14792(.A(spu_mul_op2_data[14]), .B(n9760), .Y(dpath_n491));
INVX1 mul_U14793(.A(dpath_n491), .Y(n4543));
AND2X1 mul_U14794(.A(dpath_acc_reg[14]), .B(n7196), .Y(dpath_n493));
INVX1 mul_U14795(.A(dpath_n493), .Y(n4544));
AND2X1 mul_U14796(.A(spu_mul_op2_data[13]), .B(dpath_n141), .Y(dpath_n497));
INVX1 mul_U14797(.A(dpath_n497), .Y(n4545));
AND2X1 mul_U14798(.A(dpath_acc_reg[13]), .B(n7196), .Y(dpath_n499));
INVX1 mul_U14799(.A(dpath_n499), .Y(n4546));
AND2X1 mul_U14800(.A(spu_mul_op2_data[12]), .B(dpath_n141), .Y(dpath_n503));
INVX1 mul_U14801(.A(dpath_n503), .Y(n4547));
AND2X1 mul_U14802(.A(dpath_acc_reg[12]), .B(n7196), .Y(dpath_n505));
INVX1 mul_U14803(.A(dpath_n505), .Y(n4548));
AND2X1 mul_U14804(.A(spu_mul_op2_data[11]), .B(dpath_n141), .Y(dpath_n509));
INVX1 mul_U14805(.A(dpath_n509), .Y(n4549));
AND2X1 mul_U14806(.A(dpath_acc_reg[11]), .B(n7196), .Y(dpath_n511));
INVX1 mul_U14807(.A(dpath_n511), .Y(n4550));
AND2X1 mul_U14808(.A(spu_mul_op2_data[10]), .B(n9760), .Y(dpath_n515));
INVX1 mul_U14809(.A(dpath_n515), .Y(n4551));
AND2X1 mul_U14810(.A(dpath_acc_reg[10]), .B(n7196), .Y(dpath_n517));
INVX1 mul_U14811(.A(dpath_n517), .Y(n4552));
AND2X1 mul_U14812(.A(spu_mul_op2_data[0]), .B(n9760), .Y(dpath_n521));
INVX1 mul_U14813(.A(dpath_n521), .Y(n4553));
AND2X1 mul_U14814(.A(dpath_acc_reg[0]), .B(n7196), .Y(dpath_n524));
INVX1 mul_U14815(.A(dpath_n524), .Y(n4554));
AND2X1 mul_U14816(.A(n7197), .B(dpath_acc_reg[41]), .Y(dpath_n656));
INVX1 mul_U14817(.A(dpath_n656), .Y(n4555));
AND2X1 mul_U14818(.A(dpath_n661), .B(dpath_mout[41]), .Y(dpath_n660));
INVX1 mul_U14819(.A(dpath_n660), .Y(n4556));
AND2X1 mul_U14820(.A(dpath_acc_reg[128]), .B(dpath_n665), .Y(dpath_n664));
INVX1 mul_U14821(.A(dpath_n664), .Y(n4557));
AND2X1 mul_U14822(.A(dpath_acc_reg[127]), .B(dpath_n665), .Y(dpath_n668));
INVX1 mul_U14823(.A(dpath_n668), .Y(n4558));
AND2X1 mul_U14824(.A(dpath_acc_reg[126]), .B(dpath_n665), .Y(dpath_n670));
INVX1 mul_U14825(.A(dpath_n670), .Y(n4559));
AND2X1 mul_U14826(.A(dpath_acc_reg[125]), .B(dpath_n665), .Y(dpath_n672));
INVX1 mul_U14827(.A(dpath_n672), .Y(n4560));
AND2X1 mul_U14828(.A(dpath_acc_reg[124]), .B(dpath_n665), .Y(dpath_n674));
INVX1 mul_U14829(.A(dpath_n674), .Y(n4561));
AND2X1 mul_U14830(.A(dpath_acc_reg[123]), .B(n9765), .Y(dpath_n676));
INVX1 mul_U14831(.A(dpath_n676), .Y(n4562));
AND2X1 mul_U14832(.A(dpath_acc_reg[122]), .B(n9765), .Y(dpath_n678));
INVX1 mul_U14833(.A(dpath_n678), .Y(n4563));
AND2X1 mul_U14834(.A(n7197), .B(dpath_acc_reg[40]), .Y(dpath_n682));
INVX1 mul_U14835(.A(dpath_n682), .Y(n4564));
AND2X1 mul_U14836(.A(dpath_n661), .B(dpath_mout[40]), .Y(dpath_n684));
INVX1 mul_U14837(.A(dpath_n684), .Y(n4565));
AND2X1 mul_U14838(.A(dpath_acc_reg[121]), .B(dpath_n665), .Y(dpath_n686));
INVX1 mul_U14839(.A(dpath_n686), .Y(n4566));
AND2X1 mul_U14840(.A(dpath_acc_reg[120]), .B(n9765), .Y(dpath_n688));
INVX1 mul_U14841(.A(dpath_n688), .Y(n4567));
AND2X1 mul_U14842(.A(dpath_acc_reg[119]), .B(n9765), .Y(dpath_n690));
INVX1 mul_U14843(.A(dpath_n690), .Y(n4568));
AND2X1 mul_U14844(.A(dpath_acc_reg[118]), .B(dpath_n665), .Y(dpath_n692));
INVX1 mul_U14845(.A(dpath_n692), .Y(n4569));
AND2X1 mul_U14846(.A(dpath_acc_reg[117]), .B(dpath_n665), .Y(dpath_n694));
INVX1 mul_U14847(.A(dpath_n694), .Y(n4570));
AND2X1 mul_U14848(.A(dpath_acc_reg[116]), .B(dpath_n665), .Y(dpath_n696));
INVX1 mul_U14849(.A(dpath_n696), .Y(n4571));
AND2X1 mul_U14850(.A(dpath_acc_reg[115]), .B(dpath_n665), .Y(dpath_n698));
INVX1 mul_U14851(.A(dpath_n698), .Y(n4572));
AND2X1 mul_U14852(.A(dpath_acc_reg[114]), .B(dpath_n665), .Y(dpath_n700));
INVX1 mul_U14853(.A(dpath_n700), .Y(n4573));
AND2X1 mul_U14854(.A(dpath_acc_reg[113]), .B(dpath_n665), .Y(dpath_n702));
INVX1 mul_U14855(.A(dpath_n702), .Y(n4574));
AND2X1 mul_U14856(.A(dpath_acc_reg[112]), .B(dpath_n665), .Y(dpath_n704));
INVX1 mul_U14857(.A(dpath_n704), .Y(n4575));
AND2X1 mul_U14858(.A(n7197), .B(dpath_acc_reg[39]), .Y(dpath_n708));
INVX1 mul_U14859(.A(dpath_n708), .Y(n4576));
AND2X1 mul_U14860(.A(dpath_n661), .B(dpath_mout[39]), .Y(dpath_n710));
INVX1 mul_U14861(.A(dpath_n710), .Y(n4577));
AND2X1 mul_U14862(.A(dpath_acc_reg[111]), .B(dpath_n665), .Y(dpath_n712));
INVX1 mul_U14863(.A(dpath_n712), .Y(n4578));
AND2X1 mul_U14864(.A(dpath_acc_reg[110]), .B(n9765), .Y(dpath_n714));
INVX1 mul_U14865(.A(dpath_n714), .Y(n4579));
AND2X1 mul_U14866(.A(dpath_acc_reg[109]), .B(n9765), .Y(dpath_n716));
INVX1 mul_U14867(.A(dpath_n716), .Y(n4580));
AND2X1 mul_U14868(.A(dpath_acc_reg[108]), .B(dpath_n665), .Y(dpath_n718));
INVX1 mul_U14869(.A(dpath_n718), .Y(n4581));
AND2X1 mul_U14870(.A(dpath_acc_reg[107]), .B(dpath_n665), .Y(dpath_n720));
INVX1 mul_U14871(.A(dpath_n720), .Y(n4582));
AND2X1 mul_U14872(.A(dpath_acc_reg[106]), .B(dpath_n665), .Y(dpath_n722));
INVX1 mul_U14873(.A(dpath_n722), .Y(n4583));
AND2X1 mul_U14874(.A(dpath_acc_reg[105]), .B(n9765), .Y(dpath_n724));
INVX1 mul_U14875(.A(dpath_n724), .Y(n4584));
AND2X1 mul_U14876(.A(dpath_acc_reg[104]), .B(dpath_n665), .Y(dpath_n726));
INVX1 mul_U14877(.A(dpath_n726), .Y(n4585));
AND2X1 mul_U14878(.A(dpath_acc_reg[103]), .B(n9765), .Y(dpath_n728));
INVX1 mul_U14879(.A(dpath_n728), .Y(n4586));
AND2X1 mul_U14880(.A(dpath_acc_reg[102]), .B(n9765), .Y(dpath_n730));
INVX1 mul_U14881(.A(dpath_n730), .Y(n4587));
AND2X1 mul_U14882(.A(n7197), .B(dpath_acc_reg[38]), .Y(dpath_n734));
INVX1 mul_U14883(.A(dpath_n734), .Y(n4588));
AND2X1 mul_U14884(.A(dpath_n661), .B(dpath_mout[38]), .Y(dpath_n736));
INVX1 mul_U14885(.A(dpath_n736), .Y(n4589));
AND2X1 mul_U14886(.A(dpath_acc_reg[101]), .B(n9765), .Y(dpath_n738));
INVX1 mul_U14887(.A(dpath_n738), .Y(n4590));
AND2X1 mul_U14888(.A(dpath_acc_reg[100]), .B(n9765), .Y(dpath_n740));
INVX1 mul_U14889(.A(dpath_n740), .Y(n4591));
AND2X1 mul_U14890(.A(dpath_acc_reg[99]), .B(n9765), .Y(dpath_n742));
INVX1 mul_U14891(.A(dpath_n742), .Y(n4592));
AND2X1 mul_U14892(.A(dpath_acc_reg[98]), .B(n9765), .Y(dpath_n744));
INVX1 mul_U14893(.A(dpath_n744), .Y(n4593));
AND2X1 mul_U14894(.A(dpath_acc_reg[97]), .B(n9765), .Y(dpath_n746));
INVX1 mul_U14895(.A(dpath_n746), .Y(n4594));
AND2X1 mul_U14896(.A(dpath_acc_reg[96]), .B(n9765), .Y(dpath_n748));
INVX1 mul_U14897(.A(dpath_n748), .Y(n4595));
AND2X1 mul_U14898(.A(dpath_acc_reg[95]), .B(n9765), .Y(dpath_n750));
INVX1 mul_U14899(.A(dpath_n750), .Y(n4596));
AND2X1 mul_U14900(.A(dpath_acc_reg[94]), .B(n9765), .Y(dpath_n752));
INVX1 mul_U14901(.A(dpath_n752), .Y(n4597));
AND2X1 mul_U14902(.A(dpath_acc_reg[93]), .B(n9765), .Y(dpath_n754));
INVX1 mul_U14903(.A(dpath_n754), .Y(n4598));
AND2X1 mul_U14904(.A(dpath_acc_reg[92]), .B(n9765), .Y(dpath_n756));
INVX1 mul_U14905(.A(dpath_n756), .Y(n4599));
AND2X1 mul_U14906(.A(n7197), .B(dpath_acc_reg[37]), .Y(dpath_n760));
INVX1 mul_U14907(.A(dpath_n760), .Y(n4600));
AND2X1 mul_U14908(.A(dpath_n661), .B(dpath_mout[37]), .Y(dpath_n762));
INVX1 mul_U14909(.A(dpath_n762), .Y(n4601));
AND2X1 mul_U14910(.A(dpath_acc_reg[91]), .B(n9765), .Y(dpath_n764));
INVX1 mul_U14911(.A(dpath_n764), .Y(n4602));
AND2X1 mul_U14912(.A(dpath_acc_reg[90]), .B(n9765), .Y(dpath_n766));
INVX1 mul_U14913(.A(dpath_n766), .Y(n4603));
AND2X1 mul_U14914(.A(dpath_acc_reg[89]), .B(n9765), .Y(dpath_n768));
INVX1 mul_U14915(.A(dpath_n768), .Y(n4604));
AND2X1 mul_U14916(.A(dpath_acc_reg[88]), .B(dpath_n665), .Y(dpath_n770));
INVX1 mul_U14917(.A(dpath_n770), .Y(n4605));
AND2X1 mul_U14918(.A(dpath_acc_reg[87]), .B(n9765), .Y(dpath_n772));
INVX1 mul_U14919(.A(dpath_n772), .Y(n4606));
AND2X1 mul_U14920(.A(dpath_acc_reg[86]), .B(dpath_n665), .Y(dpath_n774));
INVX1 mul_U14921(.A(dpath_n774), .Y(n4607));
AND2X1 mul_U14922(.A(dpath_acc_reg[85]), .B(n9765), .Y(dpath_n776));
INVX1 mul_U14923(.A(dpath_n776), .Y(n4608));
AND2X1 mul_U14924(.A(dpath_acc_reg[84]), .B(dpath_n665), .Y(dpath_n778));
INVX1 mul_U14925(.A(dpath_n778), .Y(n4609));
AND2X1 mul_U14926(.A(dpath_acc_reg[83]), .B(n9765), .Y(dpath_n780));
INVX1 mul_U14927(.A(dpath_n780), .Y(n4610));
AND2X1 mul_U14928(.A(dpath_acc_reg[82]), .B(dpath_n665), .Y(dpath_n782));
INVX1 mul_U14929(.A(dpath_n782), .Y(n4611));
AND2X1 mul_U14930(.A(n7197), .B(dpath_acc_reg[36]), .Y(dpath_n786));
INVX1 mul_U14931(.A(dpath_n786), .Y(n4612));
AND2X1 mul_U14932(.A(dpath_n661), .B(dpath_mout[36]), .Y(dpath_n788));
INVX1 mul_U14933(.A(dpath_n788), .Y(n4613));
AND2X1 mul_U14934(.A(dpath_acc_reg[81]), .B(n9765), .Y(dpath_n790));
INVX1 mul_U14935(.A(dpath_n790), .Y(n4614));
AND2X1 mul_U14936(.A(dpath_acc_reg[80]), .B(dpath_n665), .Y(dpath_n792));
INVX1 mul_U14937(.A(dpath_n792), .Y(n4615));
AND2X1 mul_U14938(.A(dpath_acc_reg[79]), .B(n9765), .Y(dpath_n794));
INVX1 mul_U14939(.A(dpath_n794), .Y(n4616));
AND2X1 mul_U14940(.A(dpath_acc_reg[78]), .B(dpath_n665), .Y(dpath_n796));
INVX1 mul_U14941(.A(dpath_n796), .Y(n4617));
AND2X1 mul_U14942(.A(dpath_acc_reg[77]), .B(n9765), .Y(dpath_n798));
INVX1 mul_U14943(.A(dpath_n798), .Y(n4618));
AND2X1 mul_U14944(.A(dpath_acc_reg[76]), .B(dpath_n665), .Y(dpath_n800));
INVX1 mul_U14945(.A(dpath_n800), .Y(n4619));
AND2X1 mul_U14946(.A(dpath_acc_reg[75]), .B(dpath_n665), .Y(dpath_n802));
INVX1 mul_U14947(.A(dpath_n802), .Y(n4620));
AND2X1 mul_U14948(.A(dpath_acc_reg[74]), .B(n9765), .Y(dpath_n804));
INVX1 mul_U14949(.A(dpath_n804), .Y(n4621));
AND2X1 mul_U14950(.A(dpath_acc_reg[73]), .B(dpath_n665), .Y(dpath_n806));
INVX1 mul_U14951(.A(dpath_n806), .Y(n4622));
AND2X1 mul_U14952(.A(dpath_acc_reg[72]), .B(dpath_n665), .Y(dpath_n808));
INVX1 mul_U14953(.A(dpath_n808), .Y(n4623));
AND2X1 mul_U14954(.A(n7197), .B(dpath_acc_reg[35]), .Y(dpath_n812));
INVX1 mul_U14955(.A(dpath_n812), .Y(n4624));
AND2X1 mul_U14956(.A(dpath_n661), .B(dpath_mout[35]), .Y(dpath_n814));
INVX1 mul_U14957(.A(dpath_n814), .Y(n4625));
AND2X1 mul_U14958(.A(dpath_acc_reg[71]), .B(n9765), .Y(dpath_n816));
INVX1 mul_U14959(.A(dpath_n816), .Y(n4626));
AND2X1 mul_U14960(.A(dpath_acc_reg[70]), .B(dpath_n665), .Y(dpath_n818));
INVX1 mul_U14961(.A(dpath_n818), .Y(n4627));
AND2X1 mul_U14962(.A(dpath_acc_reg[69]), .B(dpath_n665), .Y(dpath_n820));
INVX1 mul_U14963(.A(dpath_n820), .Y(n4628));
AND2X1 mul_U14964(.A(dpath_acc_reg[68]), .B(n9765), .Y(dpath_n822));
INVX1 mul_U14965(.A(dpath_n822), .Y(n4629));
AND2X1 mul_U14966(.A(dpath_acc_reg[67]), .B(dpath_n665), .Y(dpath_n824));
INVX1 mul_U14967(.A(dpath_n824), .Y(n4630));
AND2X1 mul_U14968(.A(dpath_acc_reg[66]), .B(n9765), .Y(dpath_n826));
INVX1 mul_U14969(.A(dpath_n826), .Y(n4631));
AND2X1 mul_U14970(.A(dpath_acc_reg[65]), .B(n9765), .Y(dpath_n828));
INVX1 mul_U14971(.A(dpath_n828), .Y(n4632));
AND2X1 mul_U14972(.A(dpath_acc_reg[64]), .B(dpath_n665), .Y(dpath_n830));
INVX1 mul_U14973(.A(dpath_n830), .Y(n4633));
AND2X1 mul_U14974(.A(n7197), .B(dpath_acc_reg[63]), .Y(dpath_n834));
INVX1 mul_U14975(.A(dpath_n834), .Y(n4634));
AND2X1 mul_U14976(.A(dpath_n661), .B(dpath_mout[63]), .Y(dpath_n836));
INVX1 mul_U14977(.A(dpath_n836), .Y(n4635));
AND2X1 mul_U14978(.A(n7197), .B(dpath_acc_reg[62]), .Y(dpath_n840));
INVX1 mul_U14979(.A(dpath_n840), .Y(n4636));
AND2X1 mul_U14980(.A(dpath_n661), .B(dpath_mout[62]), .Y(dpath_n842));
INVX1 mul_U14981(.A(dpath_n842), .Y(n4637));
AND2X1 mul_U14982(.A(n7197), .B(dpath_acc_reg[34]), .Y(dpath_n846));
INVX1 mul_U14983(.A(dpath_n846), .Y(n4638));
AND2X1 mul_U14984(.A(dpath_n661), .B(dpath_mout[34]), .Y(dpath_n848));
INVX1 mul_U14985(.A(dpath_n848), .Y(n4639));
AND2X1 mul_U14986(.A(n7197), .B(dpath_acc_reg[61]), .Y(dpath_n852));
INVX1 mul_U14987(.A(dpath_n852), .Y(n4640));
AND2X1 mul_U14988(.A(dpath_n661), .B(dpath_mout[61]), .Y(dpath_n854));
INVX1 mul_U14989(.A(dpath_n854), .Y(n4641));
AND2X1 mul_U14990(.A(n7197), .B(dpath_acc_reg[60]), .Y(dpath_n858));
INVX1 mul_U14991(.A(dpath_n858), .Y(n4642));
AND2X1 mul_U14992(.A(dpath_n661), .B(dpath_mout[60]), .Y(dpath_n860));
INVX1 mul_U14993(.A(dpath_n860), .Y(n4643));
AND2X1 mul_U14994(.A(n7197), .B(dpath_acc_reg[59]), .Y(dpath_n864));
INVX1 mul_U14995(.A(dpath_n864), .Y(n4644));
AND2X1 mul_U14996(.A(dpath_n661), .B(dpath_mout[59]), .Y(dpath_n866));
INVX1 mul_U14997(.A(dpath_n866), .Y(n4645));
AND2X1 mul_U14998(.A(n7197), .B(dpath_acc_reg[58]), .Y(dpath_n870));
INVX1 mul_U14999(.A(dpath_n870), .Y(n4646));
AND2X1 mul_U15000(.A(dpath_n661), .B(dpath_mout[58]), .Y(dpath_n872));
INVX1 mul_U15001(.A(dpath_n872), .Y(n4647));
AND2X1 mul_U15002(.A(n7197), .B(dpath_acc_reg[57]), .Y(dpath_n876));
INVX1 mul_U15003(.A(dpath_n876), .Y(n4648));
AND2X1 mul_U15004(.A(dpath_n661), .B(dpath_mout[57]), .Y(dpath_n878));
INVX1 mul_U15005(.A(dpath_n878), .Y(n4649));
AND2X1 mul_U15006(.A(n7197), .B(dpath_acc_reg[56]), .Y(dpath_n882));
INVX1 mul_U15007(.A(dpath_n882), .Y(n4650));
AND2X1 mul_U15008(.A(dpath_n661), .B(dpath_mout[56]), .Y(dpath_n884));
INVX1 mul_U15009(.A(dpath_n884), .Y(n4651));
AND2X1 mul_U15010(.A(n7197), .B(dpath_acc_reg[55]), .Y(dpath_n888));
INVX1 mul_U15011(.A(dpath_n888), .Y(n4652));
AND2X1 mul_U15012(.A(dpath_n661), .B(dpath_mout[55]), .Y(dpath_n890));
INVX1 mul_U15013(.A(dpath_n890), .Y(n4653));
AND2X1 mul_U15014(.A(n7197), .B(dpath_acc_reg[54]), .Y(dpath_n894));
INVX1 mul_U15015(.A(dpath_n894), .Y(n4654));
AND2X1 mul_U15016(.A(dpath_n661), .B(dpath_mout[54]), .Y(dpath_n896));
INVX1 mul_U15017(.A(dpath_n896), .Y(n4655));
AND2X1 mul_U15018(.A(n7197), .B(dpath_acc_reg[53]), .Y(dpath_n900));
INVX1 mul_U15019(.A(dpath_n900), .Y(n4656));
AND2X1 mul_U15020(.A(dpath_n661), .B(dpath_mout[53]), .Y(dpath_n902));
INVX1 mul_U15021(.A(dpath_n902), .Y(n4657));
AND2X1 mul_U15022(.A(n7197), .B(dpath_acc_reg[52]), .Y(dpath_n906));
INVX1 mul_U15023(.A(dpath_n906), .Y(n4658));
AND2X1 mul_U15024(.A(dpath_n661), .B(dpath_mout[52]), .Y(dpath_n908));
INVX1 mul_U15025(.A(dpath_n908), .Y(n4659));
AND2X1 mul_U15026(.A(n7197), .B(dpath_acc_reg[33]), .Y(dpath_n912));
INVX1 mul_U15027(.A(dpath_n912), .Y(n4660));
AND2X1 mul_U15028(.A(dpath_n661), .B(dpath_mout[33]), .Y(dpath_n914));
INVX1 mul_U15029(.A(dpath_n914), .Y(n4661));
AND2X1 mul_U15030(.A(n7197), .B(dpath_acc_reg[51]), .Y(dpath_n918));
INVX1 mul_U15031(.A(dpath_n918), .Y(n4662));
AND2X1 mul_U15032(.A(dpath_n661), .B(dpath_mout[51]), .Y(dpath_n920));
INVX1 mul_U15033(.A(dpath_n920), .Y(n4663));
AND2X1 mul_U15034(.A(n7197), .B(dpath_acc_reg[50]), .Y(dpath_n924));
INVX1 mul_U15035(.A(dpath_n924), .Y(n4664));
AND2X1 mul_U15036(.A(dpath_n661), .B(dpath_mout[50]), .Y(dpath_n926));
INVX1 mul_U15037(.A(dpath_n926), .Y(n4665));
AND2X1 mul_U15038(.A(n7197), .B(dpath_acc_reg[49]), .Y(dpath_n930));
INVX1 mul_U15039(.A(dpath_n930), .Y(n4666));
AND2X1 mul_U15040(.A(dpath_n661), .B(dpath_mout[49]), .Y(dpath_n932));
INVX1 mul_U15041(.A(dpath_n932), .Y(n4667));
AND2X1 mul_U15042(.A(n7197), .B(dpath_acc_reg[48]), .Y(dpath_n936));
INVX1 mul_U15043(.A(dpath_n936), .Y(n4668));
AND2X1 mul_U15044(.A(dpath_n661), .B(dpath_mout[48]), .Y(dpath_n938));
INVX1 mul_U15045(.A(dpath_n938), .Y(n4669));
AND2X1 mul_U15046(.A(n7197), .B(dpath_acc_reg[47]), .Y(dpath_n942));
INVX1 mul_U15047(.A(dpath_n942), .Y(n4670));
AND2X1 mul_U15048(.A(dpath_n661), .B(dpath_mout[47]), .Y(dpath_n944));
INVX1 mul_U15049(.A(dpath_n944), .Y(n4671));
AND2X1 mul_U15050(.A(n7197), .B(dpath_acc_reg[46]), .Y(dpath_n948));
INVX1 mul_U15051(.A(dpath_n948), .Y(n4672));
AND2X1 mul_U15052(.A(dpath_n661), .B(dpath_mout[46]), .Y(dpath_n950));
INVX1 mul_U15053(.A(dpath_n950), .Y(n4673));
AND2X1 mul_U15054(.A(n7197), .B(dpath_acc_reg[45]), .Y(dpath_n954));
INVX1 mul_U15055(.A(dpath_n954), .Y(n4674));
AND2X1 mul_U15056(.A(dpath_n661), .B(dpath_mout[45]), .Y(dpath_n956));
INVX1 mul_U15057(.A(dpath_n956), .Y(n4675));
AND2X1 mul_U15058(.A(n7197), .B(dpath_acc_reg[44]), .Y(dpath_n960));
INVX1 mul_U15059(.A(dpath_n960), .Y(n4676));
AND2X1 mul_U15060(.A(dpath_n661), .B(dpath_mout[44]), .Y(dpath_n962));
INVX1 mul_U15061(.A(dpath_n962), .Y(n4677));
AND2X1 mul_U15062(.A(n7197), .B(dpath_acc_reg[43]), .Y(dpath_n966));
INVX1 mul_U15063(.A(dpath_n966), .Y(n4678));
AND2X1 mul_U15064(.A(dpath_n661), .B(dpath_mout[43]), .Y(dpath_n968));
INVX1 mul_U15065(.A(dpath_n968), .Y(n4679));
AND2X1 mul_U15066(.A(n7197), .B(dpath_acc_reg[42]), .Y(dpath_n972));
INVX1 mul_U15067(.A(dpath_n972), .Y(n4680));
AND2X1 mul_U15068(.A(dpath_n661), .B(dpath_mout[42]), .Y(dpath_n974));
INVX1 mul_U15069(.A(dpath_n974), .Y(n4681));
AND2X1 mul_U15070(.A(n7197), .B(dpath_acc_reg[32]), .Y(dpath_n978));
INVX1 mul_U15071(.A(dpath_n978), .Y(n4682));
AND2X1 mul_U15072(.A(dpath_n661), .B(dpath_mout[32]), .Y(dpath_n982));
INVX1 mul_U15073(.A(dpath_n982), .Y(n4683));
AND2X1 mul_U15074(.A(byp_imm), .B(control_n10), .Y(control_n9));
INVX1 mul_U15075(.A(control_n9), .Y(n4684));
OR2X1 mul_U15076(.A(control_c3_act), .B(acc_reg_shf), .Y(control_n17));
INVX1 mul_U15077(.A(control_n17), .Y(n4685));
AND2X1 mul_U15078(.A(control_favor_e), .B(exu_mul_input_vld), .Y(control_n19));
INVX1 mul_U15079(.A(control_n19), .Y(n4686));
AND2X1 mul_U15080(.A(n8285), .B(n15172), .Y(n15174));
INVX1 mul_U15081(.A(n15174), .Y(n4687));
AND2X1 mul_U15082(.A(dpath_mulcore_ary1_a0_s_2[10]), .B(n15184), .Y(n15186));
INVX1 mul_U15083(.A(n15186), .Y(n4688));
AND2X1 mul_U15084(.A(n8057), .B(n15187), .Y(n15189));
INVX1 mul_U15085(.A(n15189), .Y(n4689));
AND2X1 mul_U15086(.A(dpath_mulcore_ary1_a0_c1[1]), .B(n15190), .Y(n15192));
INVX1 mul_U15087(.A(n15192), .Y(n4690));
AND2X1 mul_U15088(.A(n8294), .B(n15572), .Y(n15574));
INVX1 mul_U15089(.A(n15574), .Y(n4691));
AND2X1 mul_U15090(.A(dpath_mulcore_ary1_a1_s_2[10]), .B(n15584), .Y(n15586));
INVX1 mul_U15091(.A(n15586), .Y(n4692));
AND2X1 mul_U15092(.A(n8065), .B(n15587), .Y(n15589));
INVX1 mul_U15093(.A(n15589), .Y(n4693));
AND2X1 mul_U15094(.A(dpath_mulcore_ary1_a1_c1[1]), .B(n15590), .Y(n15592));
INVX1 mul_U15095(.A(n15592), .Y(n4694));
AND2X1 mul_U15096(.A(dpath_mulcore_array2_c2[96]), .B(n16028), .Y(n16030));
INVX1 mul_U15097(.A(n16030), .Y(n4695));
AND2X1 mul_U15098(.A(n8290), .B(n10023), .Y(n16590));
INVX1 mul_U15099(.A(n16590), .Y(n4696));
AND2X1 mul_U15100(.A(n8291), .B(n10020), .Y(n16594));
INVX1 mul_U15101(.A(n16594), .Y(n4697));
AND2X1 mul_U15102(.A(n8292), .B(n10017), .Y(n16598));
INVX1 mul_U15103(.A(n16598), .Y(n4698));
AND2X1 mul_U15104(.A(n8288), .B(n10014), .Y(n16602));
INVX1 mul_U15105(.A(n16602), .Y(n4699));
AND2X1 mul_U15106(.A(n8289), .B(n10027), .Y(n16605));
INVX1 mul_U15107(.A(n16605), .Y(n4700));
AND2X1 mul_U15108(.A(n8978), .B(n10008), .Y(n16610));
INVX1 mul_U15109(.A(n16610), .Y(n4701));
AND2X1 mul_U15110(.A(n8979), .B(n9819), .Y(n16617));
INVX1 mul_U15111(.A(n16617), .Y(n4702));
AND2X1 mul_U15112(.A(n8980), .B(n9820), .Y(n16624));
INVX1 mul_U15113(.A(n16624), .Y(n4703));
AND2X1 mul_U15114(.A(n8981), .B(n9821), .Y(n16631));
INVX1 mul_U15115(.A(n16631), .Y(n4704));
AND2X1 mul_U15116(.A(n8982), .B(n9822), .Y(n16638));
INVX1 mul_U15117(.A(n16638), .Y(n4705));
AND2X1 mul_U15118(.A(n8983), .B(n9823), .Y(n16645));
INVX1 mul_U15119(.A(n16645), .Y(n4706));
AND2X1 mul_U15120(.A(n8984), .B(n9995), .Y(n16652));
INVX1 mul_U15121(.A(n16652), .Y(n4707));
AND2X1 mul_U15122(.A(n8985), .B(n9992), .Y(n16659));
INVX1 mul_U15123(.A(n16659), .Y(n4708));
AND2X1 mul_U15124(.A(n8986), .B(n9989), .Y(n16666));
INVX1 mul_U15125(.A(n16666), .Y(n4709));
AND2X1 mul_U15126(.A(n8987), .B(n9986), .Y(n16673));
INVX1 mul_U15127(.A(n16673), .Y(n4710));
AND2X1 mul_U15128(.A(n8988), .B(n9983), .Y(n16680));
INVX1 mul_U15129(.A(n16680), .Y(n4711));
AND2X1 mul_U15130(.A(n8989), .B(n9980), .Y(n16687));
INVX1 mul_U15131(.A(n16687), .Y(n4712));
AND2X1 mul_U15132(.A(n8990), .B(n9977), .Y(n16694));
INVX1 mul_U15133(.A(n16694), .Y(n4713));
AND2X1 mul_U15134(.A(n8991), .B(n9974), .Y(n16701));
INVX1 mul_U15135(.A(n16701), .Y(n4714));
AND2X1 mul_U15136(.A(n8992), .B(n9971), .Y(n16708));
INVX1 mul_U15137(.A(n16708), .Y(n4715));
AND2X1 mul_U15138(.A(n8993), .B(n9968), .Y(n16715));
INVX1 mul_U15139(.A(n16715), .Y(n4716));
AND2X1 mul_U15140(.A(n8994), .B(n9965), .Y(n16722));
INVX1 mul_U15141(.A(n16722), .Y(n4717));
AND2X1 mul_U15142(.A(n8995), .B(n9962), .Y(n16729));
INVX1 mul_U15143(.A(n16729), .Y(n4718));
AND2X1 mul_U15144(.A(n8996), .B(n9959), .Y(n16736));
INVX1 mul_U15145(.A(n16736), .Y(n4719));
AND2X1 mul_U15146(.A(n8997), .B(n9956), .Y(n16743));
INVX1 mul_U15147(.A(n16743), .Y(n4720));
AND2X1 mul_U15148(.A(n8998), .B(n9953), .Y(n16750));
INVX1 mul_U15149(.A(n16750), .Y(n4721));
AND2X1 mul_U15150(.A(n8999), .B(n9950), .Y(n16757));
INVX1 mul_U15151(.A(n16757), .Y(n4722));
AND2X1 mul_U15152(.A(n9000), .B(n9947), .Y(n16764));
INVX1 mul_U15153(.A(n16764), .Y(n4723));
AND2X1 mul_U15154(.A(n9001), .B(n9944), .Y(n16771));
INVX1 mul_U15155(.A(n16771), .Y(n4724));
AND2X1 mul_U15156(.A(n9002), .B(n9941), .Y(n16778));
INVX1 mul_U15157(.A(n16778), .Y(n4725));
AND2X1 mul_U15158(.A(n9003), .B(n9938), .Y(n16785));
INVX1 mul_U15159(.A(n16785), .Y(n4726));
AND2X1 mul_U15160(.A(n9004), .B(n9935), .Y(n16792));
INVX1 mul_U15161(.A(n16792), .Y(n4727));
AND2X1 mul_U15162(.A(n9005), .B(n9932), .Y(n16799));
INVX1 mul_U15163(.A(n16799), .Y(n4728));
AND2X1 mul_U15164(.A(n9006), .B(n9929), .Y(n16806));
INVX1 mul_U15165(.A(n16806), .Y(n4729));
AND2X1 mul_U15166(.A(n9007), .B(n9926), .Y(n16813));
INVX1 mul_U15167(.A(n16813), .Y(n4730));
AND2X1 mul_U15168(.A(n9008), .B(n9923), .Y(n16820));
INVX1 mul_U15169(.A(n16820), .Y(n4731));
AND2X1 mul_U15170(.A(n9009), .B(n9920), .Y(n16827));
INVX1 mul_U15171(.A(n16827), .Y(n4732));
AND2X1 mul_U15172(.A(n9010), .B(n9917), .Y(n16834));
INVX1 mul_U15173(.A(n16834), .Y(n4733));
AND2X1 mul_U15174(.A(n9011), .B(n9914), .Y(n16841));
INVX1 mul_U15175(.A(n16841), .Y(n4734));
AND2X1 mul_U15176(.A(n9012), .B(n9911), .Y(n16848));
INVX1 mul_U15177(.A(n16848), .Y(n4735));
AND2X1 mul_U15178(.A(n9013), .B(n9908), .Y(n16855));
INVX1 mul_U15179(.A(n16855), .Y(n4736));
AND2X1 mul_U15180(.A(n9014), .B(n9905), .Y(n16862));
INVX1 mul_U15181(.A(n16862), .Y(n4737));
AND2X1 mul_U15182(.A(n9015), .B(n9902), .Y(n16869));
INVX1 mul_U15183(.A(n16869), .Y(n4738));
AND2X1 mul_U15184(.A(n9016), .B(n9899), .Y(n16876));
INVX1 mul_U15185(.A(n16876), .Y(n4739));
AND2X1 mul_U15186(.A(n9017), .B(n9896), .Y(n16883));
INVX1 mul_U15187(.A(n16883), .Y(n4740));
AND2X1 mul_U15188(.A(n9018), .B(n9893), .Y(n16890));
INVX1 mul_U15189(.A(n16890), .Y(n4741));
AND2X1 mul_U15190(.A(n9019), .B(n9890), .Y(n16897));
INVX1 mul_U15191(.A(n16897), .Y(n4742));
AND2X1 mul_U15192(.A(n9020), .B(n9887), .Y(n16904));
INVX1 mul_U15193(.A(n16904), .Y(n4743));
AND2X1 mul_U15194(.A(n9021), .B(n9884), .Y(n16911));
INVX1 mul_U15195(.A(n16911), .Y(n4744));
AND2X1 mul_U15196(.A(n9022), .B(n9881), .Y(n16918));
INVX1 mul_U15197(.A(n16918), .Y(n4745));
AND2X1 mul_U15198(.A(n9023), .B(n9878), .Y(n16925));
INVX1 mul_U15199(.A(n16925), .Y(n4746));
AND2X1 mul_U15200(.A(n9024), .B(n9875), .Y(n16932));
INVX1 mul_U15201(.A(n16932), .Y(n4747));
AND2X1 mul_U15202(.A(n9025), .B(n9872), .Y(n16939));
INVX1 mul_U15203(.A(n16939), .Y(n4748));
AND2X1 mul_U15204(.A(n9026), .B(n9869), .Y(n16946));
INVX1 mul_U15205(.A(n16946), .Y(n4749));
AND2X1 mul_U15206(.A(n9027), .B(n9866), .Y(n16953));
INVX1 mul_U15207(.A(n16953), .Y(n4750));
AND2X1 mul_U15208(.A(n9028), .B(n9863), .Y(n16960));
INVX1 mul_U15209(.A(n16960), .Y(n4751));
AND2X1 mul_U15210(.A(n9029), .B(n9860), .Y(n16967));
INVX1 mul_U15211(.A(n16967), .Y(n4752));
AND2X1 mul_U15212(.A(n9030), .B(n9857), .Y(n16974));
INVX1 mul_U15213(.A(n16974), .Y(n4753));
AND2X1 mul_U15214(.A(n9031), .B(n9849), .Y(n16981));
INVX1 mul_U15215(.A(n16981), .Y(n4754));
AND2X1 mul_U15216(.A(n9032), .B(n9850), .Y(n16988));
INVX1 mul_U15217(.A(n16988), .Y(n4755));
AND2X1 mul_U15218(.A(n9033), .B(n9851), .Y(n16995));
INVX1 mul_U15219(.A(n16995), .Y(n4756));
AND2X1 mul_U15220(.A(n9034), .B(n9852), .Y(n17002));
INVX1 mul_U15221(.A(n17002), .Y(n4757));
AND2X1 mul_U15222(.A(n9035), .B(n9846), .Y(n17009));
INVX1 mul_U15223(.A(n17009), .Y(n4758));
AND2X1 mul_U15224(.A(n9036), .B(n9847), .Y(n17016));
INVX1 mul_U15225(.A(n17016), .Y(n4759));
AND2X1 mul_U15226(.A(n9038), .B(n10007), .Y(n17029));
INVX1 mul_U15227(.A(n17029), .Y(n4760));
AND2X1 mul_U15228(.A(n8299), .B(n10019), .Y(n17034));
INVX1 mul_U15229(.A(n17034), .Y(n4761));
AND2X1 mul_U15230(.A(n8300), .B(n10016), .Y(n17038));
INVX1 mul_U15231(.A(n17038), .Y(n4762));
AND2X1 mul_U15232(.A(n8301), .B(n10013), .Y(n17042));
INVX1 mul_U15233(.A(n17042), .Y(n4763));
AND2X1 mul_U15234(.A(n8297), .B(n10010), .Y(n17046));
INVX1 mul_U15235(.A(n17046), .Y(n4764));
AND2X1 mul_U15236(.A(n8298), .B(n10022), .Y(n17049));
INVX1 mul_U15237(.A(n17049), .Y(n4765));
AND2X1 mul_U15238(.A(n9039), .B(n10005), .Y(n17054));
INVX1 mul_U15239(.A(n17054), .Y(n4766));
AND2X1 mul_U15240(.A(n9040), .B(n10003), .Y(n17061));
INVX1 mul_U15241(.A(n17061), .Y(n4767));
AND2X1 mul_U15242(.A(n9041), .B(n10001), .Y(n17068));
INVX1 mul_U15243(.A(n17068), .Y(n4768));
AND2X1 mul_U15244(.A(n9042), .B(n9999), .Y(n17075));
INVX1 mul_U15245(.A(n17075), .Y(n4769));
AND2X1 mul_U15246(.A(n9043), .B(n9997), .Y(n17082));
INVX1 mul_U15247(.A(n17082), .Y(n4770));
AND2X1 mul_U15248(.A(n9044), .B(n9994), .Y(n17089));
INVX1 mul_U15249(.A(n17089), .Y(n4771));
AND2X1 mul_U15250(.A(n9045), .B(n9991), .Y(n17096));
INVX1 mul_U15251(.A(n17096), .Y(n4772));
AND2X1 mul_U15252(.A(n9046), .B(n9988), .Y(n17103));
INVX1 mul_U15253(.A(n17103), .Y(n4773));
AND2X1 mul_U15254(.A(n9047), .B(n9985), .Y(n17110));
INVX1 mul_U15255(.A(n17110), .Y(n4774));
AND2X1 mul_U15256(.A(n9048), .B(n9982), .Y(n17117));
INVX1 mul_U15257(.A(n17117), .Y(n4775));
AND2X1 mul_U15258(.A(n9049), .B(n9979), .Y(n17124));
INVX1 mul_U15259(.A(n17124), .Y(n4776));
AND2X1 mul_U15260(.A(n9050), .B(n9976), .Y(n17131));
INVX1 mul_U15261(.A(n17131), .Y(n4777));
AND2X1 mul_U15262(.A(n9051), .B(n9973), .Y(n17138));
INVX1 mul_U15263(.A(n17138), .Y(n4778));
AND2X1 mul_U15264(.A(n9052), .B(n9970), .Y(n17145));
INVX1 mul_U15265(.A(n17145), .Y(n4779));
AND2X1 mul_U15266(.A(n9053), .B(n9967), .Y(n17152));
INVX1 mul_U15267(.A(n17152), .Y(n4780));
AND2X1 mul_U15268(.A(n9054), .B(n9964), .Y(n17159));
INVX1 mul_U15269(.A(n17159), .Y(n4781));
AND2X1 mul_U15270(.A(n9055), .B(n9961), .Y(n17166));
INVX1 mul_U15271(.A(n17166), .Y(n4782));
AND2X1 mul_U15272(.A(n9056), .B(n9958), .Y(n17173));
INVX1 mul_U15273(.A(n17173), .Y(n4783));
AND2X1 mul_U15274(.A(n9057), .B(n9955), .Y(n17180));
INVX1 mul_U15275(.A(n17180), .Y(n4784));
AND2X1 mul_U15276(.A(n9058), .B(n9952), .Y(n17187));
INVX1 mul_U15277(.A(n17187), .Y(n4785));
AND2X1 mul_U15278(.A(n9059), .B(n9949), .Y(n17194));
INVX1 mul_U15279(.A(n17194), .Y(n4786));
AND2X1 mul_U15280(.A(n9060), .B(n9946), .Y(n17201));
INVX1 mul_U15281(.A(n17201), .Y(n4787));
AND2X1 mul_U15282(.A(n9061), .B(n9943), .Y(n17208));
INVX1 mul_U15283(.A(n17208), .Y(n4788));
AND2X1 mul_U15284(.A(n9062), .B(n9940), .Y(n17215));
INVX1 mul_U15285(.A(n17215), .Y(n4789));
AND2X1 mul_U15286(.A(n9063), .B(n9937), .Y(n17222));
INVX1 mul_U15287(.A(n17222), .Y(n4790));
AND2X1 mul_U15288(.A(n9064), .B(n9934), .Y(n17229));
INVX1 mul_U15289(.A(n17229), .Y(n4791));
AND2X1 mul_U15290(.A(n9065), .B(n9931), .Y(n17236));
INVX1 mul_U15291(.A(n17236), .Y(n4792));
AND2X1 mul_U15292(.A(n9066), .B(n9928), .Y(n17243));
INVX1 mul_U15293(.A(n17243), .Y(n4793));
AND2X1 mul_U15294(.A(n9067), .B(n9925), .Y(n17250));
INVX1 mul_U15295(.A(n17250), .Y(n4794));
AND2X1 mul_U15296(.A(n9068), .B(n9922), .Y(n17257));
INVX1 mul_U15297(.A(n17257), .Y(n4795));
AND2X1 mul_U15298(.A(n9069), .B(n9919), .Y(n17264));
INVX1 mul_U15299(.A(n17264), .Y(n4796));
AND2X1 mul_U15300(.A(n9070), .B(n9916), .Y(n17271));
INVX1 mul_U15301(.A(n17271), .Y(n4797));
AND2X1 mul_U15302(.A(n9071), .B(n9913), .Y(n17278));
INVX1 mul_U15303(.A(n17278), .Y(n4798));
AND2X1 mul_U15304(.A(n9072), .B(n9910), .Y(n17285));
INVX1 mul_U15305(.A(n17285), .Y(n4799));
AND2X1 mul_U15306(.A(n9073), .B(n9907), .Y(n17292));
INVX1 mul_U15307(.A(n17292), .Y(n4800));
AND2X1 mul_U15308(.A(n9074), .B(n9904), .Y(n17299));
INVX1 mul_U15309(.A(n17299), .Y(n4801));
AND2X1 mul_U15310(.A(n9075), .B(n9901), .Y(n17306));
INVX1 mul_U15311(.A(n17306), .Y(n4802));
AND2X1 mul_U15312(.A(n9076), .B(n9898), .Y(n17313));
INVX1 mul_U15313(.A(n17313), .Y(n4803));
AND2X1 mul_U15314(.A(n9077), .B(n9895), .Y(n17320));
INVX1 mul_U15315(.A(n17320), .Y(n4804));
AND2X1 mul_U15316(.A(n9078), .B(n9892), .Y(n17327));
INVX1 mul_U15317(.A(n17327), .Y(n4805));
AND2X1 mul_U15318(.A(n9079), .B(n9889), .Y(n17334));
INVX1 mul_U15319(.A(n17334), .Y(n4806));
AND2X1 mul_U15320(.A(n9080), .B(n9886), .Y(n17341));
INVX1 mul_U15321(.A(n17341), .Y(n4807));
AND2X1 mul_U15322(.A(n9081), .B(n9883), .Y(n17348));
INVX1 mul_U15323(.A(n17348), .Y(n4808));
AND2X1 mul_U15324(.A(n9082), .B(n9880), .Y(n17355));
INVX1 mul_U15325(.A(n17355), .Y(n4809));
AND2X1 mul_U15326(.A(n9083), .B(n9877), .Y(n17362));
INVX1 mul_U15327(.A(n17362), .Y(n4810));
AND2X1 mul_U15328(.A(n9084), .B(n9874), .Y(n17369));
INVX1 mul_U15329(.A(n17369), .Y(n4811));
AND2X1 mul_U15330(.A(n9085), .B(n9871), .Y(n17376));
INVX1 mul_U15331(.A(n17376), .Y(n4812));
AND2X1 mul_U15332(.A(n9086), .B(n9868), .Y(n17383));
INVX1 mul_U15333(.A(n17383), .Y(n4813));
AND2X1 mul_U15334(.A(n9087), .B(n9865), .Y(n17390));
INVX1 mul_U15335(.A(n17390), .Y(n4814));
AND2X1 mul_U15336(.A(n9088), .B(n9862), .Y(n17397));
INVX1 mul_U15337(.A(n17397), .Y(n4815));
AND2X1 mul_U15338(.A(n9089), .B(n9859), .Y(n17404));
INVX1 mul_U15339(.A(n17404), .Y(n4816));
AND2X1 mul_U15340(.A(n9090), .B(n9856), .Y(n17411));
INVX1 mul_U15341(.A(n17411), .Y(n4817));
AND2X1 mul_U15342(.A(n9091), .B(n9826), .Y(n17418));
INVX1 mul_U15343(.A(n17418), .Y(n4818));
AND2X1 mul_U15344(.A(n9092), .B(n9824), .Y(n17425));
INVX1 mul_U15345(.A(n17425), .Y(n4819));
AND2X1 mul_U15346(.A(n9093), .B(n9825), .Y(n17432));
INVX1 mul_U15347(.A(n17432), .Y(n4820));
AND2X1 mul_U15348(.A(n9094), .B(n9836), .Y(n17439));
INVX1 mul_U15349(.A(n17439), .Y(n4821));
AND2X1 mul_U15350(.A(n9095), .B(n9837), .Y(n17446));
INVX1 mul_U15351(.A(n17446), .Y(n4822));
AND2X1 mul_U15352(.A(n9096), .B(n9833), .Y(n17453));
INVX1 mul_U15353(.A(n17453), .Y(n4823));
AND2X1 mul_U15354(.A(n9097), .B(n9834), .Y(n17460));
INVX1 mul_U15355(.A(n17460), .Y(n4824));
AND2X1 mul_U15356(.A(dpath_mulcore_booth_b1_in0[2]), .B(n9784), .Y(n17859));
INVX1 mul_U15357(.A(n17859), .Y(n4825));
AND2X1 mul_U15358(.A(n5481), .B(n9784), .Y(n17861));
INVX1 mul_U15359(.A(n17861), .Y(n4826));
AND2X1 mul_U15360(.A(n5495), .B(n9784), .Y(n17863));
INVX1 mul_U15361(.A(n17863), .Y(n4827));
AND2X1 mul_U15362(.A(dpath_mulcore_booth_b2_in0[2]), .B(n9784), .Y(n17865));
INVX1 mul_U15363(.A(n17865), .Y(n4828));
AND2X1 mul_U15364(.A(n5480), .B(n9784), .Y(n17867));
INVX1 mul_U15365(.A(n17867), .Y(n4829));
AND2X1 mul_U15366(.A(n5493), .B(n9784), .Y(n17869));
INVX1 mul_U15367(.A(n17869), .Y(n4830));
AND2X1 mul_U15368(.A(dpath_mulcore_booth_b3_in0[2]), .B(n9784), .Y(n17871));
INVX1 mul_U15369(.A(n17871), .Y(n4831));
AND2X1 mul_U15370(.A(n5479), .B(n9784), .Y(n17873));
INVX1 mul_U15371(.A(n17873), .Y(n4832));
AND2X1 mul_U15372(.A(n5491), .B(n9784), .Y(n17875));
INVX1 mul_U15373(.A(n17875), .Y(n4833));
AND2X1 mul_U15374(.A(dpath_mulcore_booth_b4_in0[2]), .B(n9784), .Y(n17877));
INVX1 mul_U15375(.A(n17877), .Y(n4834));
AND2X1 mul_U15376(.A(n5478), .B(n9784), .Y(n17879));
INVX1 mul_U15377(.A(n17879), .Y(n4835));
AND2X1 mul_U15378(.A(n5489), .B(n9784), .Y(n17881));
INVX1 mul_U15379(.A(n17881), .Y(n4836));
AND2X1 mul_U15380(.A(dpath_mulcore_booth_b5_in0[2]), .B(n9784), .Y(n17883));
INVX1 mul_U15381(.A(n17883), .Y(n4837));
AND2X1 mul_U15382(.A(n5477), .B(n9784), .Y(n17885));
INVX1 mul_U15383(.A(n17885), .Y(n4838));
AND2X1 mul_U15384(.A(n5487), .B(n9784), .Y(n17887));
INVX1 mul_U15385(.A(n17887), .Y(n4839));
AND2X1 mul_U15386(.A(dpath_mulcore_booth_b6_in0[2]), .B(n9784), .Y(n17889));
INVX1 mul_U15387(.A(n17889), .Y(n4840));
AND2X1 mul_U15388(.A(n5476), .B(n9784), .Y(n17891));
INVX1 mul_U15389(.A(n17891), .Y(n4841));
AND2X1 mul_U15390(.A(n5485), .B(n9784), .Y(n17893));
INVX1 mul_U15391(.A(n17893), .Y(n4842));
AND2X1 mul_U15392(.A(dpath_mulcore_booth_b7_in0[2]), .B(n9784), .Y(n17895));
INVX1 mul_U15393(.A(n17895), .Y(n4843));
AND2X1 mul_U15394(.A(n5475), .B(n9784), .Y(n17897));
INVX1 mul_U15395(.A(n17897), .Y(n4844));
AND2X1 mul_U15396(.A(n5482), .B(n9784), .Y(n17899));
INVX1 mul_U15397(.A(n17899), .Y(n4845));
AND2X1 mul_U15398(.A(dpath_mulcore_booth_b8_in0[2]), .B(n9784), .Y(n17901));
INVX1 mul_U15399(.A(n17901), .Y(n4846));
AND2X1 mul_U15400(.A(n5391), .B(n9784), .Y(n17903));
INVX1 mul_U15401(.A(n17903), .Y(n4847));
AND2X1 mul_U15402(.A(n5415), .B(n9784), .Y(n17905));
INVX1 mul_U15403(.A(n17905), .Y(n4848));
AND2X1 mul_U15404(.A(dpath_mulcore_booth_b9_in0[2]), .B(n9784), .Y(n17907));
INVX1 mul_U15405(.A(n17907), .Y(n4849));
AND2X1 mul_U15406(.A(n5398), .B(n9784), .Y(n17909));
INVX1 mul_U15407(.A(n17909), .Y(n4850));
AND2X1 mul_U15408(.A(n5412), .B(n9784), .Y(n17911));
INVX1 mul_U15409(.A(n17911), .Y(n4851));
AND2X1 mul_U15410(.A(dpath_mulcore_booth_b10_in0[2]), .B(n9784), .Y(n17913));
INVX1 mul_U15411(.A(n17913), .Y(n4852));
AND2X1 mul_U15412(.A(n5397), .B(n9784), .Y(n17915));
INVX1 mul_U15413(.A(n17915), .Y(n4853));
AND2X1 mul_U15414(.A(n5410), .B(n9784), .Y(n17917));
INVX1 mul_U15415(.A(n17917), .Y(n4854));
AND2X1 mul_U15416(.A(dpath_mulcore_booth_b11_in0[2]), .B(n9784), .Y(n17919));
INVX1 mul_U15417(.A(n17919), .Y(n4855));
AND2X1 mul_U15418(.A(n5396), .B(n9784), .Y(n17921));
INVX1 mul_U15419(.A(n17921), .Y(n4856));
AND2X1 mul_U15420(.A(n5408), .B(n9784), .Y(n17923));
INVX1 mul_U15421(.A(n17923), .Y(n4857));
AND2X1 mul_U15422(.A(dpath_mulcore_booth_b12_in0[2]), .B(n9784), .Y(n17925));
INVX1 mul_U15423(.A(n17925), .Y(n4858));
AND2X1 mul_U15424(.A(n5395), .B(n9784), .Y(n17927));
INVX1 mul_U15425(.A(n17927), .Y(n4859));
AND2X1 mul_U15426(.A(n5406), .B(n9784), .Y(n17929));
INVX1 mul_U15427(.A(n17929), .Y(n4860));
AND2X1 mul_U15428(.A(dpath_mulcore_booth_b13_in0[2]), .B(n9784), .Y(n17931));
INVX1 mul_U15429(.A(n17931), .Y(n4861));
AND2X1 mul_U15430(.A(n5394), .B(n9784), .Y(n17933));
INVX1 mul_U15431(.A(n17933), .Y(n4862));
AND2X1 mul_U15432(.A(n5404), .B(n9784), .Y(n17935));
INVX1 mul_U15433(.A(n17935), .Y(n4863));
AND2X1 mul_U15434(.A(dpath_mulcore_booth_b14_in0[2]), .B(n9784), .Y(n17937));
INVX1 mul_U15435(.A(n17937), .Y(n4864));
AND2X1 mul_U15436(.A(n5393), .B(n9784), .Y(n17939));
INVX1 mul_U15437(.A(n17939), .Y(n4865));
AND2X1 mul_U15438(.A(n5402), .B(n9784), .Y(n17941));
INVX1 mul_U15439(.A(n17941), .Y(n4866));
AND2X1 mul_U15440(.A(dpath_mulcore_booth_b15_in0[2]), .B(n9784), .Y(n17942));
INVX1 mul_U15441(.A(n17942), .Y(n4867));
AND2X1 mul_U15442(.A(n5392), .B(n9784), .Y(n17944));
INVX1 mul_U15443(.A(n17944), .Y(n4868));
AND2X1 mul_U15444(.A(n5399), .B(n9784), .Y(n17946));
INVX1 mul_U15445(.A(n17946), .Y(n4869));
AND2X1 mul_U15446(.A(dpath_mulcore_booth_b[32]), .B(n10082), .Y(n18012));
INVX1 mul_U15447(.A(n18012), .Y(n4870));
AND2X1 mul_U15448(.A(n18073), .B(dpath_mulcore_booth_b[32]), .Y(n18072));
INVX1 mul_U15449(.A(n18072), .Y(n4871));
AND2X1 mul_U15450(.A(n9147), .B(n10011), .Y(dpath_mulcore_ary1_a0_sc3_71__n6));
INVX1 mul_U15451(.A(dpath_mulcore_ary1_a0_sc3_71__n6), .Y(n4872));
AND2X1 mul_U15452(.A(dpath_mulcore_booth_b0_in0[2]), .B(n9784), .Y(dpath_mulcore_booth_out_mux0_n3));
INVX1 mul_U15453(.A(dpath_mulcore_booth_out_mux0_n3), .Y(n4873));
AND2X1 mul_U15454(.A(n5474), .B(n9784), .Y(dpath_mulcore_booth_out_mux0_n5));
INVX1 mul_U15455(.A(dpath_mulcore_booth_out_mux0_n5), .Y(n4874));
AND2X1 mul_U15456(.A(dpath_mulcore_booth_encode0_a_n75), .B(n9784), .Y(dpath_mulcore_booth_out_mux0_n7));
INVX1 mul_U15457(.A(dpath_mulcore_booth_out_mux0_n7), .Y(n4875));
AND2X1 mul_U15458(.A(dpath_mulcore_psum[9]), .B(n9680), .Y(dpath_mulcore_ary2_smux_n3));
INVX1 mul_U15459(.A(dpath_mulcore_ary2_smux_n3), .Y(n4876));
AND2X1 mul_U15460(.A(dpath_mulcore_psum[97]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n5));
INVX1 mul_U15461(.A(dpath_mulcore_ary2_smux_n5), .Y(n4877));
AND2X1 mul_U15462(.A(dpath_mulcore_psum[96]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n7));
INVX1 mul_U15463(.A(dpath_mulcore_ary2_smux_n7), .Y(n4878));
AND2X1 mul_U15464(.A(dpath_mulcore_psum[95]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n9));
INVX1 mul_U15465(.A(dpath_mulcore_ary2_smux_n9), .Y(n4879));
AND2X1 mul_U15466(.A(dpath_mulcore_psum[94]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n11));
INVX1 mul_U15467(.A(dpath_mulcore_ary2_smux_n11), .Y(n4880));
AND2X1 mul_U15468(.A(dpath_mulcore_psum[93]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n13));
INVX1 mul_U15469(.A(dpath_mulcore_ary2_smux_n13), .Y(n4881));
AND2X1 mul_U15470(.A(dpath_mulcore_psum[92]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n15));
INVX1 mul_U15471(.A(dpath_mulcore_ary2_smux_n15), .Y(n4882));
AND2X1 mul_U15472(.A(dpath_mulcore_psum[91]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n17));
INVX1 mul_U15473(.A(dpath_mulcore_ary2_smux_n17), .Y(n4883));
AND2X1 mul_U15474(.A(dpath_mulcore_psum[90]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n19));
INVX1 mul_U15475(.A(dpath_mulcore_ary2_smux_n19), .Y(n4884));
AND2X1 mul_U15476(.A(dpath_mulcore_psum[8]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n21));
INVX1 mul_U15477(.A(dpath_mulcore_ary2_smux_n21), .Y(n4885));
AND2X1 mul_U15478(.A(dpath_mulcore_psum[89]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n23));
INVX1 mul_U15479(.A(dpath_mulcore_ary2_smux_n23), .Y(n4886));
AND2X1 mul_U15480(.A(dpath_mulcore_psum[88]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n25));
INVX1 mul_U15481(.A(dpath_mulcore_ary2_smux_n25), .Y(n4887));
AND2X1 mul_U15482(.A(dpath_mulcore_psum[87]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n27));
INVX1 mul_U15483(.A(dpath_mulcore_ary2_smux_n27), .Y(n4888));
AND2X1 mul_U15484(.A(dpath_mulcore_psum[86]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n29));
INVX1 mul_U15485(.A(dpath_mulcore_ary2_smux_n29), .Y(n4889));
AND2X1 mul_U15486(.A(dpath_mulcore_psum[85]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n31));
INVX1 mul_U15487(.A(dpath_mulcore_ary2_smux_n31), .Y(n4890));
AND2X1 mul_U15488(.A(dpath_mulcore_psum[84]), .B(n9707), .Y(dpath_mulcore_ary2_smux_n33));
INVX1 mul_U15489(.A(dpath_mulcore_ary2_smux_n33), .Y(n4891));
AND2X1 mul_U15490(.A(dpath_mulcore_psum[83]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n35));
INVX1 mul_U15491(.A(dpath_mulcore_ary2_smux_n35), .Y(n4892));
AND2X1 mul_U15492(.A(dpath_mulcore_psum[82]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n37));
INVX1 mul_U15493(.A(dpath_mulcore_ary2_smux_n37), .Y(n4893));
AND2X1 mul_U15494(.A(dpath_mulcore_psum[81]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n39));
INVX1 mul_U15495(.A(dpath_mulcore_ary2_smux_n39), .Y(n4894));
AND2X1 mul_U15496(.A(dpath_mulcore_psum[80]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n41));
INVX1 mul_U15497(.A(dpath_mulcore_ary2_smux_n41), .Y(n4895));
AND2X1 mul_U15498(.A(dpath_mulcore_psum[7]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n43));
INVX1 mul_U15499(.A(dpath_mulcore_ary2_smux_n43), .Y(n4896));
AND2X1 mul_U15500(.A(dpath_mulcore_psum[79]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n45));
INVX1 mul_U15501(.A(dpath_mulcore_ary2_smux_n45), .Y(n4897));
AND2X1 mul_U15502(.A(dpath_mulcore_psum[78]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n47));
INVX1 mul_U15503(.A(dpath_mulcore_ary2_smux_n47), .Y(n4898));
AND2X1 mul_U15504(.A(dpath_mulcore_psum[77]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n49));
INVX1 mul_U15505(.A(dpath_mulcore_ary2_smux_n49), .Y(n4899));
AND2X1 mul_U15506(.A(dpath_mulcore_psum[76]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n51));
INVX1 mul_U15507(.A(dpath_mulcore_ary2_smux_n51), .Y(n4900));
AND2X1 mul_U15508(.A(dpath_mulcore_psum[75]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n53));
INVX1 mul_U15509(.A(dpath_mulcore_ary2_smux_n53), .Y(n4901));
AND2X1 mul_U15510(.A(dpath_mulcore_psum[74]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n55));
INVX1 mul_U15511(.A(dpath_mulcore_ary2_smux_n55), .Y(n4902));
AND2X1 mul_U15512(.A(dpath_mulcore_psum[73]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n57));
INVX1 mul_U15513(.A(dpath_mulcore_ary2_smux_n57), .Y(n4903));
AND2X1 mul_U15514(.A(dpath_mulcore_psum[72]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n59));
INVX1 mul_U15515(.A(dpath_mulcore_ary2_smux_n59), .Y(n4904));
AND2X1 mul_U15516(.A(dpath_mulcore_psum[71]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n61));
INVX1 mul_U15517(.A(dpath_mulcore_ary2_smux_n61), .Y(n4905));
AND2X1 mul_U15518(.A(dpath_mulcore_psum[70]), .B(n9708), .Y(dpath_mulcore_ary2_smux_n63));
INVX1 mul_U15519(.A(dpath_mulcore_ary2_smux_n63), .Y(n4906));
AND2X1 mul_U15520(.A(dpath_mulcore_psum[6]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n65));
INVX1 mul_U15521(.A(dpath_mulcore_ary2_smux_n65), .Y(n4907));
AND2X1 mul_U15522(.A(dpath_mulcore_psum[69]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n67));
INVX1 mul_U15523(.A(dpath_mulcore_ary2_smux_n67), .Y(n4908));
AND2X1 mul_U15524(.A(dpath_mulcore_psum[68]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n69));
INVX1 mul_U15525(.A(dpath_mulcore_ary2_smux_n69), .Y(n4909));
AND2X1 mul_U15526(.A(dpath_mulcore_psum[67]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n71));
INVX1 mul_U15527(.A(dpath_mulcore_ary2_smux_n71), .Y(n4910));
AND2X1 mul_U15528(.A(dpath_mulcore_psum[66]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n73));
INVX1 mul_U15529(.A(dpath_mulcore_ary2_smux_n73), .Y(n4911));
AND2X1 mul_U15530(.A(dpath_mulcore_psum[65]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n75));
INVX1 mul_U15531(.A(dpath_mulcore_ary2_smux_n75), .Y(n4912));
AND2X1 mul_U15532(.A(dpath_mulcore_psum[64]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n77));
INVX1 mul_U15533(.A(dpath_mulcore_ary2_smux_n77), .Y(n4913));
AND2X1 mul_U15534(.A(dpath_mulcore_psum[63]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n79));
INVX1 mul_U15535(.A(dpath_mulcore_ary2_smux_n79), .Y(n4914));
AND2X1 mul_U15536(.A(dpath_mulcore_psum[62]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n81));
INVX1 mul_U15537(.A(dpath_mulcore_ary2_smux_n81), .Y(n4915));
AND2X1 mul_U15538(.A(dpath_mulcore_psum[61]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n83));
INVX1 mul_U15539(.A(dpath_mulcore_ary2_smux_n83), .Y(n4916));
AND2X1 mul_U15540(.A(dpath_mulcore_psum[60]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n85));
INVX1 mul_U15541(.A(dpath_mulcore_ary2_smux_n85), .Y(n4917));
AND2X1 mul_U15542(.A(dpath_mulcore_psum[5]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n87));
INVX1 mul_U15543(.A(dpath_mulcore_ary2_smux_n87), .Y(n4918));
AND2X1 mul_U15544(.A(dpath_mulcore_psum[59]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n89));
INVX1 mul_U15545(.A(dpath_mulcore_ary2_smux_n89), .Y(n4919));
AND2X1 mul_U15546(.A(dpath_mulcore_psum[58]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n91));
INVX1 mul_U15547(.A(dpath_mulcore_ary2_smux_n91), .Y(n4920));
AND2X1 mul_U15548(.A(dpath_mulcore_psum[57]), .B(n9709), .Y(dpath_mulcore_ary2_smux_n93));
INVX1 mul_U15549(.A(dpath_mulcore_ary2_smux_n93), .Y(n4921));
AND2X1 mul_U15550(.A(dpath_mulcore_psum[56]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n95));
INVX1 mul_U15551(.A(dpath_mulcore_ary2_smux_n95), .Y(n4922));
AND2X1 mul_U15552(.A(dpath_mulcore_psum[55]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n97));
INVX1 mul_U15553(.A(dpath_mulcore_ary2_smux_n97), .Y(n4923));
AND2X1 mul_U15554(.A(dpath_mulcore_psum[54]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n99));
INVX1 mul_U15555(.A(dpath_mulcore_ary2_smux_n99), .Y(n4924));
AND2X1 mul_U15556(.A(dpath_mulcore_psum[53]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n101));
INVX1 mul_U15557(.A(dpath_mulcore_ary2_smux_n101), .Y(n4925));
AND2X1 mul_U15558(.A(dpath_mulcore_psum[52]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n103));
INVX1 mul_U15559(.A(dpath_mulcore_ary2_smux_n103), .Y(n4926));
AND2X1 mul_U15560(.A(dpath_mulcore_psum[51]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n105));
INVX1 mul_U15561(.A(dpath_mulcore_ary2_smux_n105), .Y(n4927));
AND2X1 mul_U15562(.A(dpath_mulcore_psum[50]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n107));
INVX1 mul_U15563(.A(dpath_mulcore_ary2_smux_n107), .Y(n4928));
AND2X1 mul_U15564(.A(dpath_mulcore_psum[4]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n109));
INVX1 mul_U15565(.A(dpath_mulcore_ary2_smux_n109), .Y(n4929));
AND2X1 mul_U15566(.A(dpath_mulcore_psum[49]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n111));
INVX1 mul_U15567(.A(dpath_mulcore_ary2_smux_n111), .Y(n4930));
AND2X1 mul_U15568(.A(dpath_mulcore_psum[48]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n113));
INVX1 mul_U15569(.A(dpath_mulcore_ary2_smux_n113), .Y(n4931));
AND2X1 mul_U15570(.A(dpath_mulcore_psum[47]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n115));
INVX1 mul_U15571(.A(dpath_mulcore_ary2_smux_n115), .Y(n4932));
AND2X1 mul_U15572(.A(dpath_mulcore_psum[46]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n117));
INVX1 mul_U15573(.A(dpath_mulcore_ary2_smux_n117), .Y(n4933));
AND2X1 mul_U15574(.A(dpath_mulcore_psum[45]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n119));
INVX1 mul_U15575(.A(dpath_mulcore_ary2_smux_n119), .Y(n4934));
AND2X1 mul_U15576(.A(dpath_mulcore_psum[44]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n121));
INVX1 mul_U15577(.A(dpath_mulcore_ary2_smux_n121), .Y(n4935));
AND2X1 mul_U15578(.A(dpath_mulcore_psum[43]), .B(n9710), .Y(dpath_mulcore_ary2_smux_n123));
INVX1 mul_U15579(.A(dpath_mulcore_ary2_smux_n123), .Y(n4936));
AND2X1 mul_U15580(.A(dpath_mulcore_psum[42]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n125));
INVX1 mul_U15581(.A(dpath_mulcore_ary2_smux_n125), .Y(n4937));
AND2X1 mul_U15582(.A(dpath_mulcore_psum[41]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n127));
INVX1 mul_U15583(.A(dpath_mulcore_ary2_smux_n127), .Y(n4938));
AND2X1 mul_U15584(.A(dpath_mulcore_psum[40]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n129));
INVX1 mul_U15585(.A(dpath_mulcore_ary2_smux_n129), .Y(n4939));
AND2X1 mul_U15586(.A(dpath_mulcore_psum[3]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n131));
INVX1 mul_U15587(.A(dpath_mulcore_ary2_smux_n131), .Y(n4940));
AND2X1 mul_U15588(.A(dpath_mulcore_psum[39]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n133));
INVX1 mul_U15589(.A(dpath_mulcore_ary2_smux_n133), .Y(n4941));
AND2X1 mul_U15590(.A(dpath_mulcore_psum[38]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n135));
INVX1 mul_U15591(.A(dpath_mulcore_ary2_smux_n135), .Y(n4942));
AND2X1 mul_U15592(.A(dpath_mulcore_psum[37]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n137));
INVX1 mul_U15593(.A(dpath_mulcore_ary2_smux_n137), .Y(n4943));
AND2X1 mul_U15594(.A(dpath_mulcore_psum[36]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n139));
INVX1 mul_U15595(.A(dpath_mulcore_ary2_smux_n139), .Y(n4944));
AND2X1 mul_U15596(.A(dpath_mulcore_psum[35]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n141));
INVX1 mul_U15597(.A(dpath_mulcore_ary2_smux_n141), .Y(n4945));
AND2X1 mul_U15598(.A(dpath_mulcore_psum[34]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n143));
INVX1 mul_U15599(.A(dpath_mulcore_ary2_smux_n143), .Y(n4946));
AND2X1 mul_U15600(.A(dpath_mulcore_psum[33]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n145));
INVX1 mul_U15601(.A(dpath_mulcore_ary2_smux_n145), .Y(n4947));
AND2X1 mul_U15602(.A(dpath_mulcore_psum[32]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n147));
INVX1 mul_U15603(.A(dpath_mulcore_ary2_smux_n147), .Y(n4948));
AND2X1 mul_U15604(.A(dpath_mulcore_psum[31]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n149));
INVX1 mul_U15605(.A(dpath_mulcore_ary2_smux_n149), .Y(n4949));
AND2X1 mul_U15606(.A(dpath_mulcore_psum[30]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n151));
INVX1 mul_U15607(.A(dpath_mulcore_ary2_smux_n151), .Y(n4950));
AND2X1 mul_U15608(.A(dpath_mulcore_psum[2]), .B(n9711), .Y(dpath_mulcore_ary2_smux_n153));
INVX1 mul_U15609(.A(dpath_mulcore_ary2_smux_n153), .Y(n4951));
AND2X1 mul_U15610(.A(dpath_mulcore_psum[29]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n155));
INVX1 mul_U15611(.A(dpath_mulcore_ary2_smux_n155), .Y(n4952));
AND2X1 mul_U15612(.A(dpath_mulcore_psum[28]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n157));
INVX1 mul_U15613(.A(dpath_mulcore_ary2_smux_n157), .Y(n4953));
AND2X1 mul_U15614(.A(dpath_mulcore_psum[27]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n159));
INVX1 mul_U15615(.A(dpath_mulcore_ary2_smux_n159), .Y(n4954));
AND2X1 mul_U15616(.A(dpath_mulcore_psum[26]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n161));
INVX1 mul_U15617(.A(dpath_mulcore_ary2_smux_n161), .Y(n4955));
AND2X1 mul_U15618(.A(dpath_mulcore_psum[25]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n163));
INVX1 mul_U15619(.A(dpath_mulcore_ary2_smux_n163), .Y(n4956));
AND2X1 mul_U15620(.A(dpath_mulcore_psum[24]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n165));
INVX1 mul_U15621(.A(dpath_mulcore_ary2_smux_n165), .Y(n4957));
AND2X1 mul_U15622(.A(dpath_mulcore_psum[23]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n167));
INVX1 mul_U15623(.A(dpath_mulcore_ary2_smux_n167), .Y(n4958));
AND2X1 mul_U15624(.A(dpath_mulcore_psum[22]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n169));
INVX1 mul_U15625(.A(dpath_mulcore_ary2_smux_n169), .Y(n4959));
AND2X1 mul_U15626(.A(dpath_mulcore_psum[21]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n171));
INVX1 mul_U15627(.A(dpath_mulcore_ary2_smux_n171), .Y(n4960));
AND2X1 mul_U15628(.A(dpath_mulcore_psum[20]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n173));
INVX1 mul_U15629(.A(dpath_mulcore_ary2_smux_n173), .Y(n4961));
AND2X1 mul_U15630(.A(dpath_mulcore_psum[1]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n175));
INVX1 mul_U15631(.A(dpath_mulcore_ary2_smux_n175), .Y(n4962));
AND2X1 mul_U15632(.A(dpath_mulcore_psum[19]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n177));
INVX1 mul_U15633(.A(dpath_mulcore_ary2_smux_n177), .Y(n4963));
AND2X1 mul_U15634(.A(dpath_mulcore_psum[18]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n179));
INVX1 mul_U15635(.A(dpath_mulcore_ary2_smux_n179), .Y(n4964));
AND2X1 mul_U15636(.A(dpath_mulcore_psum[17]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n181));
INVX1 mul_U15637(.A(dpath_mulcore_ary2_smux_n181), .Y(n4965));
AND2X1 mul_U15638(.A(dpath_mulcore_psum[16]), .B(n9712), .Y(dpath_mulcore_ary2_smux_n183));
INVX1 mul_U15639(.A(dpath_mulcore_ary2_smux_n183), .Y(n4966));
AND2X1 mul_U15640(.A(n16562), .B(n9713), .Y(dpath_mulcore_ary2_smux_n185));
INVX1 mul_U15641(.A(dpath_mulcore_ary2_smux_n185), .Y(n4967));
AND2X1 mul_U15642(.A(dpath_mulcore_psum[14]), .B(n9713), .Y(dpath_mulcore_ary2_smux_n187));
INVX1 mul_U15643(.A(dpath_mulcore_ary2_smux_n187), .Y(n4968));
AND2X1 mul_U15644(.A(dpath_mulcore_psum[13]), .B(n9713), .Y(dpath_mulcore_ary2_smux_n189));
INVX1 mul_U15645(.A(dpath_mulcore_ary2_smux_n189), .Y(n4969));
AND2X1 mul_U15646(.A(dpath_mulcore_psum[12]), .B(n9713), .Y(dpath_mulcore_ary2_smux_n191));
INVX1 mul_U15647(.A(dpath_mulcore_ary2_smux_n191), .Y(n4970));
AND2X1 mul_U15648(.A(dpath_mulcore_psum[11]), .B(n9713), .Y(dpath_mulcore_ary2_smux_n193));
INVX1 mul_U15649(.A(dpath_mulcore_ary2_smux_n193), .Y(n4971));
AND2X1 mul_U15650(.A(dpath_mulcore_psum[10]), .B(n9713), .Y(dpath_mulcore_ary2_smux_n195));
INVX1 mul_U15651(.A(dpath_mulcore_ary2_smux_n195), .Y(n4972));
AND2X1 mul_U15652(.A(dpath_mulcore_psum[0]), .B(n9713), .Y(dpath_mulcore_ary2_smux_n197));
INVX1 mul_U15653(.A(dpath_mulcore_ary2_smux_n197), .Y(n4973));
AND2X1 mul_U15654(.A(n6160), .B(n9696), .Y(dpath_mulcore_ary2_cmux_n3));
INVX1 mul_U15655(.A(dpath_mulcore_ary2_cmux_n3), .Y(n4974));
AND2X1 mul_U15656(.A(n6072), .B(n9697), .Y(dpath_mulcore_ary2_cmux_n5));
INVX1 mul_U15657(.A(dpath_mulcore_ary2_cmux_n5), .Y(n4975));
AND2X1 mul_U15658(.A(n9188), .B(n9698), .Y(dpath_mulcore_ary2_cmux_n7));
INVX1 mul_U15659(.A(dpath_mulcore_ary2_cmux_n7), .Y(n4976));
AND2X1 mul_U15660(.A(n9189), .B(n9699), .Y(dpath_mulcore_ary2_cmux_n9));
INVX1 mul_U15661(.A(dpath_mulcore_ary2_cmux_n9), .Y(n4977));
AND2X1 mul_U15662(.A(n9190), .B(n9700), .Y(dpath_mulcore_ary2_cmux_n11));
INVX1 mul_U15663(.A(dpath_mulcore_ary2_cmux_n11), .Y(n4978));
AND2X1 mul_U15664(.A(n9191), .B(n9701), .Y(dpath_mulcore_ary2_cmux_n13));
INVX1 mul_U15665(.A(dpath_mulcore_ary2_cmux_n13), .Y(n4979));
AND2X1 mul_U15666(.A(n9192), .B(n9681), .Y(dpath_mulcore_ary2_cmux_n15));
INVX1 mul_U15667(.A(dpath_mulcore_ary2_cmux_n15), .Y(n4980));
AND2X1 mul_U15668(.A(n9193), .B(n9682), .Y(dpath_mulcore_ary2_cmux_n17));
INVX1 mul_U15669(.A(dpath_mulcore_ary2_cmux_n17), .Y(n4981));
AND2X1 mul_U15670(.A(n6074), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n19));
INVX1 mul_U15671(.A(dpath_mulcore_ary2_cmux_n19), .Y(n4982));
AND2X1 mul_U15672(.A(n9194), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n21));
INVX1 mul_U15673(.A(dpath_mulcore_ary2_cmux_n21), .Y(n4983));
AND2X1 mul_U15674(.A(n9195), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n23));
INVX1 mul_U15675(.A(dpath_mulcore_ary2_cmux_n23), .Y(n4984));
AND2X1 mul_U15676(.A(n9196), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n25));
INVX1 mul_U15677(.A(dpath_mulcore_ary2_cmux_n25), .Y(n4985));
AND2X1 mul_U15678(.A(n9197), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n27));
INVX1 mul_U15679(.A(dpath_mulcore_ary2_cmux_n27), .Y(n4986));
AND2X1 mul_U15680(.A(n9198), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n29));
INVX1 mul_U15681(.A(dpath_mulcore_ary2_cmux_n29), .Y(n4987));
AND2X1 mul_U15682(.A(n9199), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n31));
INVX1 mul_U15683(.A(dpath_mulcore_ary2_cmux_n31), .Y(n4988));
AND2X1 mul_U15684(.A(n9213), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n33));
INVX1 mul_U15685(.A(dpath_mulcore_ary2_cmux_n33), .Y(n4989));
AND2X1 mul_U15686(.A(n9148), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n35));
INVX1 mul_U15687(.A(dpath_mulcore_ary2_cmux_n35), .Y(n4990));
AND2X1 mul_U15688(.A(n9200), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n37));
INVX1 mul_U15689(.A(dpath_mulcore_ary2_cmux_n37), .Y(n4991));
AND2X1 mul_U15690(.A(n9201), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n39));
INVX1 mul_U15691(.A(dpath_mulcore_ary2_cmux_n39), .Y(n4992));
AND2X1 mul_U15692(.A(n6161), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n41));
INVX1 mul_U15693(.A(dpath_mulcore_ary2_cmux_n41), .Y(n4993));
AND2X1 mul_U15694(.A(n9202), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n43));
INVX1 mul_U15695(.A(dpath_mulcore_ary2_cmux_n43), .Y(n4994));
AND2X1 mul_U15696(.A(n9203), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n45));
INVX1 mul_U15697(.A(dpath_mulcore_ary2_cmux_n45), .Y(n4995));
AND2X1 mul_U15698(.A(n9204), .B(n9702), .Y(dpath_mulcore_ary2_cmux_n47));
INVX1 mul_U15699(.A(dpath_mulcore_ary2_cmux_n47), .Y(n4996));
AND2X1 mul_U15700(.A(n9205), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n49));
INVX1 mul_U15701(.A(dpath_mulcore_ary2_cmux_n49), .Y(n4997));
AND2X1 mul_U15702(.A(n9206), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n51));
INVX1 mul_U15703(.A(dpath_mulcore_ary2_cmux_n51), .Y(n4998));
AND2X1 mul_U15704(.A(n9207), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n53));
INVX1 mul_U15705(.A(dpath_mulcore_ary2_cmux_n53), .Y(n4999));
AND2X1 mul_U15706(.A(n9208), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n55));
INVX1 mul_U15707(.A(dpath_mulcore_ary2_cmux_n55), .Y(n5000));
AND2X1 mul_U15708(.A(n9209), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n57));
INVX1 mul_U15709(.A(dpath_mulcore_ary2_cmux_n57), .Y(n5001));
AND2X1 mul_U15710(.A(n9210), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n59));
INVX1 mul_U15711(.A(dpath_mulcore_ary2_cmux_n59), .Y(n5002));
AND2X1 mul_U15712(.A(n9211), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n61));
INVX1 mul_U15713(.A(dpath_mulcore_ary2_cmux_n61), .Y(n5003));
AND2X1 mul_U15714(.A(n6162), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n63));
INVX1 mul_U15715(.A(dpath_mulcore_ary2_cmux_n63), .Y(n5004));
AND2X1 mul_U15716(.A(n9212), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n65));
INVX1 mul_U15717(.A(dpath_mulcore_ary2_cmux_n65), .Y(n5005));
AND2X1 mul_U15718(.A(n9149), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n67));
INVX1 mul_U15719(.A(dpath_mulcore_ary2_cmux_n67), .Y(n5006));
AND2X1 mul_U15720(.A(n9150), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n69));
INVX1 mul_U15721(.A(dpath_mulcore_ary2_cmux_n69), .Y(n5007));
AND2X1 mul_U15722(.A(n9151), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n71));
INVX1 mul_U15723(.A(dpath_mulcore_ary2_cmux_n71), .Y(n5008));
AND2X1 mul_U15724(.A(n9152), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n73));
INVX1 mul_U15725(.A(dpath_mulcore_ary2_cmux_n73), .Y(n5009));
AND2X1 mul_U15726(.A(n9153), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n75));
INVX1 mul_U15727(.A(dpath_mulcore_ary2_cmux_n75), .Y(n5010));
AND2X1 mul_U15728(.A(n9154), .B(n9703), .Y(dpath_mulcore_ary2_cmux_n77));
INVX1 mul_U15729(.A(dpath_mulcore_ary2_cmux_n77), .Y(n5011));
AND2X1 mul_U15730(.A(n9155), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n79));
INVX1 mul_U15731(.A(dpath_mulcore_ary2_cmux_n79), .Y(n5012));
AND2X1 mul_U15732(.A(n9156), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n81));
INVX1 mul_U15733(.A(dpath_mulcore_ary2_cmux_n81), .Y(n5013));
AND2X1 mul_U15734(.A(n9157), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n83));
INVX1 mul_U15735(.A(dpath_mulcore_ary2_cmux_n83), .Y(n5014));
AND2X1 mul_U15736(.A(n6163), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n85));
INVX1 mul_U15737(.A(dpath_mulcore_ary2_cmux_n85), .Y(n5015));
AND2X1 mul_U15738(.A(n9158), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n87));
INVX1 mul_U15739(.A(dpath_mulcore_ary2_cmux_n87), .Y(n5016));
AND2X1 mul_U15740(.A(n9159), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n89));
INVX1 mul_U15741(.A(dpath_mulcore_ary2_cmux_n89), .Y(n5017));
AND2X1 mul_U15742(.A(n9160), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n91));
INVX1 mul_U15743(.A(dpath_mulcore_ary2_cmux_n91), .Y(n5018));
AND2X1 mul_U15744(.A(n9161), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n93));
INVX1 mul_U15745(.A(dpath_mulcore_ary2_cmux_n93), .Y(n5019));
AND2X1 mul_U15746(.A(n9162), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n95));
INVX1 mul_U15747(.A(dpath_mulcore_ary2_cmux_n95), .Y(n5020));
AND2X1 mul_U15748(.A(n9163), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n97));
INVX1 mul_U15749(.A(dpath_mulcore_ary2_cmux_n97), .Y(n5021));
AND2X1 mul_U15750(.A(n9164), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n99));
INVX1 mul_U15751(.A(dpath_mulcore_ary2_cmux_n99), .Y(n5022));
AND2X1 mul_U15752(.A(n9165), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n101));
INVX1 mul_U15753(.A(dpath_mulcore_ary2_cmux_n101), .Y(n5023));
AND2X1 mul_U15754(.A(n9166), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n103));
INVX1 mul_U15755(.A(dpath_mulcore_ary2_cmux_n103), .Y(n5024));
AND2X1 mul_U15756(.A(n9167), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n105));
INVX1 mul_U15757(.A(dpath_mulcore_ary2_cmux_n105), .Y(n5025));
AND2X1 mul_U15758(.A(n6151), .B(n9704), .Y(dpath_mulcore_ary2_cmux_n107));
INVX1 mul_U15759(.A(dpath_mulcore_ary2_cmux_n107), .Y(n5026));
AND2X1 mul_U15760(.A(n9168), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n109));
INVX1 mul_U15761(.A(dpath_mulcore_ary2_cmux_n109), .Y(n5027));
AND2X1 mul_U15762(.A(n9169), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n111));
INVX1 mul_U15763(.A(dpath_mulcore_ary2_cmux_n111), .Y(n5028));
AND2X1 mul_U15764(.A(n9170), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n113));
INVX1 mul_U15765(.A(dpath_mulcore_ary2_cmux_n113), .Y(n5029));
AND2X1 mul_U15766(.A(n9171), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n115));
INVX1 mul_U15767(.A(dpath_mulcore_ary2_cmux_n115), .Y(n5030));
AND2X1 mul_U15768(.A(n9172), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n117));
INVX1 mul_U15769(.A(dpath_mulcore_ary2_cmux_n117), .Y(n5031));
AND2X1 mul_U15770(.A(n9173), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n119));
INVX1 mul_U15771(.A(dpath_mulcore_ary2_cmux_n119), .Y(n5032));
AND2X1 mul_U15772(.A(n9174), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n121));
INVX1 mul_U15773(.A(dpath_mulcore_ary2_cmux_n121), .Y(n5033));
AND2X1 mul_U15774(.A(n9175), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n123));
INVX1 mul_U15775(.A(dpath_mulcore_ary2_cmux_n123), .Y(n5034));
AND2X1 mul_U15776(.A(n9176), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n125));
INVX1 mul_U15777(.A(dpath_mulcore_ary2_cmux_n125), .Y(n5035));
AND2X1 mul_U15778(.A(n9177), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n127));
INVX1 mul_U15779(.A(dpath_mulcore_ary2_cmux_n127), .Y(n5036));
AND2X1 mul_U15780(.A(n6152), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n129));
INVX1 mul_U15781(.A(dpath_mulcore_ary2_cmux_n129), .Y(n5037));
AND2X1 mul_U15782(.A(n9178), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n131));
INVX1 mul_U15783(.A(dpath_mulcore_ary2_cmux_n131), .Y(n5038));
AND2X1 mul_U15784(.A(n9179), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n133));
INVX1 mul_U15785(.A(dpath_mulcore_ary2_cmux_n133), .Y(n5039));
AND2X1 mul_U15786(.A(n9180), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n135));
INVX1 mul_U15787(.A(dpath_mulcore_ary2_cmux_n135), .Y(n5040));
AND2X1 mul_U15788(.A(n9181), .B(n9705), .Y(dpath_mulcore_ary2_cmux_n137));
INVX1 mul_U15789(.A(dpath_mulcore_ary2_cmux_n137), .Y(n5041));
AND2X1 mul_U15790(.A(n9182), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n139));
INVX1 mul_U15791(.A(dpath_mulcore_ary2_cmux_n139), .Y(n5042));
AND2X1 mul_U15792(.A(n9183), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n141));
INVX1 mul_U15793(.A(dpath_mulcore_ary2_cmux_n141), .Y(n5043));
AND2X1 mul_U15794(.A(n9184), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n143));
INVX1 mul_U15795(.A(dpath_mulcore_ary2_cmux_n143), .Y(n5044));
AND2X1 mul_U15796(.A(n9185), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n145));
INVX1 mul_U15797(.A(dpath_mulcore_ary2_cmux_n145), .Y(n5045));
AND2X1 mul_U15798(.A(n9186), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n147));
INVX1 mul_U15799(.A(dpath_mulcore_ary2_cmux_n147), .Y(n5046));
AND2X1 mul_U15800(.A(n9187), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n149));
INVX1 mul_U15801(.A(dpath_mulcore_ary2_cmux_n149), .Y(n5047));
AND2X1 mul_U15802(.A(n6153), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n151));
INVX1 mul_U15803(.A(dpath_mulcore_ary2_cmux_n151), .Y(n5048));
AND2X1 mul_U15804(.A(n6141), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n153));
INVX1 mul_U15805(.A(dpath_mulcore_ary2_cmux_n153), .Y(n5049));
AND2X1 mul_U15806(.A(n6142), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n155));
INVX1 mul_U15807(.A(dpath_mulcore_ary2_cmux_n155), .Y(n5050));
AND2X1 mul_U15808(.A(n6143), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n157));
INVX1 mul_U15809(.A(dpath_mulcore_ary2_cmux_n157), .Y(n5051));
AND2X1 mul_U15810(.A(n6144), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n159));
INVX1 mul_U15811(.A(dpath_mulcore_ary2_cmux_n159), .Y(n5052));
AND2X1 mul_U15812(.A(n6145), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n161));
INVX1 mul_U15813(.A(dpath_mulcore_ary2_cmux_n161), .Y(n5053));
AND2X1 mul_U15814(.A(n6146), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n163));
INVX1 mul_U15815(.A(dpath_mulcore_ary2_cmux_n163), .Y(n5054));
AND2X1 mul_U15816(.A(n6147), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n165));
INVX1 mul_U15817(.A(dpath_mulcore_ary2_cmux_n165), .Y(n5055));
AND2X1 mul_U15818(.A(n6148), .B(n9706), .Y(dpath_mulcore_ary2_cmux_n167));
INVX1 mul_U15819(.A(dpath_mulcore_ary2_cmux_n167), .Y(n5056));
AND2X1 mul_U15820(.A(n6149), .B(n9680), .Y(dpath_mulcore_ary2_cmux_n169));
INVX1 mul_U15821(.A(dpath_mulcore_ary2_cmux_n169), .Y(n5057));
AND2X1 mul_U15822(.A(n6150), .B(n9680), .Y(dpath_mulcore_ary2_cmux_n171));
INVX1 mul_U15823(.A(dpath_mulcore_ary2_cmux_n171), .Y(n5058));
AND2X1 mul_U15824(.A(n6154), .B(n9680), .Y(dpath_mulcore_ary2_cmux_n173));
INVX1 mul_U15825(.A(dpath_mulcore_ary2_cmux_n173), .Y(n5059));
AND2X1 mul_U15826(.A(n6164), .B(n9700), .Y(dpath_mulcore_ary2_cmux_n175));
INVX1 mul_U15827(.A(dpath_mulcore_ary2_cmux_n175), .Y(n5060));
AND2X1 mul_U15828(.A(n6165), .B(n9696), .Y(dpath_mulcore_ary2_cmux_n177));
INVX1 mul_U15829(.A(dpath_mulcore_ary2_cmux_n177), .Y(n5061));
AND2X1 mul_U15830(.A(n6166), .B(n9681), .Y(dpath_mulcore_ary2_cmux_n179));
INVX1 mul_U15831(.A(dpath_mulcore_ary2_cmux_n179), .Y(n5062));
AND2X1 mul_U15832(.A(n6167), .B(n9701), .Y(dpath_mulcore_ary2_cmux_n181));
INVX1 mul_U15833(.A(dpath_mulcore_ary2_cmux_n181), .Y(n5063));
AND2X1 mul_U15834(.A(n16563), .B(n9698), .Y(dpath_mulcore_ary2_cmux_n183));
INVX1 mul_U15835(.A(dpath_mulcore_ary2_cmux_n183), .Y(n5064));
AND2X1 mul_U15836(.A(n6155), .B(n9682), .Y(dpath_mulcore_ary2_cmux_n185));
INVX1 mul_U15837(.A(dpath_mulcore_ary2_cmux_n185), .Y(n5065));
AND2X1 mul_U15838(.A(n6156), .B(n9680), .Y(dpath_mulcore_ary2_cmux_n187));
INVX1 mul_U15839(.A(dpath_mulcore_ary2_cmux_n187), .Y(n5066));
AND2X1 mul_U15840(.A(n6157), .B(n9699), .Y(dpath_mulcore_ary2_cmux_n189));
INVX1 mul_U15841(.A(dpath_mulcore_ary2_cmux_n189), .Y(n5067));
AND2X1 mul_U15842(.A(n6158), .B(n9700), .Y(dpath_mulcore_ary2_cmux_n191));
INVX1 mul_U15843(.A(dpath_mulcore_ary2_cmux_n191), .Y(n5068));
AND2X1 mul_U15844(.A(n6159), .B(n9696), .Y(dpath_mulcore_ary2_cmux_n193));
INVX1 mul_U15845(.A(dpath_mulcore_ary2_cmux_n193), .Y(n5069));
AND2X1 mul_U15846(.A(dpath_mulcore_pcout[0]), .B(n9681), .Y(dpath_mulcore_ary2_cmux_n195));
INVX1 mul_U15847(.A(dpath_mulcore_ary2_cmux_n195), .Y(n5070));
OR2X1 mul_U15848(.A(acc_reg_rst), .B(acc_reg_enb), .Y(dpath_ckbuf_1_enb_l));
INVX1 mul_U15849(.A(dpath_ckbuf_1_enb_l), .Y(n5071));
AND2X1 mul_U15850(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[9]), .Y(dpath_n526));
INVX1 mul_U15851(.A(dpath_n526), .Y(n5072));
AND2X1 mul_U15852(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[8]), .Y(dpath_n528));
INVX1 mul_U15853(.A(dpath_n528), .Y(n5073));
AND2X1 mul_U15854(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[7]), .Y(dpath_n530));
INVX1 mul_U15855(.A(dpath_n530), .Y(n5074));
AND2X1 mul_U15856(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[6]), .Y(dpath_n532));
INVX1 mul_U15857(.A(dpath_n532), .Y(n5075));
AND2X1 mul_U15858(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[63]), .Y(dpath_n534));
INVX1 mul_U15859(.A(dpath_n534), .Y(n5076));
AND2X1 mul_U15860(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[62]), .Y(dpath_n536));
INVX1 mul_U15861(.A(dpath_n536), .Y(n5077));
AND2X1 mul_U15862(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[61]), .Y(dpath_n538));
INVX1 mul_U15863(.A(dpath_n538), .Y(n5078));
AND2X1 mul_U15864(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[60]), .Y(dpath_n540));
INVX1 mul_U15865(.A(dpath_n540), .Y(n5079));
AND2X1 mul_U15866(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[5]), .Y(dpath_n542));
INVX1 mul_U15867(.A(dpath_n542), .Y(n5080));
AND2X1 mul_U15868(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[59]), .Y(dpath_n544));
INVX1 mul_U15869(.A(dpath_n544), .Y(n5081));
AND2X1 mul_U15870(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[58]), .Y(dpath_n546));
INVX1 mul_U15871(.A(dpath_n546), .Y(n5082));
AND2X1 mul_U15872(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[57]), .Y(dpath_n548));
INVX1 mul_U15873(.A(dpath_n548), .Y(n5083));
AND2X1 mul_U15874(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[56]), .Y(dpath_n550));
INVX1 mul_U15875(.A(dpath_n550), .Y(n5084));
AND2X1 mul_U15876(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[55]), .Y(dpath_n552));
INVX1 mul_U15877(.A(dpath_n552), .Y(n5085));
AND2X1 mul_U15878(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[54]), .Y(dpath_n554));
INVX1 mul_U15879(.A(dpath_n554), .Y(n5086));
AND2X1 mul_U15880(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[53]), .Y(dpath_n556));
INVX1 mul_U15881(.A(dpath_n556), .Y(n5087));
AND2X1 mul_U15882(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[52]), .Y(dpath_n558));
INVX1 mul_U15883(.A(dpath_n558), .Y(n5088));
AND2X1 mul_U15884(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[51]), .Y(dpath_n560));
INVX1 mul_U15885(.A(dpath_n560), .Y(n5089));
AND2X1 mul_U15886(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[50]), .Y(dpath_n562));
INVX1 mul_U15887(.A(dpath_n562), .Y(n5090));
AND2X1 mul_U15888(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[4]), .Y(dpath_n564));
INVX1 mul_U15889(.A(dpath_n564), .Y(n5091));
AND2X1 mul_U15890(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[49]), .Y(dpath_n566));
INVX1 mul_U15891(.A(dpath_n566), .Y(n5092));
AND2X1 mul_U15892(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[48]), .Y(dpath_n568));
INVX1 mul_U15893(.A(dpath_n568), .Y(n5093));
AND2X1 mul_U15894(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[47]), .Y(dpath_n570));
INVX1 mul_U15895(.A(dpath_n570), .Y(n5094));
AND2X1 mul_U15896(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[46]), .Y(dpath_n572));
INVX1 mul_U15897(.A(dpath_n572), .Y(n5095));
AND2X1 mul_U15898(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[45]), .Y(dpath_n574));
INVX1 mul_U15899(.A(dpath_n574), .Y(n5096));
AND2X1 mul_U15900(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[44]), .Y(dpath_n576));
INVX1 mul_U15901(.A(dpath_n576), .Y(n5097));
AND2X1 mul_U15902(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[43]), .Y(dpath_n578));
INVX1 mul_U15903(.A(dpath_n578), .Y(n5098));
AND2X1 mul_U15904(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[42]), .Y(dpath_n580));
INVX1 mul_U15905(.A(dpath_n580), .Y(n5099));
AND2X1 mul_U15906(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[41]), .Y(dpath_n582));
INVX1 mul_U15907(.A(dpath_n582), .Y(n5100));
AND2X1 mul_U15908(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[40]), .Y(dpath_n584));
INVX1 mul_U15909(.A(dpath_n584), .Y(n5101));
AND2X1 mul_U15910(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[3]), .Y(dpath_n586));
INVX1 mul_U15911(.A(dpath_n586), .Y(n5102));
AND2X1 mul_U15912(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[39]), .Y(dpath_n588));
INVX1 mul_U15913(.A(dpath_n588), .Y(n5103));
AND2X1 mul_U15914(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[38]), .Y(dpath_n590));
INVX1 mul_U15915(.A(dpath_n590), .Y(n5104));
AND2X1 mul_U15916(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[37]), .Y(dpath_n592));
INVX1 mul_U15917(.A(dpath_n592), .Y(n5105));
AND2X1 mul_U15918(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[36]), .Y(dpath_n594));
INVX1 mul_U15919(.A(dpath_n594), .Y(n5106));
AND2X1 mul_U15920(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[35]), .Y(dpath_n596));
INVX1 mul_U15921(.A(dpath_n596), .Y(n5107));
AND2X1 mul_U15922(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[34]), .Y(dpath_n598));
INVX1 mul_U15923(.A(dpath_n598), .Y(n5108));
AND2X1 mul_U15924(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[33]), .Y(dpath_n600));
INVX1 mul_U15925(.A(dpath_n600), .Y(n5109));
AND2X1 mul_U15926(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[32]), .Y(dpath_n602));
INVX1 mul_U15927(.A(dpath_n602), .Y(n5110));
AND2X1 mul_U15928(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[31]), .Y(dpath_n604));
INVX1 mul_U15929(.A(dpath_n604), .Y(n5111));
AND2X1 mul_U15930(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[30]), .Y(dpath_n606));
INVX1 mul_U15931(.A(dpath_n606), .Y(n5112));
AND2X1 mul_U15932(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[2]), .Y(dpath_n608));
INVX1 mul_U15933(.A(dpath_n608), .Y(n5113));
AND2X1 mul_U15934(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[29]), .Y(dpath_n610));
INVX1 mul_U15935(.A(dpath_n610), .Y(n5114));
AND2X1 mul_U15936(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[28]), .Y(dpath_n612));
INVX1 mul_U15937(.A(dpath_n612), .Y(n5115));
AND2X1 mul_U15938(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[27]), .Y(dpath_n614));
INVX1 mul_U15939(.A(dpath_n614), .Y(n5116));
AND2X1 mul_U15940(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[26]), .Y(dpath_n616));
INVX1 mul_U15941(.A(dpath_n616), .Y(n5117));
AND2X1 mul_U15942(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[25]), .Y(dpath_n618));
INVX1 mul_U15943(.A(dpath_n618), .Y(n5118));
AND2X1 mul_U15944(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[24]), .Y(dpath_n620));
INVX1 mul_U15945(.A(dpath_n620), .Y(n5119));
AND2X1 mul_U15946(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[23]), .Y(dpath_n622));
INVX1 mul_U15947(.A(dpath_n622), .Y(n5120));
AND2X1 mul_U15948(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[22]), .Y(dpath_n624));
INVX1 mul_U15949(.A(dpath_n624), .Y(n5121));
AND2X1 mul_U15950(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[21]), .Y(dpath_n626));
INVX1 mul_U15951(.A(dpath_n626), .Y(n5122));
AND2X1 mul_U15952(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[20]), .Y(dpath_n628));
INVX1 mul_U15953(.A(dpath_n628), .Y(n5123));
AND2X1 mul_U15954(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[1]), .Y(dpath_n630));
INVX1 mul_U15955(.A(dpath_n630), .Y(n5124));
AND2X1 mul_U15956(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[19]), .Y(dpath_n632));
INVX1 mul_U15957(.A(dpath_n632), .Y(n5125));
AND2X1 mul_U15958(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[18]), .Y(dpath_n634));
INVX1 mul_U15959(.A(dpath_n634), .Y(n5126));
AND2X1 mul_U15960(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[17]), .Y(dpath_n636));
INVX1 mul_U15961(.A(dpath_n636), .Y(n5127));
AND2X1 mul_U15962(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[16]), .Y(dpath_n638));
INVX1 mul_U15963(.A(dpath_n638), .Y(n5128));
AND2X1 mul_U15964(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[15]), .Y(dpath_n640));
INVX1 mul_U15965(.A(dpath_n640), .Y(n5129));
AND2X1 mul_U15966(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[14]), .Y(dpath_n642));
INVX1 mul_U15967(.A(dpath_n642), .Y(n5130));
AND2X1 mul_U15968(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[13]), .Y(dpath_n644));
INVX1 mul_U15969(.A(dpath_n644), .Y(n5131));
AND2X1 mul_U15970(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[12]), .Y(dpath_n646));
INVX1 mul_U15971(.A(dpath_n646), .Y(n5132));
AND2X1 mul_U15972(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[11]), .Y(dpath_n648));
INVX1 mul_U15973(.A(dpath_n648), .Y(n5133));
AND2X1 mul_U15974(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[10]), .Y(dpath_n650));
INVX1 mul_U15975(.A(dpath_n650), .Y(n5134));
AND2X1 mul_U15976(.A(dpath_acc_reg_shf2), .B(dpath_acc_reg[0]), .Y(dpath_n652));
INVX1 mul_U15977(.A(dpath_n652), .Y(n5135));
AND2X1 mul_U15978(.A(n9777), .B(dpath_acc_reg[73]), .Y(dpath_n986));
INVX1 mul_U15979(.A(dpath_n986), .Y(n5136));
AND2X1 mul_U15980(.A(n9777), .B(dpath_acc_reg[72]), .Y(dpath_n988));
INVX1 mul_U15981(.A(dpath_n988), .Y(n5137));
AND2X1 mul_U15982(.A(n9777), .B(dpath_acc_reg[71]), .Y(dpath_n990));
INVX1 mul_U15983(.A(dpath_n990), .Y(n5138));
AND2X1 mul_U15984(.A(dpath_acc_reg[135]), .B(acc_reg_shf), .Y(dpath_n992));
INVX1 mul_U15985(.A(dpath_n992), .Y(n5139));
AND2X1 mul_U15986(.A(dpath_acc_reg[134]), .B(acc_reg_shf), .Y(dpath_n994));
INVX1 mul_U15987(.A(dpath_n994), .Y(n5140));
AND2X1 mul_U15988(.A(n9777), .B(dpath_acc_reg[70]), .Y(dpath_n996));
INVX1 mul_U15989(.A(dpath_n996), .Y(n5141));
AND2X1 mul_U15990(.A(dpath_acc_reg[133]), .B(mul_spu_shf_ack), .Y(dpath_n998));
INVX1 mul_U15991(.A(dpath_n998), .Y(n5142));
AND2X1 mul_U15992(.A(dpath_acc_reg[132]), .B(acc_reg_shf), .Y(dpath_n1000));
INVX1 mul_U15993(.A(dpath_n1000), .Y(n5143));
AND2X1 mul_U15994(.A(dpath_acc_reg[131]), .B(acc_reg_shf), .Y(dpath_n1002));
INVX1 mul_U15995(.A(dpath_n1002), .Y(n5144));
AND2X1 mul_U15996(.A(dpath_acc_reg[130]), .B(acc_reg_shf), .Y(dpath_n1004));
INVX1 mul_U15997(.A(dpath_n1004), .Y(n5145));
AND2X1 mul_U15998(.A(dpath_acc_reg[129]), .B(mul_spu_shf_ack), .Y(dpath_n1006));
INVX1 mul_U15999(.A(dpath_n1006), .Y(n5146));
AND2X1 mul_U16000(.A(n9777), .B(dpath_acc_reg[128]), .Y(dpath_n1008));
INVX1 mul_U16001(.A(dpath_n1008), .Y(n5147));
AND2X1 mul_U16002(.A(n9777), .B(dpath_acc_reg[127]), .Y(dpath_n1010));
INVX1 mul_U16003(.A(dpath_n1010), .Y(n5148));
AND2X1 mul_U16004(.A(n9777), .B(dpath_acc_reg[126]), .Y(dpath_n1012));
INVX1 mul_U16005(.A(dpath_n1012), .Y(n5149));
AND2X1 mul_U16006(.A(n9777), .B(dpath_acc_reg[125]), .Y(dpath_n1014));
INVX1 mul_U16007(.A(dpath_n1014), .Y(n5150));
AND2X1 mul_U16008(.A(n9777), .B(dpath_acc_reg[124]), .Y(dpath_n1016));
INVX1 mul_U16009(.A(dpath_n1016), .Y(n5151));
AND2X1 mul_U16010(.A(n9777), .B(dpath_acc_reg[69]), .Y(dpath_n1018));
INVX1 mul_U16011(.A(dpath_n1018), .Y(n5152));
AND2X1 mul_U16012(.A(n9777), .B(dpath_acc_reg[123]), .Y(dpath_n1020));
INVX1 mul_U16013(.A(dpath_n1020), .Y(n5153));
AND2X1 mul_U16014(.A(n9777), .B(dpath_acc_reg[122]), .Y(dpath_n1022));
INVX1 mul_U16015(.A(dpath_n1022), .Y(n5154));
AND2X1 mul_U16016(.A(n9777), .B(dpath_acc_reg[121]), .Y(dpath_n1024));
INVX1 mul_U16017(.A(dpath_n1024), .Y(n5155));
AND2X1 mul_U16018(.A(n9777), .B(dpath_acc_reg[120]), .Y(dpath_n1026));
INVX1 mul_U16019(.A(dpath_n1026), .Y(n5156));
AND2X1 mul_U16020(.A(n9777), .B(dpath_acc_reg[119]), .Y(dpath_n1028));
INVX1 mul_U16021(.A(dpath_n1028), .Y(n5157));
AND2X1 mul_U16022(.A(n9777), .B(dpath_acc_reg[118]), .Y(dpath_n1030));
INVX1 mul_U16023(.A(dpath_n1030), .Y(n5158));
AND2X1 mul_U16024(.A(mul_spu_shf_ack), .B(dpath_acc_reg[117]), .Y(dpath_n1032));
INVX1 mul_U16025(.A(dpath_n1032), .Y(n5159));
AND2X1 mul_U16026(.A(acc_reg_shf), .B(dpath_acc_reg[116]), .Y(dpath_n1034));
INVX1 mul_U16027(.A(dpath_n1034), .Y(n5160));
AND2X1 mul_U16028(.A(n9777), .B(dpath_acc_reg[115]), .Y(dpath_n1036));
INVX1 mul_U16029(.A(dpath_n1036), .Y(n5161));
AND2X1 mul_U16030(.A(mul_spu_shf_ack), .B(dpath_acc_reg[114]), .Y(dpath_n1038));
INVX1 mul_U16031(.A(dpath_n1038), .Y(n5162));
AND2X1 mul_U16032(.A(acc_reg_shf), .B(dpath_acc_reg[68]), .Y(dpath_n1040));
INVX1 mul_U16033(.A(dpath_n1040), .Y(n5163));
AND2X1 mul_U16034(.A(n9777), .B(dpath_acc_reg[113]), .Y(dpath_n1042));
INVX1 mul_U16035(.A(dpath_n1042), .Y(n5164));
AND2X1 mul_U16036(.A(mul_spu_shf_ack), .B(dpath_acc_reg[112]), .Y(dpath_n1044));
INVX1 mul_U16037(.A(dpath_n1044), .Y(n5165));
AND2X1 mul_U16038(.A(acc_reg_shf), .B(dpath_acc_reg[111]), .Y(dpath_n1046));
INVX1 mul_U16039(.A(dpath_n1046), .Y(n5166));
AND2X1 mul_U16040(.A(n9777), .B(dpath_acc_reg[110]), .Y(dpath_n1048));
INVX1 mul_U16041(.A(dpath_n1048), .Y(n5167));
AND2X1 mul_U16042(.A(mul_spu_shf_ack), .B(dpath_acc_reg[109]), .Y(dpath_n1050));
INVX1 mul_U16043(.A(dpath_n1050), .Y(n5168));
AND2X1 mul_U16044(.A(acc_reg_shf), .B(dpath_acc_reg[108]), .Y(dpath_n1052));
INVX1 mul_U16045(.A(dpath_n1052), .Y(n5169));
AND2X1 mul_U16046(.A(n9777), .B(dpath_acc_reg[107]), .Y(dpath_n1054));
INVX1 mul_U16047(.A(dpath_n1054), .Y(n5170));
AND2X1 mul_U16048(.A(mul_spu_shf_ack), .B(dpath_acc_reg[106]), .Y(dpath_n1056));
INVX1 mul_U16049(.A(dpath_n1056), .Y(n5171));
AND2X1 mul_U16050(.A(acc_reg_shf), .B(dpath_acc_reg[105]), .Y(dpath_n1058));
INVX1 mul_U16051(.A(dpath_n1058), .Y(n5172));
AND2X1 mul_U16052(.A(n9777), .B(dpath_acc_reg[104]), .Y(dpath_n1060));
INVX1 mul_U16053(.A(dpath_n1060), .Y(n5173));
AND2X1 mul_U16054(.A(mul_spu_shf_ack), .B(dpath_acc_reg[67]), .Y(dpath_n1062));
INVX1 mul_U16055(.A(dpath_n1062), .Y(n5174));
AND2X1 mul_U16056(.A(acc_reg_shf), .B(dpath_acc_reg[103]), .Y(dpath_n1064));
INVX1 mul_U16057(.A(dpath_n1064), .Y(n5175));
AND2X1 mul_U16058(.A(n9777), .B(dpath_acc_reg[102]), .Y(dpath_n1066));
INVX1 mul_U16059(.A(dpath_n1066), .Y(n5176));
AND2X1 mul_U16060(.A(n9777), .B(dpath_acc_reg[101]), .Y(dpath_n1068));
INVX1 mul_U16061(.A(dpath_n1068), .Y(n5177));
AND2X1 mul_U16062(.A(mul_spu_shf_ack), .B(dpath_acc_reg[100]), .Y(dpath_n1070));
INVX1 mul_U16063(.A(dpath_n1070), .Y(n5178));
AND2X1 mul_U16064(.A(acc_reg_shf), .B(dpath_acc_reg[99]), .Y(dpath_n1072));
INVX1 mul_U16065(.A(dpath_n1072), .Y(n5179));
AND2X1 mul_U16066(.A(mul_spu_shf_ack), .B(dpath_acc_reg[98]), .Y(dpath_n1074));
INVX1 mul_U16067(.A(dpath_n1074), .Y(n5180));
AND2X1 mul_U16068(.A(n9777), .B(dpath_acc_reg[97]), .Y(dpath_n1076));
INVX1 mul_U16069(.A(dpath_n1076), .Y(n5181));
AND2X1 mul_U16070(.A(mul_spu_shf_ack), .B(dpath_acc_reg[96]), .Y(dpath_n1078));
INVX1 mul_U16071(.A(dpath_n1078), .Y(n5182));
AND2X1 mul_U16072(.A(acc_reg_shf), .B(dpath_acc_reg[95]), .Y(dpath_n1080));
INVX1 mul_U16073(.A(dpath_n1080), .Y(n5183));
AND2X1 mul_U16074(.A(acc_reg_shf), .B(dpath_acc_reg[94]), .Y(dpath_n1082));
INVX1 mul_U16075(.A(dpath_n1082), .Y(n5184));
AND2X1 mul_U16076(.A(n9777), .B(dpath_acc_reg[66]), .Y(dpath_n1084));
INVX1 mul_U16077(.A(dpath_n1084), .Y(n5185));
AND2X1 mul_U16078(.A(mul_spu_shf_ack), .B(dpath_acc_reg[93]), .Y(dpath_n1086));
INVX1 mul_U16079(.A(dpath_n1086), .Y(n5186));
AND2X1 mul_U16080(.A(acc_reg_shf), .B(dpath_acc_reg[92]), .Y(dpath_n1088));
INVX1 mul_U16081(.A(dpath_n1088), .Y(n5187));
AND2X1 mul_U16082(.A(mul_spu_shf_ack), .B(dpath_acc_reg[91]), .Y(dpath_n1090));
INVX1 mul_U16083(.A(dpath_n1090), .Y(n5188));
AND2X1 mul_U16084(.A(acc_reg_shf), .B(dpath_acc_reg[90]), .Y(dpath_n1092));
INVX1 mul_U16085(.A(dpath_n1092), .Y(n5189));
AND2X1 mul_U16086(.A(mul_spu_shf_ack), .B(dpath_acc_reg[89]), .Y(dpath_n1094));
INVX1 mul_U16087(.A(dpath_n1094), .Y(n5190));
AND2X1 mul_U16088(.A(acc_reg_shf), .B(dpath_acc_reg[88]), .Y(dpath_n1096));
INVX1 mul_U16089(.A(dpath_n1096), .Y(n5191));
AND2X1 mul_U16090(.A(mul_spu_shf_ack), .B(dpath_acc_reg[87]), .Y(dpath_n1098));
INVX1 mul_U16091(.A(dpath_n1098), .Y(n5192));
AND2X1 mul_U16092(.A(acc_reg_shf), .B(dpath_acc_reg[86]), .Y(dpath_n1100));
INVX1 mul_U16093(.A(dpath_n1100), .Y(n5193));
AND2X1 mul_U16094(.A(mul_spu_shf_ack), .B(dpath_acc_reg[85]), .Y(dpath_n1102));
INVX1 mul_U16095(.A(dpath_n1102), .Y(n5194));
AND2X1 mul_U16096(.A(acc_reg_shf), .B(dpath_acc_reg[84]), .Y(dpath_n1104));
INVX1 mul_U16097(.A(dpath_n1104), .Y(n5195));
AND2X1 mul_U16098(.A(mul_spu_shf_ack), .B(dpath_acc_reg[65]), .Y(dpath_n1106));
INVX1 mul_U16099(.A(dpath_n1106), .Y(n5196));
AND2X1 mul_U16100(.A(acc_reg_shf), .B(dpath_acc_reg[83]), .Y(dpath_n1108));
INVX1 mul_U16101(.A(dpath_n1108), .Y(n5197));
AND2X1 mul_U16102(.A(n9777), .B(dpath_acc_reg[82]), .Y(dpath_n1110));
INVX1 mul_U16103(.A(dpath_n1110), .Y(n5198));
AND2X1 mul_U16104(.A(n9777), .B(dpath_acc_reg[81]), .Y(dpath_n1112));
INVX1 mul_U16105(.A(dpath_n1112), .Y(n5199));
AND2X1 mul_U16106(.A(acc_reg_shf), .B(dpath_acc_reg[80]), .Y(dpath_n1114));
INVX1 mul_U16107(.A(dpath_n1114), .Y(n5200));
AND2X1 mul_U16108(.A(mul_spu_shf_ack), .B(dpath_acc_reg[79]), .Y(dpath_n1116));
INVX1 mul_U16109(.A(dpath_n1116), .Y(n5201));
AND2X1 mul_U16110(.A(acc_reg_shf), .B(dpath_acc_reg[78]), .Y(dpath_n1118));
INVX1 mul_U16111(.A(dpath_n1118), .Y(n5202));
AND2X1 mul_U16112(.A(mul_spu_shf_ack), .B(dpath_acc_reg[77]), .Y(dpath_n1120));
INVX1 mul_U16113(.A(dpath_n1120), .Y(n5203));
AND2X1 mul_U16114(.A(mul_spu_shf_ack), .B(dpath_acc_reg[76]), .Y(dpath_n1122));
INVX1 mul_U16115(.A(dpath_n1122), .Y(n5204));
AND2X1 mul_U16116(.A(mul_spu_shf_ack), .B(dpath_acc_reg[75]), .Y(dpath_n1124));
INVX1 mul_U16117(.A(dpath_n1124), .Y(n5205));
AND2X1 mul_U16118(.A(mul_spu_shf_ack), .B(dpath_acc_reg[74]), .Y(dpath_n1126));
INVX1 mul_U16119(.A(dpath_n1126), .Y(n5206));
AND2X1 mul_U16120(.A(mul_spu_shf_ack), .B(dpath_acc_reg[64]), .Y(dpath_n1128));
INVX1 mul_U16121(.A(dpath_n1128), .Y(n5207));
AND2X1 mul_U16122(.A(n5829), .B(n9818), .Y(control_n24));
INVX1 mul_U16123(.A(control_n24), .Y(n5208));
AND2X1 mul_U16124(.A(n16568), .B(n16571), .Y(n15173));
INVX1 mul_U16125(.A(n15173), .Y(n5209));
AND2X1 mul_U16126(.A(n8286), .B(dpath_mulcore_ary1_a0_s_1[10]), .Y(n15185));
INVX1 mul_U16127(.A(n15185), .Y(n5210));
AND2X1 mul_U16128(.A(n8287), .B(dpath_mulcore_ary1_a0_s_1[9]), .Y(n15188));
INVX1 mul_U16129(.A(n15188), .Y(n5211));
AND2X1 mul_U16130(.A(n8293), .B(dpath_mulcore_ary1_a0_s_1[8]), .Y(n15191));
INVX1 mul_U16131(.A(n15191), .Y(n5212));
AND2X1 mul_U16132(.A(dpath_mulcore_ary1_a1_s2[65]), .B(n8941), .Y(n15573));
INVX1 mul_U16133(.A(n15573), .Y(n5213));
AND2X1 mul_U16134(.A(n8295), .B(dpath_mulcore_ary1_a1_s_1[10]), .Y(n15585));
INVX1 mul_U16135(.A(n15585), .Y(n5214));
AND2X1 mul_U16136(.A(n8296), .B(dpath_mulcore_ary1_a1_s_1[9]), .Y(n15588));
INVX1 mul_U16137(.A(n15588), .Y(n5215));
AND2X1 mul_U16138(.A(n8302), .B(dpath_mulcore_ary1_a1_s_1[8]), .Y(n15591));
INVX1 mul_U16139(.A(n15591), .Y(n5216));
AND2X1 mul_U16140(.A(dpath_mulcore_a1s[81]), .B(dpath_mulcore_a1c[80]), .Y(n16029));
INVX1 mul_U16141(.A(n16029), .Y(n5217));
AND2X1 mul_U16142(.A(dpath_mulcore_ary1_a0_sc3_75__z), .B(n16592), .Y(n16589));
INVX1 mul_U16143(.A(n16589), .Y(n5218));
AND2X1 mul_U16144(.A(dpath_mulcore_ary1_a0_sc3_74__z), .B(n16596), .Y(n16593));
INVX1 mul_U16145(.A(n16593), .Y(n5219));
AND2X1 mul_U16146(.A(dpath_mulcore_ary1_a0_sc3_73__z), .B(n16600), .Y(n16597));
INVX1 mul_U16147(.A(n16597), .Y(n5220));
AND2X1 mul_U16148(.A(dpath_mulcore_ary1_a0_sc3_72__z), .B(n7395), .Y(n16601));
INVX1 mul_U16149(.A(n16601), .Y(n5221));
AND2X1 mul_U16150(.A(dpath_mulcore_ary1_a0_sc3_76__z), .B(n16588), .Y(n16604));
INVX1 mul_U16151(.A(n16604), .Y(n5222));
AND2X1 mul_U16152(.A(dpath_mulcore_ary1_a0_sc3_70__z), .B(n7228), .Y(n16609));
INVX1 mul_U16153(.A(n16609), .Y(n5223));
AND2X1 mul_U16154(.A(dpath_mulcore_ary1_a0_sc3_69__z), .B(n7229), .Y(n16616));
INVX1 mul_U16155(.A(n16616), .Y(n5224));
AND2X1 mul_U16156(.A(dpath_mulcore_ary1_a0_sc3_68__z), .B(n7230), .Y(n16623));
INVX1 mul_U16157(.A(n16623), .Y(n5225));
AND2X1 mul_U16158(.A(dpath_mulcore_ary1_a0_sc3_67__z), .B(n7231), .Y(n16630));
INVX1 mul_U16159(.A(n16630), .Y(n5226));
AND2X1 mul_U16160(.A(dpath_mulcore_ary1_a0_sc3_66__z), .B(n7232), .Y(n16637));
INVX1 mul_U16161(.A(n16637), .Y(n5227));
AND2X1 mul_U16162(.A(dpath_mulcore_ary1_a0_sc3_65__z), .B(n7233), .Y(n16644));
INVX1 mul_U16163(.A(n16644), .Y(n5228));
AND2X1 mul_U16164(.A(dpath_mulcore_ary1_a0_sc3_64__z), .B(n7234), .Y(n16651));
INVX1 mul_U16165(.A(n16651), .Y(n5229));
AND2X1 mul_U16166(.A(dpath_mulcore_ary1_a0_sc3_63__z), .B(n7235), .Y(n16658));
INVX1 mul_U16167(.A(n16658), .Y(n5230));
AND2X1 mul_U16168(.A(dpath_mulcore_ary1_a0_sc3_62__z), .B(n7236), .Y(n16665));
INVX1 mul_U16169(.A(n16665), .Y(n5231));
AND2X1 mul_U16170(.A(dpath_mulcore_ary1_a0_sc3_61__z), .B(n7237), .Y(n16672));
INVX1 mul_U16171(.A(n16672), .Y(n5232));
AND2X1 mul_U16172(.A(dpath_mulcore_ary1_a0_sc3_60__z), .B(n7238), .Y(n16679));
INVX1 mul_U16173(.A(n16679), .Y(n5233));
AND2X1 mul_U16174(.A(dpath_mulcore_ary1_a0_sc3_59__z), .B(n7239), .Y(n16686));
INVX1 mul_U16175(.A(n16686), .Y(n5234));
AND2X1 mul_U16176(.A(dpath_mulcore_ary1_a0_sc3_58__z), .B(n7240), .Y(n16693));
INVX1 mul_U16177(.A(n16693), .Y(n5235));
AND2X1 mul_U16178(.A(dpath_mulcore_ary1_a0_sc3_57__z), .B(n7241), .Y(n16700));
INVX1 mul_U16179(.A(n16700), .Y(n5236));
AND2X1 mul_U16180(.A(dpath_mulcore_ary1_a0_sc3_56__z), .B(n7242), .Y(n16707));
INVX1 mul_U16181(.A(n16707), .Y(n5237));
AND2X1 mul_U16182(.A(dpath_mulcore_ary1_a0_sc3_55__z), .B(n7243), .Y(n16714));
INVX1 mul_U16183(.A(n16714), .Y(n5238));
AND2X1 mul_U16184(.A(dpath_mulcore_ary1_a0_sc3_54__z), .B(n7244), .Y(n16721));
INVX1 mul_U16185(.A(n16721), .Y(n5239));
AND2X1 mul_U16186(.A(dpath_mulcore_ary1_a0_sc3_53__z), .B(n7245), .Y(n16728));
INVX1 mul_U16187(.A(n16728), .Y(n5240));
AND2X1 mul_U16188(.A(dpath_mulcore_ary1_a0_sc3_52__z), .B(n7246), .Y(n16735));
INVX1 mul_U16189(.A(n16735), .Y(n5241));
AND2X1 mul_U16190(.A(dpath_mulcore_ary1_a0_sc3_51__z), .B(n7247), .Y(n16742));
INVX1 mul_U16191(.A(n16742), .Y(n5242));
AND2X1 mul_U16192(.A(dpath_mulcore_ary1_a0_sc3_50__z), .B(n7248), .Y(n16749));
INVX1 mul_U16193(.A(n16749), .Y(n5243));
AND2X1 mul_U16194(.A(dpath_mulcore_ary1_a0_sc3_49__z), .B(n7249), .Y(n16756));
INVX1 mul_U16195(.A(n16756), .Y(n5244));
AND2X1 mul_U16196(.A(dpath_mulcore_ary1_a0_sc3_48__z), .B(n7250), .Y(n16763));
INVX1 mul_U16197(.A(n16763), .Y(n5245));
AND2X1 mul_U16198(.A(dpath_mulcore_ary1_a0_sc3_47__z), .B(n7251), .Y(n16770));
INVX1 mul_U16199(.A(n16770), .Y(n5246));
AND2X1 mul_U16200(.A(dpath_mulcore_ary1_a0_sc3_46__z), .B(n7252), .Y(n16777));
INVX1 mul_U16201(.A(n16777), .Y(n5247));
AND2X1 mul_U16202(.A(dpath_mulcore_ary1_a0_sc3_45__z), .B(n7253), .Y(n16784));
INVX1 mul_U16203(.A(n16784), .Y(n5248));
AND2X1 mul_U16204(.A(dpath_mulcore_ary1_a0_sc3_44__z), .B(n7254), .Y(n16791));
INVX1 mul_U16205(.A(n16791), .Y(n5249));
AND2X1 mul_U16206(.A(dpath_mulcore_ary1_a0_sc3_43__z), .B(n7255), .Y(n16798));
INVX1 mul_U16207(.A(n16798), .Y(n5250));
AND2X1 mul_U16208(.A(dpath_mulcore_ary1_a0_sc3_42__z), .B(n7256), .Y(n16805));
INVX1 mul_U16209(.A(n16805), .Y(n5251));
AND2X1 mul_U16210(.A(dpath_mulcore_ary1_a0_sc3_41__z), .B(n7257), .Y(n16812));
INVX1 mul_U16211(.A(n16812), .Y(n5252));
AND2X1 mul_U16212(.A(dpath_mulcore_ary1_a0_sc3_40__z), .B(n7258), .Y(n16819));
INVX1 mul_U16213(.A(n16819), .Y(n5253));
AND2X1 mul_U16214(.A(dpath_mulcore_ary1_a0_sc3_39__z), .B(n7259), .Y(n16826));
INVX1 mul_U16215(.A(n16826), .Y(n5254));
AND2X1 mul_U16216(.A(dpath_mulcore_ary1_a0_sc3_38__z), .B(n7260), .Y(n16833));
INVX1 mul_U16217(.A(n16833), .Y(n5255));
AND2X1 mul_U16218(.A(dpath_mulcore_ary1_a0_sc3_37__z), .B(n7261), .Y(n16840));
INVX1 mul_U16219(.A(n16840), .Y(n5256));
AND2X1 mul_U16220(.A(dpath_mulcore_ary1_a0_sc3_36__z), .B(n7262), .Y(n16847));
INVX1 mul_U16221(.A(n16847), .Y(n5257));
AND2X1 mul_U16222(.A(dpath_mulcore_ary1_a0_sc3_35__z), .B(n7263), .Y(n16854));
INVX1 mul_U16223(.A(n16854), .Y(n5258));
AND2X1 mul_U16224(.A(dpath_mulcore_ary1_a0_sc3_34__z), .B(n7264), .Y(n16861));
INVX1 mul_U16225(.A(n16861), .Y(n5259));
AND2X1 mul_U16226(.A(dpath_mulcore_ary1_a0_sc3_33__z), .B(n7265), .Y(n16868));
INVX1 mul_U16227(.A(n16868), .Y(n5260));
AND2X1 mul_U16228(.A(dpath_mulcore_ary1_a0_sc3_32__z), .B(n7266), .Y(n16875));
INVX1 mul_U16229(.A(n16875), .Y(n5261));
AND2X1 mul_U16230(.A(dpath_mulcore_ary1_a0_sc3_31__z), .B(n7267), .Y(n16882));
INVX1 mul_U16231(.A(n16882), .Y(n5262));
AND2X1 mul_U16232(.A(dpath_mulcore_ary1_a0_sc3_30__z), .B(n7268), .Y(n16889));
INVX1 mul_U16233(.A(n16889), .Y(n5263));
AND2X1 mul_U16234(.A(dpath_mulcore_ary1_a0_sc3_29__z), .B(n7269), .Y(n16896));
INVX1 mul_U16235(.A(n16896), .Y(n5264));
AND2X1 mul_U16236(.A(dpath_mulcore_ary1_a0_sc3_28__z), .B(n7270), .Y(n16903));
INVX1 mul_U16237(.A(n16903), .Y(n5265));
AND2X1 mul_U16238(.A(dpath_mulcore_ary1_a0_sc3_27__z), .B(n7271), .Y(n16910));
INVX1 mul_U16239(.A(n16910), .Y(n5266));
AND2X1 mul_U16240(.A(dpath_mulcore_ary1_a0_sc3_26__z), .B(n7272), .Y(n16917));
INVX1 mul_U16241(.A(n16917), .Y(n5267));
AND2X1 mul_U16242(.A(dpath_mulcore_ary1_a0_sc3_25__z), .B(n7273), .Y(n16924));
INVX1 mul_U16243(.A(n16924), .Y(n5268));
AND2X1 mul_U16244(.A(dpath_mulcore_ary1_a0_sc3_24__z), .B(n7274), .Y(n16931));
INVX1 mul_U16245(.A(n16931), .Y(n5269));
AND2X1 mul_U16246(.A(dpath_mulcore_ary1_a0_sc3_23__z), .B(n7275), .Y(n16938));
INVX1 mul_U16247(.A(n16938), .Y(n5270));
AND2X1 mul_U16248(.A(dpath_mulcore_ary1_a0_sc3_22__z), .B(n7276), .Y(n16945));
INVX1 mul_U16249(.A(n16945), .Y(n5271));
AND2X1 mul_U16250(.A(dpath_mulcore_ary1_a0_sc3_21__z), .B(n7277), .Y(n16952));
INVX1 mul_U16251(.A(n16952), .Y(n5272));
AND2X1 mul_U16252(.A(dpath_mulcore_ary1_a0_sc3_20__z), .B(n7278), .Y(n16959));
INVX1 mul_U16253(.A(n16959), .Y(n5273));
AND2X1 mul_U16254(.A(dpath_mulcore_ary1_a0_sc3_19__z), .B(n7279), .Y(n16966));
INVX1 mul_U16255(.A(n16966), .Y(n5274));
AND2X1 mul_U16256(.A(dpath_mulcore_ary1_a0_sc3_18__z), .B(n7280), .Y(n16973));
INVX1 mul_U16257(.A(n16973), .Y(n5275));
AND2X1 mul_U16258(.A(dpath_mulcore_ary1_a0_sc3_17__z), .B(n7281), .Y(n16980));
INVX1 mul_U16259(.A(n16980), .Y(n5276));
AND2X1 mul_U16260(.A(dpath_mulcore_ary1_a0_sc3_16__z), .B(n7282), .Y(n16987));
INVX1 mul_U16261(.A(n16987), .Y(n5277));
AND2X1 mul_U16262(.A(dpath_mulcore_ary1_a0_sc3_15__z), .B(n7283), .Y(n16994));
INVX1 mul_U16263(.A(n16994), .Y(n5278));
AND2X1 mul_U16264(.A(dpath_mulcore_ary1_a0_sc3_14__z), .B(n7284), .Y(n17001));
INVX1 mul_U16265(.A(n17001), .Y(n5279));
AND2X1 mul_U16266(.A(dpath_mulcore_ary1_a0_sc3_13__z), .B(n7285), .Y(n17008));
INVX1 mul_U16267(.A(n17008), .Y(n5280));
AND2X1 mul_U16268(.A(dpath_mulcore_ary1_a0_sc3_12__z), .B(n7286), .Y(n17015));
INVX1 mul_U16269(.A(n17015), .Y(n5281));
AND2X1 mul_U16270(.A(dpath_mulcore_ary1_a1_sc3_71__z), .B(n7288), .Y(n17028));
INVX1 mul_U16271(.A(n17028), .Y(n5282));
AND2X1 mul_U16272(.A(dpath_mulcore_ary1_a1_sc3_75__z), .B(n17036), .Y(n17033));
INVX1 mul_U16273(.A(n17033), .Y(n5283));
AND2X1 mul_U16274(.A(dpath_mulcore_ary1_a1_sc3_74__z), .B(n17040), .Y(n17037));
INVX1 mul_U16275(.A(n17037), .Y(n5284));
AND2X1 mul_U16276(.A(dpath_mulcore_ary1_a1_sc3_73__z), .B(n17044), .Y(n17041));
INVX1 mul_U16277(.A(n17041), .Y(n5285));
AND2X1 mul_U16278(.A(dpath_mulcore_ary1_a1_sc3_72__z), .B(n7287), .Y(n17045));
INVX1 mul_U16279(.A(n17045), .Y(n5286));
AND2X1 mul_U16280(.A(dpath_mulcore_ary1_a1_sc3_76__z), .B(n17032), .Y(n17048));
INVX1 mul_U16281(.A(n17048), .Y(n5287));
AND2X1 mul_U16282(.A(dpath_mulcore_ary1_a1_sc3_70__z), .B(n7289), .Y(n17053));
INVX1 mul_U16283(.A(n17053), .Y(n5288));
AND2X1 mul_U16284(.A(dpath_mulcore_ary1_a1_sc3_69__z), .B(n7290), .Y(n17060));
INVX1 mul_U16285(.A(n17060), .Y(n5289));
AND2X1 mul_U16286(.A(dpath_mulcore_ary1_a1_sc3_68__z), .B(n7291), .Y(n17067));
INVX1 mul_U16287(.A(n17067), .Y(n5290));
AND2X1 mul_U16288(.A(dpath_mulcore_ary1_a1_sc3_67__z), .B(n7292), .Y(n17074));
INVX1 mul_U16289(.A(n17074), .Y(n5291));
AND2X1 mul_U16290(.A(dpath_mulcore_ary1_a1_sc3_66__z), .B(n7293), .Y(n17081));
INVX1 mul_U16291(.A(n17081), .Y(n5292));
AND2X1 mul_U16292(.A(dpath_mulcore_ary1_a1_sc3_65__z), .B(n7294), .Y(n17088));
INVX1 mul_U16293(.A(n17088), .Y(n5293));
AND2X1 mul_U16294(.A(dpath_mulcore_ary1_a1_sc3_64__z), .B(n7295), .Y(n17095));
INVX1 mul_U16295(.A(n17095), .Y(n5294));
AND2X1 mul_U16296(.A(dpath_mulcore_ary1_a1_sc3_63__z), .B(n7296), .Y(n17102));
INVX1 mul_U16297(.A(n17102), .Y(n5295));
AND2X1 mul_U16298(.A(dpath_mulcore_ary1_a1_sc3_62__z), .B(n7297), .Y(n17109));
INVX1 mul_U16299(.A(n17109), .Y(n5296));
AND2X1 mul_U16300(.A(dpath_mulcore_ary1_a1_sc3_61__z), .B(n7298), .Y(n17116));
INVX1 mul_U16301(.A(n17116), .Y(n5297));
AND2X1 mul_U16302(.A(dpath_mulcore_ary1_a1_sc3_60__z), .B(n7299), .Y(n17123));
INVX1 mul_U16303(.A(n17123), .Y(n5298));
AND2X1 mul_U16304(.A(dpath_mulcore_ary1_a1_sc3_59__z), .B(n7300), .Y(n17130));
INVX1 mul_U16305(.A(n17130), .Y(n5299));
AND2X1 mul_U16306(.A(dpath_mulcore_ary1_a1_sc3_58__z), .B(n7301), .Y(n17137));
INVX1 mul_U16307(.A(n17137), .Y(n5300));
AND2X1 mul_U16308(.A(dpath_mulcore_ary1_a1_sc3_57__z), .B(n7302), .Y(n17144));
INVX1 mul_U16309(.A(n17144), .Y(n5301));
AND2X1 mul_U16310(.A(dpath_mulcore_ary1_a1_sc3_56__z), .B(n7303), .Y(n17151));
INVX1 mul_U16311(.A(n17151), .Y(n5302));
AND2X1 mul_U16312(.A(dpath_mulcore_ary1_a1_sc3_55__z), .B(n7304), .Y(n17158));
INVX1 mul_U16313(.A(n17158), .Y(n5303));
AND2X1 mul_U16314(.A(dpath_mulcore_ary1_a1_sc3_54__z), .B(n7305), .Y(n17165));
INVX1 mul_U16315(.A(n17165), .Y(n5304));
AND2X1 mul_U16316(.A(dpath_mulcore_ary1_a1_sc3_53__z), .B(n7306), .Y(n17172));
INVX1 mul_U16317(.A(n17172), .Y(n5305));
AND2X1 mul_U16318(.A(dpath_mulcore_ary1_a1_sc3_52__z), .B(n7307), .Y(n17179));
INVX1 mul_U16319(.A(n17179), .Y(n5306));
AND2X1 mul_U16320(.A(dpath_mulcore_ary1_a1_sc3_51__z), .B(n7308), .Y(n17186));
INVX1 mul_U16321(.A(n17186), .Y(n5307));
AND2X1 mul_U16322(.A(dpath_mulcore_ary1_a1_sc3_50__z), .B(n7309), .Y(n17193));
INVX1 mul_U16323(.A(n17193), .Y(n5308));
AND2X1 mul_U16324(.A(dpath_mulcore_ary1_a1_sc3_49__z), .B(n7310), .Y(n17200));
INVX1 mul_U16325(.A(n17200), .Y(n5309));
AND2X1 mul_U16326(.A(dpath_mulcore_ary1_a1_sc3_48__z), .B(n7311), .Y(n17207));
INVX1 mul_U16327(.A(n17207), .Y(n5310));
AND2X1 mul_U16328(.A(dpath_mulcore_ary1_a1_sc3_47__z), .B(n7312), .Y(n17214));
INVX1 mul_U16329(.A(n17214), .Y(n5311));
AND2X1 mul_U16330(.A(dpath_mulcore_ary1_a1_sc3_46__z), .B(n7313), .Y(n17221));
INVX1 mul_U16331(.A(n17221), .Y(n5312));
AND2X1 mul_U16332(.A(dpath_mulcore_ary1_a1_sc3_45__z), .B(n7314), .Y(n17228));
INVX1 mul_U16333(.A(n17228), .Y(n5313));
AND2X1 mul_U16334(.A(dpath_mulcore_ary1_a1_sc3_44__z), .B(n7315), .Y(n17235));
INVX1 mul_U16335(.A(n17235), .Y(n5314));
AND2X1 mul_U16336(.A(dpath_mulcore_ary1_a1_sc3_43__z), .B(n7316), .Y(n17242));
INVX1 mul_U16337(.A(n17242), .Y(n5315));
AND2X1 mul_U16338(.A(dpath_mulcore_ary1_a1_sc3_42__z), .B(n7317), .Y(n17249));
INVX1 mul_U16339(.A(n17249), .Y(n5316));
AND2X1 mul_U16340(.A(dpath_mulcore_ary1_a1_sc3_41__z), .B(n7318), .Y(n17256));
INVX1 mul_U16341(.A(n17256), .Y(n5317));
AND2X1 mul_U16342(.A(dpath_mulcore_ary1_a1_sc3_40__z), .B(n7319), .Y(n17263));
INVX1 mul_U16343(.A(n17263), .Y(n5318));
AND2X1 mul_U16344(.A(dpath_mulcore_ary1_a1_sc3_39__z), .B(n7320), .Y(n17270));
INVX1 mul_U16345(.A(n17270), .Y(n5319));
AND2X1 mul_U16346(.A(dpath_mulcore_ary1_a1_sc3_38__z), .B(n7321), .Y(n17277));
INVX1 mul_U16347(.A(n17277), .Y(n5320));
AND2X1 mul_U16348(.A(dpath_mulcore_ary1_a1_sc3_37__z), .B(n7322), .Y(n17284));
INVX1 mul_U16349(.A(n17284), .Y(n5321));
AND2X1 mul_U16350(.A(dpath_mulcore_ary1_a1_sc3_36__z), .B(n7323), .Y(n17291));
INVX1 mul_U16351(.A(n17291), .Y(n5322));
AND2X1 mul_U16352(.A(dpath_mulcore_ary1_a1_sc3_35__z), .B(n7324), .Y(n17298));
INVX1 mul_U16353(.A(n17298), .Y(n5323));
AND2X1 mul_U16354(.A(dpath_mulcore_ary1_a1_sc3_34__z), .B(n7325), .Y(n17305));
INVX1 mul_U16355(.A(n17305), .Y(n5324));
AND2X1 mul_U16356(.A(dpath_mulcore_ary1_a1_sc3_33__z), .B(n7326), .Y(n17312));
INVX1 mul_U16357(.A(n17312), .Y(n5325));
AND2X1 mul_U16358(.A(dpath_mulcore_ary1_a1_sc3_32__z), .B(n7327), .Y(n17319));
INVX1 mul_U16359(.A(n17319), .Y(n5326));
AND2X1 mul_U16360(.A(dpath_mulcore_ary1_a1_sc3_31__z), .B(n7328), .Y(n17326));
INVX1 mul_U16361(.A(n17326), .Y(n5327));
AND2X1 mul_U16362(.A(dpath_mulcore_ary1_a1_sc3_30__z), .B(n7329), .Y(n17333));
INVX1 mul_U16363(.A(n17333), .Y(n5328));
AND2X1 mul_U16364(.A(dpath_mulcore_ary1_a1_sc3_29__z), .B(n7330), .Y(n17340));
INVX1 mul_U16365(.A(n17340), .Y(n5329));
AND2X1 mul_U16366(.A(dpath_mulcore_ary1_a1_sc3_28__z), .B(n7331), .Y(n17347));
INVX1 mul_U16367(.A(n17347), .Y(n5330));
AND2X1 mul_U16368(.A(dpath_mulcore_ary1_a1_sc3_27__z), .B(n7332), .Y(n17354));
INVX1 mul_U16369(.A(n17354), .Y(n5331));
AND2X1 mul_U16370(.A(dpath_mulcore_ary1_a1_sc3_26__z), .B(n7333), .Y(n17361));
INVX1 mul_U16371(.A(n17361), .Y(n5332));
AND2X1 mul_U16372(.A(dpath_mulcore_ary1_a1_sc3_25__z), .B(n7334), .Y(n17368));
INVX1 mul_U16373(.A(n17368), .Y(n5333));
AND2X1 mul_U16374(.A(dpath_mulcore_ary1_a1_sc3_24__z), .B(n7335), .Y(n17375));
INVX1 mul_U16375(.A(n17375), .Y(n5334));
AND2X1 mul_U16376(.A(dpath_mulcore_ary1_a1_sc3_23__z), .B(n7336), .Y(n17382));
INVX1 mul_U16377(.A(n17382), .Y(n5335));
AND2X1 mul_U16378(.A(dpath_mulcore_ary1_a1_sc3_22__z), .B(n7337), .Y(n17389));
INVX1 mul_U16379(.A(n17389), .Y(n5336));
AND2X1 mul_U16380(.A(dpath_mulcore_ary1_a1_sc3_21__z), .B(n7338), .Y(n17396));
INVX1 mul_U16381(.A(n17396), .Y(n5337));
AND2X1 mul_U16382(.A(dpath_mulcore_ary1_a1_sc3_20__z), .B(n7339), .Y(n17403));
INVX1 mul_U16383(.A(n17403), .Y(n5338));
AND2X1 mul_U16384(.A(dpath_mulcore_ary1_a1_sc3_19__z), .B(n7340), .Y(n17410));
INVX1 mul_U16385(.A(n17410), .Y(n5339));
AND2X1 mul_U16386(.A(dpath_mulcore_ary1_a1_sc3_18__z), .B(n7341), .Y(n17417));
INVX1 mul_U16387(.A(n17417), .Y(n5340));
AND2X1 mul_U16388(.A(dpath_mulcore_ary1_a1_sc3_17__z), .B(n7342), .Y(n17424));
INVX1 mul_U16389(.A(n17424), .Y(n5341));
AND2X1 mul_U16390(.A(dpath_mulcore_ary1_a1_sc3_16__z), .B(n7343), .Y(n17431));
INVX1 mul_U16391(.A(n17431), .Y(n5342));
AND2X1 mul_U16392(.A(dpath_mulcore_ary1_a1_sc3_15__z), .B(n7344), .Y(n17438));
INVX1 mul_U16393(.A(n17438), .Y(n5343));
AND2X1 mul_U16394(.A(dpath_mulcore_ary1_a1_sc3_14__z), .B(n7345), .Y(n17445));
INVX1 mul_U16395(.A(n17445), .Y(n5344));
AND2X1 mul_U16396(.A(dpath_mulcore_ary1_a1_sc3_13__z), .B(n7346), .Y(n17452));
INVX1 mul_U16397(.A(n17452), .Y(n5345));
AND2X1 mul_U16398(.A(dpath_mulcore_ary1_a1_sc3_12__z), .B(n7347), .Y(n17459));
INVX1 mul_U16399(.A(n17459), .Y(n5346));
AND2X1 mul_U16400(.A(c0_act), .B(dpath_mulcore_booth_b1_in1[2]), .Y(n17858));
INVX1 mul_U16401(.A(n17858), .Y(n5347));
AND2X1 mul_U16402(.A(n5424), .B(c0_act), .Y(n17860));
INVX1 mul_U16403(.A(n17860), .Y(n5348));
AND2X1 mul_U16404(.A(n5438), .B(c0_act), .Y(n17862));
INVX1 mul_U16405(.A(n17862), .Y(n5349));
AND2X1 mul_U16406(.A(c0_act), .B(dpath_mulcore_booth_b2_in1[2]), .Y(n17864));
INVX1 mul_U16407(.A(n17864), .Y(n5350));
AND2X1 mul_U16408(.A(n5423), .B(c0_act), .Y(n17866));
INVX1 mul_U16409(.A(n17866), .Y(n5351));
AND2X1 mul_U16410(.A(n5436), .B(c0_act), .Y(n17868));
INVX1 mul_U16411(.A(n17868), .Y(n5352));
AND2X1 mul_U16412(.A(c0_act), .B(dpath_mulcore_booth_b3_in1[2]), .Y(n17870));
INVX1 mul_U16413(.A(n17870), .Y(n5353));
AND2X1 mul_U16414(.A(n5422), .B(c0_act), .Y(n17872));
INVX1 mul_U16415(.A(n17872), .Y(n5354));
AND2X1 mul_U16416(.A(n5434), .B(c0_act), .Y(n17874));
INVX1 mul_U16417(.A(n17874), .Y(n5355));
AND2X1 mul_U16418(.A(c0_act), .B(dpath_mulcore_booth_b4_in1[2]), .Y(n17876));
INVX1 mul_U16419(.A(n17876), .Y(n5356));
AND2X1 mul_U16420(.A(n5421), .B(c0_act), .Y(n17878));
INVX1 mul_U16421(.A(n17878), .Y(n5357));
AND2X1 mul_U16422(.A(n5432), .B(c0_act), .Y(n17880));
INVX1 mul_U16423(.A(n17880), .Y(n5358));
AND2X1 mul_U16424(.A(c0_act), .B(dpath_mulcore_booth_b5_in1[2]), .Y(n17882));
INVX1 mul_U16425(.A(n17882), .Y(n5359));
AND2X1 mul_U16426(.A(n5420), .B(c0_act), .Y(n17884));
INVX1 mul_U16427(.A(n17884), .Y(n5360));
AND2X1 mul_U16428(.A(n5430), .B(c0_act), .Y(n17886));
INVX1 mul_U16429(.A(n17886), .Y(n5361));
AND2X1 mul_U16430(.A(c0_act), .B(dpath_mulcore_booth_b6_in1[2]), .Y(n17888));
INVX1 mul_U16431(.A(n17888), .Y(n5362));
AND2X1 mul_U16432(.A(n5419), .B(c0_act), .Y(n17890));
INVX1 mul_U16433(.A(n17890), .Y(n5363));
AND2X1 mul_U16434(.A(n5428), .B(c0_act), .Y(n17892));
INVX1 mul_U16435(.A(n17892), .Y(n5364));
AND2X1 mul_U16436(.A(c0_act), .B(dpath_mulcore_booth_b7_in1[2]), .Y(n17894));
INVX1 mul_U16437(.A(n17894), .Y(n5365));
AND2X1 mul_U16438(.A(n5418), .B(c0_act), .Y(n17896));
INVX1 mul_U16439(.A(n17896), .Y(n5366));
AND2X1 mul_U16440(.A(n5425), .B(c0_act), .Y(n17898));
INVX1 mul_U16441(.A(n17898), .Y(n5367));
AND2X1 mul_U16442(.A(c0_act), .B(dpath_mulcore_booth_b8_in1[2]), .Y(n17900));
INVX1 mul_U16443(.A(n17900), .Y(n5368));
AND2X1 mul_U16444(.A(n5443), .B(c0_act), .Y(n17902));
INVX1 mul_U16445(.A(n17902), .Y(n5369));
AND2X1 mul_U16446(.A(n5467), .B(c0_act), .Y(n17904));
INVX1 mul_U16447(.A(n17904), .Y(n5370));
AND2X1 mul_U16448(.A(c0_act), .B(dpath_mulcore_booth_b9_in1[2]), .Y(n17906));
INVX1 mul_U16449(.A(n17906), .Y(n5371));
AND2X1 mul_U16450(.A(n5450), .B(c0_act), .Y(n17908));
INVX1 mul_U16451(.A(n17908), .Y(n5372));
AND2X1 mul_U16452(.A(n5464), .B(c0_act), .Y(n17910));
INVX1 mul_U16453(.A(n17910), .Y(n5373));
AND2X1 mul_U16454(.A(c0_act), .B(dpath_mulcore_booth_b10_in1[2]), .Y(n17912));
INVX1 mul_U16455(.A(n17912), .Y(n5374));
AND2X1 mul_U16456(.A(n5449), .B(c0_act), .Y(n17914));
INVX1 mul_U16457(.A(n17914), .Y(n5375));
AND2X1 mul_U16458(.A(n5462), .B(c0_act), .Y(n17916));
INVX1 mul_U16459(.A(n17916), .Y(n5376));
AND2X1 mul_U16460(.A(c0_act), .B(dpath_mulcore_booth_b11_in1[2]), .Y(n17918));
INVX1 mul_U16461(.A(n17918), .Y(n5377));
AND2X1 mul_U16462(.A(n5448), .B(c0_act), .Y(n17920));
INVX1 mul_U16463(.A(n17920), .Y(n5378));
AND2X1 mul_U16464(.A(n5460), .B(c0_act), .Y(n17922));
INVX1 mul_U16465(.A(n17922), .Y(n5379));
AND2X1 mul_U16466(.A(c0_act), .B(dpath_mulcore_booth_b12_in1[2]), .Y(n17924));
INVX1 mul_U16467(.A(n17924), .Y(n5380));
AND2X1 mul_U16468(.A(n5447), .B(c0_act), .Y(n17926));
INVX1 mul_U16469(.A(n17926), .Y(n5381));
AND2X1 mul_U16470(.A(n5458), .B(c0_act), .Y(n17928));
INVX1 mul_U16471(.A(n17928), .Y(n5382));
AND2X1 mul_U16472(.A(c0_act), .B(dpath_mulcore_booth_b13_in1[2]), .Y(n17930));
INVX1 mul_U16473(.A(n17930), .Y(n5383));
AND2X1 mul_U16474(.A(n5446), .B(c0_act), .Y(n17932));
INVX1 mul_U16475(.A(n17932), .Y(n5384));
AND2X1 mul_U16476(.A(n5456), .B(c0_act), .Y(n17934));
INVX1 mul_U16477(.A(n17934), .Y(n5385));
AND2X1 mul_U16478(.A(c0_act), .B(dpath_mulcore_booth_b14_in1[2]), .Y(n17936));
INVX1 mul_U16479(.A(n17936), .Y(n5386));
AND2X1 mul_U16480(.A(n5445), .B(c0_act), .Y(n17938));
INVX1 mul_U16481(.A(n17938), .Y(n5387));
AND2X1 mul_U16482(.A(n5454), .B(c0_act), .Y(n17940));
INVX1 mul_U16483(.A(n17940), .Y(n5388));
AND2X1 mul_U16484(.A(n5444), .B(c0_act), .Y(n17943));
INVX1 mul_U16485(.A(n17943), .Y(n5389));
AND2X1 mul_U16486(.A(n5451), .B(c0_act), .Y(n17945));
INVX1 mul_U16487(.A(n17945), .Y(n5390));
INVX1 mul_U16488(.A(dpath_mulcore_booth_b8_in0[1]), .Y(n5391));
INVX1 mul_U16489(.A(dpath_mulcore_booth_b15_in0[1]), .Y(n5392));
INVX1 mul_U16490(.A(dpath_mulcore_booth_b14_in0[1]), .Y(n5393));
INVX1 mul_U16491(.A(dpath_mulcore_booth_b13_in0[1]), .Y(n5394));
INVX1 mul_U16492(.A(dpath_mulcore_booth_b12_in0[1]), .Y(n5395));
INVX1 mul_U16493(.A(dpath_mulcore_booth_b11_in0[1]), .Y(n5396));
INVX1 mul_U16494(.A(dpath_mulcore_booth_b10_in0[1]), .Y(n5397));
AND2X1 mul_U16495(.A(n17975), .B(n17976), .Y(dpath_mulcore_booth_b9_in0[1]));
INVX1 mul_U16496(.A(dpath_mulcore_booth_b9_in0[1]), .Y(n5398));
INVX1 mul_U16497(.A(dpath_mulcore_booth_b15_in0[0]), .Y(n5399));
AND2X1 mul_U16498(.A(n5401), .B(dpath_mulcore_booth_b14_in0[2]), .Y(n17979));
INVX1 mul_U16499(.A(n17979), .Y(n5400));
OR2X1 mul_U16500(.A(dpath_mulcore_booth_b15_in0[2]), .B(n9806), .Y(n17982));
INVX1 mul_U16501(.A(n17982), .Y(n5401));
INVX1 mul_U16502(.A(dpath_mulcore_booth_b14_in0[0]), .Y(n5402));
AND2X1 mul_U16503(.A(n17986), .B(dpath_mulcore_booth_b13_in0[2]), .Y(n17983));
INVX1 mul_U16504(.A(n17983), .Y(n5403));
INVX1 mul_U16505(.A(dpath_mulcore_booth_b13_in0[0]), .Y(n5404));
AND2X1 mul_U16506(.A(n17990), .B(dpath_mulcore_booth_b12_in0[2]), .Y(n17987));
INVX1 mul_U16507(.A(n17987), .Y(n5405));
INVX1 mul_U16508(.A(dpath_mulcore_booth_b12_in0[0]), .Y(n5406));
AND2X1 mul_U16509(.A(n17994), .B(dpath_mulcore_booth_b11_in0[2]), .Y(n17991));
INVX1 mul_U16510(.A(n17991), .Y(n5407));
INVX1 mul_U16511(.A(dpath_mulcore_booth_b11_in0[0]), .Y(n5408));
AND2X1 mul_U16512(.A(n17998), .B(dpath_mulcore_booth_b10_in0[2]), .Y(n17995));
INVX1 mul_U16513(.A(n17995), .Y(n5409));
INVX1 mul_U16514(.A(dpath_mulcore_booth_b10_in0[0]), .Y(n5410));
AND2X1 mul_U16515(.A(n18002), .B(dpath_mulcore_booth_b9_in0[2]), .Y(n17999));
INVX1 mul_U16516(.A(n17999), .Y(n5411));
INVX1 mul_U16517(.A(dpath_mulcore_booth_b9_in0[0]), .Y(n5412));
OR2X1 mul_U16518(.A(dpath_mul_op2_d[18]), .B(dpath_mulcore_booth_b8_in0[2]), .Y(n18005));
INVX1 mul_U16519(.A(n18005), .Y(n5413));
AND2X1 mul_U16520(.A(n18006), .B(dpath_mul_op2_d[18]), .Y(n18003));
INVX1 mul_U16521(.A(n18003), .Y(n5414));
INVX1 mul_U16522(.A(dpath_mulcore_booth_b8_in0[0]), .Y(n5415));
AND2X1 mul_U16523(.A(n5417), .B(dpath_mulcore_booth_b8_in0[2]), .Y(n18007));
INVX1 mul_U16524(.A(n18007), .Y(n5416));
OR2X1 mul_U16525(.A(dpath_mulcore_booth_b7_in0[2]), .B(dpath_mul_op2_d[16]), .Y(n18010));
INVX1 mul_U16526(.A(n18010), .Y(n5417));
INVX1 mul_U16527(.A(dpath_mulcore_booth_b7_in1[1]), .Y(n5418));
INVX1 mul_U16528(.A(dpath_mulcore_booth_b6_in1[1]), .Y(n5419));
INVX1 mul_U16529(.A(dpath_mulcore_booth_b5_in1[1]), .Y(n5420));
INVX1 mul_U16530(.A(dpath_mulcore_booth_b4_in1[1]), .Y(n5421));
INVX1 mul_U16531(.A(dpath_mulcore_booth_b3_in1[1]), .Y(n5422));
INVX1 mul_U16532(.A(dpath_mulcore_booth_b2_in1[1]), .Y(n5423));
AND2X1 mul_U16533(.A(n18039), .B(n18040), .Y(dpath_mulcore_booth_b1_in1[1]));
INVX1 mul_U16534(.A(dpath_mulcore_booth_b1_in1[1]), .Y(n5424));
INVX1 mul_U16535(.A(dpath_mulcore_booth_b7_in1[0]), .Y(n5425));
AND2X1 mul_U16536(.A(n5427), .B(dpath_mulcore_booth_b6_in1[2]), .Y(n18043));
INVX1 mul_U16537(.A(n18043), .Y(n5426));
OR2X1 mul_U16538(.A(dpath_mulcore_booth_b7_in1[2]), .B(n10095), .Y(n18046));
INVX1 mul_U16539(.A(n18046), .Y(n5427));
INVX1 mul_U16540(.A(dpath_mulcore_booth_b6_in1[0]), .Y(n5428));
AND2X1 mul_U16541(.A(n18050), .B(dpath_mulcore_booth_b5_in1[2]), .Y(n18047));
INVX1 mul_U16542(.A(n18047), .Y(n5429));
INVX1 mul_U16543(.A(dpath_mulcore_booth_b5_in1[0]), .Y(n5430));
AND2X1 mul_U16544(.A(n18054), .B(dpath_mulcore_booth_b4_in1[2]), .Y(n18051));
INVX1 mul_U16545(.A(n18051), .Y(n5431));
INVX1 mul_U16546(.A(dpath_mulcore_booth_b4_in1[0]), .Y(n5432));
AND2X1 mul_U16547(.A(n18058), .B(dpath_mulcore_booth_b3_in1[2]), .Y(n18055));
INVX1 mul_U16548(.A(n18055), .Y(n5433));
INVX1 mul_U16549(.A(dpath_mulcore_booth_b3_in1[0]), .Y(n5434));
AND2X1 mul_U16550(.A(n18062), .B(dpath_mulcore_booth_b2_in1[2]), .Y(n18059));
INVX1 mul_U16551(.A(n18059), .Y(n5435));
INVX1 mul_U16552(.A(dpath_mulcore_booth_b2_in1[0]), .Y(n5436));
AND2X1 mul_U16553(.A(n18066), .B(dpath_mulcore_booth_b1_in1[2]), .Y(n18063));
INVX1 mul_U16554(.A(n18063), .Y(n5437));
INVX1 mul_U16555(.A(dpath_mulcore_booth_b1_in1[0]), .Y(n5438));
OR2X1 mul_U16556(.A(dpath_mulcore_booth_b[34]), .B(dpath_mulcore_booth_b0_in1[2]), .Y(n18069));
INVX1 mul_U16557(.A(n18069), .Y(n5439));
AND2X1 mul_U16558(.A(n18070), .B(dpath_mulcore_booth_b[34]), .Y(n18067));
INVX1 mul_U16559(.A(n18067), .Y(n5440));
AND2X1 mul_U16560(.A(n5442), .B(dpath_mulcore_booth_b0_in1[2]), .Y(n18071));
INVX1 mul_U16561(.A(n18071), .Y(n5441));
OR2X1 mul_U16562(.A(dpath_mulcore_booth_b[31]), .B(dpath_mulcore_booth_b[32]), .Y(n18074));
INVX1 mul_U16563(.A(n18074), .Y(n5442));
INVX1 mul_U16564(.A(dpath_mulcore_booth_b8_in1[1]), .Y(n5443));
INVX1 mul_U16565(.A(dpath_mulcore_booth_b15_in1[1]), .Y(n5444));
INVX1 mul_U16566(.A(dpath_mulcore_booth_b14_in1[1]), .Y(n5445));
INVX1 mul_U16567(.A(dpath_mulcore_booth_b13_in1[1]), .Y(n5446));
INVX1 mul_U16568(.A(dpath_mulcore_booth_b12_in1[1]), .Y(n5447));
INVX1 mul_U16569(.A(dpath_mulcore_booth_b11_in1[1]), .Y(n5448));
INVX1 mul_U16570(.A(dpath_mulcore_booth_b10_in1[1]), .Y(n5449));
AND2X1 mul_U16571(.A(n18103), .B(n18104), .Y(dpath_mulcore_booth_b9_in1[1]));
INVX1 mul_U16572(.A(dpath_mulcore_booth_b9_in1[1]), .Y(n5450));
INVX1 mul_U16573(.A(dpath_mulcore_booth_b15_in1[0]), .Y(n5451));
AND2X1 mul_U16574(.A(n5453), .B(dpath_mulcore_booth_b14_in1[2]), .Y(n18107));
INVX1 mul_U16575(.A(n18107), .Y(n5452));
OR2X1 mul_U16576(.A(dpath_mulcore_booth_b15_in1[2]), .B(n10109), .Y(n18110));
INVX1 mul_U16577(.A(n18110), .Y(n5453));
INVX1 mul_U16578(.A(dpath_mulcore_booth_b14_in1[0]), .Y(n5454));
AND2X1 mul_U16579(.A(n18114), .B(dpath_mulcore_booth_b13_in1[2]), .Y(n18111));
INVX1 mul_U16580(.A(n18111), .Y(n5455));
INVX1 mul_U16581(.A(dpath_mulcore_booth_b13_in1[0]), .Y(n5456));
AND2X1 mul_U16582(.A(n18118), .B(dpath_mulcore_booth_b12_in1[2]), .Y(n18115));
INVX1 mul_U16583(.A(n18115), .Y(n5457));
INVX1 mul_U16584(.A(dpath_mulcore_booth_b12_in1[0]), .Y(n5458));
AND2X1 mul_U16585(.A(n18122), .B(dpath_mulcore_booth_b11_in1[2]), .Y(n18119));
INVX1 mul_U16586(.A(n18119), .Y(n5459));
INVX1 mul_U16587(.A(dpath_mulcore_booth_b11_in1[0]), .Y(n5460));
AND2X1 mul_U16588(.A(n18126), .B(dpath_mulcore_booth_b10_in1[2]), .Y(n18123));
INVX1 mul_U16589(.A(n18123), .Y(n5461));
INVX1 mul_U16590(.A(dpath_mulcore_booth_b10_in1[0]), .Y(n5462));
AND2X1 mul_U16591(.A(n18130), .B(dpath_mulcore_booth_b9_in1[2]), .Y(n18127));
INVX1 mul_U16592(.A(n18127), .Y(n5463));
INVX1 mul_U16593(.A(dpath_mulcore_booth_b9_in1[0]), .Y(n5464));
OR2X1 mul_U16594(.A(dpath_mulcore_booth_b[50]), .B(dpath_mulcore_booth_b8_in1[2]), .Y(n18133));
INVX1 mul_U16595(.A(n18133), .Y(n5465));
AND2X1 mul_U16596(.A(n18134), .B(dpath_mulcore_booth_b[50]), .Y(n18131));
INVX1 mul_U16597(.A(n18131), .Y(n5466));
INVX1 mul_U16598(.A(dpath_mulcore_booth_b8_in1[0]), .Y(n5467));
AND2X1 mul_U16599(.A(n5469), .B(dpath_mulcore_booth_b8_in1[2]), .Y(n18135));
INVX1 mul_U16600(.A(n18135), .Y(n5468));
OR2X1 mul_U16601(.A(dpath_mulcore_booth_b7_in1[2]), .B(dpath_mulcore_booth_b[48]), .Y(n18138));
INVX1 mul_U16602(.A(n18138), .Y(n5469));
AND2X1 mul_U16603(.A(dpath_mulcore_ary1_a0_sc3_71__z), .B(n7227), .Y(dpath_mulcore_ary1_a0_sc3_71__n5));
INVX1 mul_U16604(.A(dpath_mulcore_ary1_a0_sc3_71__n5), .Y(n5470));
AND2X1 mul_U16605(.A(c0_act), .B(dpath_mulcore_booth_b0_in1[2]), .Y(dpath_mulcore_booth_out_mux0_n2));
INVX1 mul_U16606(.A(dpath_mulcore_booth_out_mux0_n2), .Y(n5471));
INVX1 mul_U16607(.A(dpath_mulcore_booth_out_mux0_n4), .Y(n5472));
INVX1 mul_U16608(.A(dpath_mulcore_booth_out_mux0_n6), .Y(n5473));
AND2X1 mul_U16609(.A(dpath_mulcore_booth_encode0_a_n17), .B(n9786), .Y(dpath_mulcore_booth_b0_in0[1]));
INVX1 mul_U16610(.A(dpath_mulcore_booth_b0_in0[1]), .Y(n5474));
INVX1 mul_U16611(.A(dpath_mulcore_booth_b7_in0[1]), .Y(n5475));
INVX1 mul_U16612(.A(dpath_mulcore_booth_b6_in0[1]), .Y(n5476));
INVX1 mul_U16613(.A(dpath_mulcore_booth_b5_in0[1]), .Y(n5477));
INVX1 mul_U16614(.A(dpath_mulcore_booth_b4_in0[1]), .Y(n5478));
INVX1 mul_U16615(.A(dpath_mulcore_booth_b3_in0[1]), .Y(n5479));
INVX1 mul_U16616(.A(dpath_mulcore_booth_b2_in0[1]), .Y(n5480));
AND2X1 mul_U16617(.A(dpath_mulcore_booth_encode0_a_n43), .B(dpath_mulcore_booth_encode0_a_n44), .Y(dpath_mulcore_booth_b1_in0[1]));
INVX1 mul_U16618(.A(dpath_mulcore_booth_b1_in0[1]), .Y(n5481));
INVX1 mul_U16619(.A(dpath_mulcore_booth_b7_in0[0]), .Y(n5482));
AND2X1 mul_U16620(.A(n5484), .B(dpath_mulcore_booth_b6_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n47));
INVX1 mul_U16621(.A(dpath_mulcore_booth_encode0_a_n47), .Y(n5483));
OR2X1 mul_U16622(.A(dpath_mulcore_booth_b7_in0[2]), .B(n9791), .Y(dpath_mulcore_booth_encode0_a_n50));
INVX1 mul_U16623(.A(dpath_mulcore_booth_encode0_a_n50), .Y(n5484));
INVX1 mul_U16624(.A(dpath_mulcore_booth_b6_in0[0]), .Y(n5485));
AND2X1 mul_U16625(.A(dpath_mulcore_booth_encode0_a_n54), .B(dpath_mulcore_booth_b5_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n51));
INVX1 mul_U16626(.A(dpath_mulcore_booth_encode0_a_n51), .Y(n5486));
INVX1 mul_U16627(.A(dpath_mulcore_booth_b5_in0[0]), .Y(n5487));
AND2X1 mul_U16628(.A(dpath_mulcore_booth_encode0_a_n58), .B(dpath_mulcore_booth_b4_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n55));
INVX1 mul_U16629(.A(dpath_mulcore_booth_encode0_a_n55), .Y(n5488));
INVX1 mul_U16630(.A(dpath_mulcore_booth_b4_in0[0]), .Y(n5489));
AND2X1 mul_U16631(.A(dpath_mulcore_booth_encode0_a_n62), .B(dpath_mulcore_booth_b3_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n59));
INVX1 mul_U16632(.A(dpath_mulcore_booth_encode0_a_n59), .Y(n5490));
INVX1 mul_U16633(.A(dpath_mulcore_booth_b3_in0[0]), .Y(n5491));
AND2X1 mul_U16634(.A(dpath_mulcore_booth_encode0_a_n66), .B(dpath_mulcore_booth_b2_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n63));
INVX1 mul_U16635(.A(dpath_mulcore_booth_encode0_a_n63), .Y(n5492));
INVX1 mul_U16636(.A(dpath_mulcore_booth_b2_in0[0]), .Y(n5493));
AND2X1 mul_U16637(.A(dpath_mulcore_booth_encode0_a_n70), .B(dpath_mulcore_booth_b1_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n67));
INVX1 mul_U16638(.A(dpath_mulcore_booth_encode0_a_n67), .Y(n5494));
INVX1 mul_U16639(.A(dpath_mulcore_booth_b1_in0[0]), .Y(n5495));
OR2X1 mul_U16640(.A(dpath_mul_op2_d[2]), .B(dpath_mulcore_booth_b0_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n73));
INVX1 mul_U16641(.A(dpath_mulcore_booth_encode0_a_n73), .Y(n5496));
AND2X1 mul_U16642(.A(dpath_mulcore_booth_encode0_a_n74), .B(dpath_mul_op2_d[2]), .Y(dpath_mulcore_booth_encode0_a_n71));
INVX1 mul_U16643(.A(dpath_mulcore_booth_encode0_a_n71), .Y(n5497));
AND2X1 mul_U16644(.A(n9683), .B(dpath_mulcore_psum[8]), .Y(dpath_mulcore_ary2_smux_n2));
INVX1 mul_U16645(.A(dpath_mulcore_ary2_smux_n2), .Y(n5498));
AND2X1 mul_U16646(.A(dpath_mulcore_psum[96]), .B(n9691), .Y(dpath_mulcore_ary2_smux_n4));
INVX1 mul_U16647(.A(dpath_mulcore_ary2_smux_n4), .Y(n5499));
AND2X1 mul_U16648(.A(dpath_mulcore_psum[95]), .B(n9691), .Y(dpath_mulcore_ary2_smux_n6));
INVX1 mul_U16649(.A(dpath_mulcore_ary2_smux_n6), .Y(n5500));
AND2X1 mul_U16650(.A(dpath_mulcore_psum[94]), .B(n9691), .Y(dpath_mulcore_ary2_smux_n8));
INVX1 mul_U16651(.A(dpath_mulcore_ary2_smux_n8), .Y(n5501));
AND2X1 mul_U16652(.A(dpath_mulcore_psum[93]), .B(n9691), .Y(dpath_mulcore_ary2_smux_n10));
INVX1 mul_U16653(.A(dpath_mulcore_ary2_smux_n10), .Y(n5502));
AND2X1 mul_U16654(.A(dpath_mulcore_psum[92]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n12));
INVX1 mul_U16655(.A(dpath_mulcore_ary2_smux_n12), .Y(n5503));
AND2X1 mul_U16656(.A(dpath_mulcore_psum[91]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n14));
INVX1 mul_U16657(.A(dpath_mulcore_ary2_smux_n14), .Y(n5504));
AND2X1 mul_U16658(.A(dpath_mulcore_psum[90]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n16));
INVX1 mul_U16659(.A(dpath_mulcore_ary2_smux_n16), .Y(n5505));
AND2X1 mul_U16660(.A(dpath_mulcore_psum[89]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n18));
INVX1 mul_U16661(.A(dpath_mulcore_ary2_smux_n18), .Y(n5506));
AND2X1 mul_U16662(.A(dpath_mulcore_psum[7]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n20));
INVX1 mul_U16663(.A(dpath_mulcore_ary2_smux_n20), .Y(n5507));
AND2X1 mul_U16664(.A(dpath_mulcore_psum[88]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n22));
INVX1 mul_U16665(.A(dpath_mulcore_ary2_smux_n22), .Y(n5508));
AND2X1 mul_U16666(.A(dpath_mulcore_psum[87]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n24));
INVX1 mul_U16667(.A(dpath_mulcore_ary2_smux_n24), .Y(n5509));
AND2X1 mul_U16668(.A(dpath_mulcore_psum[86]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n26));
INVX1 mul_U16669(.A(dpath_mulcore_ary2_smux_n26), .Y(n5510));
AND2X1 mul_U16670(.A(dpath_mulcore_psum[85]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n28));
INVX1 mul_U16671(.A(dpath_mulcore_ary2_smux_n28), .Y(n5511));
AND2X1 mul_U16672(.A(dpath_mulcore_psum[84]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n30));
INVX1 mul_U16673(.A(dpath_mulcore_ary2_smux_n30), .Y(n5512));
AND2X1 mul_U16674(.A(dpath_mulcore_psum[83]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n32));
INVX1 mul_U16675(.A(dpath_mulcore_ary2_smux_n32), .Y(n5513));
AND2X1 mul_U16676(.A(dpath_mulcore_psum[82]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n34));
INVX1 mul_U16677(.A(dpath_mulcore_ary2_smux_n34), .Y(n5514));
AND2X1 mul_U16678(.A(dpath_mulcore_psum[81]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n36));
INVX1 mul_U16679(.A(dpath_mulcore_ary2_smux_n36), .Y(n5515));
AND2X1 mul_U16680(.A(dpath_mulcore_psum[80]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n38));
INVX1 mul_U16681(.A(dpath_mulcore_ary2_smux_n38), .Y(n5516));
AND2X1 mul_U16682(.A(dpath_mulcore_psum[79]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n40));
INVX1 mul_U16683(.A(dpath_mulcore_ary2_smux_n40), .Y(n5517));
AND2X1 mul_U16684(.A(dpath_mulcore_psum[6]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n42));
INVX1 mul_U16685(.A(dpath_mulcore_ary2_smux_n42), .Y(n5518));
AND2X1 mul_U16686(.A(dpath_mulcore_psum[78]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n44));
INVX1 mul_U16687(.A(dpath_mulcore_ary2_smux_n44), .Y(n5519));
AND2X1 mul_U16688(.A(dpath_mulcore_psum[77]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n46));
INVX1 mul_U16689(.A(dpath_mulcore_ary2_smux_n46), .Y(n5520));
AND2X1 mul_U16690(.A(dpath_mulcore_psum[76]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n48));
INVX1 mul_U16691(.A(dpath_mulcore_ary2_smux_n48), .Y(n5521));
AND2X1 mul_U16692(.A(dpath_mulcore_psum[75]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n50));
INVX1 mul_U16693(.A(dpath_mulcore_ary2_smux_n50), .Y(n5522));
AND2X1 mul_U16694(.A(dpath_mulcore_psum[74]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n52));
INVX1 mul_U16695(.A(dpath_mulcore_ary2_smux_n52), .Y(n5523));
AND2X1 mul_U16696(.A(dpath_mulcore_psum[73]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n54));
INVX1 mul_U16697(.A(dpath_mulcore_ary2_smux_n54), .Y(n5524));
AND2X1 mul_U16698(.A(dpath_mulcore_psum[72]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n56));
INVX1 mul_U16699(.A(dpath_mulcore_ary2_smux_n56), .Y(n5525));
AND2X1 mul_U16700(.A(dpath_mulcore_psum[71]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n58));
INVX1 mul_U16701(.A(dpath_mulcore_ary2_smux_n58), .Y(n5526));
AND2X1 mul_U16702(.A(dpath_mulcore_psum[70]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n60));
INVX1 mul_U16703(.A(dpath_mulcore_ary2_smux_n60), .Y(n5527));
AND2X1 mul_U16704(.A(dpath_mulcore_psum[69]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n62));
INVX1 mul_U16705(.A(dpath_mulcore_ary2_smux_n62), .Y(n5528));
AND2X1 mul_U16706(.A(dpath_mulcore_psum[5]), .B(n9686), .Y(dpath_mulcore_ary2_smux_n64));
INVX1 mul_U16707(.A(dpath_mulcore_ary2_smux_n64), .Y(n5529));
AND2X1 mul_U16708(.A(dpath_mulcore_psum[68]), .B(n9674), .Y(dpath_mulcore_ary2_smux_n66));
INVX1 mul_U16709(.A(dpath_mulcore_ary2_smux_n66), .Y(n5530));
AND2X1 mul_U16710(.A(dpath_mulcore_psum[67]), .B(n9676), .Y(dpath_mulcore_ary2_smux_n68));
INVX1 mul_U16711(.A(dpath_mulcore_ary2_smux_n68), .Y(n5531));
AND2X1 mul_U16712(.A(dpath_mulcore_psum[66]), .B(n9677), .Y(dpath_mulcore_ary2_smux_n70));
INVX1 mul_U16713(.A(dpath_mulcore_ary2_smux_n70), .Y(n5532));
AND2X1 mul_U16714(.A(dpath_mulcore_psum[65]), .B(n9690), .Y(dpath_mulcore_ary2_smux_n72));
INVX1 mul_U16715(.A(dpath_mulcore_ary2_smux_n72), .Y(n5533));
AND2X1 mul_U16716(.A(dpath_mulcore_psum[64]), .B(n9689), .Y(dpath_mulcore_ary2_smux_n74));
INVX1 mul_U16717(.A(dpath_mulcore_ary2_smux_n74), .Y(n5534));
AND2X1 mul_U16718(.A(dpath_mulcore_psum[63]), .B(n9687), .Y(dpath_mulcore_ary2_smux_n76));
INVX1 mul_U16719(.A(dpath_mulcore_ary2_smux_n76), .Y(n5535));
AND2X1 mul_U16720(.A(dpath_mulcore_psum[62]), .B(n9688), .Y(dpath_mulcore_ary2_smux_n78));
INVX1 mul_U16721(.A(dpath_mulcore_ary2_smux_n78), .Y(n5536));
AND2X1 mul_U16722(.A(dpath_mulcore_psum[61]), .B(n9692), .Y(dpath_mulcore_ary2_smux_n80));
INVX1 mul_U16723(.A(dpath_mulcore_ary2_smux_n80), .Y(n5537));
AND2X1 mul_U16724(.A(dpath_mulcore_psum[60]), .B(n9691), .Y(dpath_mulcore_ary2_smux_n82));
INVX1 mul_U16725(.A(dpath_mulcore_ary2_smux_n82), .Y(n5538));
AND2X1 mul_U16726(.A(dpath_mulcore_psum[59]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n84));
INVX1 mul_U16727(.A(dpath_mulcore_ary2_smux_n84), .Y(n5539));
AND2X1 mul_U16728(.A(dpath_mulcore_psum[4]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n86));
INVX1 mul_U16729(.A(dpath_mulcore_ary2_smux_n86), .Y(n5540));
AND2X1 mul_U16730(.A(dpath_mulcore_psum[58]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n88));
INVX1 mul_U16731(.A(dpath_mulcore_ary2_smux_n88), .Y(n5541));
AND2X1 mul_U16732(.A(dpath_mulcore_psum[57]), .B(n9691), .Y(dpath_mulcore_ary2_smux_n90));
INVX1 mul_U16733(.A(dpath_mulcore_ary2_smux_n90), .Y(n5542));
AND2X1 mul_U16734(.A(dpath_mulcore_psum[56]), .B(n9693), .Y(dpath_mulcore_ary2_smux_n92));
INVX1 mul_U16735(.A(dpath_mulcore_ary2_smux_n92), .Y(n5543));
AND2X1 mul_U16736(.A(dpath_mulcore_psum[55]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n94));
INVX1 mul_U16737(.A(dpath_mulcore_ary2_smux_n94), .Y(n5544));
AND2X1 mul_U16738(.A(dpath_mulcore_psum[54]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n96));
INVX1 mul_U16739(.A(dpath_mulcore_ary2_smux_n96), .Y(n5545));
AND2X1 mul_U16740(.A(dpath_mulcore_psum[53]), .B(n9673), .Y(dpath_mulcore_ary2_smux_n98));
INVX1 mul_U16741(.A(dpath_mulcore_ary2_smux_n98), .Y(n5546));
AND2X1 mul_U16742(.A(dpath_mulcore_psum[52]), .B(n9675), .Y(dpath_mulcore_ary2_smux_n100));
INVX1 mul_U16743(.A(dpath_mulcore_ary2_smux_n100), .Y(n5547));
AND2X1 mul_U16744(.A(dpath_mulcore_psum[51]), .B(n9678), .Y(dpath_mulcore_ary2_smux_n102));
INVX1 mul_U16745(.A(dpath_mulcore_ary2_smux_n102), .Y(n5548));
AND2X1 mul_U16746(.A(dpath_mulcore_psum[50]), .B(n9679), .Y(dpath_mulcore_ary2_smux_n104));
INVX1 mul_U16747(.A(dpath_mulcore_ary2_smux_n104), .Y(n5549));
AND2X1 mul_U16748(.A(dpath_mulcore_psum[49]), .B(n9684), .Y(dpath_mulcore_ary2_smux_n106));
INVX1 mul_U16749(.A(dpath_mulcore_ary2_smux_n106), .Y(n5550));
AND2X1 mul_U16750(.A(dpath_mulcore_psum[3]), .B(n9683), .Y(dpath_mulcore_ary2_smux_n108));
INVX1 mul_U16751(.A(dpath_mulcore_ary2_smux_n108), .Y(n5551));
AND2X1 mul_U16752(.A(dpath_mulcore_psum[48]), .B(n9685), .Y(dpath_mulcore_ary2_smux_n110));
INVX1 mul_U16753(.A(dpath_mulcore_ary2_smux_n110), .Y(n5552));
AND2X1 mul_U16754(.A(dpath_mulcore_psum[47]), .B(n9671), .Y(dpath_mulcore_ary2_smux_n112));
INVX1 mul_U16755(.A(dpath_mulcore_ary2_smux_n112), .Y(n5553));
AND2X1 mul_U16756(.A(dpath_mulcore_psum[46]), .B(n9672), .Y(dpath_mulcore_ary2_smux_n114));
INVX1 mul_U16757(.A(dpath_mulcore_ary2_smux_n114), .Y(n5554));
AND2X1 mul_U16758(.A(dpath_mulcore_psum[45]), .B(dpath_mulcore_x2_c2c3), .Y(dpath_mulcore_ary2_smux_n116));
INVX1 mul_U16759(.A(dpath_mulcore_ary2_smux_n116), .Y(n5555));
AND2X1 mul_U16760(.A(dpath_mulcore_psum[44]), .B(dpath_mulcore_x2_c2c3), .Y(dpath_mulcore_ary2_smux_n118));
INVX1 mul_U16761(.A(dpath_mulcore_ary2_smux_n118), .Y(n5556));
AND2X1 mul_U16762(.A(dpath_mulcore_psum[43]), .B(dpath_mulcore_x2_c2c3), .Y(dpath_mulcore_ary2_smux_n120));
INVX1 mul_U16763(.A(dpath_mulcore_ary2_smux_n120), .Y(n5557));
AND2X1 mul_U16764(.A(dpath_mulcore_psum[42]), .B(n9671), .Y(dpath_mulcore_ary2_smux_n122));
INVX1 mul_U16765(.A(dpath_mulcore_ary2_smux_n122), .Y(n5558));
AND2X1 mul_U16766(.A(dpath_mulcore_psum[41]), .B(n9675), .Y(dpath_mulcore_ary2_smux_n124));
INVX1 mul_U16767(.A(dpath_mulcore_ary2_smux_n124), .Y(n5559));
AND2X1 mul_U16768(.A(dpath_mulcore_psum[40]), .B(n9678), .Y(dpath_mulcore_ary2_smux_n126));
INVX1 mul_U16769(.A(dpath_mulcore_ary2_smux_n126), .Y(n5560));
AND2X1 mul_U16770(.A(dpath_mulcore_psum[39]), .B(n9679), .Y(dpath_mulcore_ary2_smux_n128));
INVX1 mul_U16771(.A(dpath_mulcore_ary2_smux_n128), .Y(n5561));
AND2X1 mul_U16772(.A(dpath_mulcore_psum[2]), .B(n9672), .Y(dpath_mulcore_ary2_smux_n130));
INVX1 mul_U16773(.A(dpath_mulcore_ary2_smux_n130), .Y(n5562));
AND2X1 mul_U16774(.A(dpath_mulcore_psum[38]), .B(dpath_mulcore_x2_c2c3), .Y(dpath_mulcore_ary2_smux_n132));
INVX1 mul_U16775(.A(dpath_mulcore_ary2_smux_n132), .Y(n5563));
AND2X1 mul_U16776(.A(dpath_mulcore_psum[37]), .B(n9671), .Y(dpath_mulcore_ary2_smux_n134));
INVX1 mul_U16777(.A(dpath_mulcore_ary2_smux_n134), .Y(n5564));
AND2X1 mul_U16778(.A(dpath_mulcore_psum[36]), .B(n9675), .Y(dpath_mulcore_ary2_smux_n136));
INVX1 mul_U16779(.A(dpath_mulcore_ary2_smux_n136), .Y(n5565));
AND2X1 mul_U16780(.A(dpath_mulcore_psum[35]), .B(n9678), .Y(dpath_mulcore_ary2_smux_n138));
INVX1 mul_U16781(.A(dpath_mulcore_ary2_smux_n138), .Y(n5566));
AND2X1 mul_U16782(.A(dpath_mulcore_psum[34]), .B(n9679), .Y(dpath_mulcore_ary2_smux_n140));
INVX1 mul_U16783(.A(dpath_mulcore_ary2_smux_n140), .Y(n5567));
AND2X1 mul_U16784(.A(dpath_mulcore_psum[33]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n142));
INVX1 mul_U16785(.A(dpath_mulcore_ary2_smux_n142), .Y(n5568));
AND2X1 mul_U16786(.A(dpath_mulcore_psum[32]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n144));
INVX1 mul_U16787(.A(dpath_mulcore_ary2_smux_n144), .Y(n5569));
AND2X1 mul_U16788(.A(dpath_mulcore_psum[31]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n146));
INVX1 mul_U16789(.A(dpath_mulcore_ary2_smux_n146), .Y(n5570));
AND2X1 mul_U16790(.A(dpath_mulcore_psum[30]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n148));
INVX1 mul_U16791(.A(dpath_mulcore_ary2_smux_n148), .Y(n5571));
AND2X1 mul_U16792(.A(dpath_mulcore_psum[29]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n150));
INVX1 mul_U16793(.A(dpath_mulcore_ary2_smux_n150), .Y(n5572));
AND2X1 mul_U16794(.A(dpath_mulcore_psum[1]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n152));
INVX1 mul_U16795(.A(dpath_mulcore_ary2_smux_n152), .Y(n5573));
AND2X1 mul_U16796(.A(dpath_mulcore_psum[28]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n154));
INVX1 mul_U16797(.A(dpath_mulcore_ary2_smux_n154), .Y(n5574));
AND2X1 mul_U16798(.A(dpath_mulcore_psum[27]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n156));
INVX1 mul_U16799(.A(dpath_mulcore_ary2_smux_n156), .Y(n5575));
AND2X1 mul_U16800(.A(dpath_mulcore_psum[26]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n158));
INVX1 mul_U16801(.A(dpath_mulcore_ary2_smux_n158), .Y(n5576));
AND2X1 mul_U16802(.A(dpath_mulcore_psum[25]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n160));
INVX1 mul_U16803(.A(dpath_mulcore_ary2_smux_n160), .Y(n5577));
AND2X1 mul_U16804(.A(dpath_mulcore_psum[24]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n162));
INVX1 mul_U16805(.A(dpath_mulcore_ary2_smux_n162), .Y(n5578));
AND2X1 mul_U16806(.A(dpath_mulcore_psum[23]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n164));
INVX1 mul_U16807(.A(dpath_mulcore_ary2_smux_n164), .Y(n5579));
AND2X1 mul_U16808(.A(dpath_mulcore_psum[22]), .B(n9694), .Y(dpath_mulcore_ary2_smux_n166));
INVX1 mul_U16809(.A(dpath_mulcore_ary2_smux_n166), .Y(n5580));
AND2X1 mul_U16810(.A(dpath_mulcore_psum[21]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n168));
INVX1 mul_U16811(.A(dpath_mulcore_ary2_smux_n168), .Y(n5581));
AND2X1 mul_U16812(.A(dpath_mulcore_psum[20]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n170));
INVX1 mul_U16813(.A(dpath_mulcore_ary2_smux_n170), .Y(n5582));
AND2X1 mul_U16814(.A(dpath_mulcore_psum[19]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n172));
INVX1 mul_U16815(.A(dpath_mulcore_ary2_smux_n172), .Y(n5583));
AND2X1 mul_U16816(.A(dpath_mulcore_psum[0]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n174));
INVX1 mul_U16817(.A(dpath_mulcore_ary2_smux_n174), .Y(n5584));
AND2X1 mul_U16818(.A(dpath_mulcore_psum[18]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n176));
INVX1 mul_U16819(.A(dpath_mulcore_ary2_smux_n176), .Y(n5585));
AND2X1 mul_U16820(.A(dpath_mulcore_psum[17]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n178));
INVX1 mul_U16821(.A(dpath_mulcore_ary2_smux_n178), .Y(n5586));
AND2X1 mul_U16822(.A(dpath_mulcore_psum[16]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n180));
INVX1 mul_U16823(.A(dpath_mulcore_ary2_smux_n180), .Y(n5587));
AND2X1 mul_U16824(.A(n16562), .B(n9695), .Y(dpath_mulcore_ary2_smux_n182));
INVX1 mul_U16825(.A(dpath_mulcore_ary2_smux_n182), .Y(n5588));
AND2X1 mul_U16826(.A(dpath_mulcore_psum[14]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n184));
INVX1 mul_U16827(.A(dpath_mulcore_ary2_smux_n184), .Y(n5589));
AND2X1 mul_U16828(.A(dpath_mulcore_psum[13]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n186));
INVX1 mul_U16829(.A(dpath_mulcore_ary2_smux_n186), .Y(n5590));
AND2X1 mul_U16830(.A(dpath_mulcore_psum[12]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n188));
INVX1 mul_U16831(.A(dpath_mulcore_ary2_smux_n188), .Y(n5591));
AND2X1 mul_U16832(.A(dpath_mulcore_psum[11]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n190));
INVX1 mul_U16833(.A(dpath_mulcore_ary2_smux_n190), .Y(n5592));
AND2X1 mul_U16834(.A(dpath_mulcore_psum[10]), .B(n9695), .Y(dpath_mulcore_ary2_smux_n192));
INVX1 mul_U16835(.A(dpath_mulcore_ary2_smux_n192), .Y(n5593));
AND2X1 mul_U16836(.A(dpath_mulcore_psum[9]), .B(n9685), .Y(dpath_mulcore_ary2_smux_n194));
INVX1 mul_U16837(.A(dpath_mulcore_ary2_smux_n194), .Y(n5594));
AND2X1 mul_U16838(.A(dpath_mulcore_psumx2), .B(n9686), .Y(dpath_mulcore_ary2_smux_n196));
INVX1 mul_U16839(.A(dpath_mulcore_ary2_smux_n196), .Y(n5595));
AND2X1 mul_U16840(.A(n9683), .B(n6074), .Y(dpath_mulcore_ary2_cmux_n2));
INVX1 mul_U16841(.A(dpath_mulcore_ary2_cmux_n2), .Y(n5596));
AND2X1 mul_U16842(.A(n9188), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n4));
INVX1 mul_U16843(.A(dpath_mulcore_ary2_cmux_n4), .Y(n5597));
AND2X1 mul_U16844(.A(n9189), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n6));
INVX1 mul_U16845(.A(dpath_mulcore_ary2_cmux_n6), .Y(n5598));
AND2X1 mul_U16846(.A(n9190), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n8));
INVX1 mul_U16847(.A(dpath_mulcore_ary2_cmux_n8), .Y(n5599));
AND2X1 mul_U16848(.A(n9191), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n10));
INVX1 mul_U16849(.A(dpath_mulcore_ary2_cmux_n10), .Y(n5600));
AND2X1 mul_U16850(.A(n9192), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n12));
INVX1 mul_U16851(.A(dpath_mulcore_ary2_cmux_n12), .Y(n5601));
AND2X1 mul_U16852(.A(n9193), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n14));
INVX1 mul_U16853(.A(dpath_mulcore_ary2_cmux_n14), .Y(n5602));
AND2X1 mul_U16854(.A(n9194), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n16));
INVX1 mul_U16855(.A(dpath_mulcore_ary2_cmux_n16), .Y(n5603));
AND2X1 mul_U16856(.A(n6161), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n18));
INVX1 mul_U16857(.A(dpath_mulcore_ary2_cmux_n18), .Y(n5604));
AND2X1 mul_U16858(.A(n9195), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n20));
INVX1 mul_U16859(.A(dpath_mulcore_ary2_cmux_n20), .Y(n5605));
AND2X1 mul_U16860(.A(n9196), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n22));
INVX1 mul_U16861(.A(dpath_mulcore_ary2_cmux_n22), .Y(n5606));
AND2X1 mul_U16862(.A(n9197), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n24));
INVX1 mul_U16863(.A(dpath_mulcore_ary2_cmux_n24), .Y(n5607));
AND2X1 mul_U16864(.A(n9198), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n26));
INVX1 mul_U16865(.A(dpath_mulcore_ary2_cmux_n26), .Y(n5608));
AND2X1 mul_U16866(.A(n9199), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n28));
INVX1 mul_U16867(.A(dpath_mulcore_ary2_cmux_n28), .Y(n5609));
AND2X1 mul_U16868(.A(n9213), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n30));
INVX1 mul_U16869(.A(dpath_mulcore_ary2_cmux_n30), .Y(n5610));
AND2X1 mul_U16870(.A(n9148), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n32));
INVX1 mul_U16871(.A(dpath_mulcore_ary2_cmux_n32), .Y(n5611));
AND2X1 mul_U16872(.A(n9200), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n34));
INVX1 mul_U16873(.A(dpath_mulcore_ary2_cmux_n34), .Y(n5612));
AND2X1 mul_U16874(.A(n9201), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n36));
INVX1 mul_U16875(.A(dpath_mulcore_ary2_cmux_n36), .Y(n5613));
AND2X1 mul_U16876(.A(n9202), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n38));
INVX1 mul_U16877(.A(dpath_mulcore_ary2_cmux_n38), .Y(n5614));
AND2X1 mul_U16878(.A(n6162), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n40));
INVX1 mul_U16879(.A(dpath_mulcore_ary2_cmux_n40), .Y(n5615));
AND2X1 mul_U16880(.A(n9203), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n42));
INVX1 mul_U16881(.A(dpath_mulcore_ary2_cmux_n42), .Y(n5616));
AND2X1 mul_U16882(.A(n9204), .B(n9690), .Y(dpath_mulcore_ary2_cmux_n44));
INVX1 mul_U16883(.A(dpath_mulcore_ary2_cmux_n44), .Y(n5617));
AND2X1 mul_U16884(.A(n9205), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n46));
INVX1 mul_U16885(.A(dpath_mulcore_ary2_cmux_n46), .Y(n5618));
AND2X1 mul_U16886(.A(n9206), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n48));
INVX1 mul_U16887(.A(dpath_mulcore_ary2_cmux_n48), .Y(n5619));
AND2X1 mul_U16888(.A(n9207), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n50));
INVX1 mul_U16889(.A(dpath_mulcore_ary2_cmux_n50), .Y(n5620));
AND2X1 mul_U16890(.A(n9208), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n52));
INVX1 mul_U16891(.A(dpath_mulcore_ary2_cmux_n52), .Y(n5621));
AND2X1 mul_U16892(.A(n9209), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n54));
INVX1 mul_U16893(.A(dpath_mulcore_ary2_cmux_n54), .Y(n5622));
AND2X1 mul_U16894(.A(n9210), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n56));
INVX1 mul_U16895(.A(dpath_mulcore_ary2_cmux_n56), .Y(n5623));
AND2X1 mul_U16896(.A(n9211), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n58));
INVX1 mul_U16897(.A(dpath_mulcore_ary2_cmux_n58), .Y(n5624));
AND2X1 mul_U16898(.A(n9212), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n60));
INVX1 mul_U16899(.A(dpath_mulcore_ary2_cmux_n60), .Y(n5625));
AND2X1 mul_U16900(.A(n6163), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n62));
INVX1 mul_U16901(.A(dpath_mulcore_ary2_cmux_n62), .Y(n5626));
AND2X1 mul_U16902(.A(n9149), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n64));
INVX1 mul_U16903(.A(dpath_mulcore_ary2_cmux_n64), .Y(n5627));
AND2X1 mul_U16904(.A(n9150), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n66));
INVX1 mul_U16905(.A(dpath_mulcore_ary2_cmux_n66), .Y(n5628));
AND2X1 mul_U16906(.A(n9151), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n68));
INVX1 mul_U16907(.A(dpath_mulcore_ary2_cmux_n68), .Y(n5629));
AND2X1 mul_U16908(.A(n9152), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n70));
INVX1 mul_U16909(.A(dpath_mulcore_ary2_cmux_n70), .Y(n5630));
AND2X1 mul_U16910(.A(n9153), .B(n9672), .Y(dpath_mulcore_ary2_cmux_n72));
INVX1 mul_U16911(.A(dpath_mulcore_ary2_cmux_n72), .Y(n5631));
AND2X1 mul_U16912(.A(n9154), .B(n9672), .Y(dpath_mulcore_ary2_cmux_n74));
INVX1 mul_U16913(.A(dpath_mulcore_ary2_cmux_n74), .Y(n5632));
AND2X1 mul_U16914(.A(n9155), .B(n9672), .Y(dpath_mulcore_ary2_cmux_n76));
INVX1 mul_U16915(.A(dpath_mulcore_ary2_cmux_n76), .Y(n5633));
AND2X1 mul_U16916(.A(n9156), .B(n9672), .Y(dpath_mulcore_ary2_cmux_n78));
INVX1 mul_U16917(.A(dpath_mulcore_ary2_cmux_n78), .Y(n5634));
AND2X1 mul_U16918(.A(n9157), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n80));
INVX1 mul_U16919(.A(dpath_mulcore_ary2_cmux_n80), .Y(n5635));
AND2X1 mul_U16920(.A(n9158), .B(n9692), .Y(dpath_mulcore_ary2_cmux_n82));
INVX1 mul_U16921(.A(dpath_mulcore_ary2_cmux_n82), .Y(n5636));
AND2X1 mul_U16922(.A(n6151), .B(n9693), .Y(dpath_mulcore_ary2_cmux_n84));
INVX1 mul_U16923(.A(dpath_mulcore_ary2_cmux_n84), .Y(n5637));
AND2X1 mul_U16924(.A(n9159), .B(dpath_mulcore_x2_c2c3), .Y(dpath_mulcore_ary2_cmux_n86));
INVX1 mul_U16925(.A(dpath_mulcore_ary2_cmux_n86), .Y(n5638));
AND2X1 mul_U16926(.A(n9160), .B(n9692), .Y(dpath_mulcore_ary2_cmux_n88));
INVX1 mul_U16927(.A(dpath_mulcore_ary2_cmux_n88), .Y(n5639));
AND2X1 mul_U16928(.A(n9161), .B(dpath_mulcore_x2_c2c3), .Y(dpath_mulcore_ary2_cmux_n90));
INVX1 mul_U16929(.A(dpath_mulcore_ary2_cmux_n90), .Y(n5640));
AND2X1 mul_U16930(.A(n9162), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n92));
INVX1 mul_U16931(.A(dpath_mulcore_ary2_cmux_n92), .Y(n5641));
AND2X1 mul_U16932(.A(n9163), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n94));
INVX1 mul_U16933(.A(dpath_mulcore_ary2_cmux_n94), .Y(n5642));
AND2X1 mul_U16934(.A(n9164), .B(n9689), .Y(dpath_mulcore_ary2_cmux_n96));
INVX1 mul_U16935(.A(dpath_mulcore_ary2_cmux_n96), .Y(n5643));
AND2X1 mul_U16936(.A(n9165), .B(n9673), .Y(dpath_mulcore_ary2_cmux_n98));
INVX1 mul_U16937(.A(dpath_mulcore_ary2_cmux_n98), .Y(n5644));
AND2X1 mul_U16938(.A(n9166), .B(dpath_mulcore_x2_c2c3), .Y(dpath_mulcore_ary2_cmux_n100));
INVX1 mul_U16939(.A(dpath_mulcore_ary2_cmux_n100), .Y(n5645));
AND2X1 mul_U16940(.A(n9167), .B(n9673), .Y(dpath_mulcore_ary2_cmux_n102));
INVX1 mul_U16941(.A(dpath_mulcore_ary2_cmux_n102), .Y(n5646));
AND2X1 mul_U16942(.A(n9168), .B(dpath_mulcore_x2_c2c3), .Y(dpath_mulcore_ary2_cmux_n104));
INVX1 mul_U16943(.A(dpath_mulcore_ary2_cmux_n104), .Y(n5647));
AND2X1 mul_U16944(.A(n6152), .B(n9673), .Y(dpath_mulcore_ary2_cmux_n106));
INVX1 mul_U16945(.A(dpath_mulcore_ary2_cmux_n106), .Y(n5648));
AND2X1 mul_U16946(.A(n9169), .B(dpath_mulcore_x2_c2c3), .Y(dpath_mulcore_ary2_cmux_n108));
INVX1 mul_U16947(.A(dpath_mulcore_ary2_cmux_n108), .Y(n5649));
AND2X1 mul_U16948(.A(n9170), .B(n9673), .Y(dpath_mulcore_ary2_cmux_n110));
INVX1 mul_U16949(.A(dpath_mulcore_ary2_cmux_n110), .Y(n5650));
AND2X1 mul_U16950(.A(n9171), .B(n9676), .Y(dpath_mulcore_ary2_cmux_n112));
INVX1 mul_U16951(.A(dpath_mulcore_ary2_cmux_n112), .Y(n5651));
AND2X1 mul_U16952(.A(n9172), .B(n9677), .Y(dpath_mulcore_ary2_cmux_n114));
INVX1 mul_U16953(.A(dpath_mulcore_ary2_cmux_n114), .Y(n5652));
AND2X1 mul_U16954(.A(n9173), .B(n9678), .Y(dpath_mulcore_ary2_cmux_n116));
INVX1 mul_U16955(.A(dpath_mulcore_ary2_cmux_n116), .Y(n5653));
AND2X1 mul_U16956(.A(n9174), .B(n9679), .Y(dpath_mulcore_ary2_cmux_n118));
INVX1 mul_U16957(.A(dpath_mulcore_ary2_cmux_n118), .Y(n5654));
AND2X1 mul_U16958(.A(n9175), .B(n9694), .Y(dpath_mulcore_ary2_cmux_n120));
INVX1 mul_U16959(.A(dpath_mulcore_ary2_cmux_n120), .Y(n5655));
AND2X1 mul_U16960(.A(n9176), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n122));
INVX1 mul_U16961(.A(dpath_mulcore_ary2_cmux_n122), .Y(n5656));
AND2X1 mul_U16962(.A(n9177), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n124));
INVX1 mul_U16963(.A(dpath_mulcore_ary2_cmux_n124), .Y(n5657));
AND2X1 mul_U16964(.A(n9178), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n126));
INVX1 mul_U16965(.A(dpath_mulcore_ary2_cmux_n126), .Y(n5658));
AND2X1 mul_U16966(.A(n6153), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n128));
INVX1 mul_U16967(.A(dpath_mulcore_ary2_cmux_n128), .Y(n5659));
AND2X1 mul_U16968(.A(n9179), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n130));
INVX1 mul_U16969(.A(dpath_mulcore_ary2_cmux_n130), .Y(n5660));
AND2X1 mul_U16970(.A(n9180), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n132));
INVX1 mul_U16971(.A(dpath_mulcore_ary2_cmux_n132), .Y(n5661));
AND2X1 mul_U16972(.A(n9181), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n134));
INVX1 mul_U16973(.A(dpath_mulcore_ary2_cmux_n134), .Y(n5662));
AND2X1 mul_U16974(.A(n9182), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n136));
INVX1 mul_U16975(.A(dpath_mulcore_ary2_cmux_n136), .Y(n5663));
AND2X1 mul_U16976(.A(n9183), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n138));
INVX1 mul_U16977(.A(dpath_mulcore_ary2_cmux_n138), .Y(n5664));
AND2X1 mul_U16978(.A(n9184), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n140));
INVX1 mul_U16979(.A(dpath_mulcore_ary2_cmux_n140), .Y(n5665));
AND2X1 mul_U16980(.A(n9185), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n142));
INVX1 mul_U16981(.A(dpath_mulcore_ary2_cmux_n142), .Y(n5666));
AND2X1 mul_U16982(.A(n9186), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n144));
INVX1 mul_U16983(.A(dpath_mulcore_ary2_cmux_n144), .Y(n5667));
AND2X1 mul_U16984(.A(n9187), .B(n9691), .Y(dpath_mulcore_ary2_cmux_n146));
INVX1 mul_U16985(.A(dpath_mulcore_ary2_cmux_n146), .Y(n5668));
AND2X1 mul_U16986(.A(n6141), .B(n9688), .Y(dpath_mulcore_ary2_cmux_n148));
INVX1 mul_U16987(.A(dpath_mulcore_ary2_cmux_n148), .Y(n5669));
AND2X1 mul_U16988(.A(n6154), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n150));
INVX1 mul_U16989(.A(dpath_mulcore_ary2_cmux_n150), .Y(n5670));
AND2X1 mul_U16990(.A(n6142), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n152));
INVX1 mul_U16991(.A(dpath_mulcore_ary2_cmux_n152), .Y(n5671));
AND2X1 mul_U16992(.A(n6143), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n154));
INVX1 mul_U16993(.A(dpath_mulcore_ary2_cmux_n154), .Y(n5672));
AND2X1 mul_U16994(.A(n6144), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n156));
INVX1 mul_U16995(.A(dpath_mulcore_ary2_cmux_n156), .Y(n5673));
AND2X1 mul_U16996(.A(n6145), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n158));
INVX1 mul_U16997(.A(dpath_mulcore_ary2_cmux_n158), .Y(n5674));
AND2X1 mul_U16998(.A(n6146), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n160));
INVX1 mul_U16999(.A(dpath_mulcore_ary2_cmux_n160), .Y(n5675));
AND2X1 mul_U17000(.A(n6147), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n162));
INVX1 mul_U17001(.A(dpath_mulcore_ary2_cmux_n162), .Y(n5676));
AND2X1 mul_U17002(.A(n6148), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n164));
INVX1 mul_U17003(.A(dpath_mulcore_ary2_cmux_n164), .Y(n5677));
AND2X1 mul_U17004(.A(n6149), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n166));
INVX1 mul_U17005(.A(dpath_mulcore_ary2_cmux_n166), .Y(n5678));
AND2X1 mul_U17006(.A(n6150), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n168));
INVX1 mul_U17007(.A(dpath_mulcore_ary2_cmux_n168), .Y(n5679));
AND2X1 mul_U17008(.A(n6164), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n170));
INVX1 mul_U17009(.A(dpath_mulcore_ary2_cmux_n170), .Y(n5680));
AND2X1 mul_U17010(.A(dpath_mulcore_pcout[0]), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n172));
INVX1 mul_U17011(.A(dpath_mulcore_ary2_cmux_n172), .Y(n5681));
AND2X1 mul_U17012(.A(n6165), .B(n9687), .Y(dpath_mulcore_ary2_cmux_n174));
INVX1 mul_U17013(.A(dpath_mulcore_ary2_cmux_n174), .Y(n5682));
AND2X1 mul_U17014(.A(n6166), .B(n9686), .Y(dpath_mulcore_ary2_cmux_n176));
INVX1 mul_U17015(.A(dpath_mulcore_ary2_cmux_n176), .Y(n5683));
AND2X1 mul_U17016(.A(n6167), .B(n9686), .Y(dpath_mulcore_ary2_cmux_n178));
INVX1 mul_U17017(.A(dpath_mulcore_ary2_cmux_n178), .Y(n5684));
AND2X1 mul_U17018(.A(n16563), .B(n9686), .Y(dpath_mulcore_ary2_cmux_n180));
INVX1 mul_U17019(.A(dpath_mulcore_ary2_cmux_n180), .Y(n5685));
AND2X1 mul_U17020(.A(n6155), .B(n9686), .Y(dpath_mulcore_ary2_cmux_n182));
INVX1 mul_U17021(.A(dpath_mulcore_ary2_cmux_n182), .Y(n5686));
AND2X1 mul_U17022(.A(n6156), .B(n9686), .Y(dpath_mulcore_ary2_cmux_n184));
INVX1 mul_U17023(.A(dpath_mulcore_ary2_cmux_n184), .Y(n5687));
AND2X1 mul_U17024(.A(n6157), .B(n9695), .Y(dpath_mulcore_ary2_cmux_n186));
INVX1 mul_U17025(.A(dpath_mulcore_ary2_cmux_n186), .Y(n5688));
AND2X1 mul_U17026(.A(n6158), .B(n9686), .Y(dpath_mulcore_ary2_cmux_n188));
INVX1 mul_U17027(.A(dpath_mulcore_ary2_cmux_n188), .Y(n5689));
AND2X1 mul_U17028(.A(n6159), .B(n9686), .Y(dpath_mulcore_ary2_cmux_n190));
INVX1 mul_U17029(.A(dpath_mulcore_ary2_cmux_n190), .Y(n5690));
AND2X1 mul_U17030(.A(n6160), .B(n9686), .Y(dpath_mulcore_ary2_cmux_n192));
INVX1 mul_U17031(.A(dpath_mulcore_ary2_cmux_n192), .Y(n5691));
AND2X1 mul_U17032(.A(dpath_mulcore_pcoutx2), .B(n9686), .Y(dpath_mulcore_ary2_cmux_n194));
INVX1 mul_U17033(.A(dpath_mulcore_ary2_cmux_n194), .Y(n5692));
AND2X1 mul_U17034(.A(dpath_mout[9]), .B(n9753), .Y(dpath_n525));
INVX1 mul_U17035(.A(dpath_n525), .Y(n5693));
AND2X1 mul_U17036(.A(dpath_mout[8]), .B(n9753), .Y(dpath_n527));
INVX1 mul_U17037(.A(dpath_n527), .Y(n5694));
AND2X1 mul_U17038(.A(dpath_mout[7]), .B(n9753), .Y(dpath_n529));
INVX1 mul_U17039(.A(dpath_n529), .Y(n5695));
AND2X1 mul_U17040(.A(dpath_mout[6]), .B(n9753), .Y(dpath_n531));
INVX1 mul_U17041(.A(dpath_n531), .Y(n5696));
AND2X1 mul_U17042(.A(dpath_mout[63]), .B(n9753), .Y(dpath_n533));
INVX1 mul_U17043(.A(dpath_n533), .Y(n5697));
AND2X1 mul_U17044(.A(dpath_mout[62]), .B(n9753), .Y(dpath_n535));
INVX1 mul_U17045(.A(dpath_n535), .Y(n5698));
AND2X1 mul_U17046(.A(dpath_mout[61]), .B(n9753), .Y(dpath_n537));
INVX1 mul_U17047(.A(dpath_n537), .Y(n5699));
AND2X1 mul_U17048(.A(dpath_mout[60]), .B(n9753), .Y(dpath_n539));
INVX1 mul_U17049(.A(dpath_n539), .Y(n5700));
AND2X1 mul_U17050(.A(dpath_mout[5]), .B(n9753), .Y(dpath_n541));
INVX1 mul_U17051(.A(dpath_n541), .Y(n5701));
AND2X1 mul_U17052(.A(dpath_mout[59]), .B(n9753), .Y(dpath_n543));
INVX1 mul_U17053(.A(dpath_n543), .Y(n5702));
AND2X1 mul_U17054(.A(dpath_mout[58]), .B(n9753), .Y(dpath_n545));
INVX1 mul_U17055(.A(dpath_n545), .Y(n5703));
AND2X1 mul_U17056(.A(dpath_mout[57]), .B(n9753), .Y(dpath_n547));
INVX1 mul_U17057(.A(dpath_n547), .Y(n5704));
AND2X1 mul_U17058(.A(dpath_mout[56]), .B(n9753), .Y(dpath_n549));
INVX1 mul_U17059(.A(dpath_n549), .Y(n5705));
AND2X1 mul_U17060(.A(dpath_mout[55]), .B(n9753), .Y(dpath_n551));
INVX1 mul_U17061(.A(dpath_n551), .Y(n5706));
AND2X1 mul_U17062(.A(dpath_mout[54]), .B(n9753), .Y(dpath_n553));
INVX1 mul_U17063(.A(dpath_n553), .Y(n5707));
AND2X1 mul_U17064(.A(dpath_mout[53]), .B(n9753), .Y(dpath_n555));
INVX1 mul_U17065(.A(dpath_n555), .Y(n5708));
AND2X1 mul_U17066(.A(dpath_mout[52]), .B(n9753), .Y(dpath_n557));
INVX1 mul_U17067(.A(dpath_n557), .Y(n5709));
AND2X1 mul_U17068(.A(dpath_mout[51]), .B(n9753), .Y(dpath_n559));
INVX1 mul_U17069(.A(dpath_n559), .Y(n5710));
AND2X1 mul_U17070(.A(dpath_mout[50]), .B(n9753), .Y(dpath_n561));
INVX1 mul_U17071(.A(dpath_n561), .Y(n5711));
AND2X1 mul_U17072(.A(dpath_mout[4]), .B(n9753), .Y(dpath_n563));
INVX1 mul_U17073(.A(dpath_n563), .Y(n5712));
AND2X1 mul_U17074(.A(dpath_mout[49]), .B(n9753), .Y(dpath_n565));
INVX1 mul_U17075(.A(dpath_n565), .Y(n5713));
AND2X1 mul_U17076(.A(dpath_mout[48]), .B(n9753), .Y(dpath_n567));
INVX1 mul_U17077(.A(dpath_n567), .Y(n5714));
AND2X1 mul_U17078(.A(dpath_mout[47]), .B(n9753), .Y(dpath_n569));
INVX1 mul_U17079(.A(dpath_n569), .Y(n5715));
AND2X1 mul_U17080(.A(dpath_mout[46]), .B(n9753), .Y(dpath_n571));
INVX1 mul_U17081(.A(dpath_n571), .Y(n5716));
AND2X1 mul_U17082(.A(dpath_mout[45]), .B(n9753), .Y(dpath_n573));
INVX1 mul_U17083(.A(dpath_n573), .Y(n5717));
AND2X1 mul_U17084(.A(dpath_mout[44]), .B(n9753), .Y(dpath_n575));
INVX1 mul_U17085(.A(dpath_n575), .Y(n5718));
AND2X1 mul_U17086(.A(dpath_mout[43]), .B(n9753), .Y(dpath_n577));
INVX1 mul_U17087(.A(dpath_n577), .Y(n5719));
AND2X1 mul_U17088(.A(dpath_mout[42]), .B(n9753), .Y(dpath_n579));
INVX1 mul_U17089(.A(dpath_n579), .Y(n5720));
AND2X1 mul_U17090(.A(dpath_mout[41]), .B(n9753), .Y(dpath_n581));
INVX1 mul_U17091(.A(dpath_n581), .Y(n5721));
AND2X1 mul_U17092(.A(dpath_mout[40]), .B(n9753), .Y(dpath_n583));
INVX1 mul_U17093(.A(dpath_n583), .Y(n5722));
AND2X1 mul_U17094(.A(dpath_mout[3]), .B(n9753), .Y(dpath_n585));
INVX1 mul_U17095(.A(dpath_n585), .Y(n5723));
AND2X1 mul_U17096(.A(dpath_mout[39]), .B(n9753), .Y(dpath_n587));
INVX1 mul_U17097(.A(dpath_n587), .Y(n5724));
AND2X1 mul_U17098(.A(dpath_mout[38]), .B(n9753), .Y(dpath_n589));
INVX1 mul_U17099(.A(dpath_n589), .Y(n5725));
AND2X1 mul_U17100(.A(dpath_mout[37]), .B(n9753), .Y(dpath_n591));
INVX1 mul_U17101(.A(dpath_n591), .Y(n5726));
AND2X1 mul_U17102(.A(dpath_mout[36]), .B(n9753), .Y(dpath_n593));
INVX1 mul_U17103(.A(dpath_n593), .Y(n5727));
AND2X1 mul_U17104(.A(dpath_mout[35]), .B(n9753), .Y(dpath_n595));
INVX1 mul_U17105(.A(dpath_n595), .Y(n5728));
AND2X1 mul_U17106(.A(dpath_mout[34]), .B(n9753), .Y(dpath_n597));
INVX1 mul_U17107(.A(dpath_n597), .Y(n5729));
AND2X1 mul_U17108(.A(dpath_mout[33]), .B(n9753), .Y(dpath_n599));
INVX1 mul_U17109(.A(dpath_n599), .Y(n5730));
AND2X1 mul_U17110(.A(dpath_mout[32]), .B(n9753), .Y(dpath_n601));
INVX1 mul_U17111(.A(dpath_n601), .Y(n5731));
AND2X1 mul_U17112(.A(dpath_mout[31]), .B(n9753), .Y(dpath_n603));
INVX1 mul_U17113(.A(dpath_n603), .Y(n5732));
AND2X1 mul_U17114(.A(dpath_mout[30]), .B(n9753), .Y(dpath_n605));
INVX1 mul_U17115(.A(dpath_n605), .Y(n5733));
AND2X1 mul_U17116(.A(dpath_mout[2]), .B(n9753), .Y(dpath_n607));
INVX1 mul_U17117(.A(dpath_n607), .Y(n5734));
AND2X1 mul_U17118(.A(dpath_mout[29]), .B(n9753), .Y(dpath_n609));
INVX1 mul_U17119(.A(dpath_n609), .Y(n5735));
AND2X1 mul_U17120(.A(dpath_mout[28]), .B(n9753), .Y(dpath_n611));
INVX1 mul_U17121(.A(dpath_n611), .Y(n5736));
AND2X1 mul_U17122(.A(dpath_mout[27]), .B(n9753), .Y(dpath_n613));
INVX1 mul_U17123(.A(dpath_n613), .Y(n5737));
AND2X1 mul_U17124(.A(dpath_mout[26]), .B(n9753), .Y(dpath_n615));
INVX1 mul_U17125(.A(dpath_n615), .Y(n5738));
AND2X1 mul_U17126(.A(dpath_mout[25]), .B(n9753), .Y(dpath_n617));
INVX1 mul_U17127(.A(dpath_n617), .Y(n5739));
AND2X1 mul_U17128(.A(dpath_mout[24]), .B(n9753), .Y(dpath_n619));
INVX1 mul_U17129(.A(dpath_n619), .Y(n5740));
AND2X1 mul_U17130(.A(dpath_mout[23]), .B(n9753), .Y(dpath_n621));
INVX1 mul_U17131(.A(dpath_n621), .Y(n5741));
AND2X1 mul_U17132(.A(dpath_mout[22]), .B(n9753), .Y(dpath_n623));
INVX1 mul_U17133(.A(dpath_n623), .Y(n5742));
AND2X1 mul_U17134(.A(dpath_mout[21]), .B(n9753), .Y(dpath_n625));
INVX1 mul_U17135(.A(dpath_n625), .Y(n5743));
AND2X1 mul_U17136(.A(dpath_mout[20]), .B(n9753), .Y(dpath_n627));
INVX1 mul_U17137(.A(dpath_n627), .Y(n5744));
AND2X1 mul_U17138(.A(dpath_mout[1]), .B(n9753), .Y(dpath_n629));
INVX1 mul_U17139(.A(dpath_n629), .Y(n5745));
AND2X1 mul_U17140(.A(dpath_mout[19]), .B(n9753), .Y(dpath_n631));
INVX1 mul_U17141(.A(dpath_n631), .Y(n5746));
AND2X1 mul_U17142(.A(dpath_mout[18]), .B(n9753), .Y(dpath_n633));
INVX1 mul_U17143(.A(dpath_n633), .Y(n5747));
AND2X1 mul_U17144(.A(dpath_mout[17]), .B(n9753), .Y(dpath_n635));
INVX1 mul_U17145(.A(dpath_n635), .Y(n5748));
AND2X1 mul_U17146(.A(dpath_mout[16]), .B(n9753), .Y(dpath_n637));
INVX1 mul_U17147(.A(dpath_n637), .Y(n5749));
AND2X1 mul_U17148(.A(dpath_mout[15]), .B(n9753), .Y(dpath_n639));
INVX1 mul_U17149(.A(dpath_n639), .Y(n5750));
AND2X1 mul_U17150(.A(dpath_mout[14]), .B(n9753), .Y(dpath_n641));
INVX1 mul_U17151(.A(dpath_n641), .Y(n5751));
AND2X1 mul_U17152(.A(dpath_mout[13]), .B(n9753), .Y(dpath_n643));
INVX1 mul_U17153(.A(dpath_n643), .Y(n5752));
AND2X1 mul_U17154(.A(dpath_mout[12]), .B(n9753), .Y(dpath_n645));
INVX1 mul_U17155(.A(dpath_n645), .Y(n5753));
AND2X1 mul_U17156(.A(dpath_mout[11]), .B(n9753), .Y(dpath_n647));
INVX1 mul_U17157(.A(dpath_n647), .Y(n5754));
AND2X1 mul_U17158(.A(dpath_mout[10]), .B(n9753), .Y(dpath_n649));
INVX1 mul_U17159(.A(dpath_n649), .Y(n5755));
AND2X1 mul_U17160(.A(dpath_mout[0]), .B(n9753), .Y(dpath_n651));
INVX1 mul_U17161(.A(dpath_n651), .Y(n5756));
AND2X1 mul_U17162(.A(dpath_mout[9]), .B(n9782), .Y(dpath_n985));
INVX1 mul_U17163(.A(dpath_n985), .Y(n5757));
AND2X1 mul_U17164(.A(dpath_mout[8]), .B(n9783), .Y(dpath_n987));
INVX1 mul_U17165(.A(dpath_n987), .Y(n5758));
AND2X1 mul_U17166(.A(dpath_mout[7]), .B(n9781), .Y(dpath_n989));
INVX1 mul_U17167(.A(dpath_n989), .Y(n5759));
AND2X1 mul_U17168(.A(dpath_mout[71]), .B(n9778), .Y(dpath_n991));
INVX1 mul_U17169(.A(dpath_n991), .Y(n5760));
AND2X1 mul_U17170(.A(dpath_mout[70]), .B(n9779), .Y(dpath_n993));
INVX1 mul_U17171(.A(dpath_n993), .Y(n5761));
AND2X1 mul_U17172(.A(dpath_mout[6]), .B(n9780), .Y(dpath_n995));
INVX1 mul_U17173(.A(dpath_n995), .Y(n5762));
AND2X1 mul_U17174(.A(dpath_mout[69]), .B(n9779), .Y(dpath_n997));
INVX1 mul_U17175(.A(dpath_n997), .Y(n5763));
AND2X1 mul_U17176(.A(dpath_mout[68]), .B(n9779), .Y(dpath_n999));
INVX1 mul_U17177(.A(dpath_n999), .Y(n5764));
AND2X1 mul_U17178(.A(dpath_mout[67]), .B(n9779), .Y(dpath_n1001));
INVX1 mul_U17179(.A(dpath_n1001), .Y(n5765));
AND2X1 mul_U17180(.A(dpath_mout[66]), .B(n9779), .Y(dpath_n1003));
INVX1 mul_U17181(.A(dpath_n1003), .Y(n5766));
AND2X1 mul_U17182(.A(dpath_mout[65]), .B(n9778), .Y(dpath_n1005));
INVX1 mul_U17183(.A(dpath_n1005), .Y(n5767));
AND2X1 mul_U17184(.A(dpath_mout[64]), .B(n9780), .Y(dpath_n1007));
INVX1 mul_U17185(.A(dpath_n1007), .Y(n5768));
AND2X1 mul_U17186(.A(dpath_mout[63]), .B(n9779), .Y(dpath_n1009));
INVX1 mul_U17187(.A(dpath_n1009), .Y(n5769));
AND2X1 mul_U17188(.A(dpath_mout[62]), .B(n9781), .Y(dpath_n1011));
INVX1 mul_U17189(.A(dpath_n1011), .Y(n5770));
AND2X1 mul_U17190(.A(dpath_mout[61]), .B(n9778), .Y(dpath_n1013));
INVX1 mul_U17191(.A(dpath_n1013), .Y(n5771));
AND2X1 mul_U17192(.A(dpath_mout[60]), .B(n9783), .Y(dpath_n1015));
INVX1 mul_U17193(.A(dpath_n1015), .Y(n5772));
AND2X1 mul_U17194(.A(dpath_mout[5]), .B(n9782), .Y(dpath_n1017));
INVX1 mul_U17195(.A(dpath_n1017), .Y(n5773));
AND2X1 mul_U17196(.A(dpath_mout[59]), .B(n9781), .Y(dpath_n1019));
INVX1 mul_U17197(.A(dpath_n1019), .Y(n5774));
AND2X1 mul_U17198(.A(dpath_mout[58]), .B(n9778), .Y(dpath_n1021));
INVX1 mul_U17199(.A(dpath_n1021), .Y(n5775));
AND2X1 mul_U17200(.A(dpath_mout[57]), .B(n9779), .Y(dpath_n1023));
INVX1 mul_U17201(.A(dpath_n1023), .Y(n5776));
AND2X1 mul_U17202(.A(dpath_mout[56]), .B(n9778), .Y(dpath_n1025));
INVX1 mul_U17203(.A(dpath_n1025), .Y(n5777));
AND2X1 mul_U17204(.A(dpath_mout[55]), .B(n9780), .Y(dpath_n1027));
INVX1 mul_U17205(.A(dpath_n1027), .Y(n5778));
AND2X1 mul_U17206(.A(dpath_mout[54]), .B(n9782), .Y(dpath_n1029));
INVX1 mul_U17207(.A(dpath_n1029), .Y(n5779));
AND2X1 mul_U17208(.A(dpath_mout[53]), .B(n9783), .Y(dpath_n1031));
INVX1 mul_U17209(.A(dpath_n1031), .Y(n5780));
AND2X1 mul_U17210(.A(dpath_mout[52]), .B(n9781), .Y(dpath_n1033));
INVX1 mul_U17211(.A(dpath_n1033), .Y(n5781));
AND2X1 mul_U17212(.A(dpath_mout[51]), .B(n9778), .Y(dpath_n1035));
INVX1 mul_U17213(.A(dpath_n1035), .Y(n5782));
AND2X1 mul_U17214(.A(dpath_mout[50]), .B(n9778), .Y(dpath_n1037));
INVX1 mul_U17215(.A(dpath_n1037), .Y(n5783));
AND2X1 mul_U17216(.A(dpath_mout[4]), .B(n9779), .Y(dpath_n1039));
INVX1 mul_U17217(.A(dpath_n1039), .Y(n5784));
AND2X1 mul_U17218(.A(dpath_mout[49]), .B(n9778), .Y(dpath_n1041));
INVX1 mul_U17219(.A(dpath_n1041), .Y(n5785));
AND2X1 mul_U17220(.A(dpath_mout[48]), .B(n9780), .Y(dpath_n1043));
INVX1 mul_U17221(.A(dpath_n1043), .Y(n5786));
AND2X1 mul_U17222(.A(dpath_mout[47]), .B(n9782), .Y(dpath_n1045));
INVX1 mul_U17223(.A(dpath_n1045), .Y(n5787));
AND2X1 mul_U17224(.A(dpath_mout[46]), .B(n9783), .Y(dpath_n1047));
INVX1 mul_U17225(.A(dpath_n1047), .Y(n5788));
AND2X1 mul_U17226(.A(dpath_mout[45]), .B(n9779), .Y(dpath_n1049));
INVX1 mul_U17227(.A(dpath_n1049), .Y(n5789));
AND2X1 mul_U17228(.A(dpath_mout[44]), .B(n9779), .Y(dpath_n1051));
INVX1 mul_U17229(.A(dpath_n1051), .Y(n5790));
AND2X1 mul_U17230(.A(dpath_mout[43]), .B(n9782), .Y(dpath_n1053));
INVX1 mul_U17231(.A(dpath_n1053), .Y(n5791));
AND2X1 mul_U17232(.A(dpath_mout[42]), .B(n9783), .Y(dpath_n1055));
INVX1 mul_U17233(.A(dpath_n1055), .Y(n5792));
AND2X1 mul_U17234(.A(dpath_mout[41]), .B(n9781), .Y(dpath_n1057));
INVX1 mul_U17235(.A(dpath_n1057), .Y(n5793));
AND2X1 mul_U17236(.A(dpath_mout[40]), .B(n9778), .Y(dpath_n1059));
INVX1 mul_U17237(.A(dpath_n1059), .Y(n5794));
AND2X1 mul_U17238(.A(dpath_mout[3]), .B(n9779), .Y(dpath_n1061));
INVX1 mul_U17239(.A(dpath_n1061), .Y(n5795));
AND2X1 mul_U17240(.A(dpath_mout[39]), .B(n9779), .Y(dpath_n1063));
INVX1 mul_U17241(.A(dpath_n1063), .Y(n5796));
AND2X1 mul_U17242(.A(dpath_mout[38]), .B(n9778), .Y(dpath_n1065));
INVX1 mul_U17243(.A(dpath_n1065), .Y(n5797));
AND2X1 mul_U17244(.A(dpath_mout[37]), .B(n9780), .Y(dpath_n1067));
INVX1 mul_U17245(.A(dpath_n1067), .Y(n5798));
AND2X1 mul_U17246(.A(dpath_mout[36]), .B(n9781), .Y(dpath_n1069));
INVX1 mul_U17247(.A(dpath_n1069), .Y(n5799));
AND2X1 mul_U17248(.A(dpath_mout[35]), .B(n9782), .Y(dpath_n1071));
INVX1 mul_U17249(.A(dpath_n1071), .Y(n5800));
AND2X1 mul_U17250(.A(dpath_mout[34]), .B(n9783), .Y(dpath_n1073));
INVX1 mul_U17251(.A(dpath_n1073), .Y(n5801));
AND2X1 mul_U17252(.A(dpath_mout[33]), .B(n9779), .Y(dpath_n1075));
INVX1 mul_U17253(.A(dpath_n1075), .Y(n5802));
AND2X1 mul_U17254(.A(dpath_mout[32]), .B(n9778), .Y(dpath_n1077));
INVX1 mul_U17255(.A(dpath_n1077), .Y(n5803));
AND2X1 mul_U17256(.A(dpath_mout[31]), .B(n9779), .Y(dpath_n1079));
INVX1 mul_U17257(.A(dpath_n1079), .Y(n5804));
AND2X1 mul_U17258(.A(dpath_mout[30]), .B(n9778), .Y(dpath_n1081));
INVX1 mul_U17259(.A(dpath_n1081), .Y(n5805));
AND2X1 mul_U17260(.A(dpath_mout[2]), .B(n9779), .Y(dpath_n1083));
INVX1 mul_U17261(.A(dpath_n1083), .Y(n5806));
AND2X1 mul_U17262(.A(dpath_mout[29]), .B(n9778), .Y(dpath_n1085));
INVX1 mul_U17263(.A(dpath_n1085), .Y(n5807));
AND2X1 mul_U17264(.A(dpath_mout[28]), .B(n9779), .Y(dpath_n1087));
INVX1 mul_U17265(.A(dpath_n1087), .Y(n5808));
AND2X1 mul_U17266(.A(dpath_mout[27]), .B(n9780), .Y(dpath_n1089));
INVX1 mul_U17267(.A(dpath_n1089), .Y(n5809));
AND2X1 mul_U17268(.A(dpath_mout[26]), .B(n9778), .Y(dpath_n1091));
INVX1 mul_U17269(.A(dpath_n1091), .Y(n5810));
AND2X1 mul_U17270(.A(dpath_mout[25]), .B(n9779), .Y(dpath_n1093));
INVX1 mul_U17271(.A(dpath_n1093), .Y(n5811));
AND2X1 mul_U17272(.A(dpath_mout[24]), .B(n9780), .Y(dpath_n1095));
INVX1 mul_U17273(.A(dpath_n1095), .Y(n5812));
AND2X1 mul_U17274(.A(dpath_mout[23]), .B(n9779), .Y(dpath_n1097));
INVX1 mul_U17275(.A(dpath_n1097), .Y(n5813));
AND2X1 mul_U17276(.A(dpath_mout[22]), .B(n9778), .Y(dpath_n1099));
INVX1 mul_U17277(.A(dpath_n1099), .Y(n5814));
AND2X1 mul_U17278(.A(dpath_mout[21]), .B(n9780), .Y(dpath_n1101));
INVX1 mul_U17279(.A(dpath_n1101), .Y(n5815));
AND2X1 mul_U17280(.A(dpath_mout[20]), .B(n9780), .Y(dpath_n1103));
INVX1 mul_U17281(.A(dpath_n1103), .Y(n5816));
AND2X1 mul_U17282(.A(dpath_mout[1]), .B(n9780), .Y(dpath_n1105));
INVX1 mul_U17283(.A(dpath_n1105), .Y(n5817));
AND2X1 mul_U17284(.A(dpath_mout[19]), .B(n9780), .Y(dpath_n1107));
INVX1 mul_U17285(.A(dpath_n1107), .Y(n5818));
AND2X1 mul_U17286(.A(dpath_mout[18]), .B(n9780), .Y(dpath_n1109));
INVX1 mul_U17287(.A(dpath_n1109), .Y(n5819));
AND2X1 mul_U17288(.A(dpath_mout[17]), .B(n9780), .Y(dpath_n1111));
INVX1 mul_U17289(.A(dpath_n1111), .Y(n5820));
AND2X1 mul_U17290(.A(dpath_mout[16]), .B(n9780), .Y(dpath_n1113));
INVX1 mul_U17291(.A(dpath_n1113), .Y(n5821));
AND2X1 mul_U17292(.A(dpath_mout[15]), .B(n9780), .Y(dpath_n1115));
INVX1 mul_U17293(.A(dpath_n1115), .Y(n5822));
AND2X1 mul_U17294(.A(dpath_mout[14]), .B(n9780), .Y(dpath_n1117));
INVX1 mul_U17295(.A(dpath_n1117), .Y(n5823));
AND2X1 mul_U17296(.A(dpath_mout[13]), .B(n9780), .Y(dpath_n1119));
INVX1 mul_U17297(.A(dpath_n1119), .Y(n5824));
AND2X1 mul_U17298(.A(dpath_mout[12]), .B(n9780), .Y(dpath_n1121));
INVX1 mul_U17299(.A(dpath_n1121), .Y(n5825));
AND2X1 mul_U17300(.A(dpath_mout[11]), .B(n9780), .Y(dpath_n1123));
INVX1 mul_U17301(.A(dpath_n1123), .Y(n5826));
AND2X1 mul_U17302(.A(dpath_mout[10]), .B(n9780), .Y(dpath_n1125));
INVX1 mul_U17303(.A(dpath_n1125), .Y(n5827));
AND2X1 mul_U17304(.A(dpath_mout[0]), .B(n9782), .Y(dpath_n1127));
INVX1 mul_U17305(.A(dpath_n1127), .Y(n5828));
OR2X1 mul_U17306(.A(control_acc_actc4), .B(acc_actc3), .Y(control_n25));
INVX1 mul_U17307(.A(control_n25), .Y(n5829));
AND2X1 mul_U17308(.A(dpath_acc_reg[134]), .B(dpath_acc_reg[133]), .Y(n10600));
INVX1 mul_U17309(.A(n10600), .Y(n5830));
INVX1 mul_U17310(.A(control_n13), .Y(n5831));
INVX1 mul_U17311(.A(dpath_n137), .Y(n5832));
INVX1 mul_U17312(.A(dpath_n146), .Y(n5833));
INVX1 mul_U17313(.A(dpath_n152), .Y(n5834));
INVX1 mul_U17314(.A(dpath_n158), .Y(n5835));
INVX1 mul_U17315(.A(dpath_n164), .Y(n5836));
INVX1 mul_U17316(.A(dpath_n170), .Y(n5837));
INVX1 mul_U17317(.A(dpath_n176), .Y(n5838));
INVX1 mul_U17318(.A(dpath_n182), .Y(n5839));
INVX1 mul_U17319(.A(dpath_n188), .Y(n5840));
INVX1 mul_U17320(.A(dpath_n194), .Y(n5841));
INVX1 mul_U17321(.A(dpath_n200), .Y(n5842));
INVX1 mul_U17322(.A(dpath_n206), .Y(n5843));
INVX1 mul_U17323(.A(dpath_n212), .Y(n5844));
INVX1 mul_U17324(.A(dpath_n218), .Y(n5845));
INVX1 mul_U17325(.A(dpath_n224), .Y(n5846));
INVX1 mul_U17326(.A(dpath_n230), .Y(n5847));
INVX1 mul_U17327(.A(dpath_n236), .Y(n5848));
INVX1 mul_U17328(.A(dpath_n242), .Y(n5849));
INVX1 mul_U17329(.A(dpath_n248), .Y(n5850));
INVX1 mul_U17330(.A(dpath_n254), .Y(n5851));
INVX1 mul_U17331(.A(dpath_n260), .Y(n5852));
INVX1 mul_U17332(.A(dpath_n266), .Y(n5853));
INVX1 mul_U17333(.A(dpath_n272), .Y(n5854));
INVX1 mul_U17334(.A(dpath_n278), .Y(n5855));
INVX1 mul_U17335(.A(dpath_n284), .Y(n5856));
INVX1 mul_U17336(.A(dpath_n290), .Y(n5857));
INVX1 mul_U17337(.A(dpath_n296), .Y(n5858));
INVX1 mul_U17338(.A(dpath_n302), .Y(n5859));
INVX1 mul_U17339(.A(dpath_n308), .Y(n5860));
INVX1 mul_U17340(.A(dpath_n314), .Y(n5861));
INVX1 mul_U17341(.A(dpath_n320), .Y(n5862));
INVX1 mul_U17342(.A(dpath_n326), .Y(n5863));
INVX1 mul_U17343(.A(dpath_n332), .Y(n5864));
INVX1 mul_U17344(.A(dpath_n338), .Y(n5865));
INVX1 mul_U17345(.A(dpath_n344), .Y(n5866));
INVX1 mul_U17346(.A(dpath_n350), .Y(n5867));
INVX1 mul_U17347(.A(dpath_n356), .Y(n5868));
INVX1 mul_U17348(.A(dpath_n362), .Y(n5869));
INVX1 mul_U17349(.A(dpath_n368), .Y(n5870));
INVX1 mul_U17350(.A(dpath_n374), .Y(n5871));
INVX1 mul_U17351(.A(dpath_n380), .Y(n5872));
INVX1 mul_U17352(.A(dpath_n386), .Y(n5873));
INVX1 mul_U17353(.A(dpath_n392), .Y(n5874));
INVX1 mul_U17354(.A(dpath_n398), .Y(n5875));
INVX1 mul_U17355(.A(dpath_n404), .Y(n5876));
INVX1 mul_U17356(.A(dpath_n410), .Y(n5877));
INVX1 mul_U17357(.A(dpath_n416), .Y(n5878));
INVX1 mul_U17358(.A(dpath_n422), .Y(n5879));
INVX1 mul_U17359(.A(dpath_n428), .Y(n5880));
INVX1 mul_U17360(.A(dpath_n434), .Y(n5881));
INVX1 mul_U17361(.A(dpath_n440), .Y(n5882));
INVX1 mul_U17362(.A(dpath_n446), .Y(n5883));
INVX1 mul_U17363(.A(dpath_n452), .Y(n5884));
INVX1 mul_U17364(.A(dpath_n458), .Y(n5885));
INVX1 mul_U17365(.A(dpath_n464), .Y(n5886));
INVX1 mul_U17366(.A(dpath_n470), .Y(n5887));
INVX1 mul_U17367(.A(dpath_n476), .Y(n5888));
INVX1 mul_U17368(.A(dpath_n482), .Y(n5889));
INVX1 mul_U17369(.A(dpath_n488), .Y(n5890));
INVX1 mul_U17370(.A(dpath_n494), .Y(n5891));
INVX1 mul_U17371(.A(dpath_n500), .Y(n5892));
INVX1 mul_U17372(.A(dpath_n506), .Y(n5893));
INVX1 mul_U17373(.A(dpath_n512), .Y(n5894));
INVX1 mul_U17374(.A(dpath_n518), .Y(n5895));
INVX1 mul_U17375(.A(dpath_n653), .Y(n5896));
INVX1 mul_U17376(.A(dpath_n679), .Y(n5897));
INVX1 mul_U17377(.A(dpath_n705), .Y(n5898));
INVX1 mul_U17378(.A(dpath_n731), .Y(n5899));
INVX1 mul_U17379(.A(dpath_n757), .Y(n5900));
INVX1 mul_U17380(.A(dpath_n783), .Y(n5901));
INVX1 mul_U17381(.A(dpath_n809), .Y(n5902));
INVX1 mul_U17382(.A(dpath_n831), .Y(n5903));
INVX1 mul_U17383(.A(dpath_n837), .Y(n5904));
INVX1 mul_U17384(.A(dpath_n843), .Y(n5905));
INVX1 mul_U17385(.A(dpath_n849), .Y(n5906));
INVX1 mul_U17386(.A(dpath_n855), .Y(n5907));
INVX1 mul_U17387(.A(dpath_n861), .Y(n5908));
INVX1 mul_U17388(.A(dpath_n867), .Y(n5909));
INVX1 mul_U17389(.A(dpath_n873), .Y(n5910));
INVX1 mul_U17390(.A(dpath_n879), .Y(n5911));
INVX1 mul_U17391(.A(dpath_n885), .Y(n5912));
INVX1 mul_U17392(.A(dpath_n891), .Y(n5913));
INVX1 mul_U17393(.A(dpath_n897), .Y(n5914));
INVX1 mul_U17394(.A(dpath_n903), .Y(n5915));
INVX1 mul_U17395(.A(dpath_n909), .Y(n5916));
INVX1 mul_U17396(.A(dpath_n915), .Y(n5917));
INVX1 mul_U17397(.A(dpath_n921), .Y(n5918));
INVX1 mul_U17398(.A(dpath_n927), .Y(n5919));
INVX1 mul_U17399(.A(dpath_n933), .Y(n5920));
INVX1 mul_U17400(.A(dpath_n939), .Y(n5921));
INVX1 mul_U17401(.A(dpath_n945), .Y(n5922));
INVX1 mul_U17402(.A(dpath_n951), .Y(n5923));
INVX1 mul_U17403(.A(dpath_n957), .Y(n5924));
INVX1 mul_U17404(.A(dpath_n963), .Y(n5925));
INVX1 mul_U17405(.A(dpath_n969), .Y(n5926));
INVX1 mul_U17406(.A(dpath_n975), .Y(n5927));
AND2X1 mul_U17407(.A(dpath_mulcore_b4[1]), .B(n9730), .Y(n13691));
INVX1 mul_U17408(.A(n13691), .Y(n5928));
AND2X1 mul_U17409(.A(dpath_mulcore_b4[1]), .B(dpath_mulcore_b4[0]), .Y(n13692));
INVX1 mul_U17410(.A(n13692), .Y(n5929));
AND2X1 mul_U17411(.A(dpath_mulcore_b3[1]), .B(n9728), .Y(n13693));
INVX1 mul_U17412(.A(n13693), .Y(n5930));
OR2X1 mul_U17413(.A(n9727), .B(n6057), .Y(dpath_mulcore_ary1_a0_I1_I0_b0n_1));
INVX1 mul_U17414(.A(dpath_mulcore_ary1_a0_I1_I0_b0n_1), .Y(n5931));
AND2X1 mul_U17415(.A(dpath_mulcore_b1[1]), .B(n9724), .Y(n13702));
INVX1 mul_U17416(.A(n13702), .Y(n5932));
AND2X1 mul_U17417(.A(dpath_mulcore_b1[1]), .B(dpath_mulcore_b1[0]), .Y(n13703));
INVX1 mul_U17418(.A(n13703), .Y(n5933));
AND2X1 mul_U17419(.A(dpath_mulcore_b0[1]), .B(n9722), .Y(n13704));
INVX1 mul_U17420(.A(n13704), .Y(n5934));
OR2X1 mul_U17421(.A(n9721), .B(n6058), .Y(dpath_mulcore_ary1_a0_I0_I0_b0n_1));
INVX1 mul_U17422(.A(dpath_mulcore_ary1_a0_I0_I0_b0n_1), .Y(n5935));
AND2X1 mul_U17423(.A(dpath_mulcore_b15[1]), .B(n9752), .Y(n13713));
INVX1 mul_U17424(.A(n13713), .Y(n5936));
AND2X1 mul_U17425(.A(dpath_mulcore_b15[1]), .B(dpath_mulcore_b15[0]), .Y(n13714));
INVX1 mul_U17426(.A(n13714), .Y(n5937));
AND2X1 mul_U17427(.A(dpath_mulcore_b14[1]), .B(n9750), .Y(n13715));
INVX1 mul_U17428(.A(n13715), .Y(n5938));
OR2X1 mul_U17429(.A(n9749), .B(n6059), .Y(dpath_mulcore_ary1_a1_I2_I0_b0n_1));
INVX1 mul_U17430(.A(dpath_mulcore_ary1_a1_I2_I0_b0n_1), .Y(n5939));
AND2X1 mul_U17431(.A(dpath_mulcore_b12[1]), .B(n9746), .Y(n13724));
INVX1 mul_U17432(.A(n13724), .Y(n5940));
AND2X1 mul_U17433(.A(dpath_mulcore_b12[1]), .B(dpath_mulcore_b12[0]), .Y(n13725));
INVX1 mul_U17434(.A(n13725), .Y(n5941));
AND2X1 mul_U17435(.A(dpath_mulcore_b11[1]), .B(n9744), .Y(n13726));
INVX1 mul_U17436(.A(n13726), .Y(n5942));
OR2X1 mul_U17437(.A(n9743), .B(n6060), .Y(dpath_mulcore_ary1_a1_I1_I0_b0n_1));
INVX1 mul_U17438(.A(dpath_mulcore_ary1_a1_I1_I0_b0n_1), .Y(n5943));
AND2X1 mul_U17439(.A(dpath_mulcore_b9[1]), .B(n9740), .Y(n13735));
INVX1 mul_U17440(.A(n13735), .Y(n5944));
AND2X1 mul_U17441(.A(dpath_mulcore_b9[1]), .B(dpath_mulcore_b9[0]), .Y(n13736));
INVX1 mul_U17442(.A(n13736), .Y(n5945));
AND2X1 mul_U17443(.A(dpath_mulcore_b8[1]), .B(n9738), .Y(n13737));
INVX1 mul_U17444(.A(n13737), .Y(n5946));
OR2X1 mul_U17445(.A(n9737), .B(n6061), .Y(dpath_mulcore_ary1_a1_I0_I0_b0n_1));
INVX1 mul_U17446(.A(dpath_mulcore_ary1_a1_I0_I0_b0n_1), .Y(n5947));
AND2X1 mul_U17447(.A(dpath_mulcore_b2[1]), .B(dpath_mulcore_b2[0]), .Y(n17803));
INVX1 mul_U17448(.A(n17803), .Y(n5948));
AND2X1 mul_U17449(.A(dpath_mulcore_b2[1]), .B(n9726), .Y(n17804));
INVX1 mul_U17450(.A(n17804), .Y(n5949));
AND2X1 mul_U17451(.A(dpath_mulcore_b13[1]), .B(dpath_mulcore_b13[0]), .Y(n17805));
INVX1 mul_U17452(.A(n17805), .Y(n5950));
AND2X1 mul_U17453(.A(dpath_mulcore_b13[1]), .B(n9748), .Y(n17806));
INVX1 mul_U17454(.A(n17806), .Y(n5951));
AND2X1 mul_U17455(.A(dpath_mulcore_b10[1]), .B(dpath_mulcore_b10[0]), .Y(n17807));
INVX1 mul_U17456(.A(n17807), .Y(n5952));
AND2X1 mul_U17457(.A(dpath_mulcore_b10[1]), .B(n9742), .Y(n17808));
INVX1 mul_U17458(.A(n17808), .Y(n5953));
OR2X1 mul_U17459(.A(n9733), .B(n6062), .Y(dpath_mulcore_ary1_a0_I2_I0_b0n_1));
INVX1 mul_U17460(.A(dpath_mulcore_ary1_a0_I2_I0_b0n_1), .Y(n5954));
AND2X1 mul_U17461(.A(dpath_mulcore_b6[1]), .B(n9734), .Y(n17810));
INVX1 mul_U17462(.A(n17810), .Y(n5955));
AND2X1 mul_U17463(.A(dpath_mulcore_b7[1]), .B(dpath_mulcore_b7[0]), .Y(n17811));
INVX1 mul_U17464(.A(n17811), .Y(n5956));
AND2X1 mul_U17465(.A(dpath_mulcore_b7[1]), .B(n9736), .Y(n17812));
INVX1 mul_U17466(.A(n17812), .Y(n5957));
AND2X1 mul_U17467(.A(dpath_mulcore_b5[1]), .B(dpath_mulcore_b5[0]), .Y(dpath_mulcore_ary1_a0_p1n_n4));
INVX1 mul_U17468(.A(dpath_mulcore_ary1_a0_p1n_n4), .Y(n5958));
AND2X1 mul_U17469(.A(dpath_mulcore_b5[1]), .B(n9732), .Y(dpath_mulcore_ary1_a0_p1n_n5));
INVX1 mul_U17470(.A(dpath_mulcore_ary1_a0_p1n_n5), .Y(n5959));
INVX1 mul_U17471(.A(dpath_n138), .Y(n5960));
INVX1 mul_U17472(.A(dpath_n147), .Y(n5961));
INVX1 mul_U17473(.A(dpath_n153), .Y(n5962));
INVX1 mul_U17474(.A(dpath_n159), .Y(n5963));
INVX1 mul_U17475(.A(dpath_n165), .Y(n5964));
INVX1 mul_U17476(.A(dpath_n171), .Y(n5965));
INVX1 mul_U17477(.A(dpath_n177), .Y(n5966));
INVX1 mul_U17478(.A(dpath_n183), .Y(n5967));
INVX1 mul_U17479(.A(dpath_n189), .Y(n5968));
INVX1 mul_U17480(.A(dpath_n195), .Y(n5969));
INVX1 mul_U17481(.A(dpath_n201), .Y(n5970));
INVX1 mul_U17482(.A(dpath_n207), .Y(n5971));
INVX1 mul_U17483(.A(dpath_n213), .Y(n5972));
INVX1 mul_U17484(.A(dpath_n219), .Y(n5973));
INVX1 mul_U17485(.A(dpath_n225), .Y(n5974));
INVX1 mul_U17486(.A(dpath_n231), .Y(n5975));
INVX1 mul_U17487(.A(dpath_n237), .Y(n5976));
INVX1 mul_U17488(.A(dpath_n243), .Y(n5977));
INVX1 mul_U17489(.A(dpath_n249), .Y(n5978));
INVX1 mul_U17490(.A(dpath_n255), .Y(n5979));
INVX1 mul_U17491(.A(dpath_n261), .Y(n5980));
INVX1 mul_U17492(.A(dpath_n267), .Y(n5981));
INVX1 mul_U17493(.A(dpath_n273), .Y(n5982));
INVX1 mul_U17494(.A(dpath_n279), .Y(n5983));
INVX1 mul_U17495(.A(dpath_n285), .Y(n5984));
INVX1 mul_U17496(.A(dpath_n291), .Y(n5985));
INVX1 mul_U17497(.A(dpath_n297), .Y(n5986));
INVX1 mul_U17498(.A(dpath_n303), .Y(n5987));
INVX1 mul_U17499(.A(dpath_n309), .Y(n5988));
INVX1 mul_U17500(.A(dpath_n315), .Y(n5989));
INVX1 mul_U17501(.A(dpath_n321), .Y(n5990));
INVX1 mul_U17502(.A(dpath_n327), .Y(n5991));
INVX1 mul_U17503(.A(dpath_n333), .Y(n5992));
INVX1 mul_U17504(.A(dpath_n339), .Y(n5993));
INVX1 mul_U17505(.A(dpath_n345), .Y(n5994));
INVX1 mul_U17506(.A(dpath_n351), .Y(n5995));
INVX1 mul_U17507(.A(dpath_n357), .Y(n5996));
INVX1 mul_U17508(.A(dpath_n363), .Y(n5997));
INVX1 mul_U17509(.A(dpath_n369), .Y(n5998));
INVX1 mul_U17510(.A(dpath_n375), .Y(n5999));
INVX1 mul_U17511(.A(dpath_n381), .Y(n6000));
INVX1 mul_U17512(.A(dpath_n387), .Y(n6001));
INVX1 mul_U17513(.A(dpath_n393), .Y(n6002));
INVX1 mul_U17514(.A(dpath_n399), .Y(n6003));
INVX1 mul_U17515(.A(dpath_n405), .Y(n6004));
INVX1 mul_U17516(.A(dpath_n411), .Y(n6005));
INVX1 mul_U17517(.A(dpath_n417), .Y(n6006));
INVX1 mul_U17518(.A(dpath_n423), .Y(n6007));
INVX1 mul_U17519(.A(dpath_n429), .Y(n6008));
INVX1 mul_U17520(.A(dpath_n435), .Y(n6009));
INVX1 mul_U17521(.A(dpath_n441), .Y(n6010));
INVX1 mul_U17522(.A(dpath_n447), .Y(n6011));
INVX1 mul_U17523(.A(dpath_n453), .Y(n6012));
INVX1 mul_U17524(.A(dpath_n459), .Y(n6013));
INVX1 mul_U17525(.A(dpath_n465), .Y(n6014));
INVX1 mul_U17526(.A(dpath_n471), .Y(n6015));
INVX1 mul_U17527(.A(dpath_n477), .Y(n6016));
INVX1 mul_U17528(.A(dpath_n483), .Y(n6017));
INVX1 mul_U17529(.A(dpath_n489), .Y(n6018));
INVX1 mul_U17530(.A(dpath_n495), .Y(n6019));
INVX1 mul_U17531(.A(dpath_n501), .Y(n6020));
INVX1 mul_U17532(.A(dpath_n507), .Y(n6021));
INVX1 mul_U17533(.A(dpath_n513), .Y(n6022));
INVX1 mul_U17534(.A(dpath_n519), .Y(n6023));
INVX1 mul_U17535(.A(dpath_n654), .Y(n6024));
INVX1 mul_U17536(.A(dpath_n680), .Y(n6025));
INVX1 mul_U17537(.A(dpath_n706), .Y(n6026));
INVX1 mul_U17538(.A(dpath_n732), .Y(n6027));
INVX1 mul_U17539(.A(dpath_n758), .Y(n6028));
INVX1 mul_U17540(.A(dpath_n784), .Y(n6029));
INVX1 mul_U17541(.A(dpath_n810), .Y(n6030));
INVX1 mul_U17542(.A(dpath_n832), .Y(n6031));
INVX1 mul_U17543(.A(dpath_n838), .Y(n6032));
INVX1 mul_U17544(.A(dpath_n844), .Y(n6033));
INVX1 mul_U17545(.A(dpath_n850), .Y(n6034));
INVX1 mul_U17546(.A(dpath_n856), .Y(n6035));
INVX1 mul_U17547(.A(dpath_n862), .Y(n6036));
INVX1 mul_U17548(.A(dpath_n868), .Y(n6037));
INVX1 mul_U17549(.A(dpath_n874), .Y(n6038));
INVX1 mul_U17550(.A(dpath_n880), .Y(n6039));
INVX1 mul_U17551(.A(dpath_n886), .Y(n6040));
INVX1 mul_U17552(.A(dpath_n892), .Y(n6041));
INVX1 mul_U17553(.A(dpath_n898), .Y(n6042));
INVX1 mul_U17554(.A(dpath_n904), .Y(n6043));
INVX1 mul_U17555(.A(dpath_n910), .Y(n6044));
INVX1 mul_U17556(.A(dpath_n916), .Y(n6045));
INVX1 mul_U17557(.A(dpath_n922), .Y(n6046));
INVX1 mul_U17558(.A(dpath_n928), .Y(n6047));
INVX1 mul_U17559(.A(dpath_n934), .Y(n6048));
INVX1 mul_U17560(.A(dpath_n940), .Y(n6049));
INVX1 mul_U17561(.A(dpath_n946), .Y(n6050));
INVX1 mul_U17562(.A(dpath_n952), .Y(n6051));
INVX1 mul_U17563(.A(dpath_n958), .Y(n6052));
INVX1 mul_U17564(.A(dpath_n964), .Y(n6053));
INVX1 mul_U17565(.A(dpath_n970), .Y(n6054));
INVX1 mul_U17566(.A(dpath_n976), .Y(n6055));
AND2X1 mul_U17567(.A(dpath_acc_reg[131]), .B(dpath_acc_reg[130]), .Y(n10599));
INVX1 mul_U17568(.A(n10599), .Y(n6056));
AND2X1 mul_U17569(.A(dpath_mulcore_b3[1]), .B(dpath_mulcore_b3[0]), .Y(n13694));
INVX1 mul_U17570(.A(n13694), .Y(n6057));
AND2X1 mul_U17571(.A(dpath_mulcore_b0[1]), .B(dpath_mulcore_b0[0]), .Y(n13705));
INVX1 mul_U17572(.A(n13705), .Y(n6058));
AND2X1 mul_U17573(.A(dpath_mulcore_b14[1]), .B(dpath_mulcore_b14[0]), .Y(n13716));
INVX1 mul_U17574(.A(n13716), .Y(n6059));
AND2X1 mul_U17575(.A(dpath_mulcore_b11[1]), .B(dpath_mulcore_b11[0]), .Y(n13727));
INVX1 mul_U17576(.A(n13727), .Y(n6060));
AND2X1 mul_U17577(.A(dpath_mulcore_b8[1]), .B(dpath_mulcore_b8[0]), .Y(n13738));
INVX1 mul_U17578(.A(n13738), .Y(n6061));
AND2X1 mul_U17579(.A(dpath_mulcore_b6[1]), .B(dpath_mulcore_b6[0]), .Y(n17809));
INVX1 mul_U17580(.A(n17809), .Y(n6062));
INVX1 mul_U17581(.A(control_n14), .Y(n6063));
AND2X1 mul_U17582(.A(dpath_mulcore_b16), .B(n10032), .Y(dpath_mulcore_ary1_a1_I2_I2_p2_l_67));
AND2X1 mul_U17583(.A(dpath_mulcore_b16), .B(n10031), .Y(dpath_mulcore_ary1_a1_I2_I2_p2_l_66));
AND2X1 mul_U17584(.A(dpath_mulcore_b16), .B(n10030), .Y(dpath_mulcore_ary1_a1_I2_I2_p2_l_65));
AND2X1 mul_U17585(.A(dpath_mulcore_b16), .B(n10029), .Y(dpath_mulcore_ary1_a1_I2_I2_p2_l_64));
AND2X1 mul_U17586(.A(dpath_mulcore_b16), .B(n10028), .Y(dpath_mulcore_ary1_a1_I2_p2_l[63]));
AND2X1 mul_U17587(.A(dpath_mulcore_b16), .B(n10024), .Y(dpath_mulcore_ary1_a1_I2_p2_l[62]));
AND2X1 mul_U17588(.A(dpath_mulcore_b16), .B(n10021), .Y(dpath_mulcore_ary1_a1_I2_p2_l[61]));
AND2X1 mul_U17589(.A(dpath_mulcore_b16), .B(n10018), .Y(dpath_mulcore_ary1_a1_I2_p2_l[60]));
AND2X1 mul_U17590(.A(dpath_mulcore_b16), .B(n10015), .Y(dpath_mulcore_ary1_a1_I2_p2_l[59]));
AND2X1 mul_U17591(.A(dpath_mulcore_b16), .B(n10012), .Y(dpath_mulcore_ary1_a1_I2_p2_l[58]));
AND2X1 mul_U17592(.A(dpath_mulcore_b16), .B(n10009), .Y(dpath_mulcore_ary1_a1_I2_p2_l[57]));
AND2X1 mul_U17593(.A(dpath_mulcore_b16), .B(n10006), .Y(dpath_mulcore_ary1_a1_I2_p2_l[56]));
AND2X1 mul_U17594(.A(dpath_mulcore_b16), .B(n10004), .Y(dpath_mulcore_ary1_a1_I2_p2_l[55]));
AND2X1 mul_U17595(.A(dpath_mulcore_b16), .B(n10002), .Y(dpath_mulcore_ary1_a1_I2_p2_l[54]));
AND2X1 mul_U17596(.A(dpath_mulcore_b16), .B(n10000), .Y(dpath_mulcore_ary1_a1_I2_p2_l[53]));
AND2X1 mul_U17597(.A(dpath_mulcore_b16), .B(n9998), .Y(dpath_mulcore_ary1_a1_I2_p2_l[52]));
AND2X1 mul_U17598(.A(dpath_mulcore_b16), .B(n9996), .Y(dpath_mulcore_ary1_a1_I2_p2_l[51]));
AND2X1 mul_U17599(.A(dpath_mulcore_b16), .B(n9993), .Y(dpath_mulcore_ary1_a1_I2_p2_l[50]));
AND2X1 mul_U17600(.A(dpath_mulcore_b16), .B(n9990), .Y(dpath_mulcore_ary1_a1_I2_p2_l[49]));
AND2X1 mul_U17601(.A(dpath_mulcore_b16), .B(n9987), .Y(dpath_mulcore_ary1_a1_I2_p2_l[48]));
AND2X1 mul_U17602(.A(dpath_mulcore_b16), .B(n9984), .Y(dpath_mulcore_ary1_a1_I2_p2_l[47]));
AND2X1 mul_U17603(.A(dpath_mulcore_b16), .B(n9981), .Y(dpath_mulcore_ary1_a1_I2_p2_l[46]));
AND2X1 mul_U17604(.A(dpath_mulcore_b16), .B(n9978), .Y(dpath_mulcore_ary1_a1_I2_p2_l[45]));
AND2X1 mul_U17605(.A(dpath_mulcore_b16), .B(n9975), .Y(dpath_mulcore_ary1_a1_I2_p2_l[44]));
AND2X1 mul_U17606(.A(dpath_mulcore_b16), .B(n9972), .Y(dpath_mulcore_ary1_a1_I2_p2_l[43]));
AND2X1 mul_U17607(.A(dpath_mulcore_b16), .B(n9969), .Y(dpath_mulcore_ary1_a1_I2_p2_l[42]));
AND2X1 mul_U17608(.A(dpath_mulcore_b16), .B(n9966), .Y(dpath_mulcore_ary1_a1_I2_p2_l[41]));
AND2X1 mul_U17609(.A(dpath_mulcore_b16), .B(n9963), .Y(dpath_mulcore_ary1_a1_I2_p2_l[40]));
AND2X1 mul_U17610(.A(dpath_mulcore_b16), .B(n9960), .Y(dpath_mulcore_ary1_a1_I2_p2_l[39]));
AND2X1 mul_U17611(.A(dpath_mulcore_b16), .B(n9957), .Y(dpath_mulcore_ary1_a1_I2_p2_l[38]));
AND2X1 mul_U17612(.A(dpath_mulcore_b16), .B(n9954), .Y(dpath_mulcore_ary1_a1_I2_p2_l[37]));
AND2X1 mul_U17613(.A(dpath_mulcore_b16), .B(n9951), .Y(dpath_mulcore_ary1_a1_I2_p2_l[36]));
AND2X1 mul_U17614(.A(dpath_mulcore_b16), .B(n9948), .Y(dpath_mulcore_ary1_a1_I2_p2_l[35]));
AND2X1 mul_U17615(.A(dpath_mulcore_b16), .B(n9945), .Y(dpath_mulcore_ary1_a1_I2_p2_l[34]));
AND2X1 mul_U17616(.A(dpath_mulcore_b16), .B(n9942), .Y(dpath_mulcore_ary1_a1_I2_p2_l[33]));
AND2X1 mul_U17617(.A(dpath_mulcore_b16), .B(n9939), .Y(dpath_mulcore_ary1_a1_I2_p2_l[32]));
AND2X1 mul_U17618(.A(dpath_mulcore_b16), .B(n9936), .Y(dpath_mulcore_ary1_a1_I2_p2_l[31]));
AND2X1 mul_U17619(.A(dpath_mulcore_b16), .B(n9933), .Y(dpath_mulcore_ary1_a1_I2_p2_l[30]));
AND2X1 mul_U17620(.A(dpath_mulcore_b16), .B(n9930), .Y(dpath_mulcore_ary1_a1_I2_p2_l[29]));
AND2X1 mul_U17621(.A(dpath_mulcore_b16), .B(n9927), .Y(dpath_mulcore_ary1_a1_I2_p2_l[28]));
AND2X1 mul_U17622(.A(dpath_mulcore_b16), .B(n9924), .Y(dpath_mulcore_ary1_a1_I2_p2_l[27]));
AND2X1 mul_U17623(.A(dpath_mulcore_b16), .B(n9921), .Y(dpath_mulcore_ary1_a1_I2_p2_l[26]));
AND2X1 mul_U17624(.A(dpath_mulcore_b16), .B(n9918), .Y(dpath_mulcore_ary1_a1_I2_p2_l[25]));
AND2X1 mul_U17625(.A(dpath_mulcore_b16), .B(n9915), .Y(dpath_mulcore_ary1_a1_I2_p2_l[24]));
AND2X1 mul_U17626(.A(dpath_mulcore_b16), .B(n9912), .Y(dpath_mulcore_ary1_a1_I2_p2_l[23]));
AND2X1 mul_U17627(.A(dpath_mulcore_b16), .B(n9909), .Y(dpath_mulcore_ary1_a1_I2_p2_l[22]));
AND2X1 mul_U17628(.A(dpath_mulcore_b16), .B(n9906), .Y(dpath_mulcore_ary1_a1_I2_p2_l[21]));
AND2X1 mul_U17629(.A(dpath_mulcore_b16), .B(n9903), .Y(dpath_mulcore_ary1_a1_I2_p2_l[20]));
AND2X1 mul_U17630(.A(dpath_mulcore_b16), .B(n9900), .Y(dpath_mulcore_ary1_a1_I2_p2_l[19]));
AND2X1 mul_U17631(.A(dpath_mulcore_b16), .B(n9897), .Y(dpath_mulcore_ary1_a1_I2_p2_l[18]));
AND2X1 mul_U17632(.A(dpath_mulcore_b16), .B(n9894), .Y(dpath_mulcore_ary1_a1_I2_p2_l[17]));
AND2X1 mul_U17633(.A(dpath_mulcore_b16), .B(n9891), .Y(dpath_mulcore_ary1_a1_I2_p2_l[16]));
AND2X1 mul_U17634(.A(dpath_mulcore_b16), .B(n9888), .Y(dpath_mulcore_ary1_a1_I2_p2_l[15]));
AND2X1 mul_U17635(.A(dpath_mulcore_b16), .B(n9885), .Y(dpath_mulcore_ary1_a1_I2_p2_l[14]));
AND2X1 mul_U17636(.A(dpath_mulcore_b16), .B(n9882), .Y(dpath_mulcore_ary1_a1_I2_p2_l[13]));
AND2X1 mul_U17637(.A(dpath_mulcore_b16), .B(n9879), .Y(dpath_mulcore_ary1_a1_I2_p2_l[12]));
AND2X1 mul_U17638(.A(dpath_mulcore_b16), .B(n9876), .Y(dpath_mulcore_ary1_a1_I2_p2_l[11]));
AND2X1 mul_U17639(.A(dpath_mulcore_b16), .B(n9873), .Y(dpath_mulcore_ary1_a1_I2_p2_l[10]));
AND2X1 mul_U17640(.A(dpath_mulcore_b16), .B(n9870), .Y(dpath_mulcore_ary1_a1_I2_p2_l[9]));
AND2X1 mul_U17641(.A(dpath_mulcore_b16), .B(n9867), .Y(dpath_mulcore_ary1_a1_I2_p2_l[8]));
AND2X1 mul_U17642(.A(dpath_mulcore_b16), .B(n9864), .Y(dpath_mulcore_ary1_a1_I2_p2_l[7]));
AND2X1 mul_U17643(.A(dpath_mulcore_b16), .B(n9861), .Y(dpath_mulcore_ary1_a1_I2_p2_l[6]));
AND2X1 mul_U17644(.A(dpath_mulcore_b16), .B(n9858), .Y(dpath_mulcore_ary1_a1_I2_p2_l[5]));
AND2X1 mul_U17645(.A(dpath_mulcore_b16), .B(n9855), .Y(dpath_mulcore_ary1_a1_I2_p2_l[4]));
AND2X1 mul_U17646(.A(n7420), .B(n8389), .Y(n13745));
AND2X1 mul_U17647(.A(n7421), .B(n8390), .Y(n13747));
AND2X1 mul_U17648(.A(n7422), .B(n8391), .Y(n13749));
AND2X1 mul_U17649(.A(n7423), .B(n8392), .Y(n13751));
AND2X1 mul_U17650(.A(n7424), .B(n8393), .Y(n13753));
AND2X1 mul_U17651(.A(n7425), .B(n8394), .Y(n13755));
AND2X1 mul_U17652(.A(n7426), .B(n8395), .Y(n13757));
AND2X1 mul_U17653(.A(n7427), .B(n8396), .Y(n13759));
AND2X1 mul_U17654(.A(n7428), .B(n8397), .Y(n13761));
AND2X1 mul_U17655(.A(n7429), .B(n8398), .Y(n13763));
AND2X1 mul_U17656(.A(n7430), .B(n8399), .Y(n13765));
AND2X1 mul_U17657(.A(n7431), .B(n8400), .Y(n13767));
AND2X1 mul_U17658(.A(n7432), .B(n8401), .Y(n13769));
AND2X1 mul_U17659(.A(n7433), .B(n8402), .Y(n13771));
AND2X1 mul_U17660(.A(n7434), .B(n8403), .Y(n13773));
AND2X1 mul_U17661(.A(n7435), .B(n8404), .Y(n13775));
AND2X1 mul_U17662(.A(n7436), .B(n8405), .Y(n13777));
AND2X1 mul_U17663(.A(n7437), .B(n8406), .Y(n13779));
AND2X1 mul_U17664(.A(n7438), .B(n8407), .Y(n13781));
AND2X1 mul_U17665(.A(n7439), .B(n8408), .Y(n13783));
AND2X1 mul_U17666(.A(n7440), .B(n8409), .Y(n13785));
AND2X1 mul_U17667(.A(n7441), .B(n8410), .Y(n13787));
AND2X1 mul_U17668(.A(n7442), .B(n8411), .Y(n13789));
AND2X1 mul_U17669(.A(n7443), .B(n8412), .Y(n13791));
AND2X1 mul_U17670(.A(n7444), .B(n8413), .Y(n13793));
AND2X1 mul_U17671(.A(n7445), .B(n8414), .Y(n13795));
AND2X1 mul_U17672(.A(n7446), .B(n8415), .Y(n13797));
AND2X1 mul_U17673(.A(n7447), .B(n8416), .Y(n13799));
AND2X1 mul_U17674(.A(n7448), .B(n8417), .Y(n13801));
AND2X1 mul_U17675(.A(n7449), .B(n8418), .Y(n13803));
AND2X1 mul_U17676(.A(n7450), .B(n8419), .Y(n13805));
AND2X1 mul_U17677(.A(n7451), .B(n8420), .Y(n13807));
AND2X1 mul_U17678(.A(n7452), .B(n8421), .Y(n13809));
AND2X1 mul_U17679(.A(n7453), .B(n8422), .Y(n13811));
AND2X1 mul_U17680(.A(n7454), .B(n8423), .Y(n13813));
AND2X1 mul_U17681(.A(n7455), .B(n8424), .Y(n13815));
AND2X1 mul_U17682(.A(n7456), .B(n8425), .Y(n13817));
AND2X1 mul_U17683(.A(n7457), .B(n8426), .Y(n13819));
AND2X1 mul_U17684(.A(n7458), .B(n8427), .Y(n13821));
AND2X1 mul_U17685(.A(n7459), .B(n8428), .Y(n13823));
AND2X1 mul_U17686(.A(n7460), .B(n8429), .Y(n13825));
AND2X1 mul_U17687(.A(n7461), .B(n8430), .Y(n13827));
AND2X1 mul_U17688(.A(n7462), .B(n8431), .Y(n13829));
AND2X1 mul_U17689(.A(n7463), .B(n8432), .Y(n13831));
AND2X1 mul_U17690(.A(n7464), .B(n8433), .Y(n13833));
AND2X1 mul_U17691(.A(n7465), .B(n8434), .Y(n13835));
AND2X1 mul_U17692(.A(n7466), .B(n8435), .Y(n13837));
AND2X1 mul_U17693(.A(n7467), .B(n8436), .Y(n13839));
AND2X1 mul_U17694(.A(n7468), .B(n8437), .Y(n13841));
AND2X1 mul_U17695(.A(n7469), .B(n8438), .Y(n13843));
AND2X1 mul_U17696(.A(n7470), .B(n8439), .Y(n13845));
AND2X1 mul_U17697(.A(n7471), .B(n8440), .Y(n13847));
AND2X1 mul_U17698(.A(n7472), .B(n8441), .Y(n13849));
AND2X1 mul_U17699(.A(n7473), .B(n8442), .Y(n13851));
AND2X1 mul_U17700(.A(n7474), .B(n8443), .Y(n13853));
AND2X1 mul_U17701(.A(n7475), .B(n8444), .Y(n13855));
AND2X1 mul_U17702(.A(n7476), .B(n8445), .Y(n13857));
AND2X1 mul_U17703(.A(n7477), .B(n8446), .Y(n13859));
AND2X1 mul_U17704(.A(n7478), .B(n8447), .Y(n13861));
AND2X1 mul_U17705(.A(n7799), .B(n9480), .Y(n14790));
AND2X1 mul_U17706(.A(n7926), .B(n9482), .Y(n14798));
AND2X1 mul_U17707(.A(n6075), .B(n9699), .Y(n14897));
AND2X1 mul_U17708(.A(n9684), .B(dpath_areg[0]), .Y(n14968));
AND2X1 mul_U17709(.A(dpath_mulcore_ps[47]), .B(dpath_mulcore_pc[46]), .Y(n16044));
AND2X1 mul_U17710(.A(dpath_mulcore_a0c[19]), .B(dpath_mulcore_a0s[20]), .Y(n16368));
AND2X1 mul_U17711(.A(n8269), .B(dpath_mulcore_array2_s3[15]), .Y(n16563));
AND2X1 mul_U17712(.A(n7417), .B(n9483), .Y(n16569));
AND2X1 mul_U17713(.A(n7418), .B(n8977), .Y(n16571));
AND2X1 mul_U17714(.A(n7419), .B(n8388), .Y(n16573));
AND2X1 mul_U17715(.A(n7481), .B(n9476), .Y(n16580));
AND2X1 mul_U17716(.A(n9484), .B(dpath_mulcore_ary1_a0_s_2[75]), .Y(n16588));
AND2X1 mul_U17717(.A(dpath_mulcore_ary1_a0_I1_I2_net073), .B(dpath_mulcore_ary1_a0_s_2[74]), .Y(n16592));
AND2X1 mul_U17718(.A(dpath_mulcore_ary1_a0_s1[67]), .B(dpath_mulcore_ary1_a0_s_2[73]), .Y(n16596));
AND2X1 mul_U17719(.A(dpath_mulcore_ary1_a0_s1[66]), .B(dpath_mulcore_ary1_a0_s_2[72]), .Y(n16600));
AND2X1 mul_U17720(.A(n9485), .B(dpath_mulcore_ary1_a1_s_2[75]), .Y(n17032));
AND2X1 mul_U17721(.A(dpath_mulcore_ary1_a1_I1_I2_net073), .B(dpath_mulcore_ary1_a1_s_2[74]), .Y(n17036));
AND2X1 mul_U17722(.A(dpath_mulcore_ary1_a1_s1[67]), .B(dpath_mulcore_ary1_a1_s_2[73]), .Y(n17040));
AND2X1 mul_U17723(.A(dpath_mulcore_ary1_a1_s1[66]), .B(dpath_mulcore_ary1_a1_s_2[72]), .Y(n17044));
AND2X1 mul_U17724(.A(n9100), .B(dpath_mulcore_array2_s1[67]), .Y(n17471));
AND2X1 mul_U17725(.A(dpath_mulcore_array2_s2[20]), .B(n10033), .Y(n17800));
AND2X1 mul_U17726(.A(dpath_mulcore_a1sum[6]), .B(n9531), .Y(n18139));
AND2X1 mul_U17727(.A(dpath_mulcore_cyc2), .B(n9531), .Y(n18140));
AND2X1 mul_U17728(.A(n6168), .B(n9531), .Y(n18141));
AND2X1 mul_U17729(.A(dpath_mulcore_a1sum[79]), .B(n9531), .Y(n18142));
AND2X1 mul_U17730(.A(dpath_mulcore_a1sum[78]), .B(n9531), .Y(n18143));
AND2X1 mul_U17731(.A(dpath_mulcore_a1sum[77]), .B(n9531), .Y(n18144));
AND2X1 mul_U17732(.A(dpath_mulcore_a1sum[5]), .B(n9531), .Y(n18145));
AND2X1 mul_U17733(.A(dpath_mulcore_a1sum[76]), .B(n9531), .Y(n18146));
AND2X1 mul_U17734(.A(dpath_mulcore_a1sum[75]), .B(n9531), .Y(n18147));
AND2X1 mul_U17735(.A(dpath_mulcore_a1sum[74]), .B(n9532), .Y(n18148));
AND2X1 mul_U17736(.A(dpath_mulcore_a1sum[73]), .B(n9520), .Y(n18149));
AND2X1 mul_U17737(.A(dpath_mulcore_a1sum[72]), .B(n9517), .Y(n18150));
AND2X1 mul_U17738(.A(dpath_mulcore_a1sum[71]), .B(n9517), .Y(n18151));
AND2X1 mul_U17739(.A(dpath_mulcore_a1sum[70]), .B(n9517), .Y(n18152));
AND2X1 mul_U17740(.A(dpath_mulcore_a1sum[69]), .B(n9517), .Y(n18153));
AND2X1 mul_U17741(.A(dpath_mulcore_a1sum[68]), .B(n9517), .Y(n18154));
AND2X1 mul_U17742(.A(dpath_mulcore_a1sum[67]), .B(n9517), .Y(n18155));
AND2X1 mul_U17743(.A(dpath_mulcore_a1sum[4]), .B(n9517), .Y(n18156));
AND2X1 mul_U17744(.A(dpath_mulcore_a1sum[66]), .B(n9517), .Y(n18157));
AND2X1 mul_U17745(.A(dpath_mulcore_a1sum[65]), .B(n9517), .Y(n18158));
AND2X1 mul_U17746(.A(dpath_mulcore_a1sum[64]), .B(n9517), .Y(n18159));
AND2X1 mul_U17747(.A(dpath_mulcore_a1sum[63]), .B(n9518), .Y(n18160));
AND2X1 mul_U17748(.A(dpath_mulcore_a1sum[62]), .B(n9518), .Y(n18161));
AND2X1 mul_U17749(.A(dpath_mulcore_a1sum[61]), .B(n9518), .Y(n18162));
AND2X1 mul_U17750(.A(dpath_mulcore_a1sum[60]), .B(n9518), .Y(n18163));
AND2X1 mul_U17751(.A(dpath_mulcore_a1sum[59]), .B(n9518), .Y(n18164));
AND2X1 mul_U17752(.A(dpath_mulcore_a1sum[58]), .B(n9518), .Y(n18165));
AND2X1 mul_U17753(.A(dpath_mulcore_a1sum[57]), .B(n9518), .Y(n18166));
AND2X1 mul_U17754(.A(dpath_mulcore_a1sum[3]), .B(n9518), .Y(n18167));
AND2X1 mul_U17755(.A(dpath_mulcore_a1sum[56]), .B(n9518), .Y(n18168));
AND2X1 mul_U17756(.A(dpath_mulcore_a1sum[55]), .B(n9518), .Y(n18169));
AND2X1 mul_U17757(.A(dpath_mulcore_a1sum[54]), .B(n9518), .Y(n18170));
AND2X1 mul_U17758(.A(dpath_mulcore_a1sum[53]), .B(n9518), .Y(n18171));
AND2X1 mul_U17759(.A(dpath_mulcore_a1sum[52]), .B(n9518), .Y(n18172));
AND2X1 mul_U17760(.A(dpath_mulcore_a1sum[51]), .B(n9496), .Y(n18173));
AND2X1 mul_U17761(.A(dpath_mulcore_a1sum[50]), .B(n9496), .Y(n18174));
AND2X1 mul_U17762(.A(dpath_mulcore_a1sum[49]), .B(n9496), .Y(n18175));
AND2X1 mul_U17763(.A(dpath_mulcore_a1sum[48]), .B(n9528), .Y(n18176));
AND2X1 mul_U17764(.A(dpath_mulcore_a1sum[47]), .B(n9525), .Y(n18177));
AND2X1 mul_U17765(.A(dpath_mulcore_a1sum[2]), .B(n9526), .Y(n18178));
AND2X1 mul_U17766(.A(dpath_mulcore_a1sum[46]), .B(n9529), .Y(n18179));
AND2X1 mul_U17767(.A(dpath_mulcore_a1sum[45]), .B(n9531), .Y(n18180));
AND2X1 mul_U17768(.A(dpath_mulcore_a1sum[44]), .B(n9536), .Y(n18181));
AND2X1 mul_U17769(.A(dpath_mulcore_a1sum[43]), .B(n9537), .Y(n18182));
AND2X1 mul_U17770(.A(dpath_mulcore_a1sum[42]), .B(n9538), .Y(n18183));
AND2X1 mul_U17771(.A(dpath_mulcore_a1sum[41]), .B(n9499), .Y(n18184));
AND2X1 mul_U17772(.A(dpath_mulcore_a1sum[40]), .B(n9493), .Y(n18185));
AND2X1 mul_U17773(.A(dpath_mulcore_a1sum[39]), .B(n9519), .Y(n18186));
AND2X1 mul_U17774(.A(dpath_mulcore_a1sum[38]), .B(n9519), .Y(n18187));
AND2X1 mul_U17775(.A(dpath_mulcore_a1sum[37]), .B(n9519), .Y(n18188));
AND2X1 mul_U17776(.A(dpath_mulcore_a1sum[1]), .B(n9519), .Y(n18189));
AND2X1 mul_U17777(.A(dpath_mulcore_a1sum[36]), .B(n9519), .Y(n18190));
AND2X1 mul_U17778(.A(dpath_mulcore_a1sum[35]), .B(n9519), .Y(n18191));
AND2X1 mul_U17779(.A(dpath_mulcore_a1sum[34]), .B(n9519), .Y(n18192));
AND2X1 mul_U17780(.A(dpath_mulcore_a1sum[33]), .B(n9519), .Y(n18193));
AND2X1 mul_U17781(.A(dpath_mulcore_a1sum[32]), .B(n9519), .Y(n18194));
AND2X1 mul_U17782(.A(dpath_mulcore_a1sum[31]), .B(n9519), .Y(n18195));
AND2X1 mul_U17783(.A(dpath_mulcore_a1sum[30]), .B(n9519), .Y(n18196));
AND2X1 mul_U17784(.A(dpath_mulcore_a1sum[29]), .B(n9519), .Y(n18197));
AND2X1 mul_U17785(.A(dpath_mulcore_a1sum[28]), .B(n9519), .Y(n18198));
AND2X1 mul_U17786(.A(dpath_mulcore_a1sum[27]), .B(n9520), .Y(n18199));
AND2X1 mul_U17787(.A(dpath_mulcore_a1sum[0]), .B(n9520), .Y(n18200));
AND2X1 mul_U17788(.A(dpath_mulcore_a1sum[26]), .B(n9520), .Y(n18201));
AND2X1 mul_U17789(.A(dpath_mulcore_a1sum[25]), .B(n9520), .Y(n18202));
AND2X1 mul_U17790(.A(dpath_mulcore_a1sum[24]), .B(n9520), .Y(n18203));
AND2X1 mul_U17791(.A(dpath_mulcore_a1sum[23]), .B(n9520), .Y(n18204));
AND2X1 mul_U17792(.A(dpath_mulcore_a1sum[22]), .B(n9520), .Y(n18205));
AND2X1 mul_U17793(.A(dpath_mulcore_a1sum[21]), .B(n9520), .Y(n18206));
AND2X1 mul_U17794(.A(dpath_mulcore_a1sum[20]), .B(n9520), .Y(n18207));
AND2X1 mul_U17795(.A(dpath_mulcore_a1sum[19]), .B(n9520), .Y(n18208));
AND2X1 mul_U17796(.A(dpath_mulcore_a1sum[18]), .B(n9520), .Y(n18209));
AND2X1 mul_U17797(.A(dpath_mulcore_a1sum[17]), .B(n9520), .Y(n18210));
AND2X1 mul_U17798(.A(dpath_mulcore_a1sum[16]), .B(n9521), .Y(n18211));
AND2X1 mul_U17799(.A(dpath_mulcore_a1sum[15]), .B(n9521), .Y(n18212));
AND2X1 mul_U17800(.A(dpath_mulcore_a1sum[14]), .B(n9521), .Y(n18213));
AND2X1 mul_U17801(.A(dpath_mulcore_a1sum[13]), .B(n9521), .Y(n18214));
AND2X1 mul_U17802(.A(dpath_mulcore_a1sum[12]), .B(n9521), .Y(n18215));
AND2X1 mul_U17803(.A(dpath_mulcore_ary1_a1_sc3_11__z), .B(n9521), .Y(n18216));
AND2X1 mul_U17804(.A(dpath_mulcore_a1sum[10]), .B(n9521), .Y(n18217));
AND2X1 mul_U17805(.A(dpath_mulcore_a1sum[9]), .B(n9521), .Y(n18218));
AND2X1 mul_U17806(.A(dpath_mulcore_a1sum[8]), .B(n9521), .Y(n18219));
AND2X1 mul_U17807(.A(dpath_mulcore_a1sum[7]), .B(n9521), .Y(n18220));
AND2X1 mul_U17808(.A(n14782), .B(n9518), .Y(n18223));
AND2X1 mul_U17809(.A(dpath_mulcore_a1cout[79]), .B(n9496), .Y(n18224));
AND2X1 mul_U17810(.A(dpath_mulcore_a1cout[78]), .B(n9519), .Y(n18225));
AND2X1 mul_U17811(.A(dpath_mulcore_a1cout[7]), .B(n9535), .Y(n18244));
AND2X1 mul_U17812(.A(dpath_mulcore_a1cout[6]), .B(n9528), .Y(n18255));
AND2X1 mul_U17813(.A(dpath_mulcore_a1cout[5]), .B(n9528), .Y(n18266));
AND2X1 mul_U17814(.A(dpath_mulcore_a1cout[4]), .B(n9529), .Y(n18277));
AND2X1 mul_U17815(.A(n17466), .B(n9531), .Y(n18297));
AND2X1 mul_U17816(.A(dpath_mul_op2_d[38]), .B(n9510), .Y(n18303));
AND2X1 mul_U17817(.A(dpath_mul_op2_d[37]), .B(n9510), .Y(n18304));
AND2X1 mul_U17818(.A(dpath_mul_op2_d[36]), .B(n9510), .Y(n18305));
AND2X1 mul_U17819(.A(dpath_mul_op2_d[35]), .B(n9533), .Y(n18306));
AND2X1 mul_U17820(.A(dpath_mul_op2_d[34]), .B(n9525), .Y(n18307));
AND2X1 mul_U17821(.A(dpath_mul_op2_d[33]), .B(n9525), .Y(n18308));
AND2X1 mul_U17822(.A(dpath_mul_op2_d[63]), .B(n9525), .Y(n18309));
AND2X1 mul_U17823(.A(dpath_mul_op2_d[62]), .B(n9525), .Y(n18310));
AND2X1 mul_U17824(.A(dpath_mul_op2_d[61]), .B(n9525), .Y(n18311));
AND2X1 mul_U17825(.A(dpath_mul_op2_d[60]), .B(n9525), .Y(n18312));
AND2X1 mul_U17826(.A(dpath_mul_op2_d[59]), .B(n9525), .Y(n18313));
AND2X1 mul_U17827(.A(dpath_mul_op2_d[32]), .B(n9525), .Y(n18314));
AND2X1 mul_U17828(.A(dpath_mul_op2_d[58]), .B(n9525), .Y(n18315));
AND2X1 mul_U17829(.A(dpath_mul_op2_d[57]), .B(n9525), .Y(n18316));
AND2X1 mul_U17830(.A(dpath_mul_op2_d[56]), .B(n9525), .Y(n18317));
AND2X1 mul_U17831(.A(dpath_mul_op2_d[55]), .B(n9526), .Y(n18318));
AND2X1 mul_U17832(.A(dpath_mul_op2_d[54]), .B(n9526), .Y(n18319));
AND2X1 mul_U17833(.A(dpath_mul_op2_d[53]), .B(n9526), .Y(n18320));
AND2X1 mul_U17834(.A(dpath_mul_op2_d[52]), .B(n9526), .Y(n18321));
AND2X1 mul_U17835(.A(dpath_mul_op2_d[51]), .B(n9526), .Y(n18322));
AND2X1 mul_U17836(.A(dpath_mul_op2_d[50]), .B(n9526), .Y(n18323));
AND2X1 mul_U17837(.A(dpath_mul_op2_d[49]), .B(n9526), .Y(n18324));
AND2X1 mul_U17838(.A(dpath_mul_op2_d[48]), .B(n9526), .Y(n18325));
AND2X1 mul_U17839(.A(dpath_mul_op2_d[47]), .B(n9526), .Y(n18326));
AND2X1 mul_U17840(.A(dpath_mul_op2_d[46]), .B(n9526), .Y(n18327));
AND2X1 mul_U17841(.A(dpath_mul_op2_d[45]), .B(n9526), .Y(n18328));
AND2X1 mul_U17842(.A(dpath_mul_op2_d[44]), .B(n9526), .Y(n18329));
AND2X1 mul_U17843(.A(dpath_mul_op2_d[43]), .B(n9526), .Y(n18330));
AND2X1 mul_U17844(.A(dpath_mul_op2_d[42]), .B(n9520), .Y(n18331));
AND2X1 mul_U17845(.A(dpath_mul_op2_d[41]), .B(n9521), .Y(n18332));
AND2X1 mul_U17846(.A(dpath_mul_op2_d[40]), .B(n9510), .Y(n18333));
AND2X1 mul_U17847(.A(dpath_mul_op2_d[39]), .B(n9511), .Y(n18334));
AND2X1 mul_U17848(.A(dpath_mulcore_add_cin), .B(n9509), .Y(n18335));
AND2X1 mul_U17849(.A(dpath_mulcore_booth_b15_in0[2]), .B(n9509), .Y(n18336));
AND2X1 mul_U17850(.A(dpath_mulcore_booth_out_mux16_n2), .B(n9509), .Y(n18337));
AND2X1 mul_U17851(.A(c0_act), .B(dpath_mulcore_booth_b15_in1[2]), .Y(dpath_mulcore_booth_out_mux16_n2));
INVX1 mul_U17852(.A(dpath_mulcore_booth_out_mux16_n2), .Y(n6064));
AND2X1 mul_U17853(.A(n9786), .B(dpath_mulcore_booth_b0_in0[2]), .Y(dpath_mulcore_booth_encode0_a_n75));
AND2X1 mul_U17854(.A(dpath_mout[38]), .B(n9507), .Y(dpath_mulcore_pip_dff_n3));
AND2X1 mul_U17855(.A(dpath_mout[37]), .B(n9507), .Y(dpath_mulcore_pip_dff_n5));
AND2X1 mul_U17856(.A(dpath_mout[36]), .B(n9507), .Y(dpath_mulcore_pip_dff_n7));
AND2X1 mul_U17857(.A(dpath_mout[35]), .B(n9507), .Y(dpath_mulcore_pip_dff_n9));
AND2X1 mul_U17858(.A(dpath_mout[34]), .B(n9507), .Y(dpath_mulcore_pip_dff_n11));
AND2X1 mul_U17859(.A(dpath_mout[33]), .B(n9507), .Y(dpath_mulcore_pip_dff_n13));
AND2X1 mul_U17860(.A(dpath_mout[63]), .B(n9507), .Y(dpath_mulcore_pip_dff_n15));
AND2X1 mul_U17861(.A(dpath_mout[62]), .B(n9507), .Y(dpath_mulcore_pip_dff_n17));
AND2X1 mul_U17862(.A(dpath_mout[61]), .B(n9507), .Y(dpath_mulcore_pip_dff_n19));
AND2X1 mul_U17863(.A(dpath_mout[60]), .B(n9507), .Y(dpath_mulcore_pip_dff_n21));
AND2X1 mul_U17864(.A(dpath_mout[59]), .B(n9507), .Y(dpath_mulcore_pip_dff_n23));
AND2X1 mul_U17865(.A(dpath_mout[32]), .B(n9507), .Y(dpath_mulcore_pip_dff_n25));
AND2X1 mul_U17866(.A(dpath_mout[58]), .B(n9508), .Y(dpath_mulcore_pip_dff_n27));
AND2X1 mul_U17867(.A(dpath_mout[57]), .B(n9508), .Y(dpath_mulcore_pip_dff_n29));
AND2X1 mul_U17868(.A(dpath_mout[56]), .B(n9508), .Y(dpath_mulcore_pip_dff_n31));
AND2X1 mul_U17869(.A(dpath_mout[55]), .B(n9508), .Y(dpath_mulcore_pip_dff_n33));
AND2X1 mul_U17870(.A(dpath_mout[54]), .B(n9508), .Y(dpath_mulcore_pip_dff_n35));
AND2X1 mul_U17871(.A(dpath_mout[53]), .B(n9508), .Y(dpath_mulcore_pip_dff_n37));
AND2X1 mul_U17872(.A(dpath_mout[52]), .B(n9508), .Y(dpath_mulcore_pip_dff_n39));
AND2X1 mul_U17873(.A(dpath_mout[51]), .B(n9508), .Y(dpath_mulcore_pip_dff_n41));
AND2X1 mul_U17874(.A(dpath_mout[50]), .B(n9508), .Y(dpath_mulcore_pip_dff_n43));
AND2X1 mul_U17875(.A(dpath_mout[49]), .B(n9508), .Y(dpath_mulcore_pip_dff_n45));
AND2X1 mul_U17876(.A(dpath_mout[48]), .B(n9508), .Y(dpath_mulcore_pip_dff_n47));
AND2X1 mul_U17877(.A(dpath_mout[47]), .B(n9508), .Y(dpath_mulcore_pip_dff_n49));
AND2X1 mul_U17878(.A(dpath_mout[46]), .B(n9508), .Y(dpath_mulcore_pip_dff_n51));
AND2X1 mul_U17879(.A(dpath_mout[45]), .B(n9509), .Y(dpath_mulcore_pip_dff_n53));
AND2X1 mul_U17880(.A(dpath_mout[44]), .B(n9509), .Y(dpath_mulcore_pip_dff_n55));
AND2X1 mul_U17881(.A(dpath_mout[43]), .B(n9509), .Y(dpath_mulcore_pip_dff_n57));
AND2X1 mul_U17882(.A(dpath_mout[42]), .B(n9509), .Y(dpath_mulcore_pip_dff_n59));
AND2X1 mul_U17883(.A(dpath_mout[41]), .B(n9509), .Y(dpath_mulcore_pip_dff_n61));
AND2X1 mul_U17884(.A(dpath_mout[40]), .B(n9509), .Y(dpath_mulcore_pip_dff_n63));
AND2X1 mul_U17885(.A(dpath_mout[39]), .B(n9509), .Y(dpath_mulcore_pip_dff_n65));
AND2X1 mul_U17886(.A(dpath_mulcore_addout[96]), .B(n9514), .Y(dpath_mulcore_out_dff_n3));
AND2X1 mul_U17887(.A(dpath_mulcore_addout[95]), .B(n9515), .Y(dpath_mulcore_out_dff_n5));
AND2X1 mul_U17888(.A(dpath_mulcore_addout[94]), .B(n9515), .Y(dpath_mulcore_out_dff_n7));
AND2X1 mul_U17889(.A(dpath_mulcore_addout[93]), .B(n9515), .Y(dpath_mulcore_out_dff_n9));
AND2X1 mul_U17890(.A(dpath_mulcore_addout[92]), .B(n9515), .Y(dpath_mulcore_out_dff_n11));
AND2X1 mul_U17891(.A(dpath_mulcore_addout[91]), .B(n9515), .Y(dpath_mulcore_out_dff_n13));
AND2X1 mul_U17892(.A(dpath_mulcore_addout[90]), .B(n9515), .Y(dpath_mulcore_out_dff_n15));
AND2X1 mul_U17893(.A(dpath_mulcore_addout[89]), .B(n9515), .Y(dpath_mulcore_out_dff_n17));
AND2X1 mul_U17894(.A(dpath_mulcore_addout[88]), .B(n9515), .Y(dpath_mulcore_out_dff_n19));
AND2X1 mul_U17895(.A(dpath_mulcore_addout[87]), .B(n9515), .Y(dpath_mulcore_out_dff_n21));
AND2X1 mul_U17896(.A(dpath_mulcore_addout[6]), .B(n9515), .Y(dpath_mulcore_out_dff_n23));
AND2X1 mul_U17897(.A(dpath_mulcore_addout[86]), .B(n9515), .Y(dpath_mulcore_out_dff_n25));
AND2X1 mul_U17898(.A(dpath_mulcore_addout[85]), .B(n9515), .Y(dpath_mulcore_out_dff_n27));
AND2X1 mul_U17899(.A(dpath_mulcore_addout[84]), .B(n9515), .Y(dpath_mulcore_out_dff_n29));
AND2X1 mul_U17900(.A(dpath_mulcore_addout[83]), .B(n9516), .Y(dpath_mulcore_out_dff_n31));
AND2X1 mul_U17901(.A(dpath_mulcore_addout[82]), .B(n9516), .Y(dpath_mulcore_out_dff_n33));
AND2X1 mul_U17902(.A(dpath_mulcore_addout[81]), .B(n9516), .Y(dpath_mulcore_out_dff_n35));
AND2X1 mul_U17903(.A(dpath_mulcore_addout[80]), .B(n9516), .Y(dpath_mulcore_out_dff_n37));
AND2X1 mul_U17904(.A(dpath_mulcore_addout[79]), .B(n9516), .Y(dpath_mulcore_out_dff_n39));
AND2X1 mul_U17905(.A(dpath_mulcore_addout[78]), .B(n9516), .Y(dpath_mulcore_out_dff_n41));
AND2X1 mul_U17906(.A(dpath_mulcore_addout[77]), .B(n9516), .Y(dpath_mulcore_out_dff_n43));
AND2X1 mul_U17907(.A(dpath_mulcore_addout[5]), .B(n9516), .Y(dpath_mulcore_out_dff_n45));
AND2X1 mul_U17908(.A(dpath_mulcore_addout[76]), .B(n9516), .Y(dpath_mulcore_out_dff_n47));
AND2X1 mul_U17909(.A(dpath_mulcore_addout[75]), .B(n9516), .Y(dpath_mulcore_out_dff_n49));
AND2X1 mul_U17910(.A(dpath_mulcore_addout[74]), .B(n9516), .Y(dpath_mulcore_out_dff_n51));
AND2X1 mul_U17911(.A(dpath_mulcore_addout[73]), .B(n9516), .Y(dpath_mulcore_out_dff_n53));
AND2X1 mul_U17912(.A(dpath_mulcore_addout[72]), .B(n9516), .Y(dpath_mulcore_out_dff_n55));
AND2X1 mul_U17913(.A(dpath_mulcore_addout[71]), .B(n9517), .Y(dpath_mulcore_out_dff_n57));
AND2X1 mul_U17914(.A(dpath_mulcore_addout[70]), .B(n9517), .Y(dpath_mulcore_out_dff_n59));
AND2X1 mul_U17915(.A(dpath_mulcore_addout[69]), .B(n9505), .Y(dpath_mulcore_out_dff_n61));
AND2X1 mul_U17916(.A(dpath_mulcore_addout[68]), .B(n9494), .Y(dpath_mulcore_out_dff_n63));
AND2X1 mul_U17917(.A(dpath_mulcore_addout[67]), .B(n9492), .Y(dpath_mulcore_out_dff_n65));
AND2X1 mul_U17918(.A(dpath_mulcore_addout[4]), .B(n9494), .Y(dpath_mulcore_out_dff_n67));
AND2X1 mul_U17919(.A(dpath_mulcore_addout[66]), .B(n9492), .Y(dpath_mulcore_out_dff_n69));
AND2X1 mul_U17920(.A(dpath_mulcore_addout[65]), .B(n9494), .Y(dpath_mulcore_out_dff_n71));
AND2X1 mul_U17921(.A(dpath_mulcore_addout[64]), .B(n9492), .Y(dpath_mulcore_out_dff_n73));
AND2X1 mul_U17922(.A(dpath_mulcore_addout[63]), .B(n9494), .Y(dpath_mulcore_out_dff_n75));
AND2X1 mul_U17923(.A(dpath_mulcore_addout[62]), .B(n9511), .Y(dpath_mulcore_out_dff_n77));
AND2X1 mul_U17924(.A(dpath_mulcore_addout[61]), .B(n9492), .Y(dpath_mulcore_out_dff_n79));
AND2X1 mul_U17925(.A(dpath_mulcore_addout[60]), .B(n9502), .Y(dpath_mulcore_out_dff_n81));
AND2X1 mul_U17926(.A(dpath_mulcore_addout[59]), .B(n9502), .Y(dpath_mulcore_out_dff_n83));
AND2X1 mul_U17927(.A(dpath_mulcore_addout[58]), .B(n9502), .Y(dpath_mulcore_out_dff_n85));
AND2X1 mul_U17928(.A(dpath_mulcore_addout[57]), .B(n9502), .Y(dpath_mulcore_out_dff_n87));
AND2X1 mul_U17929(.A(dpath_mulcore_addout[3]), .B(n9502), .Y(dpath_mulcore_out_dff_n89));
AND2X1 mul_U17930(.A(dpath_mulcore_addout[56]), .B(n9502), .Y(dpath_mulcore_out_dff_n91));
AND2X1 mul_U17931(.A(dpath_mulcore_addout[55]), .B(n9502), .Y(dpath_mulcore_out_dff_n93));
AND2X1 mul_U17932(.A(dpath_mulcore_addout[54]), .B(n9502), .Y(dpath_mulcore_out_dff_n95));
AND2X1 mul_U17933(.A(dpath_mulcore_addout[53]), .B(n9502), .Y(dpath_mulcore_out_dff_n97));
AND2X1 mul_U17934(.A(dpath_mulcore_addout[52]), .B(n9502), .Y(dpath_mulcore_out_dff_n99));
AND2X1 mul_U17935(.A(dpath_mulcore_addout[51]), .B(n9502), .Y(dpath_mulcore_out_dff_n101));
AND2X1 mul_U17936(.A(dpath_mulcore_addout[50]), .B(n9502), .Y(dpath_mulcore_out_dff_n103));
AND2X1 mul_U17937(.A(dpath_mulcore_addout[49]), .B(n9502), .Y(dpath_mulcore_out_dff_n105));
AND2X1 mul_U17938(.A(dpath_mulcore_addout[48]), .B(n9503), .Y(dpath_mulcore_out_dff_n107));
AND2X1 mul_U17939(.A(dpath_mulcore_addout[47]), .B(n9503), .Y(dpath_mulcore_out_dff_n109));
AND2X1 mul_U17940(.A(dpath_mulcore_addout[2]), .B(n9503), .Y(dpath_mulcore_out_dff_n111));
AND2X1 mul_U17941(.A(dpath_mulcore_addout[46]), .B(n9503), .Y(dpath_mulcore_out_dff_n113));
AND2X1 mul_U17942(.A(dpath_mulcore_addout[45]), .B(n9503), .Y(dpath_mulcore_out_dff_n115));
AND2X1 mul_U17943(.A(dpath_mulcore_addout[44]), .B(n9503), .Y(dpath_mulcore_out_dff_n117));
AND2X1 mul_U17944(.A(dpath_mulcore_addout[43]), .B(n9503), .Y(dpath_mulcore_out_dff_n119));
AND2X1 mul_U17945(.A(dpath_mulcore_addout[42]), .B(n9503), .Y(dpath_mulcore_out_dff_n121));
AND2X1 mul_U17946(.A(dpath_mulcore_addout[41]), .B(n9503), .Y(dpath_mulcore_out_dff_n123));
AND2X1 mul_U17947(.A(dpath_mulcore_addout[40]), .B(n9503), .Y(dpath_mulcore_out_dff_n125));
AND2X1 mul_U17948(.A(dpath_mulcore_addout[39]), .B(n9503), .Y(dpath_mulcore_out_dff_n127));
AND2X1 mul_U17949(.A(dpath_mulcore_addout[38]), .B(n9503), .Y(dpath_mulcore_out_dff_n129));
AND2X1 mul_U17950(.A(dpath_mulcore_addout[37]), .B(n9503), .Y(dpath_mulcore_out_dff_n131));
AND2X1 mul_U17951(.A(dpath_mulcore_addout[1]), .B(n9504), .Y(dpath_mulcore_out_dff_n133));
AND2X1 mul_U17952(.A(dpath_mulcore_addout[36]), .B(n9504), .Y(dpath_mulcore_out_dff_n135));
AND2X1 mul_U17953(.A(dpath_mulcore_addout[35]), .B(n9504), .Y(dpath_mulcore_out_dff_n137));
AND2X1 mul_U17954(.A(dpath_mulcore_addout[34]), .B(n9504), .Y(dpath_mulcore_out_dff_n139));
AND2X1 mul_U17955(.A(dpath_mulcore_addout[33]), .B(n9504), .Y(dpath_mulcore_out_dff_n141));
AND2X1 mul_U17956(.A(dpath_mulcore_addout[32]), .B(n9504), .Y(dpath_mulcore_out_dff_n143));
AND2X1 mul_U17957(.A(dpath_mulcore_addout[31]), .B(n9504), .Y(dpath_mulcore_out_dff_n145));
AND2X1 mul_U17958(.A(dpath_mulcore_addout[30]), .B(n9504), .Y(dpath_mulcore_out_dff_n147));
AND2X1 mul_U17959(.A(dpath_mulcore_addout[29]), .B(n9504), .Y(dpath_mulcore_out_dff_n149));
AND2X1 mul_U17960(.A(dpath_mulcore_addout[28]), .B(n9504), .Y(dpath_mulcore_out_dff_n151));
AND2X1 mul_U17961(.A(dpath_mulcore_addout[27]), .B(n9504), .Y(dpath_mulcore_out_dff_n153));
AND2X1 mul_U17962(.A(dpath_mulcore_addout[0]), .B(n9504), .Y(dpath_mulcore_out_dff_n155));
AND2X1 mul_U17963(.A(dpath_mulcore_addout[26]), .B(n9504), .Y(dpath_mulcore_out_dff_n157));
AND2X1 mul_U17964(.A(dpath_mulcore_addout[25]), .B(n9505), .Y(dpath_mulcore_out_dff_n159));
AND2X1 mul_U17965(.A(dpath_mulcore_addout[24]), .B(n9505), .Y(dpath_mulcore_out_dff_n161));
AND2X1 mul_U17966(.A(dpath_mulcore_addout[23]), .B(n9505), .Y(dpath_mulcore_out_dff_n163));
AND2X1 mul_U17967(.A(dpath_mulcore_addout[22]), .B(n9505), .Y(dpath_mulcore_out_dff_n165));
AND2X1 mul_U17968(.A(dpath_mulcore_addout[21]), .B(n9505), .Y(dpath_mulcore_out_dff_n167));
AND2X1 mul_U17969(.A(dpath_mulcore_addout[20]), .B(n9505), .Y(dpath_mulcore_out_dff_n169));
AND2X1 mul_U17970(.A(dpath_mulcore_addout[19]), .B(n9505), .Y(dpath_mulcore_out_dff_n171));
AND2X1 mul_U17971(.A(dpath_mulcore_addout[18]), .B(n9505), .Y(dpath_mulcore_out_dff_n173));
AND2X1 mul_U17972(.A(dpath_mulcore_addout[17]), .B(n9505), .Y(dpath_mulcore_out_dff_n175));
AND2X1 mul_U17973(.A(dpath_mulcore_addout[16]), .B(n9505), .Y(dpath_mulcore_out_dff_n177));
AND2X1 mul_U17974(.A(dpath_mulcore_addout[15]), .B(n9505), .Y(dpath_mulcore_out_dff_n179));
AND2X1 mul_U17975(.A(dpath_mulcore_addout[14]), .B(n9505), .Y(dpath_mulcore_out_dff_n181));
AND2X1 mul_U17976(.A(dpath_mulcore_addout[13]), .B(n9506), .Y(dpath_mulcore_out_dff_n183));
AND2X1 mul_U17977(.A(dpath_mulcore_addout[12]), .B(n9506), .Y(dpath_mulcore_out_dff_n185));
AND2X1 mul_U17978(.A(dpath_mulcore_addout[11]), .B(n9506), .Y(dpath_mulcore_out_dff_n187));
AND2X1 mul_U17979(.A(dpath_mulcore_addout[10]), .B(n9506), .Y(dpath_mulcore_out_dff_n189));
AND2X1 mul_U17980(.A(dpath_mulcore_addout[9]), .B(n9506), .Y(dpath_mulcore_out_dff_n191));
AND2X1 mul_U17981(.A(dpath_mulcore_addout[8]), .B(n9506), .Y(dpath_mulcore_out_dff_n193));
AND2X1 mul_U17982(.A(dpath_mulcore_addout[103]), .B(n9506), .Y(dpath_mulcore_out_dff_n195));
AND2X1 mul_U17983(.A(dpath_mulcore_addout[102]), .B(n9506), .Y(dpath_mulcore_out_dff_n197));
AND2X1 mul_U17984(.A(dpath_mulcore_addout[101]), .B(n9506), .Y(dpath_mulcore_out_dff_n199));
AND2X1 mul_U17985(.A(dpath_mulcore_addout[100]), .B(n9506), .Y(dpath_mulcore_out_dff_n201));
AND2X1 mul_U17986(.A(dpath_mulcore_addout[99]), .B(n9506), .Y(dpath_mulcore_out_dff_n203));
AND2X1 mul_U17987(.A(dpath_mulcore_addout[98]), .B(n9506), .Y(dpath_mulcore_out_dff_n205));
AND2X1 mul_U17988(.A(dpath_mulcore_addout[97]), .B(n9506), .Y(dpath_mulcore_out_dff_n207));
AND2X1 mul_U17989(.A(dpath_mulcore_addout[7]), .B(n9507), .Y(dpath_mulcore_out_dff_n209));
AND2X1 mul_U17990(.A(dpath_mulcore_pcout_in[36]), .B(n9511), .Y(dpath_mulcore_pcout_dff_n3));
AND2X1 mul_U17991(.A(dpath_mulcore_pcout_in[35]), .B(n9511), .Y(dpath_mulcore_pcout_dff_n5));
AND2X1 mul_U17992(.A(dpath_mulcore_pcout_in[97]), .B(n9511), .Y(dpath_mulcore_pcout_dff_n9));
AND2X1 mul_U17993(.A(dpath_mulcore_pcout_in[34]), .B(n9511), .Y(dpath_mulcore_pcout_dff_n11));
AND2X1 mul_U17994(.A(dpath_mulcore_pcout_in[96]), .B(n9511), .Y(dpath_mulcore_pcout_dff_n13));
AND2X1 mul_U17995(.A(dpath_mulcore_pcout_in[95]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n15));
AND2X1 mul_U17996(.A(dpath_mulcore_pcout_in[94]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n17));
AND2X1 mul_U17997(.A(dpath_mulcore_pcout_in[93]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n19));
AND2X1 mul_U17998(.A(dpath_mulcore_pcout_in[92]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n21));
AND2X1 mul_U17999(.A(dpath_mulcore_pcout_in[91]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n23));
AND2X1 mul_U18000(.A(dpath_mulcore_pcout_in[90]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n25));
AND2X1 mul_U18001(.A(dpath_mulcore_pcout_in[89]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n27));
AND2X1 mul_U18002(.A(dpath_mulcore_pcout_in[88]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n29));
AND2X1 mul_U18003(.A(dpath_mulcore_pcout_in[87]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n31));
AND2X1 mul_U18004(.A(dpath_mulcore_pcout_in[33]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n33));
AND2X1 mul_U18005(.A(dpath_mulcore_pcout_in[86]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n35));
AND2X1 mul_U18006(.A(dpath_mulcore_pcout_in[85]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n37));
AND2X1 mul_U18007(.A(dpath_mulcore_pcout_in[84]), .B(n9512), .Y(dpath_mulcore_pcout_dff_n39));
AND2X1 mul_U18008(.A(dpath_mulcore_pcout_in[83]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n41));
AND2X1 mul_U18009(.A(dpath_mulcore_pcout_in[82]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n43));
AND2X1 mul_U18010(.A(dpath_mulcore_pcout_in[81]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n45));
AND2X1 mul_U18011(.A(dpath_mulcore_pcout_in[80]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n47));
AND2X1 mul_U18012(.A(dpath_mulcore_pcout_in[79]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n49));
AND2X1 mul_U18013(.A(dpath_mulcore_pcout_in[78]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n51));
AND2X1 mul_U18014(.A(dpath_mulcore_pcout_in[77]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n53));
AND2X1 mul_U18015(.A(dpath_mulcore_pcout_in[32]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n55));
AND2X1 mul_U18016(.A(dpath_mulcore_pcout_in[76]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n57));
AND2X1 mul_U18017(.A(dpath_mulcore_pcout_in[75]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n59));
AND2X1 mul_U18018(.A(dpath_mulcore_pcout_in[74]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n61));
AND2X1 mul_U18019(.A(dpath_mulcore_pcout_in[73]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n63));
AND2X1 mul_U18020(.A(dpath_mulcore_pcout_in[72]), .B(n9513), .Y(dpath_mulcore_pcout_dff_n65));
AND2X1 mul_U18021(.A(dpath_mulcore_pcout_in[71]), .B(n9498), .Y(dpath_mulcore_pcout_dff_n67));
AND2X1 mul_U18022(.A(dpath_mulcore_pcout_in[70]), .B(n9498), .Y(dpath_mulcore_pcout_dff_n69));
AND2X1 mul_U18023(.A(dpath_mulcore_pcout_in[69]), .B(n9497), .Y(dpath_mulcore_pcout_dff_n71));
AND2X1 mul_U18024(.A(dpath_mulcore_pcout_in[68]), .B(n9498), .Y(dpath_mulcore_pcout_dff_n73));
AND2X1 mul_U18025(.A(dpath_mulcore_pcout_in[67]), .B(n9497), .Y(dpath_mulcore_pcout_dff_n75));
AND2X1 mul_U18026(.A(dpath_mulcore_pcout_in[31]), .B(n9492), .Y(dpath_mulcore_pcout_dff_n77));
AND2X1 mul_U18027(.A(dpath_mulcore_pcout_in[66]), .B(n9498), .Y(dpath_mulcore_pcout_dff_n79));
AND2X1 mul_U18028(.A(dpath_mulcore_pcout_in[65]), .B(n9494), .Y(dpath_mulcore_pcout_dff_n81));
AND2X1 mul_U18029(.A(dpath_mulcore_pcout_in[64]), .B(n9496), .Y(dpath_mulcore_pcout_dff_n83));
AND2X1 mul_U18030(.A(dpath_mulcore_pcout_in[63]), .B(n9495), .Y(dpath_mulcore_pcout_dff_n85));
AND2X1 mul_U18031(.A(dpath_mulcore_pcout_in[62]), .B(n9550), .Y(dpath_mulcore_pcout_dff_n87));
AND2X1 mul_U18032(.A(dpath_mulcore_pcout_in[61]), .B(n9497), .Y(dpath_mulcore_pcout_dff_n89));
AND2X1 mul_U18033(.A(dpath_mulcore_pcout_in[60]), .B(n9498), .Y(dpath_mulcore_pcout_dff_n91));
AND2X1 mul_U18034(.A(dpath_mulcore_pcout_in[59]), .B(n9498), .Y(dpath_mulcore_pcout_dff_n93));
AND2X1 mul_U18035(.A(dpath_mulcore_pcout_in[58]), .B(n9498), .Y(dpath_mulcore_pcout_dff_n95));
AND2X1 mul_U18036(.A(dpath_mulcore_pcout_in[57]), .B(n9541), .Y(dpath_mulcore_pcout_dff_n97));
AND2X1 mul_U18037(.A(dpath_mulcore_pcout_in[30]), .B(n9540), .Y(dpath_mulcore_pcout_dff_n99));
AND2X1 mul_U18038(.A(dpath_mulcore_pcout_in[56]), .B(n9539), .Y(dpath_mulcore_pcout_dff_n101));
AND2X1 mul_U18039(.A(dpath_mulcore_pcout_in[55]), .B(n9511), .Y(dpath_mulcore_pcout_dff_n103));
AND2X1 mul_U18040(.A(dpath_mulcore_pcout_in[54]), .B(n9518), .Y(dpath_mulcore_pcout_dff_n105));
AND2X1 mul_U18041(.A(dpath_mulcore_pcout_in[53]), .B(n9517), .Y(dpath_mulcore_pcout_dff_n107));
AND2X1 mul_U18042(.A(dpath_mulcore_pcout_in[52]), .B(n9548), .Y(dpath_mulcore_pcout_dff_n109));
AND2X1 mul_U18043(.A(dpath_mulcore_pcout_in[51]), .B(n9549), .Y(dpath_mulcore_pcout_dff_n111));
AND2X1 mul_U18044(.A(dpath_mulcore_pcout_in[50]), .B(n9552), .Y(dpath_mulcore_pcout_dff_n113));
AND2X1 mul_U18045(.A(dpath_mulcore_pcout_in[49]), .B(n9551), .Y(dpath_mulcore_pcout_dff_n115));
AND2X1 mul_U18046(.A(dpath_mulcore_pcout_in[48]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n117));
AND2X1 mul_U18047(.A(dpath_mulcore_pcout_in[47]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n119));
AND2X1 mul_U18048(.A(dpath_mulcore_pcout_in[46]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n121));
AND2X1 mul_U18049(.A(dpath_mulcore_pcout_in[45]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n123));
AND2X1 mul_U18050(.A(dpath_mulcore_pcout_in[44]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n125));
AND2X1 mul_U18051(.A(dpath_mulcore_pcout_in[43]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n127));
AND2X1 mul_U18052(.A(dpath_mulcore_pcout_in[42]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n129));
AND2X1 mul_U18053(.A(dpath_mulcore_pcout_in[41]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n131));
AND2X1 mul_U18054(.A(dpath_mulcore_pcout_in[40]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n133));
AND2X1 mul_U18055(.A(dpath_mulcore_pcout_in[39]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n135));
AND2X1 mul_U18056(.A(dpath_mulcore_pcout_in[38]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n137));
AND2X1 mul_U18057(.A(dpath_mulcore_pcout_in[37]), .B(n9514), .Y(dpath_mulcore_pcout_dff_n139));
AND2X1 mul_U18058(.A(dpath_mulcore_psum_in[37]), .B(n9552), .Y(dpath_mulcore_psum_dff_n3));
AND2X1 mul_U18059(.A(dpath_mulcore_psum_in[36]), .B(n9552), .Y(dpath_mulcore_psum_dff_n5));
AND2X1 mul_U18060(.A(dpath_mulcore_psum_in[98]), .B(n9552), .Y(dpath_mulcore_psum_dff_n7));
AND2X1 mul_U18061(.A(dpath_mulcore_psum_in[35]), .B(n9552), .Y(dpath_mulcore_psum_dff_n9));
AND2X1 mul_U18062(.A(dpath_mulcore_psum_in[97]), .B(n9552), .Y(dpath_mulcore_psum_dff_n11));
AND2X1 mul_U18063(.A(dpath_mulcore_psum_in[96]), .B(n9552), .Y(dpath_mulcore_psum_dff_n13));
AND2X1 mul_U18064(.A(dpath_mulcore_psum_in[95]), .B(n9552), .Y(dpath_mulcore_psum_dff_n15));
AND2X1 mul_U18065(.A(dpath_mulcore_psum_in[94]), .B(n9552), .Y(dpath_mulcore_psum_dff_n17));
AND2X1 mul_U18066(.A(dpath_mulcore_psum_in[93]), .B(n9552), .Y(dpath_mulcore_psum_dff_n19));
AND2X1 mul_U18067(.A(dpath_mulcore_psum_in[92]), .B(n9553), .Y(dpath_mulcore_psum_dff_n21));
AND2X1 mul_U18068(.A(dpath_mulcore_psum_in[91]), .B(n9553), .Y(dpath_mulcore_psum_dff_n23));
AND2X1 mul_U18069(.A(dpath_mulcore_psum_in[90]), .B(n9553), .Y(dpath_mulcore_psum_dff_n25));
AND2X1 mul_U18070(.A(dpath_mulcore_psum_in[89]), .B(n9553), .Y(dpath_mulcore_psum_dff_n27));
AND2X1 mul_U18071(.A(dpath_mulcore_psum_in[88]), .B(n9553), .Y(dpath_mulcore_psum_dff_n29));
AND2X1 mul_U18072(.A(dpath_mulcore_psum_in[34]), .B(n9553), .Y(dpath_mulcore_psum_dff_n31));
AND2X1 mul_U18073(.A(dpath_mulcore_psum_in[87]), .B(n9553), .Y(dpath_mulcore_psum_dff_n33));
AND2X1 mul_U18074(.A(dpath_mulcore_psum_in[86]), .B(n9553), .Y(dpath_mulcore_psum_dff_n35));
AND2X1 mul_U18075(.A(dpath_mulcore_psum_in[85]), .B(n9553), .Y(dpath_mulcore_psum_dff_n37));
AND2X1 mul_U18076(.A(dpath_mulcore_psum_in[84]), .B(n9553), .Y(dpath_mulcore_psum_dff_n39));
AND2X1 mul_U18077(.A(dpath_mulcore_psum_in[83]), .B(n9553), .Y(dpath_mulcore_psum_dff_n41));
AND2X1 mul_U18078(.A(dpath_mulcore_psum_in[82]), .B(n9553), .Y(dpath_mulcore_psum_dff_n43));
AND2X1 mul_U18079(.A(dpath_mulcore_psum_in[81]), .B(n9553), .Y(dpath_mulcore_psum_dff_n45));
AND2X1 mul_U18080(.A(dpath_mulcore_psum_in[80]), .B(n9554), .Y(dpath_mulcore_psum_dff_n47));
AND2X1 mul_U18081(.A(dpath_mulcore_psum_in[79]), .B(n9554), .Y(dpath_mulcore_psum_dff_n49));
AND2X1 mul_U18082(.A(dpath_mulcore_psum_in[78]), .B(n9554), .Y(dpath_mulcore_psum_dff_n51));
AND2X1 mul_U18083(.A(dpath_mulcore_psum_in[33]), .B(n9554), .Y(dpath_mulcore_psum_dff_n53));
AND2X1 mul_U18084(.A(dpath_mulcore_psum_in[77]), .B(n9554), .Y(dpath_mulcore_psum_dff_n55));
AND2X1 mul_U18085(.A(dpath_mulcore_psum_in[76]), .B(n9554), .Y(dpath_mulcore_psum_dff_n57));
AND2X1 mul_U18086(.A(dpath_mulcore_psum_in[75]), .B(n9554), .Y(dpath_mulcore_psum_dff_n59));
AND2X1 mul_U18087(.A(dpath_mulcore_psum_in[74]), .B(n9554), .Y(dpath_mulcore_psum_dff_n61));
AND2X1 mul_U18088(.A(dpath_mulcore_psum_in[73]), .B(n9554), .Y(dpath_mulcore_psum_dff_n63));
AND2X1 mul_U18089(.A(dpath_mulcore_psum_in[72]), .B(n9554), .Y(dpath_mulcore_psum_dff_n65));
AND2X1 mul_U18090(.A(dpath_mulcore_psum_in[71]), .B(n9554), .Y(dpath_mulcore_psum_dff_n67));
AND2X1 mul_U18091(.A(dpath_mulcore_psum_in[70]), .B(n9554), .Y(dpath_mulcore_psum_dff_n69));
AND2X1 mul_U18092(.A(dpath_mulcore_psum_in[69]), .B(n9554), .Y(dpath_mulcore_psum_dff_n71));
AND2X1 mul_U18093(.A(dpath_mulcore_psum_in[68]), .B(n9555), .Y(dpath_mulcore_psum_dff_n73));
AND2X1 mul_U18094(.A(dpath_mulcore_psum_in[32]), .B(n9555), .Y(dpath_mulcore_psum_dff_n75));
AND2X1 mul_U18095(.A(dpath_mulcore_psum_in[67]), .B(n9555), .Y(dpath_mulcore_psum_dff_n77));
AND2X1 mul_U18096(.A(dpath_mulcore_psum_in[66]), .B(n9555), .Y(dpath_mulcore_psum_dff_n79));
AND2X1 mul_U18097(.A(dpath_mulcore_psum_in[65]), .B(n9555), .Y(dpath_mulcore_psum_dff_n81));
AND2X1 mul_U18098(.A(dpath_mulcore_psum_in[64]), .B(n9555), .Y(dpath_mulcore_psum_dff_n83));
AND2X1 mul_U18099(.A(dpath_mulcore_psum_in[63]), .B(n9555), .Y(dpath_mulcore_psum_dff_n85));
AND2X1 mul_U18100(.A(dpath_mulcore_psum_in[62]), .B(n9555), .Y(dpath_mulcore_psum_dff_n87));
AND2X1 mul_U18101(.A(dpath_mulcore_psum_in[61]), .B(n9555), .Y(dpath_mulcore_psum_dff_n89));
AND2X1 mul_U18102(.A(dpath_mulcore_psum_in[60]), .B(n9555), .Y(dpath_mulcore_psum_dff_n91));
AND2X1 mul_U18103(.A(dpath_mulcore_psum_in[59]), .B(n9555), .Y(dpath_mulcore_psum_dff_n93));
AND2X1 mul_U18104(.A(dpath_mulcore_psum_in[58]), .B(n9555), .Y(dpath_mulcore_psum_dff_n95));
AND2X1 mul_U18105(.A(dpath_mulcore_psum_in[31]), .B(n9555), .Y(dpath_mulcore_psum_dff_n97));
AND2X1 mul_U18106(.A(dpath_mulcore_psum_in[57]), .B(n9556), .Y(dpath_mulcore_psum_dff_n99));
AND2X1 mul_U18107(.A(dpath_mulcore_psum_in[56]), .B(n9517), .Y(dpath_mulcore_psum_dff_n101));
AND2X1 mul_U18108(.A(dpath_mulcore_psum_in[55]), .B(n9512), .Y(dpath_mulcore_psum_dff_n103));
AND2X1 mul_U18109(.A(dpath_mulcore_psum_in[54]), .B(n9510), .Y(dpath_mulcore_psum_dff_n105));
AND2X1 mul_U18110(.A(dpath_mulcore_psum_in[53]), .B(n9510), .Y(dpath_mulcore_psum_dff_n107));
AND2X1 mul_U18111(.A(dpath_mulcore_psum_in[52]), .B(n9510), .Y(dpath_mulcore_psum_dff_n109));
AND2X1 mul_U18112(.A(dpath_mulcore_psum_in[51]), .B(n9510), .Y(dpath_mulcore_psum_dff_n111));
AND2X1 mul_U18113(.A(dpath_mulcore_psum_in[50]), .B(n9510), .Y(dpath_mulcore_psum_dff_n113));
AND2X1 mul_U18114(.A(dpath_mulcore_psum_in[49]), .B(n9510), .Y(dpath_mulcore_psum_dff_n115));
AND2X1 mul_U18115(.A(dpath_mulcore_psum_in[48]), .B(n9510), .Y(dpath_mulcore_psum_dff_n117));
AND2X1 mul_U18116(.A(dpath_mulcore_psum_in[47]), .B(n9510), .Y(dpath_mulcore_psum_dff_n119));
AND2X1 mul_U18117(.A(dpath_mulcore_psum_in[46]), .B(n9510), .Y(dpath_mulcore_psum_dff_n121));
AND2X1 mul_U18118(.A(dpath_mulcore_psum_in[45]), .B(n9510), .Y(dpath_mulcore_psum_dff_n123));
AND2X1 mul_U18119(.A(dpath_mulcore_psum_in[44]), .B(n9511), .Y(dpath_mulcore_psum_dff_n125));
AND2X1 mul_U18120(.A(dpath_mulcore_psum_in[43]), .B(n9511), .Y(dpath_mulcore_psum_dff_n127));
AND2X1 mul_U18121(.A(dpath_mulcore_psum_in[42]), .B(n9511), .Y(dpath_mulcore_psum_dff_n129));
AND2X1 mul_U18122(.A(dpath_mulcore_psum_in[41]), .B(n9511), .Y(dpath_mulcore_psum_dff_n131));
AND2X1 mul_U18123(.A(dpath_mulcore_psum_in[40]), .B(n9511), .Y(dpath_mulcore_psum_dff_n133));
AND2X1 mul_U18124(.A(dpath_mulcore_psum_in[39]), .B(n9511), .Y(dpath_mulcore_psum_dff_n135));
AND2X1 mul_U18125(.A(dpath_mulcore_psum_in[38]), .B(n9511), .Y(dpath_mulcore_psum_dff_n137));
AND2X1 mul_U18126(.A(dpath_mulcore_a0sum[6]), .B(n9557), .Y(dpath_mulcore_a0sum_dff_n3));
AND2X1 mul_U18127(.A(dpath_mulcore_a0sum[79]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n9));
AND2X1 mul_U18128(.A(dpath_mulcore_a0sum[78]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n11));
AND2X1 mul_U18129(.A(dpath_mulcore_a0sum[77]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n13));
AND2X1 mul_U18130(.A(dpath_mulcore_a0sum[5]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n15));
AND2X1 mul_U18131(.A(dpath_mulcore_a0sum[76]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n17));
AND2X1 mul_U18132(.A(dpath_mulcore_a0sum[75]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n19));
AND2X1 mul_U18133(.A(dpath_mulcore_a0sum[74]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n21));
AND2X1 mul_U18134(.A(dpath_mulcore_a0sum[73]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n23));
AND2X1 mul_U18135(.A(dpath_mulcore_a0sum[72]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n25));
AND2X1 mul_U18136(.A(dpath_mulcore_a0sum[71]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n27));
AND2X1 mul_U18137(.A(dpath_mulcore_a0sum[70]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n29));
AND2X1 mul_U18138(.A(dpath_mulcore_a0sum[69]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n31));
AND2X1 mul_U18139(.A(dpath_mulcore_a0sum[68]), .B(n9533), .Y(dpath_mulcore_a0sum_dff_n33));
AND2X1 mul_U18140(.A(dpath_mulcore_a0sum[67]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n35));
AND2X1 mul_U18141(.A(dpath_mulcore_a0sum[4]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n37));
AND2X1 mul_U18142(.A(dpath_mulcore_a0sum[66]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n39));
AND2X1 mul_U18143(.A(dpath_mulcore_a0sum[65]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n41));
AND2X1 mul_U18144(.A(dpath_mulcore_a0sum[64]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n43));
AND2X1 mul_U18145(.A(dpath_mulcore_a0sum[63]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n45));
AND2X1 mul_U18146(.A(dpath_mulcore_a0sum[62]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n47));
AND2X1 mul_U18147(.A(dpath_mulcore_a0sum[61]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n49));
AND2X1 mul_U18148(.A(dpath_mulcore_a0sum[60]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n51));
AND2X1 mul_U18149(.A(dpath_mulcore_a0sum[59]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n53));
AND2X1 mul_U18150(.A(dpath_mulcore_a0sum[58]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n55));
AND2X1 mul_U18151(.A(dpath_mulcore_a0sum[57]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n57));
AND2X1 mul_U18152(.A(dpath_mulcore_a0sum[3]), .B(n9534), .Y(dpath_mulcore_a0sum_dff_n59));
AND2X1 mul_U18153(.A(dpath_mulcore_a0sum[56]), .B(n9495), .Y(dpath_mulcore_a0sum_dff_n61));
AND2X1 mul_U18154(.A(dpath_mulcore_a0sum[55]), .B(n9495), .Y(dpath_mulcore_a0sum_dff_n63));
AND2X1 mul_U18155(.A(dpath_mulcore_a0sum[54]), .B(n9559), .Y(dpath_mulcore_a0sum_dff_n65));
AND2X1 mul_U18156(.A(dpath_mulcore_a0sum[53]), .B(n9560), .Y(dpath_mulcore_a0sum_dff_n67));
AND2X1 mul_U18157(.A(dpath_mulcore_a0sum[52]), .B(n9561), .Y(dpath_mulcore_a0sum_dff_n69));
AND2X1 mul_U18158(.A(dpath_mulcore_a0sum[51]), .B(n9502), .Y(dpath_mulcore_a0sum_dff_n71));
AND2X1 mul_U18159(.A(dpath_mulcore_a0sum[50]), .B(n9503), .Y(dpath_mulcore_a0sum_dff_n73));
AND2X1 mul_U18160(.A(dpath_mulcore_a0sum[49]), .B(n9504), .Y(dpath_mulcore_a0sum_dff_n75));
AND2X1 mul_U18161(.A(dpath_mulcore_a0sum[48]), .B(n9505), .Y(dpath_mulcore_a0sum_dff_n77));
AND2X1 mul_U18162(.A(dpath_mulcore_a0sum[47]), .B(n9506), .Y(dpath_mulcore_a0sum_dff_n79));
AND2X1 mul_U18163(.A(dpath_mulcore_a0sum[2]), .B(n9507), .Y(dpath_mulcore_a0sum_dff_n81));
AND2X1 mul_U18164(.A(dpath_mulcore_a0sum[46]), .B(n9508), .Y(dpath_mulcore_a0sum_dff_n83));
AND2X1 mul_U18165(.A(dpath_mulcore_a0sum[45]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n85));
AND2X1 mul_U18166(.A(dpath_mulcore_a0sum[44]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n87));
AND2X1 mul_U18167(.A(dpath_mulcore_a0sum[43]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n89));
AND2X1 mul_U18168(.A(dpath_mulcore_a0sum[42]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n91));
AND2X1 mul_U18169(.A(dpath_mulcore_a0sum[41]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n93));
AND2X1 mul_U18170(.A(dpath_mulcore_a0sum[40]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n95));
AND2X1 mul_U18171(.A(dpath_mulcore_a0sum[39]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n97));
AND2X1 mul_U18172(.A(dpath_mulcore_a0sum[38]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n99));
AND2X1 mul_U18173(.A(dpath_mulcore_a0sum[37]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n101));
AND2X1 mul_U18174(.A(dpath_mulcore_a0sum[1]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n103));
AND2X1 mul_U18175(.A(dpath_mulcore_a0sum[36]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n105));
AND2X1 mul_U18176(.A(dpath_mulcore_a0sum[35]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n107));
AND2X1 mul_U18177(.A(dpath_mulcore_a0sum[34]), .B(n9535), .Y(dpath_mulcore_a0sum_dff_n109));
AND2X1 mul_U18178(.A(dpath_mulcore_a0sum[33]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n111));
AND2X1 mul_U18179(.A(dpath_mulcore_a0sum[32]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n113));
AND2X1 mul_U18180(.A(dpath_mulcore_a0sum[31]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n115));
AND2X1 mul_U18181(.A(dpath_mulcore_a0sum[30]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n117));
AND2X1 mul_U18182(.A(dpath_mulcore_a0sum[29]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n119));
AND2X1 mul_U18183(.A(dpath_mulcore_a0sum[28]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n121));
AND2X1 mul_U18184(.A(dpath_mulcore_a0sum[27]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n123));
AND2X1 mul_U18185(.A(dpath_mulcore_a0sum[0]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n125));
AND2X1 mul_U18186(.A(dpath_mulcore_a0sum[26]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n127));
AND2X1 mul_U18187(.A(dpath_mulcore_a0sum[25]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n129));
AND2X1 mul_U18188(.A(dpath_mulcore_a0sum[24]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n131));
AND2X1 mul_U18189(.A(dpath_mulcore_a0sum[23]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n133));
AND2X1 mul_U18190(.A(dpath_mulcore_a0sum[22]), .B(n9536), .Y(dpath_mulcore_a0sum_dff_n135));
AND2X1 mul_U18191(.A(dpath_mulcore_a0sum[21]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n137));
AND2X1 mul_U18192(.A(dpath_mulcore_a0sum[20]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n139));
AND2X1 mul_U18193(.A(dpath_mulcore_a0sum[19]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n141));
AND2X1 mul_U18194(.A(dpath_mulcore_a0sum[18]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n143));
AND2X1 mul_U18195(.A(dpath_mulcore_a0sum[17]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n145));
AND2X1 mul_U18196(.A(dpath_mulcore_a0sum[16]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n147));
AND2X1 mul_U18197(.A(dpath_mulcore_a0sum[15]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n149));
AND2X1 mul_U18198(.A(dpath_mulcore_a0sum[14]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n151));
AND2X1 mul_U18199(.A(dpath_mulcore_a0sum[13]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n153));
AND2X1 mul_U18200(.A(dpath_mulcore_a0sum[12]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n155));
AND2X1 mul_U18201(.A(dpath_mulcore_ary1_a0_sc3_11__z), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n157));
AND2X1 mul_U18202(.A(dpath_mulcore_a0sum[10]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n159));
AND2X1 mul_U18203(.A(dpath_mulcore_a0sum[9]), .B(n9537), .Y(dpath_mulcore_a0sum_dff_n161));
AND2X1 mul_U18204(.A(dpath_mulcore_a0sum[8]), .B(n9538), .Y(dpath_mulcore_a0sum_dff_n163));
AND2X1 mul_U18205(.A(dpath_mulcore_a0sum[7]), .B(n9538), .Y(dpath_mulcore_a0sum_dff_n165));
AND2X1 mul_U18206(.A(dpath_mulcore_a0cout[79]), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n11));
AND2X1 mul_U18207(.A(dpath_mulcore_a0cout[78]), .B(n9544), .Y(dpath_mulcore_a0cot_dff_n13));
AND2X1 mul_U18208(.A(dpath_mulcore_a0cout[7]), .B(n9545), .Y(dpath_mulcore_a0cot_dff_n51));
AND2X1 mul_U18209(.A(dpath_mulcore_a0cout[6]), .B(n9546), .Y(dpath_mulcore_a0cot_dff_n73));
AND2X1 mul_U18210(.A(dpath_mulcore_a0cout[5]), .B(n9547), .Y(dpath_mulcore_a0cot_dff_n95));
AND2X1 mul_U18211(.A(dpath_mulcore_a0cout[4]), .B(n9532), .Y(dpath_mulcore_a0cot_dff_n117));
AND2X1 mul_U18212(.A(n17022), .B(n9558), .Y(dpath_mulcore_a0cot_dff_n157));
AND2X1 mul_U18213(.A(dpath_acc_reg_in[135]), .B(n7195), .Y(dpath_accum_n2));
AND2X1 mul_U18214(.A(dpath_acc_reg_in[134]), .B(n7195), .Y(dpath_accum_n5));
AND2X1 mul_U18215(.A(dpath_acc_reg_in[133]), .B(n7195), .Y(dpath_accum_n7));
AND2X1 mul_U18216(.A(dpath_acc_reg_in[132]), .B(n7195), .Y(dpath_accum_n9));
AND2X1 mul_U18217(.A(dpath_acc_reg_in[131]), .B(n7195), .Y(dpath_accum_n11));
AND2X1 mul_U18218(.A(dpath_acc_reg_in[130]), .B(n7195), .Y(dpath_accum_n13));
AND2X1 mul_U18219(.A(dpath_acc_reg_in[129]), .B(n7195), .Y(dpath_accum_n15));
AND2X1 mul_U18220(.A(dpath_acc_reg_in[128]), .B(n7195), .Y(dpath_accum_n17));
AND2X1 mul_U18221(.A(dpath_acc_reg_in[127]), .B(n7195), .Y(dpath_accum_n19));
AND2X1 mul_U18222(.A(dpath_acc_reg_in[126]), .B(n9592), .Y(dpath_accum_n21));
AND2X1 mul_U18223(.A(dpath_acc_reg_in[125]), .B(n7195), .Y(dpath_accum_n23));
AND2X1 mul_U18224(.A(dpath_acc_reg_in[124]), .B(n7195), .Y(dpath_accum_n25));
AND2X1 mul_U18225(.A(dpath_acc_reg_in[123]), .B(n7195), .Y(dpath_accum_n27));
AND2X1 mul_U18226(.A(dpath_acc_reg_in[122]), .B(n9592), .Y(dpath_accum_n29));
AND2X1 mul_U18227(.A(dpath_acc_reg_in[121]), .B(n9592), .Y(dpath_accum_n31));
AND2X1 mul_U18228(.A(dpath_acc_reg_in[120]), .B(n9592), .Y(dpath_accum_n33));
AND2X1 mul_U18229(.A(dpath_acc_reg_in[119]), .B(n9592), .Y(dpath_accum_n35));
AND2X1 mul_U18230(.A(dpath_acc_reg_in[118]), .B(n9592), .Y(dpath_accum_n37));
AND2X1 mul_U18231(.A(dpath_acc_reg_in[117]), .B(n9592), .Y(dpath_accum_n39));
AND2X1 mul_U18232(.A(dpath_acc_reg_in[116]), .B(n9592), .Y(dpath_accum_n41));
AND2X1 mul_U18233(.A(dpath_acc_reg_in[115]), .B(n9592), .Y(dpath_accum_n43));
AND2X1 mul_U18234(.A(dpath_acc_reg_in[114]), .B(n7195), .Y(dpath_accum_n45));
AND2X1 mul_U18235(.A(dpath_acc_reg_in[113]), .B(n9592), .Y(dpath_accum_n47));
AND2X1 mul_U18236(.A(dpath_acc_reg_in[112]), .B(n7195), .Y(dpath_accum_n49));
AND2X1 mul_U18237(.A(dpath_acc_reg_in[111]), .B(n7195), .Y(dpath_accum_n51));
AND2X1 mul_U18238(.A(dpath_acc_reg_in[110]), .B(n9592), .Y(dpath_accum_n53));
AND2X1 mul_U18239(.A(dpath_acc_reg_in[109]), .B(n9592), .Y(dpath_accum_n55));
AND2X1 mul_U18240(.A(dpath_acc_reg_in[108]), .B(n7195), .Y(dpath_accum_n57));
AND2X1 mul_U18241(.A(dpath_acc_reg_in[107]), .B(n9592), .Y(dpath_accum_n59));
AND2X1 mul_U18242(.A(dpath_acc_reg_in[106]), .B(n7195), .Y(dpath_accum_n61));
AND2X1 mul_U18243(.A(dpath_acc_reg_in[105]), .B(n7195), .Y(dpath_accum_n63));
AND2X1 mul_U18244(.A(dpath_acc_reg_in[104]), .B(n9592), .Y(dpath_accum_n65));
AND2X1 mul_U18245(.A(dpath_acc_reg_in[103]), .B(n9592), .Y(dpath_accum_n67));
AND2X1 mul_U18246(.A(dpath_acc_reg_in[102]), .B(n7195), .Y(dpath_accum_n69));
AND2X1 mul_U18247(.A(dpath_acc_reg_in[101]), .B(n9592), .Y(dpath_accum_n71));
AND2X1 mul_U18248(.A(dpath_acc_reg_in[100]), .B(n9592), .Y(dpath_accum_n73));
AND2X1 mul_U18249(.A(dpath_acc_reg_in[99]), .B(n7195), .Y(dpath_accum_n75));
AND2X1 mul_U18250(.A(dpath_acc_reg_in[98]), .B(n7195), .Y(dpath_accum_n77));
AND2X1 mul_U18251(.A(dpath_acc_reg_in[97]), .B(n7195), .Y(dpath_accum_n79));
AND2X1 mul_U18252(.A(dpath_acc_reg_in[96]), .B(n9592), .Y(dpath_accum_n81));
AND2X1 mul_U18253(.A(dpath_acc_reg_in[95]), .B(n9592), .Y(dpath_accum_n83));
AND2X1 mul_U18254(.A(dpath_acc_reg_in[94]), .B(n7195), .Y(dpath_accum_n85));
AND2X1 mul_U18255(.A(dpath_acc_reg_in[93]), .B(n9592), .Y(dpath_accum_n87));
AND2X1 mul_U18256(.A(dpath_acc_reg_in[92]), .B(n7195), .Y(dpath_accum_n89));
AND2X1 mul_U18257(.A(dpath_acc_reg_in[91]), .B(n9592), .Y(dpath_accum_n91));
AND2X1 mul_U18258(.A(dpath_acc_reg_in[90]), .B(n7195), .Y(dpath_accum_n93));
AND2X1 mul_U18259(.A(dpath_acc_reg_in[89]), .B(n9592), .Y(dpath_accum_n95));
AND2X1 mul_U18260(.A(dpath_acc_reg_in[88]), .B(n9592), .Y(dpath_accum_n97));
AND2X1 mul_U18261(.A(dpath_acc_reg_in[87]), .B(n9592), .Y(dpath_accum_n99));
AND2X1 mul_U18262(.A(dpath_acc_reg_in[86]), .B(n7195), .Y(dpath_accum_n101));
AND2X1 mul_U18263(.A(dpath_acc_reg_in[85]), .B(n9592), .Y(dpath_accum_n103));
AND2X1 mul_U18264(.A(dpath_acc_reg_in[84]), .B(n7195), .Y(dpath_accum_n105));
AND2X1 mul_U18265(.A(dpath_acc_reg_in[83]), .B(n9592), .Y(dpath_accum_n107));
AND2X1 mul_U18266(.A(dpath_acc_reg_in[82]), .B(n9592), .Y(dpath_accum_n109));
AND2X1 mul_U18267(.A(dpath_acc_reg_in[81]), .B(n7195), .Y(dpath_accum_n111));
AND2X1 mul_U18268(.A(dpath_acc_reg_in[80]), .B(n7195), .Y(dpath_accum_n113));
AND2X1 mul_U18269(.A(dpath_acc_reg_in[79]), .B(n7195), .Y(dpath_accum_n115));
AND2X1 mul_U18270(.A(dpath_acc_reg_in[78]), .B(n7195), .Y(dpath_accum_n117));
AND2X1 mul_U18271(.A(dpath_acc_reg_in[77]), .B(n9592), .Y(dpath_accum_n119));
AND2X1 mul_U18272(.A(dpath_acc_reg_in[76]), .B(n9592), .Y(dpath_accum_n121));
AND2X1 mul_U18273(.A(dpath_acc_reg_in[75]), .B(n7195), .Y(dpath_accum_n123));
AND2X1 mul_U18274(.A(dpath_acc_reg_in[74]), .B(n9592), .Y(dpath_accum_n125));
AND2X1 mul_U18275(.A(dpath_acc_reg_in[73]), .B(n9592), .Y(dpath_accum_n127));
AND2X1 mul_U18276(.A(dpath_acc_reg_in[72]), .B(n9592), .Y(dpath_accum_n129));
AND2X1 mul_U18277(.A(mul_spu_shf_ack), .B(n9532), .Y(dpath_dffshf_n3));
AND2X1 mul_U18278(.A(grst_l), .B(n9494), .Y(rstff_n4));
OR2X1 mul_U18279(.A(n6073), .B(n9815), .Y(n18338));
INVX1 mul_U18280(.A(n18338), .Y(mul_exu_ack));
INVX1 mul_U18281(.A(n10582), .Y(n6066));
AND2X1 mul_U18282(.A(dpath_acc_reg[129]), .B(dpath_mulcore_add_co96), .Y(n10591));
INVX1 mul_U18283(.A(n10591), .Y(n6067));
AND2X1 mul_U18284(.A(n10594), .B(dpath_acc_reg[131]), .Y(n10593));
INVX1 mul_U18285(.A(n10593), .Y(n6068));
AND2X1 mul_U18286(.A(n10596), .B(dpath_acc_reg[133]), .Y(n10597));
INVX1 mul_U18287(.A(n10597), .Y(n6069));
INVX1 mul_U18288(.A(n10603), .Y(n6070));
INVX1 mul_U18289(.A(dpath_mulcore_array2_c2[67]), .Y(n6071));
INVX1 mul_U18290(.A(dpath_mulcore_pcout[96]), .Y(n6072));
AND2X1 mul_U18291(.A(control_n20), .B(exu_mul_input_vld), .Y(control_n12));
INVX1 mul_U18292(.A(control_n12), .Y(n6073));
INVX1 mul_U18293(.A(dpath_mulcore_pcout[8]), .Y(n6074));
INVX1 mul_U18294(.A(dpath_areg[96]), .Y(n6075));
INVX1 mul_U18295(.A(dpath_areg[95]), .Y(n6076));
INVX1 mul_U18296(.A(dpath_areg[94]), .Y(n6077));
INVX1 mul_U18297(.A(dpath_areg[93]), .Y(n6078));
INVX1 mul_U18298(.A(dpath_areg[92]), .Y(n6079));
INVX1 mul_U18299(.A(dpath_areg[91]), .Y(n6080));
INVX1 mul_U18300(.A(dpath_areg[90]), .Y(n6081));
INVX1 mul_U18301(.A(dpath_areg[89]), .Y(n6082));
INVX1 mul_U18302(.A(dpath_areg[88]), .Y(n6083));
INVX1 mul_U18303(.A(dpath_areg[87]), .Y(n6084));
INVX1 mul_U18304(.A(dpath_areg[86]), .Y(n6085));
INVX1 mul_U18305(.A(dpath_areg[85]), .Y(n6086));
INVX1 mul_U18306(.A(dpath_areg[84]), .Y(n6087));
INVX1 mul_U18307(.A(dpath_areg[83]), .Y(n6088));
INVX1 mul_U18308(.A(dpath_areg[82]), .Y(n6089));
INVX1 mul_U18309(.A(dpath_areg[81]), .Y(n6090));
INVX1 mul_U18310(.A(dpath_areg[80]), .Y(n6091));
INVX1 mul_U18311(.A(dpath_areg[79]), .Y(n6092));
INVX1 mul_U18312(.A(dpath_areg[78]), .Y(n6093));
INVX1 mul_U18313(.A(dpath_areg[77]), .Y(n6094));
INVX1 mul_U18314(.A(dpath_areg[76]), .Y(n6095));
INVX1 mul_U18315(.A(dpath_areg[75]), .Y(n6096));
INVX1 mul_U18316(.A(dpath_areg[74]), .Y(n6097));
INVX1 mul_U18317(.A(dpath_areg[73]), .Y(n6098));
INVX1 mul_U18318(.A(dpath_areg[72]), .Y(n6099));
INVX1 mul_U18319(.A(dpath_areg[71]), .Y(n6100));
INVX1 mul_U18320(.A(dpath_areg[70]), .Y(n6101));
INVX1 mul_U18321(.A(dpath_areg[69]), .Y(n6102));
INVX1 mul_U18322(.A(dpath_areg[68]), .Y(n6103));
INVX1 mul_U18323(.A(dpath_areg[67]), .Y(n6104));
INVX1 mul_U18324(.A(dpath_areg[66]), .Y(n6105));
INVX1 mul_U18325(.A(dpath_areg[65]), .Y(n6106));
INVX1 mul_U18326(.A(dpath_areg[64]), .Y(n6107));
INVX1 mul_U18327(.A(dpath_areg[63]), .Y(n6108));
INVX1 mul_U18328(.A(dpath_areg[62]), .Y(n6109));
INVX1 mul_U18329(.A(dpath_areg[61]), .Y(n6110));
INVX1 mul_U18330(.A(dpath_areg[60]), .Y(n6111));
INVX1 mul_U18331(.A(dpath_areg[59]), .Y(n6112));
INVX1 mul_U18332(.A(dpath_areg[58]), .Y(n6113));
INVX1 mul_U18333(.A(dpath_areg[57]), .Y(n6114));
INVX1 mul_U18334(.A(dpath_areg[56]), .Y(n6115));
INVX1 mul_U18335(.A(dpath_areg[55]), .Y(n6116));
INVX1 mul_U18336(.A(dpath_areg[54]), .Y(n6117));
INVX1 mul_U18337(.A(dpath_areg[53]), .Y(n6118));
INVX1 mul_U18338(.A(dpath_areg[52]), .Y(n6119));
INVX1 mul_U18339(.A(dpath_areg[51]), .Y(n6120));
INVX1 mul_U18340(.A(dpath_areg[50]), .Y(n6121));
INVX1 mul_U18341(.A(dpath_areg[49]), .Y(n6122));
INVX1 mul_U18342(.A(dpath_areg[48]), .Y(n6123));
INVX1 mul_U18343(.A(dpath_areg[47]), .Y(n6124));
INVX1 mul_U18344(.A(dpath_areg[46]), .Y(n6125));
INVX1 mul_U18345(.A(dpath_areg[45]), .Y(n6126));
INVX1 mul_U18346(.A(dpath_areg[44]), .Y(n6127));
INVX1 mul_U18347(.A(dpath_areg[43]), .Y(n6128));
INVX1 mul_U18348(.A(dpath_areg[42]), .Y(n6129));
INVX1 mul_U18349(.A(dpath_areg[41]), .Y(n6130));
INVX1 mul_U18350(.A(dpath_areg[40]), .Y(n6131));
INVX1 mul_U18351(.A(dpath_areg[39]), .Y(n6132));
INVX1 mul_U18352(.A(dpath_areg[38]), .Y(n6133));
INVX1 mul_U18353(.A(dpath_areg[37]), .Y(n6134));
INVX1 mul_U18354(.A(dpath_areg[36]), .Y(n6135));
INVX1 mul_U18355(.A(dpath_areg[35]), .Y(n6136));
INVX1 mul_U18356(.A(dpath_areg[34]), .Y(n6137));
INVX1 mul_U18357(.A(dpath_areg[33]), .Y(n6138));
INVX1 mul_U18358(.A(dpath_areg[32]), .Y(n6139));
AND2X1 mul_U18359(.A(byp_imm), .B(acc_actc2), .Y(dpath_n983));
INVX1 mul_U18360(.A(dpath_n983), .Y(n6140));
INVX1 mul_U18361(.A(dpath_mulcore_pcout[29]), .Y(n6141));
INVX1 mul_U18362(.A(dpath_mulcore_pcout[28]), .Y(n6142));
INVX1 mul_U18363(.A(dpath_mulcore_pcout[27]), .Y(n6143));
INVX1 mul_U18364(.A(dpath_mulcore_pcout[26]), .Y(n6144));
INVX1 mul_U18365(.A(dpath_mulcore_pcout[25]), .Y(n6145));
INVX1 mul_U18366(.A(dpath_mulcore_pcout[24]), .Y(n6146));
INVX1 mul_U18367(.A(dpath_mulcore_pcout[23]), .Y(n6147));
INVX1 mul_U18368(.A(dpath_mulcore_pcout[22]), .Y(n6148));
INVX1 mul_U18369(.A(dpath_mulcore_pcout[21]), .Y(n6149));
INVX1 mul_U18370(.A(dpath_mulcore_pcout[20]), .Y(n6150));
INVX1 mul_U18371(.A(dpath_mulcore_pcout[4]), .Y(n6151));
INVX1 mul_U18372(.A(dpath_mulcore_pcout[3]), .Y(n6152));
INVX1 mul_U18373(.A(dpath_mulcore_pcout[2]), .Y(n6153));
INVX1 mul_U18374(.A(dpath_mulcore_pcout[1]), .Y(n6154));
INVX1 mul_U18375(.A(dpath_mulcore_pcout[14]), .Y(n6155));
INVX1 mul_U18376(.A(dpath_mulcore_pcout[13]), .Y(n6156));
INVX1 mul_U18377(.A(dpath_mulcore_pcout[12]), .Y(n6157));
INVX1 mul_U18378(.A(dpath_mulcore_pcout[11]), .Y(n6158));
INVX1 mul_U18379(.A(dpath_mulcore_pcout[10]), .Y(n6159));
INVX1 mul_U18380(.A(dpath_mulcore_pcout[9]), .Y(n6160));
INVX1 mul_U18381(.A(dpath_mulcore_pcout[7]), .Y(n6161));
INVX1 mul_U18382(.A(dpath_mulcore_pcout[6]), .Y(n6162));
INVX1 mul_U18383(.A(dpath_mulcore_pcout[5]), .Y(n6163));
INVX1 mul_U18384(.A(dpath_mulcore_pcout[19]), .Y(n6164));
INVX1 mul_U18385(.A(dpath_mulcore_pcout[18]), .Y(n6165));
INVX1 mul_U18386(.A(dpath_mulcore_pcout[17]), .Y(n6166));
INVX1 mul_U18387(.A(dpath_mulcore_pcout[16]), .Y(n6167));
AND2X1 mul_U18388(.A(dpath_mulcore_ary1_a1_I2_I2_p2_l_67), .B(n9478), .Y(n14782));
INVX1 mul_U18389(.A(n14782), .Y(n6168));
AND2X1 mul_U18390(.A(dpath_mulcore_b7[1]), .B(n10606), .Y(dpath_mulcore_ary1_a0_I2_I2_p1_l_65));
INVX1 mul_U18391(.A(dpath_mulcore_ary1_a0_I2_I2_p1_l_65), .Y(n6169));
AND2X1 mul_U18392(.A(dpath_mulcore_b7[1]), .B(n10609), .Y(dpath_mulcore_ary1_a0_I2_I2_p1_l_64));
INVX1 mul_U18393(.A(dpath_mulcore_ary1_a0_I2_I2_p1_l_64), .Y(n6170));
AND2X1 mul_U18394(.A(dpath_mulcore_b7[1]), .B(n10612), .Y(dpath_mulcore_ary1_a0_I2_p1_l[63]));
INVX1 mul_U18395(.A(dpath_mulcore_ary1_a0_I2_p1_l[63]), .Y(n6171));
AND2X1 mul_U18396(.A(dpath_mulcore_b6[1]), .B(n10615), .Y(dpath_mulcore_ary1_a0_I2_p0_l[63]));
INVX1 mul_U18397(.A(dpath_mulcore_ary1_a0_I2_p0_l[63]), .Y(n6172));
AND2X1 mul_U18398(.A(dpath_mulcore_b7[1]), .B(n10618), .Y(dpath_mulcore_ary1_a0_I2_p1_l[62]));
INVX1 mul_U18399(.A(dpath_mulcore_ary1_a0_I2_p1_l[62]), .Y(n6173));
AND2X1 mul_U18400(.A(dpath_mulcore_b6[1]), .B(n10621), .Y(dpath_mulcore_ary1_a0_I2_p0_l[62]));
INVX1 mul_U18401(.A(dpath_mulcore_ary1_a0_I2_p0_l[62]), .Y(n6174));
AND2X1 mul_U18402(.A(dpath_mulcore_b7[1]), .B(n10624), .Y(dpath_mulcore_ary1_a0_I2_p1_l[61]));
INVX1 mul_U18403(.A(dpath_mulcore_ary1_a0_I2_p1_l[61]), .Y(n6175));
AND2X1 mul_U18404(.A(dpath_mulcore_b6[1]), .B(n10627), .Y(dpath_mulcore_ary1_a0_I2_p0_l[61]));
INVX1 mul_U18405(.A(dpath_mulcore_ary1_a0_I2_p0_l[61]), .Y(n6176));
AND2X1 mul_U18406(.A(dpath_mulcore_b7[1]), .B(n10630), .Y(dpath_mulcore_ary1_a0_I2_p1_l[60]));
INVX1 mul_U18407(.A(dpath_mulcore_ary1_a0_I2_p1_l[60]), .Y(n6177));
AND2X1 mul_U18408(.A(dpath_mulcore_b6[1]), .B(n10633), .Y(dpath_mulcore_ary1_a0_I2_p0_l[60]));
INVX1 mul_U18409(.A(dpath_mulcore_ary1_a0_I2_p0_l[60]), .Y(n6178));
AND2X1 mul_U18410(.A(dpath_mulcore_b7[1]), .B(n10636), .Y(dpath_mulcore_ary1_a0_I2_p1_l[59]));
INVX1 mul_U18411(.A(dpath_mulcore_ary1_a0_I2_p1_l[59]), .Y(n6179));
AND2X1 mul_U18412(.A(dpath_mulcore_b6[1]), .B(n10639), .Y(dpath_mulcore_ary1_a0_I2_p0_l[59]));
INVX1 mul_U18413(.A(dpath_mulcore_ary1_a0_I2_p0_l[59]), .Y(n6180));
AND2X1 mul_U18414(.A(dpath_mulcore_b7[1]), .B(n10642), .Y(dpath_mulcore_ary1_a0_I2_p1_l[58]));
INVX1 mul_U18415(.A(dpath_mulcore_ary1_a0_I2_p1_l[58]), .Y(n6181));
AND2X1 mul_U18416(.A(dpath_mulcore_b6[1]), .B(n10645), .Y(dpath_mulcore_ary1_a0_I2_p0_l[58]));
INVX1 mul_U18417(.A(dpath_mulcore_ary1_a0_I2_p0_l[58]), .Y(n6182));
AND2X1 mul_U18418(.A(dpath_mulcore_b7[1]), .B(n10648), .Y(dpath_mulcore_ary1_a0_I2_p1_l[57]));
INVX1 mul_U18419(.A(dpath_mulcore_ary1_a0_I2_p1_l[57]), .Y(n6183));
AND2X1 mul_U18420(.A(dpath_mulcore_b6[1]), .B(n10651), .Y(dpath_mulcore_ary1_a0_I2_p0_l[57]));
INVX1 mul_U18421(.A(dpath_mulcore_ary1_a0_I2_p0_l[57]), .Y(n6184));
AND2X1 mul_U18422(.A(dpath_mulcore_b7[1]), .B(n10654), .Y(dpath_mulcore_ary1_a0_I2_p1_l[56]));
INVX1 mul_U18423(.A(dpath_mulcore_ary1_a0_I2_p1_l[56]), .Y(n6185));
AND2X1 mul_U18424(.A(dpath_mulcore_b6[1]), .B(n10657), .Y(dpath_mulcore_ary1_a0_I2_p0_l[56]));
INVX1 mul_U18425(.A(dpath_mulcore_ary1_a0_I2_p0_l[56]), .Y(n6186));
AND2X1 mul_U18426(.A(dpath_mulcore_b7[1]), .B(n10660), .Y(dpath_mulcore_ary1_a0_I2_p1_l[55]));
INVX1 mul_U18427(.A(dpath_mulcore_ary1_a0_I2_p1_l[55]), .Y(n6187));
AND2X1 mul_U18428(.A(dpath_mulcore_b6[1]), .B(n10663), .Y(dpath_mulcore_ary1_a0_I2_p0_l[55]));
INVX1 mul_U18429(.A(dpath_mulcore_ary1_a0_I2_p0_l[55]), .Y(n6188));
AND2X1 mul_U18430(.A(dpath_mulcore_b7[1]), .B(n10666), .Y(dpath_mulcore_ary1_a0_I2_p1_l[54]));
INVX1 mul_U18431(.A(dpath_mulcore_ary1_a0_I2_p1_l[54]), .Y(n6189));
AND2X1 mul_U18432(.A(dpath_mulcore_b6[1]), .B(n10669), .Y(dpath_mulcore_ary1_a0_I2_p0_l[54]));
INVX1 mul_U18433(.A(dpath_mulcore_ary1_a0_I2_p0_l[54]), .Y(n6190));
AND2X1 mul_U18434(.A(dpath_mulcore_b7[1]), .B(n10672), .Y(dpath_mulcore_ary1_a0_I2_p1_l[53]));
INVX1 mul_U18435(.A(dpath_mulcore_ary1_a0_I2_p1_l[53]), .Y(n6191));
AND2X1 mul_U18436(.A(dpath_mulcore_b6[1]), .B(n10675), .Y(dpath_mulcore_ary1_a0_I2_p0_l[53]));
INVX1 mul_U18437(.A(dpath_mulcore_ary1_a0_I2_p0_l[53]), .Y(n6192));
AND2X1 mul_U18438(.A(dpath_mulcore_b7[1]), .B(n10678), .Y(dpath_mulcore_ary1_a0_I2_p1_l[52]));
INVX1 mul_U18439(.A(dpath_mulcore_ary1_a0_I2_p1_l[52]), .Y(n6193));
AND2X1 mul_U18440(.A(dpath_mulcore_b6[1]), .B(n10681), .Y(dpath_mulcore_ary1_a0_I2_p0_l[52]));
INVX1 mul_U18441(.A(dpath_mulcore_ary1_a0_I2_p0_l[52]), .Y(n6194));
AND2X1 mul_U18442(.A(dpath_mulcore_b7[1]), .B(n10684), .Y(dpath_mulcore_ary1_a0_I2_p1_l[51]));
INVX1 mul_U18443(.A(dpath_mulcore_ary1_a0_I2_p1_l[51]), .Y(n6195));
AND2X1 mul_U18444(.A(dpath_mulcore_b6[1]), .B(n10687), .Y(dpath_mulcore_ary1_a0_I2_p0_l[51]));
INVX1 mul_U18445(.A(dpath_mulcore_ary1_a0_I2_p0_l[51]), .Y(n6196));
AND2X1 mul_U18446(.A(dpath_mulcore_b7[1]), .B(n10690), .Y(dpath_mulcore_ary1_a0_I2_p1_l[50]));
INVX1 mul_U18447(.A(dpath_mulcore_ary1_a0_I2_p1_l[50]), .Y(n6197));
AND2X1 mul_U18448(.A(dpath_mulcore_b6[1]), .B(n10693), .Y(dpath_mulcore_ary1_a0_I2_p0_l[50]));
INVX1 mul_U18449(.A(dpath_mulcore_ary1_a0_I2_p0_l[50]), .Y(n6198));
AND2X1 mul_U18450(.A(dpath_mulcore_b7[1]), .B(n10696), .Y(dpath_mulcore_ary1_a0_I2_p1_l[49]));
INVX1 mul_U18451(.A(dpath_mulcore_ary1_a0_I2_p1_l[49]), .Y(n6199));
AND2X1 mul_U18452(.A(dpath_mulcore_b6[1]), .B(n10699), .Y(dpath_mulcore_ary1_a0_I2_p0_l[49]));
INVX1 mul_U18453(.A(dpath_mulcore_ary1_a0_I2_p0_l[49]), .Y(n6200));
AND2X1 mul_U18454(.A(dpath_mulcore_b7[1]), .B(n10702), .Y(dpath_mulcore_ary1_a0_I2_p1_l[48]));
INVX1 mul_U18455(.A(dpath_mulcore_ary1_a0_I2_p1_l[48]), .Y(n6201));
AND2X1 mul_U18456(.A(dpath_mulcore_b6[1]), .B(n10705), .Y(dpath_mulcore_ary1_a0_I2_p0_l[48]));
INVX1 mul_U18457(.A(dpath_mulcore_ary1_a0_I2_p0_l[48]), .Y(n6202));
AND2X1 mul_U18458(.A(dpath_mulcore_b7[1]), .B(n10708), .Y(dpath_mulcore_ary1_a0_I2_p1_l[47]));
INVX1 mul_U18459(.A(dpath_mulcore_ary1_a0_I2_p1_l[47]), .Y(n6203));
AND2X1 mul_U18460(.A(dpath_mulcore_b6[1]), .B(n10711), .Y(dpath_mulcore_ary1_a0_I2_p0_l[47]));
INVX1 mul_U18461(.A(dpath_mulcore_ary1_a0_I2_p0_l[47]), .Y(n6204));
AND2X1 mul_U18462(.A(dpath_mulcore_b7[1]), .B(n10714), .Y(dpath_mulcore_ary1_a0_I2_p1_l[46]));
INVX1 mul_U18463(.A(dpath_mulcore_ary1_a0_I2_p1_l[46]), .Y(n6205));
AND2X1 mul_U18464(.A(dpath_mulcore_b6[1]), .B(n10717), .Y(dpath_mulcore_ary1_a0_I2_p0_l[46]));
INVX1 mul_U18465(.A(dpath_mulcore_ary1_a0_I2_p0_l[46]), .Y(n6206));
AND2X1 mul_U18466(.A(dpath_mulcore_b7[1]), .B(n10720), .Y(dpath_mulcore_ary1_a0_I2_p1_l[45]));
INVX1 mul_U18467(.A(dpath_mulcore_ary1_a0_I2_p1_l[45]), .Y(n6207));
AND2X1 mul_U18468(.A(dpath_mulcore_b6[1]), .B(n10723), .Y(dpath_mulcore_ary1_a0_I2_p0_l[45]));
INVX1 mul_U18469(.A(dpath_mulcore_ary1_a0_I2_p0_l[45]), .Y(n6208));
AND2X1 mul_U18470(.A(dpath_mulcore_b7[1]), .B(n10726), .Y(dpath_mulcore_ary1_a0_I2_p1_l[44]));
INVX1 mul_U18471(.A(dpath_mulcore_ary1_a0_I2_p1_l[44]), .Y(n6209));
AND2X1 mul_U18472(.A(dpath_mulcore_b6[1]), .B(n10729), .Y(dpath_mulcore_ary1_a0_I2_p0_l[44]));
INVX1 mul_U18473(.A(dpath_mulcore_ary1_a0_I2_p0_l[44]), .Y(n6210));
AND2X1 mul_U18474(.A(dpath_mulcore_b7[1]), .B(n10732), .Y(dpath_mulcore_ary1_a0_I2_p1_l[43]));
INVX1 mul_U18475(.A(dpath_mulcore_ary1_a0_I2_p1_l[43]), .Y(n6211));
AND2X1 mul_U18476(.A(dpath_mulcore_b6[1]), .B(n10735), .Y(dpath_mulcore_ary1_a0_I2_p0_l[43]));
INVX1 mul_U18477(.A(dpath_mulcore_ary1_a0_I2_p0_l[43]), .Y(n6212));
AND2X1 mul_U18478(.A(dpath_mulcore_b7[1]), .B(n10738), .Y(dpath_mulcore_ary1_a0_I2_p1_l[42]));
INVX1 mul_U18479(.A(dpath_mulcore_ary1_a0_I2_p1_l[42]), .Y(n6213));
AND2X1 mul_U18480(.A(dpath_mulcore_b6[1]), .B(n10741), .Y(dpath_mulcore_ary1_a0_I2_p0_l[42]));
INVX1 mul_U18481(.A(dpath_mulcore_ary1_a0_I2_p0_l[42]), .Y(n6214));
AND2X1 mul_U18482(.A(dpath_mulcore_b7[1]), .B(n10744), .Y(dpath_mulcore_ary1_a0_I2_p1_l[41]));
INVX1 mul_U18483(.A(dpath_mulcore_ary1_a0_I2_p1_l[41]), .Y(n6215));
AND2X1 mul_U18484(.A(dpath_mulcore_b6[1]), .B(n10747), .Y(dpath_mulcore_ary1_a0_I2_p0_l[41]));
INVX1 mul_U18485(.A(dpath_mulcore_ary1_a0_I2_p0_l[41]), .Y(n6216));
AND2X1 mul_U18486(.A(dpath_mulcore_b7[1]), .B(n10750), .Y(dpath_mulcore_ary1_a0_I2_p1_l[40]));
INVX1 mul_U18487(.A(dpath_mulcore_ary1_a0_I2_p1_l[40]), .Y(n6217));
AND2X1 mul_U18488(.A(dpath_mulcore_b6[1]), .B(n10753), .Y(dpath_mulcore_ary1_a0_I2_p0_l[40]));
INVX1 mul_U18489(.A(dpath_mulcore_ary1_a0_I2_p0_l[40]), .Y(n6218));
AND2X1 mul_U18490(.A(dpath_mulcore_b7[1]), .B(n10756), .Y(dpath_mulcore_ary1_a0_I2_p1_l[39]));
INVX1 mul_U18491(.A(dpath_mulcore_ary1_a0_I2_p1_l[39]), .Y(n6219));
AND2X1 mul_U18492(.A(dpath_mulcore_b6[1]), .B(n10759), .Y(dpath_mulcore_ary1_a0_I2_p0_l[39]));
INVX1 mul_U18493(.A(dpath_mulcore_ary1_a0_I2_p0_l[39]), .Y(n6220));
AND2X1 mul_U18494(.A(dpath_mulcore_b7[1]), .B(n10762), .Y(dpath_mulcore_ary1_a0_I2_p1_l[38]));
INVX1 mul_U18495(.A(dpath_mulcore_ary1_a0_I2_p1_l[38]), .Y(n6221));
AND2X1 mul_U18496(.A(dpath_mulcore_b6[1]), .B(n10765), .Y(dpath_mulcore_ary1_a0_I2_p0_l[38]));
INVX1 mul_U18497(.A(dpath_mulcore_ary1_a0_I2_p0_l[38]), .Y(n6222));
AND2X1 mul_U18498(.A(dpath_mulcore_b7[1]), .B(n10768), .Y(dpath_mulcore_ary1_a0_I2_p1_l[37]));
INVX1 mul_U18499(.A(dpath_mulcore_ary1_a0_I2_p1_l[37]), .Y(n6223));
AND2X1 mul_U18500(.A(dpath_mulcore_b6[1]), .B(n10771), .Y(dpath_mulcore_ary1_a0_I2_p0_l[37]));
INVX1 mul_U18501(.A(dpath_mulcore_ary1_a0_I2_p0_l[37]), .Y(n6224));
AND2X1 mul_U18502(.A(dpath_mulcore_b7[1]), .B(n10774), .Y(dpath_mulcore_ary1_a0_I2_p1_l[36]));
INVX1 mul_U18503(.A(dpath_mulcore_ary1_a0_I2_p1_l[36]), .Y(n6225));
AND2X1 mul_U18504(.A(dpath_mulcore_b6[1]), .B(n10777), .Y(dpath_mulcore_ary1_a0_I2_p0_l[36]));
INVX1 mul_U18505(.A(dpath_mulcore_ary1_a0_I2_p0_l[36]), .Y(n6226));
AND2X1 mul_U18506(.A(dpath_mulcore_b7[1]), .B(n10780), .Y(dpath_mulcore_ary1_a0_I2_p1_l[35]));
INVX1 mul_U18507(.A(dpath_mulcore_ary1_a0_I2_p1_l[35]), .Y(n6227));
AND2X1 mul_U18508(.A(dpath_mulcore_b6[1]), .B(n10783), .Y(dpath_mulcore_ary1_a0_I2_p0_l[35]));
INVX1 mul_U18509(.A(dpath_mulcore_ary1_a0_I2_p0_l[35]), .Y(n6228));
AND2X1 mul_U18510(.A(dpath_mulcore_b7[1]), .B(n10786), .Y(dpath_mulcore_ary1_a0_I2_p1_l[34]));
INVX1 mul_U18511(.A(dpath_mulcore_ary1_a0_I2_p1_l[34]), .Y(n6229));
AND2X1 mul_U18512(.A(dpath_mulcore_b6[1]), .B(n10789), .Y(dpath_mulcore_ary1_a0_I2_p0_l[34]));
INVX1 mul_U18513(.A(dpath_mulcore_ary1_a0_I2_p0_l[34]), .Y(n6230));
AND2X1 mul_U18514(.A(dpath_mulcore_b7[1]), .B(n10792), .Y(dpath_mulcore_ary1_a0_I2_p1_l[33]));
INVX1 mul_U18515(.A(dpath_mulcore_ary1_a0_I2_p1_l[33]), .Y(n6231));
AND2X1 mul_U18516(.A(dpath_mulcore_b6[1]), .B(n10795), .Y(dpath_mulcore_ary1_a0_I2_p0_l[33]));
INVX1 mul_U18517(.A(dpath_mulcore_ary1_a0_I2_p0_l[33]), .Y(n6232));
AND2X1 mul_U18518(.A(dpath_mulcore_b7[1]), .B(n10798), .Y(dpath_mulcore_ary1_a0_I2_p1_l[32]));
INVX1 mul_U18519(.A(dpath_mulcore_ary1_a0_I2_p1_l[32]), .Y(n6233));
AND2X1 mul_U18520(.A(dpath_mulcore_b6[1]), .B(n10801), .Y(dpath_mulcore_ary1_a0_I2_p0_l[32]));
INVX1 mul_U18521(.A(dpath_mulcore_ary1_a0_I2_p0_l[32]), .Y(n6234));
AND2X1 mul_U18522(.A(dpath_mulcore_b7[1]), .B(n10804), .Y(dpath_mulcore_ary1_a0_I2_p1_l[31]));
INVX1 mul_U18523(.A(dpath_mulcore_ary1_a0_I2_p1_l[31]), .Y(n6235));
AND2X1 mul_U18524(.A(dpath_mulcore_b6[1]), .B(n10807), .Y(dpath_mulcore_ary1_a0_I2_p0_l[31]));
INVX1 mul_U18525(.A(dpath_mulcore_ary1_a0_I2_p0_l[31]), .Y(n6236));
AND2X1 mul_U18526(.A(dpath_mulcore_b7[1]), .B(n10810), .Y(dpath_mulcore_ary1_a0_I2_p1_l[30]));
INVX1 mul_U18527(.A(dpath_mulcore_ary1_a0_I2_p1_l[30]), .Y(n6237));
AND2X1 mul_U18528(.A(dpath_mulcore_b6[1]), .B(n10813), .Y(dpath_mulcore_ary1_a0_I2_p0_l[30]));
INVX1 mul_U18529(.A(dpath_mulcore_ary1_a0_I2_p0_l[30]), .Y(n6238));
AND2X1 mul_U18530(.A(dpath_mulcore_b7[1]), .B(n10816), .Y(dpath_mulcore_ary1_a0_I2_p1_l[29]));
INVX1 mul_U18531(.A(dpath_mulcore_ary1_a0_I2_p1_l[29]), .Y(n6239));
AND2X1 mul_U18532(.A(dpath_mulcore_b6[1]), .B(n10819), .Y(dpath_mulcore_ary1_a0_I2_p0_l[29]));
INVX1 mul_U18533(.A(dpath_mulcore_ary1_a0_I2_p0_l[29]), .Y(n6240));
AND2X1 mul_U18534(.A(dpath_mulcore_b7[1]), .B(n10822), .Y(dpath_mulcore_ary1_a0_I2_p1_l[28]));
INVX1 mul_U18535(.A(dpath_mulcore_ary1_a0_I2_p1_l[28]), .Y(n6241));
AND2X1 mul_U18536(.A(dpath_mulcore_b6[1]), .B(n10825), .Y(dpath_mulcore_ary1_a0_I2_p0_l[28]));
INVX1 mul_U18537(.A(dpath_mulcore_ary1_a0_I2_p0_l[28]), .Y(n6242));
AND2X1 mul_U18538(.A(dpath_mulcore_b7[1]), .B(n10828), .Y(dpath_mulcore_ary1_a0_I2_p1_l[27]));
INVX1 mul_U18539(.A(dpath_mulcore_ary1_a0_I2_p1_l[27]), .Y(n6243));
AND2X1 mul_U18540(.A(dpath_mulcore_b6[1]), .B(n10831), .Y(dpath_mulcore_ary1_a0_I2_p0_l[27]));
INVX1 mul_U18541(.A(dpath_mulcore_ary1_a0_I2_p0_l[27]), .Y(n6244));
AND2X1 mul_U18542(.A(dpath_mulcore_b7[1]), .B(n10834), .Y(dpath_mulcore_ary1_a0_I2_p1_l[26]));
INVX1 mul_U18543(.A(dpath_mulcore_ary1_a0_I2_p1_l[26]), .Y(n6245));
AND2X1 mul_U18544(.A(dpath_mulcore_b6[1]), .B(n10837), .Y(dpath_mulcore_ary1_a0_I2_p0_l[26]));
INVX1 mul_U18545(.A(dpath_mulcore_ary1_a0_I2_p0_l[26]), .Y(n6246));
AND2X1 mul_U18546(.A(dpath_mulcore_b7[1]), .B(n10840), .Y(dpath_mulcore_ary1_a0_I2_p1_l[25]));
INVX1 mul_U18547(.A(dpath_mulcore_ary1_a0_I2_p1_l[25]), .Y(n6247));
AND2X1 mul_U18548(.A(dpath_mulcore_b6[1]), .B(n10843), .Y(dpath_mulcore_ary1_a0_I2_p0_l[25]));
INVX1 mul_U18549(.A(dpath_mulcore_ary1_a0_I2_p0_l[25]), .Y(n6248));
AND2X1 mul_U18550(.A(dpath_mulcore_b7[1]), .B(n10846), .Y(dpath_mulcore_ary1_a0_I2_p1_l[24]));
INVX1 mul_U18551(.A(dpath_mulcore_ary1_a0_I2_p1_l[24]), .Y(n6249));
AND2X1 mul_U18552(.A(dpath_mulcore_b6[1]), .B(n10849), .Y(dpath_mulcore_ary1_a0_I2_p0_l[24]));
INVX1 mul_U18553(.A(dpath_mulcore_ary1_a0_I2_p0_l[24]), .Y(n6250));
AND2X1 mul_U18554(.A(dpath_mulcore_b7[1]), .B(n10852), .Y(dpath_mulcore_ary1_a0_I2_p1_l[23]));
INVX1 mul_U18555(.A(dpath_mulcore_ary1_a0_I2_p1_l[23]), .Y(n6251));
AND2X1 mul_U18556(.A(dpath_mulcore_b6[1]), .B(n10855), .Y(dpath_mulcore_ary1_a0_I2_p0_l[23]));
INVX1 mul_U18557(.A(dpath_mulcore_ary1_a0_I2_p0_l[23]), .Y(n6252));
AND2X1 mul_U18558(.A(dpath_mulcore_b7[1]), .B(n10858), .Y(dpath_mulcore_ary1_a0_I2_p1_l[22]));
INVX1 mul_U18559(.A(dpath_mulcore_ary1_a0_I2_p1_l[22]), .Y(n6253));
AND2X1 mul_U18560(.A(dpath_mulcore_b6[1]), .B(n10861), .Y(dpath_mulcore_ary1_a0_I2_p0_l[22]));
INVX1 mul_U18561(.A(dpath_mulcore_ary1_a0_I2_p0_l[22]), .Y(n6254));
AND2X1 mul_U18562(.A(dpath_mulcore_b7[1]), .B(n10864), .Y(dpath_mulcore_ary1_a0_I2_p1_l[21]));
INVX1 mul_U18563(.A(dpath_mulcore_ary1_a0_I2_p1_l[21]), .Y(n6255));
AND2X1 mul_U18564(.A(dpath_mulcore_b6[1]), .B(n10867), .Y(dpath_mulcore_ary1_a0_I2_p0_l[21]));
INVX1 mul_U18565(.A(dpath_mulcore_ary1_a0_I2_p0_l[21]), .Y(n6256));
AND2X1 mul_U18566(.A(dpath_mulcore_b7[1]), .B(n10870), .Y(dpath_mulcore_ary1_a0_I2_p1_l[20]));
INVX1 mul_U18567(.A(dpath_mulcore_ary1_a0_I2_p1_l[20]), .Y(n6257));
AND2X1 mul_U18568(.A(dpath_mulcore_b6[1]), .B(n10873), .Y(dpath_mulcore_ary1_a0_I2_p0_l[20]));
INVX1 mul_U18569(.A(dpath_mulcore_ary1_a0_I2_p0_l[20]), .Y(n6258));
AND2X1 mul_U18570(.A(dpath_mulcore_b7[1]), .B(n10876), .Y(dpath_mulcore_ary1_a0_I2_p1_l[19]));
INVX1 mul_U18571(.A(dpath_mulcore_ary1_a0_I2_p1_l[19]), .Y(n6259));
AND2X1 mul_U18572(.A(dpath_mulcore_b6[1]), .B(n10879), .Y(dpath_mulcore_ary1_a0_I2_p0_l[19]));
INVX1 mul_U18573(.A(dpath_mulcore_ary1_a0_I2_p0_l[19]), .Y(n6260));
AND2X1 mul_U18574(.A(dpath_mulcore_b7[1]), .B(n10882), .Y(dpath_mulcore_ary1_a0_I2_p1_l[18]));
INVX1 mul_U18575(.A(dpath_mulcore_ary1_a0_I2_p1_l[18]), .Y(n6261));
AND2X1 mul_U18576(.A(dpath_mulcore_b6[1]), .B(n10885), .Y(dpath_mulcore_ary1_a0_I2_p0_l[18]));
INVX1 mul_U18577(.A(dpath_mulcore_ary1_a0_I2_p0_l[18]), .Y(n6262));
AND2X1 mul_U18578(.A(dpath_mulcore_b7[1]), .B(n10888), .Y(dpath_mulcore_ary1_a0_I2_p1_l[17]));
INVX1 mul_U18579(.A(dpath_mulcore_ary1_a0_I2_p1_l[17]), .Y(n6263));
AND2X1 mul_U18580(.A(dpath_mulcore_b6[1]), .B(n10891), .Y(dpath_mulcore_ary1_a0_I2_p0_l[17]));
INVX1 mul_U18581(.A(dpath_mulcore_ary1_a0_I2_p0_l[17]), .Y(n6264));
AND2X1 mul_U18582(.A(dpath_mulcore_b7[1]), .B(n10894), .Y(dpath_mulcore_ary1_a0_I2_p1_l[16]));
INVX1 mul_U18583(.A(dpath_mulcore_ary1_a0_I2_p1_l[16]), .Y(n6265));
AND2X1 mul_U18584(.A(dpath_mulcore_b6[1]), .B(n10897), .Y(dpath_mulcore_ary1_a0_I2_p0_l[16]));
INVX1 mul_U18585(.A(dpath_mulcore_ary1_a0_I2_p0_l[16]), .Y(n6266));
AND2X1 mul_U18586(.A(dpath_mulcore_b7[1]), .B(n10900), .Y(dpath_mulcore_ary1_a0_I2_p1_l[15]));
INVX1 mul_U18587(.A(dpath_mulcore_ary1_a0_I2_p1_l[15]), .Y(n6267));
AND2X1 mul_U18588(.A(dpath_mulcore_b6[1]), .B(n10903), .Y(dpath_mulcore_ary1_a0_I2_p0_l[15]));
INVX1 mul_U18589(.A(dpath_mulcore_ary1_a0_I2_p0_l[15]), .Y(n6268));
AND2X1 mul_U18590(.A(dpath_mulcore_b7[1]), .B(n10906), .Y(dpath_mulcore_ary1_a0_I2_p1_l[14]));
INVX1 mul_U18591(.A(dpath_mulcore_ary1_a0_I2_p1_l[14]), .Y(n6269));
AND2X1 mul_U18592(.A(dpath_mulcore_b6[1]), .B(n10909), .Y(dpath_mulcore_ary1_a0_I2_p0_l[14]));
INVX1 mul_U18593(.A(dpath_mulcore_ary1_a0_I2_p0_l[14]), .Y(n6270));
AND2X1 mul_U18594(.A(dpath_mulcore_b7[1]), .B(n10912), .Y(dpath_mulcore_ary1_a0_I2_p1_l[13]));
INVX1 mul_U18595(.A(dpath_mulcore_ary1_a0_I2_p1_l[13]), .Y(n6271));
AND2X1 mul_U18596(.A(dpath_mulcore_b6[1]), .B(n10915), .Y(dpath_mulcore_ary1_a0_I2_p0_l[13]));
INVX1 mul_U18597(.A(dpath_mulcore_ary1_a0_I2_p0_l[13]), .Y(n6272));
AND2X1 mul_U18598(.A(dpath_mulcore_b7[1]), .B(n10918), .Y(dpath_mulcore_ary1_a0_I2_p1_l[12]));
INVX1 mul_U18599(.A(dpath_mulcore_ary1_a0_I2_p1_l[12]), .Y(n6273));
AND2X1 mul_U18600(.A(dpath_mulcore_b6[1]), .B(n10921), .Y(dpath_mulcore_ary1_a0_I2_p0_l[12]));
INVX1 mul_U18601(.A(dpath_mulcore_ary1_a0_I2_p0_l[12]), .Y(n6274));
AND2X1 mul_U18602(.A(dpath_mulcore_b7[1]), .B(n10924), .Y(dpath_mulcore_ary1_a0_I2_p1_l[11]));
INVX1 mul_U18603(.A(dpath_mulcore_ary1_a0_I2_p1_l[11]), .Y(n6275));
AND2X1 mul_U18604(.A(dpath_mulcore_b6[1]), .B(n10927), .Y(dpath_mulcore_ary1_a0_I2_p0_l[11]));
INVX1 mul_U18605(.A(dpath_mulcore_ary1_a0_I2_p0_l[11]), .Y(n6276));
AND2X1 mul_U18606(.A(dpath_mulcore_b7[1]), .B(n10930), .Y(dpath_mulcore_ary1_a0_I2_p1_l[10]));
INVX1 mul_U18607(.A(dpath_mulcore_ary1_a0_I2_p1_l[10]), .Y(n6277));
AND2X1 mul_U18608(.A(dpath_mulcore_b6[1]), .B(n10933), .Y(dpath_mulcore_ary1_a0_I2_p0_l[10]));
INVX1 mul_U18609(.A(dpath_mulcore_ary1_a0_I2_p0_l[10]), .Y(n6278));
AND2X1 mul_U18610(.A(dpath_mulcore_b7[1]), .B(n10936), .Y(dpath_mulcore_ary1_a0_I2_p1_l[9]));
INVX1 mul_U18611(.A(dpath_mulcore_ary1_a0_I2_p1_l[9]), .Y(n6279));
AND2X1 mul_U18612(.A(dpath_mulcore_b6[1]), .B(n10939), .Y(dpath_mulcore_ary1_a0_I2_p0_l[9]));
INVX1 mul_U18613(.A(dpath_mulcore_ary1_a0_I2_p0_l[9]), .Y(n6280));
AND2X1 mul_U18614(.A(dpath_mulcore_b7[1]), .B(n10942), .Y(dpath_mulcore_ary1_a0_I2_p1_l[8]));
INVX1 mul_U18615(.A(dpath_mulcore_ary1_a0_I2_p1_l[8]), .Y(n6281));
AND2X1 mul_U18616(.A(dpath_mulcore_b6[1]), .B(n10945), .Y(dpath_mulcore_ary1_a0_I2_p0_l[8]));
INVX1 mul_U18617(.A(dpath_mulcore_ary1_a0_I2_p0_l[8]), .Y(n6282));
AND2X1 mul_U18618(.A(dpath_mulcore_b7[1]), .B(n10948), .Y(dpath_mulcore_ary1_a0_I2_p1_l[7]));
INVX1 mul_U18619(.A(dpath_mulcore_ary1_a0_I2_p1_l[7]), .Y(n6283));
AND2X1 mul_U18620(.A(dpath_mulcore_b6[1]), .B(n10951), .Y(dpath_mulcore_ary1_a0_I2_p0_l[7]));
INVX1 mul_U18621(.A(dpath_mulcore_ary1_a0_I2_p0_l[7]), .Y(n6284));
AND2X1 mul_U18622(.A(dpath_mulcore_b7[1]), .B(n10954), .Y(dpath_mulcore_ary1_a0_I2_p1_l[6]));
INVX1 mul_U18623(.A(dpath_mulcore_ary1_a0_I2_p1_l[6]), .Y(n6285));
AND2X1 mul_U18624(.A(dpath_mulcore_b6[1]), .B(n10957), .Y(dpath_mulcore_ary1_a0_I2_p0_l[6]));
INVX1 mul_U18625(.A(dpath_mulcore_ary1_a0_I2_p0_l[6]), .Y(n6286));
AND2X1 mul_U18626(.A(dpath_mulcore_b7[1]), .B(n10960), .Y(dpath_mulcore_ary1_a0_I2_p1_l[5]));
INVX1 mul_U18627(.A(dpath_mulcore_ary1_a0_I2_p1_l[5]), .Y(n6287));
AND2X1 mul_U18628(.A(dpath_mulcore_b6[1]), .B(n10963), .Y(dpath_mulcore_ary1_a0_I2_p0_l[5]));
INVX1 mul_U18629(.A(dpath_mulcore_ary1_a0_I2_p0_l[5]), .Y(n6288));
AND2X1 mul_U18630(.A(dpath_mulcore_b7[1]), .B(n10966), .Y(dpath_mulcore_ary1_a0_I2_p1_l[4]));
INVX1 mul_U18631(.A(dpath_mulcore_ary1_a0_I2_p1_l[4]), .Y(n6289));
AND2X1 mul_U18632(.A(dpath_mulcore_b6[1]), .B(n10969), .Y(dpath_mulcore_ary1_a0_I2_p0_l[4]));
INVX1 mul_U18633(.A(dpath_mulcore_ary1_a0_I2_p0_l[4]), .Y(n6290));
AND2X1 mul_U18634(.A(dpath_mulcore_b6[1]), .B(n10972), .Y(dpath_mulcore_ary1_a0_I2_p0_l[3]));
INVX1 mul_U18635(.A(dpath_mulcore_ary1_a0_I2_p0_l[3]), .Y(n6291));
AND2X1 mul_U18636(.A(dpath_mulcore_b7[1]), .B(n10975), .Y(dpath_mulcore_ary1_a0_I2_p1_l[3]));
INVX1 mul_U18637(.A(dpath_mulcore_ary1_a0_I2_p1_l[3]), .Y(n6292));
AND2X1 mul_U18638(.A(dpath_mulcore_b6[1]), .B(n10978), .Y(dpath_mulcore_ary1_a0_I2_I0_p0_l_2));
INVX1 mul_U18639(.A(dpath_mulcore_ary1_a0_I2_I0_p0_l_2), .Y(n6293));
AND2X1 mul_U18640(.A(dpath_mulcore_b6[1]), .B(n10981), .Y(dpath_mulcore_ary1_a0_I2_I0_p0_l_1));
INVX1 mul_U18641(.A(dpath_mulcore_ary1_a0_I2_I0_p0_l_1), .Y(n6294));
AND2X1 mul_U18642(.A(dpath_mulcore_b6[1]), .B(n10983), .Y(dpath_mulcore_ary1_a0_I2_I0_p0_l_0));
INVX1 mul_U18643(.A(dpath_mulcore_ary1_a0_I2_I0_p0_l_0), .Y(n6295));
AND2X1 mul_U18644(.A(dpath_mulcore_b7[1]), .B(n10985), .Y(dpath_mulcore_ary1_a0_I2_I0_p1_l_2));
INVX1 mul_U18645(.A(dpath_mulcore_ary1_a0_I2_I0_p1_l_2), .Y(n6296));
AND2X1 mul_U18646(.A(dpath_mulcore_b5[1]), .B(n10988), .Y(dpath_mulcore_ary1_a0_I1_I2_p2_l_67));
INVX1 mul_U18647(.A(dpath_mulcore_ary1_a0_I1_I2_p2_l_67), .Y(n6297));
AND2X1 mul_U18648(.A(dpath_mulcore_b5[1]), .B(n10991), .Y(dpath_mulcore_ary1_a0_I1_I2_p2_l_66));
INVX1 mul_U18649(.A(dpath_mulcore_ary1_a0_I1_I2_p2_l_66), .Y(n6298));
AND2X1 mul_U18650(.A(dpath_mulcore_b5[1]), .B(n10994), .Y(dpath_mulcore_ary1_a0_I1_I2_p2_l_65));
INVX1 mul_U18651(.A(dpath_mulcore_ary1_a0_I1_I2_p2_l_65), .Y(n6299));
AND2X1 mul_U18652(.A(dpath_mulcore_b4[1]), .B(n10997), .Y(dpath_mulcore_ary1_a0_I1_I2_p1_l_65));
INVX1 mul_U18653(.A(dpath_mulcore_ary1_a0_I1_I2_p1_l_65), .Y(n6300));
AND2X1 mul_U18654(.A(dpath_mulcore_b4[1]), .B(n11000), .Y(dpath_mulcore_ary1_a0_I1_I2_p1_l_64));
INVX1 mul_U18655(.A(dpath_mulcore_ary1_a0_I1_I2_p1_l_64), .Y(n6301));
AND2X1 mul_U18656(.A(dpath_mulcore_b5[1]), .B(n11003), .Y(dpath_mulcore_ary1_a0_I1_I2_p2_l_64));
INVX1 mul_U18657(.A(dpath_mulcore_ary1_a0_I1_I2_p2_l_64), .Y(n6302));
AND2X1 mul_U18658(.A(dpath_mulcore_b5[1]), .B(n11006), .Y(dpath_mulcore_ary1_a0_I1_p2_l[63]));
INVX1 mul_U18659(.A(dpath_mulcore_ary1_a0_I1_p2_l[63]), .Y(n6303));
AND2X1 mul_U18660(.A(dpath_mulcore_b4[1]), .B(n11009), .Y(dpath_mulcore_ary1_a0_I1_p1_l[63]));
INVX1 mul_U18661(.A(dpath_mulcore_ary1_a0_I1_p1_l[63]), .Y(n6304));
AND2X1 mul_U18662(.A(dpath_mulcore_b3[1]), .B(n11012), .Y(dpath_mulcore_ary1_a0_I1_p0_l[63]));
INVX1 mul_U18663(.A(dpath_mulcore_ary1_a0_I1_p0_l[63]), .Y(n6305));
AND2X1 mul_U18664(.A(dpath_mulcore_b5[1]), .B(n11015), .Y(dpath_mulcore_ary1_a0_I1_p2_l[62]));
INVX1 mul_U18665(.A(dpath_mulcore_ary1_a0_I1_p2_l[62]), .Y(n6306));
AND2X1 mul_U18666(.A(dpath_mulcore_b4[1]), .B(n11018), .Y(dpath_mulcore_ary1_a0_I1_p1_l[62]));
INVX1 mul_U18667(.A(dpath_mulcore_ary1_a0_I1_p1_l[62]), .Y(n6307));
AND2X1 mul_U18668(.A(dpath_mulcore_b3[1]), .B(n11021), .Y(dpath_mulcore_ary1_a0_I1_p0_l[62]));
INVX1 mul_U18669(.A(dpath_mulcore_ary1_a0_I1_p0_l[62]), .Y(n6308));
AND2X1 mul_U18670(.A(dpath_mulcore_b5[1]), .B(n11024), .Y(dpath_mulcore_ary1_a0_I1_p2_l[61]));
INVX1 mul_U18671(.A(dpath_mulcore_ary1_a0_I1_p2_l[61]), .Y(n6309));
AND2X1 mul_U18672(.A(dpath_mulcore_b4[1]), .B(n11027), .Y(dpath_mulcore_ary1_a0_I1_p1_l[61]));
INVX1 mul_U18673(.A(dpath_mulcore_ary1_a0_I1_p1_l[61]), .Y(n6310));
AND2X1 mul_U18674(.A(dpath_mulcore_b3[1]), .B(n11030), .Y(dpath_mulcore_ary1_a0_I1_p0_l[61]));
INVX1 mul_U18675(.A(dpath_mulcore_ary1_a0_I1_p0_l[61]), .Y(n6311));
AND2X1 mul_U18676(.A(dpath_mulcore_b5[1]), .B(n11033), .Y(dpath_mulcore_ary1_a0_I1_p2_l[60]));
INVX1 mul_U18677(.A(dpath_mulcore_ary1_a0_I1_p2_l[60]), .Y(n6312));
AND2X1 mul_U18678(.A(dpath_mulcore_b4[1]), .B(n11036), .Y(dpath_mulcore_ary1_a0_I1_p1_l[60]));
INVX1 mul_U18679(.A(dpath_mulcore_ary1_a0_I1_p1_l[60]), .Y(n6313));
AND2X1 mul_U18680(.A(dpath_mulcore_b3[1]), .B(n11039), .Y(dpath_mulcore_ary1_a0_I1_p0_l[60]));
INVX1 mul_U18681(.A(dpath_mulcore_ary1_a0_I1_p0_l[60]), .Y(n6314));
AND2X1 mul_U18682(.A(dpath_mulcore_b5[1]), .B(n11042), .Y(dpath_mulcore_ary1_a0_I1_p2_l[59]));
INVX1 mul_U18683(.A(dpath_mulcore_ary1_a0_I1_p2_l[59]), .Y(n6315));
AND2X1 mul_U18684(.A(dpath_mulcore_b4[1]), .B(n11045), .Y(dpath_mulcore_ary1_a0_I1_p1_l[59]));
INVX1 mul_U18685(.A(dpath_mulcore_ary1_a0_I1_p1_l[59]), .Y(n6316));
AND2X1 mul_U18686(.A(dpath_mulcore_b3[1]), .B(n11048), .Y(dpath_mulcore_ary1_a0_I1_p0_l[59]));
INVX1 mul_U18687(.A(dpath_mulcore_ary1_a0_I1_p0_l[59]), .Y(n6317));
AND2X1 mul_U18688(.A(dpath_mulcore_b5[1]), .B(n11051), .Y(dpath_mulcore_ary1_a0_I1_p2_l[58]));
INVX1 mul_U18689(.A(dpath_mulcore_ary1_a0_I1_p2_l[58]), .Y(n6318));
AND2X1 mul_U18690(.A(dpath_mulcore_b4[1]), .B(n11054), .Y(dpath_mulcore_ary1_a0_I1_p1_l[58]));
INVX1 mul_U18691(.A(dpath_mulcore_ary1_a0_I1_p1_l[58]), .Y(n6319));
AND2X1 mul_U18692(.A(dpath_mulcore_b3[1]), .B(n11057), .Y(dpath_mulcore_ary1_a0_I1_p0_l[58]));
INVX1 mul_U18693(.A(dpath_mulcore_ary1_a0_I1_p0_l[58]), .Y(n6320));
AND2X1 mul_U18694(.A(dpath_mulcore_b5[1]), .B(n11060), .Y(dpath_mulcore_ary1_a0_I1_p2_l[57]));
INVX1 mul_U18695(.A(dpath_mulcore_ary1_a0_I1_p2_l[57]), .Y(n6321));
AND2X1 mul_U18696(.A(dpath_mulcore_b4[1]), .B(n11063), .Y(dpath_mulcore_ary1_a0_I1_p1_l[57]));
INVX1 mul_U18697(.A(dpath_mulcore_ary1_a0_I1_p1_l[57]), .Y(n6322));
AND2X1 mul_U18698(.A(dpath_mulcore_b3[1]), .B(n11066), .Y(dpath_mulcore_ary1_a0_I1_p0_l[57]));
INVX1 mul_U18699(.A(dpath_mulcore_ary1_a0_I1_p0_l[57]), .Y(n6323));
AND2X1 mul_U18700(.A(dpath_mulcore_b5[1]), .B(n11069), .Y(dpath_mulcore_ary1_a0_I1_p2_l[56]));
INVX1 mul_U18701(.A(dpath_mulcore_ary1_a0_I1_p2_l[56]), .Y(n6324));
AND2X1 mul_U18702(.A(dpath_mulcore_b4[1]), .B(n11072), .Y(dpath_mulcore_ary1_a0_I1_p1_l[56]));
INVX1 mul_U18703(.A(dpath_mulcore_ary1_a0_I1_p1_l[56]), .Y(n6325));
AND2X1 mul_U18704(.A(dpath_mulcore_b3[1]), .B(n11075), .Y(dpath_mulcore_ary1_a0_I1_p0_l[56]));
INVX1 mul_U18705(.A(dpath_mulcore_ary1_a0_I1_p0_l[56]), .Y(n6326));
AND2X1 mul_U18706(.A(dpath_mulcore_b5[1]), .B(n11078), .Y(dpath_mulcore_ary1_a0_I1_p2_l[55]));
INVX1 mul_U18707(.A(dpath_mulcore_ary1_a0_I1_p2_l[55]), .Y(n6327));
AND2X1 mul_U18708(.A(dpath_mulcore_b4[1]), .B(n11081), .Y(dpath_mulcore_ary1_a0_I1_p1_l[55]));
INVX1 mul_U18709(.A(dpath_mulcore_ary1_a0_I1_p1_l[55]), .Y(n6328));
AND2X1 mul_U18710(.A(dpath_mulcore_b3[1]), .B(n11084), .Y(dpath_mulcore_ary1_a0_I1_p0_l[55]));
INVX1 mul_U18711(.A(dpath_mulcore_ary1_a0_I1_p0_l[55]), .Y(n6329));
AND2X1 mul_U18712(.A(dpath_mulcore_b5[1]), .B(n11087), .Y(dpath_mulcore_ary1_a0_I1_p2_l[54]));
INVX1 mul_U18713(.A(dpath_mulcore_ary1_a0_I1_p2_l[54]), .Y(n6330));
AND2X1 mul_U18714(.A(dpath_mulcore_b4[1]), .B(n11090), .Y(dpath_mulcore_ary1_a0_I1_p1_l[54]));
INVX1 mul_U18715(.A(dpath_mulcore_ary1_a0_I1_p1_l[54]), .Y(n6331));
AND2X1 mul_U18716(.A(dpath_mulcore_b3[1]), .B(n11093), .Y(dpath_mulcore_ary1_a0_I1_p0_l[54]));
INVX1 mul_U18717(.A(dpath_mulcore_ary1_a0_I1_p0_l[54]), .Y(n6332));
AND2X1 mul_U18718(.A(dpath_mulcore_b5[1]), .B(n11096), .Y(dpath_mulcore_ary1_a0_I1_p2_l[53]));
INVX1 mul_U18719(.A(dpath_mulcore_ary1_a0_I1_p2_l[53]), .Y(n6333));
AND2X1 mul_U18720(.A(dpath_mulcore_b4[1]), .B(n11099), .Y(dpath_mulcore_ary1_a0_I1_p1_l[53]));
INVX1 mul_U18721(.A(dpath_mulcore_ary1_a0_I1_p1_l[53]), .Y(n6334));
AND2X1 mul_U18722(.A(dpath_mulcore_b3[1]), .B(n11102), .Y(dpath_mulcore_ary1_a0_I1_p0_l[53]));
INVX1 mul_U18723(.A(dpath_mulcore_ary1_a0_I1_p0_l[53]), .Y(n6335));
AND2X1 mul_U18724(.A(dpath_mulcore_b5[1]), .B(n11105), .Y(dpath_mulcore_ary1_a0_I1_p2_l[52]));
INVX1 mul_U18725(.A(dpath_mulcore_ary1_a0_I1_p2_l[52]), .Y(n6336));
AND2X1 mul_U18726(.A(dpath_mulcore_b4[1]), .B(n11108), .Y(dpath_mulcore_ary1_a0_I1_p1_l[52]));
INVX1 mul_U18727(.A(dpath_mulcore_ary1_a0_I1_p1_l[52]), .Y(n6337));
AND2X1 mul_U18728(.A(dpath_mulcore_b3[1]), .B(n11111), .Y(dpath_mulcore_ary1_a0_I1_p0_l[52]));
INVX1 mul_U18729(.A(dpath_mulcore_ary1_a0_I1_p0_l[52]), .Y(n6338));
AND2X1 mul_U18730(.A(dpath_mulcore_b5[1]), .B(n11114), .Y(dpath_mulcore_ary1_a0_I1_p2_l[51]));
INVX1 mul_U18731(.A(dpath_mulcore_ary1_a0_I1_p2_l[51]), .Y(n6339));
AND2X1 mul_U18732(.A(dpath_mulcore_b4[1]), .B(n11117), .Y(dpath_mulcore_ary1_a0_I1_p1_l[51]));
INVX1 mul_U18733(.A(dpath_mulcore_ary1_a0_I1_p1_l[51]), .Y(n6340));
AND2X1 mul_U18734(.A(dpath_mulcore_b3[1]), .B(n11120), .Y(dpath_mulcore_ary1_a0_I1_p0_l[51]));
INVX1 mul_U18735(.A(dpath_mulcore_ary1_a0_I1_p0_l[51]), .Y(n6341));
AND2X1 mul_U18736(.A(dpath_mulcore_b5[1]), .B(n11123), .Y(dpath_mulcore_ary1_a0_I1_p2_l[50]));
INVX1 mul_U18737(.A(dpath_mulcore_ary1_a0_I1_p2_l[50]), .Y(n6342));
AND2X1 mul_U18738(.A(dpath_mulcore_b4[1]), .B(n11126), .Y(dpath_mulcore_ary1_a0_I1_p1_l[50]));
INVX1 mul_U18739(.A(dpath_mulcore_ary1_a0_I1_p1_l[50]), .Y(n6343));
AND2X1 mul_U18740(.A(dpath_mulcore_b3[1]), .B(n11129), .Y(dpath_mulcore_ary1_a0_I1_p0_l[50]));
INVX1 mul_U18741(.A(dpath_mulcore_ary1_a0_I1_p0_l[50]), .Y(n6344));
AND2X1 mul_U18742(.A(dpath_mulcore_b5[1]), .B(n11132), .Y(dpath_mulcore_ary1_a0_I1_p2_l[49]));
INVX1 mul_U18743(.A(dpath_mulcore_ary1_a0_I1_p2_l[49]), .Y(n6345));
AND2X1 mul_U18744(.A(dpath_mulcore_b4[1]), .B(n11135), .Y(dpath_mulcore_ary1_a0_I1_p1_l[49]));
INVX1 mul_U18745(.A(dpath_mulcore_ary1_a0_I1_p1_l[49]), .Y(n6346));
AND2X1 mul_U18746(.A(dpath_mulcore_b3[1]), .B(n11138), .Y(dpath_mulcore_ary1_a0_I1_p0_l[49]));
INVX1 mul_U18747(.A(dpath_mulcore_ary1_a0_I1_p0_l[49]), .Y(n6347));
AND2X1 mul_U18748(.A(dpath_mulcore_b5[1]), .B(n11141), .Y(dpath_mulcore_ary1_a0_I1_p2_l[48]));
INVX1 mul_U18749(.A(dpath_mulcore_ary1_a0_I1_p2_l[48]), .Y(n6348));
AND2X1 mul_U18750(.A(dpath_mulcore_b4[1]), .B(n11144), .Y(dpath_mulcore_ary1_a0_I1_p1_l[48]));
INVX1 mul_U18751(.A(dpath_mulcore_ary1_a0_I1_p1_l[48]), .Y(n6349));
AND2X1 mul_U18752(.A(dpath_mulcore_b3[1]), .B(n11147), .Y(dpath_mulcore_ary1_a0_I1_p0_l[48]));
INVX1 mul_U18753(.A(dpath_mulcore_ary1_a0_I1_p0_l[48]), .Y(n6350));
AND2X1 mul_U18754(.A(dpath_mulcore_b5[1]), .B(n11150), .Y(dpath_mulcore_ary1_a0_I1_p2_l[47]));
INVX1 mul_U18755(.A(dpath_mulcore_ary1_a0_I1_p2_l[47]), .Y(n6351));
AND2X1 mul_U18756(.A(dpath_mulcore_b4[1]), .B(n11153), .Y(dpath_mulcore_ary1_a0_I1_p1_l[47]));
INVX1 mul_U18757(.A(dpath_mulcore_ary1_a0_I1_p1_l[47]), .Y(n6352));
AND2X1 mul_U18758(.A(dpath_mulcore_b3[1]), .B(n11156), .Y(dpath_mulcore_ary1_a0_I1_p0_l[47]));
INVX1 mul_U18759(.A(dpath_mulcore_ary1_a0_I1_p0_l[47]), .Y(n6353));
AND2X1 mul_U18760(.A(dpath_mulcore_b5[1]), .B(n11159), .Y(dpath_mulcore_ary1_a0_I1_p2_l[46]));
INVX1 mul_U18761(.A(dpath_mulcore_ary1_a0_I1_p2_l[46]), .Y(n6354));
AND2X1 mul_U18762(.A(dpath_mulcore_b4[1]), .B(n11162), .Y(dpath_mulcore_ary1_a0_I1_p1_l[46]));
INVX1 mul_U18763(.A(dpath_mulcore_ary1_a0_I1_p1_l[46]), .Y(n6355));
AND2X1 mul_U18764(.A(dpath_mulcore_b3[1]), .B(n11165), .Y(dpath_mulcore_ary1_a0_I1_p0_l[46]));
INVX1 mul_U18765(.A(dpath_mulcore_ary1_a0_I1_p0_l[46]), .Y(n6356));
AND2X1 mul_U18766(.A(dpath_mulcore_b5[1]), .B(n11168), .Y(dpath_mulcore_ary1_a0_I1_p2_l[45]));
INVX1 mul_U18767(.A(dpath_mulcore_ary1_a0_I1_p2_l[45]), .Y(n6357));
AND2X1 mul_U18768(.A(dpath_mulcore_b4[1]), .B(n11171), .Y(dpath_mulcore_ary1_a0_I1_p1_l[45]));
INVX1 mul_U18769(.A(dpath_mulcore_ary1_a0_I1_p1_l[45]), .Y(n6358));
AND2X1 mul_U18770(.A(dpath_mulcore_b3[1]), .B(n11174), .Y(dpath_mulcore_ary1_a0_I1_p0_l[45]));
INVX1 mul_U18771(.A(dpath_mulcore_ary1_a0_I1_p0_l[45]), .Y(n6359));
AND2X1 mul_U18772(.A(dpath_mulcore_b5[1]), .B(n11177), .Y(dpath_mulcore_ary1_a0_I1_p2_l[44]));
INVX1 mul_U18773(.A(dpath_mulcore_ary1_a0_I1_p2_l[44]), .Y(n6360));
AND2X1 mul_U18774(.A(dpath_mulcore_b4[1]), .B(n11180), .Y(dpath_mulcore_ary1_a0_I1_p1_l[44]));
INVX1 mul_U18775(.A(dpath_mulcore_ary1_a0_I1_p1_l[44]), .Y(n6361));
AND2X1 mul_U18776(.A(dpath_mulcore_b3[1]), .B(n11183), .Y(dpath_mulcore_ary1_a0_I1_p0_l[44]));
INVX1 mul_U18777(.A(dpath_mulcore_ary1_a0_I1_p0_l[44]), .Y(n6362));
AND2X1 mul_U18778(.A(dpath_mulcore_b5[1]), .B(n11186), .Y(dpath_mulcore_ary1_a0_I1_p2_l[43]));
INVX1 mul_U18779(.A(dpath_mulcore_ary1_a0_I1_p2_l[43]), .Y(n6363));
AND2X1 mul_U18780(.A(dpath_mulcore_b4[1]), .B(n11189), .Y(dpath_mulcore_ary1_a0_I1_p1_l[43]));
INVX1 mul_U18781(.A(dpath_mulcore_ary1_a0_I1_p1_l[43]), .Y(n6364));
AND2X1 mul_U18782(.A(dpath_mulcore_b3[1]), .B(n11192), .Y(dpath_mulcore_ary1_a0_I1_p0_l[43]));
INVX1 mul_U18783(.A(dpath_mulcore_ary1_a0_I1_p0_l[43]), .Y(n6365));
AND2X1 mul_U18784(.A(dpath_mulcore_b5[1]), .B(n11195), .Y(dpath_mulcore_ary1_a0_I1_p2_l[42]));
INVX1 mul_U18785(.A(dpath_mulcore_ary1_a0_I1_p2_l[42]), .Y(n6366));
AND2X1 mul_U18786(.A(dpath_mulcore_b4[1]), .B(n11198), .Y(dpath_mulcore_ary1_a0_I1_p1_l[42]));
INVX1 mul_U18787(.A(dpath_mulcore_ary1_a0_I1_p1_l[42]), .Y(n6367));
AND2X1 mul_U18788(.A(dpath_mulcore_b3[1]), .B(n11201), .Y(dpath_mulcore_ary1_a0_I1_p0_l[42]));
INVX1 mul_U18789(.A(dpath_mulcore_ary1_a0_I1_p0_l[42]), .Y(n6368));
AND2X1 mul_U18790(.A(dpath_mulcore_b5[1]), .B(n11204), .Y(dpath_mulcore_ary1_a0_I1_p2_l[41]));
INVX1 mul_U18791(.A(dpath_mulcore_ary1_a0_I1_p2_l[41]), .Y(n6369));
AND2X1 mul_U18792(.A(dpath_mulcore_b4[1]), .B(n11207), .Y(dpath_mulcore_ary1_a0_I1_p1_l[41]));
INVX1 mul_U18793(.A(dpath_mulcore_ary1_a0_I1_p1_l[41]), .Y(n6370));
AND2X1 mul_U18794(.A(dpath_mulcore_b3[1]), .B(n11210), .Y(dpath_mulcore_ary1_a0_I1_p0_l[41]));
INVX1 mul_U18795(.A(dpath_mulcore_ary1_a0_I1_p0_l[41]), .Y(n6371));
AND2X1 mul_U18796(.A(dpath_mulcore_b5[1]), .B(n11213), .Y(dpath_mulcore_ary1_a0_I1_p2_l[40]));
INVX1 mul_U18797(.A(dpath_mulcore_ary1_a0_I1_p2_l[40]), .Y(n6372));
AND2X1 mul_U18798(.A(dpath_mulcore_b4[1]), .B(n11216), .Y(dpath_mulcore_ary1_a0_I1_p1_l[40]));
INVX1 mul_U18799(.A(dpath_mulcore_ary1_a0_I1_p1_l[40]), .Y(n6373));
AND2X1 mul_U18800(.A(dpath_mulcore_b3[1]), .B(n11219), .Y(dpath_mulcore_ary1_a0_I1_p0_l[40]));
INVX1 mul_U18801(.A(dpath_mulcore_ary1_a0_I1_p0_l[40]), .Y(n6374));
AND2X1 mul_U18802(.A(dpath_mulcore_b5[1]), .B(n11222), .Y(dpath_mulcore_ary1_a0_I1_p2_l[39]));
INVX1 mul_U18803(.A(dpath_mulcore_ary1_a0_I1_p2_l[39]), .Y(n6375));
AND2X1 mul_U18804(.A(dpath_mulcore_b4[1]), .B(n11225), .Y(dpath_mulcore_ary1_a0_I1_p1_l[39]));
INVX1 mul_U18805(.A(dpath_mulcore_ary1_a0_I1_p1_l[39]), .Y(n6376));
AND2X1 mul_U18806(.A(dpath_mulcore_b3[1]), .B(n11228), .Y(dpath_mulcore_ary1_a0_I1_p0_l[39]));
INVX1 mul_U18807(.A(dpath_mulcore_ary1_a0_I1_p0_l[39]), .Y(n6377));
AND2X1 mul_U18808(.A(dpath_mulcore_b5[1]), .B(n11231), .Y(dpath_mulcore_ary1_a0_I1_p2_l[38]));
INVX1 mul_U18809(.A(dpath_mulcore_ary1_a0_I1_p2_l[38]), .Y(n6378));
AND2X1 mul_U18810(.A(dpath_mulcore_b4[1]), .B(n11234), .Y(dpath_mulcore_ary1_a0_I1_p1_l[38]));
INVX1 mul_U18811(.A(dpath_mulcore_ary1_a0_I1_p1_l[38]), .Y(n6379));
AND2X1 mul_U18812(.A(dpath_mulcore_b3[1]), .B(n11237), .Y(dpath_mulcore_ary1_a0_I1_p0_l[38]));
INVX1 mul_U18813(.A(dpath_mulcore_ary1_a0_I1_p0_l[38]), .Y(n6380));
AND2X1 mul_U18814(.A(dpath_mulcore_b5[1]), .B(n11240), .Y(dpath_mulcore_ary1_a0_I1_p2_l[37]));
INVX1 mul_U18815(.A(dpath_mulcore_ary1_a0_I1_p2_l[37]), .Y(n6381));
AND2X1 mul_U18816(.A(dpath_mulcore_b4[1]), .B(n11243), .Y(dpath_mulcore_ary1_a0_I1_p1_l[37]));
INVX1 mul_U18817(.A(dpath_mulcore_ary1_a0_I1_p1_l[37]), .Y(n6382));
AND2X1 mul_U18818(.A(dpath_mulcore_b3[1]), .B(n11246), .Y(dpath_mulcore_ary1_a0_I1_p0_l[37]));
INVX1 mul_U18819(.A(dpath_mulcore_ary1_a0_I1_p0_l[37]), .Y(n6383));
AND2X1 mul_U18820(.A(dpath_mulcore_b5[1]), .B(n11249), .Y(dpath_mulcore_ary1_a0_I1_p2_l[36]));
INVX1 mul_U18821(.A(dpath_mulcore_ary1_a0_I1_p2_l[36]), .Y(n6384));
AND2X1 mul_U18822(.A(dpath_mulcore_b4[1]), .B(n11252), .Y(dpath_mulcore_ary1_a0_I1_p1_l[36]));
INVX1 mul_U18823(.A(dpath_mulcore_ary1_a0_I1_p1_l[36]), .Y(n6385));
AND2X1 mul_U18824(.A(dpath_mulcore_b3[1]), .B(n11255), .Y(dpath_mulcore_ary1_a0_I1_p0_l[36]));
INVX1 mul_U18825(.A(dpath_mulcore_ary1_a0_I1_p0_l[36]), .Y(n6386));
AND2X1 mul_U18826(.A(dpath_mulcore_b5[1]), .B(n11258), .Y(dpath_mulcore_ary1_a0_I1_p2_l[35]));
INVX1 mul_U18827(.A(dpath_mulcore_ary1_a0_I1_p2_l[35]), .Y(n6387));
AND2X1 mul_U18828(.A(dpath_mulcore_b4[1]), .B(n11261), .Y(dpath_mulcore_ary1_a0_I1_p1_l[35]));
INVX1 mul_U18829(.A(dpath_mulcore_ary1_a0_I1_p1_l[35]), .Y(n6388));
AND2X1 mul_U18830(.A(dpath_mulcore_b3[1]), .B(n11264), .Y(dpath_mulcore_ary1_a0_I1_p0_l[35]));
INVX1 mul_U18831(.A(dpath_mulcore_ary1_a0_I1_p0_l[35]), .Y(n6389));
AND2X1 mul_U18832(.A(dpath_mulcore_b5[1]), .B(n11267), .Y(dpath_mulcore_ary1_a0_I1_p2_l[34]));
INVX1 mul_U18833(.A(dpath_mulcore_ary1_a0_I1_p2_l[34]), .Y(n6390));
AND2X1 mul_U18834(.A(dpath_mulcore_b4[1]), .B(n11270), .Y(dpath_mulcore_ary1_a0_I1_p1_l[34]));
INVX1 mul_U18835(.A(dpath_mulcore_ary1_a0_I1_p1_l[34]), .Y(n6391));
AND2X1 mul_U18836(.A(dpath_mulcore_b3[1]), .B(n11273), .Y(dpath_mulcore_ary1_a0_I1_p0_l[34]));
INVX1 mul_U18837(.A(dpath_mulcore_ary1_a0_I1_p0_l[34]), .Y(n6392));
AND2X1 mul_U18838(.A(dpath_mulcore_b5[1]), .B(n11276), .Y(dpath_mulcore_ary1_a0_I1_p2_l[33]));
INVX1 mul_U18839(.A(dpath_mulcore_ary1_a0_I1_p2_l[33]), .Y(n6393));
AND2X1 mul_U18840(.A(dpath_mulcore_b4[1]), .B(n11279), .Y(dpath_mulcore_ary1_a0_I1_p1_l[33]));
INVX1 mul_U18841(.A(dpath_mulcore_ary1_a0_I1_p1_l[33]), .Y(n6394));
AND2X1 mul_U18842(.A(dpath_mulcore_b3[1]), .B(n11282), .Y(dpath_mulcore_ary1_a0_I1_p0_l[33]));
INVX1 mul_U18843(.A(dpath_mulcore_ary1_a0_I1_p0_l[33]), .Y(n6395));
AND2X1 mul_U18844(.A(dpath_mulcore_b5[1]), .B(n11285), .Y(dpath_mulcore_ary1_a0_I1_p2_l[32]));
INVX1 mul_U18845(.A(dpath_mulcore_ary1_a0_I1_p2_l[32]), .Y(n6396));
AND2X1 mul_U18846(.A(dpath_mulcore_b4[1]), .B(n11288), .Y(dpath_mulcore_ary1_a0_I1_p1_l[32]));
INVX1 mul_U18847(.A(dpath_mulcore_ary1_a0_I1_p1_l[32]), .Y(n6397));
AND2X1 mul_U18848(.A(dpath_mulcore_b3[1]), .B(n11291), .Y(dpath_mulcore_ary1_a0_I1_p0_l[32]));
INVX1 mul_U18849(.A(dpath_mulcore_ary1_a0_I1_p0_l[32]), .Y(n6398));
AND2X1 mul_U18850(.A(dpath_mulcore_b5[1]), .B(n11294), .Y(dpath_mulcore_ary1_a0_I1_p2_l[31]));
INVX1 mul_U18851(.A(dpath_mulcore_ary1_a0_I1_p2_l[31]), .Y(n6399));
AND2X1 mul_U18852(.A(dpath_mulcore_b4[1]), .B(n11297), .Y(dpath_mulcore_ary1_a0_I1_p1_l[31]));
INVX1 mul_U18853(.A(dpath_mulcore_ary1_a0_I1_p1_l[31]), .Y(n6400));
AND2X1 mul_U18854(.A(dpath_mulcore_b3[1]), .B(n11300), .Y(dpath_mulcore_ary1_a0_I1_p0_l[31]));
INVX1 mul_U18855(.A(dpath_mulcore_ary1_a0_I1_p0_l[31]), .Y(n6401));
AND2X1 mul_U18856(.A(dpath_mulcore_b5[1]), .B(n11303), .Y(dpath_mulcore_ary1_a0_I1_p2_l[30]));
INVX1 mul_U18857(.A(dpath_mulcore_ary1_a0_I1_p2_l[30]), .Y(n6402));
AND2X1 mul_U18858(.A(dpath_mulcore_b4[1]), .B(n11306), .Y(dpath_mulcore_ary1_a0_I1_p1_l[30]));
INVX1 mul_U18859(.A(dpath_mulcore_ary1_a0_I1_p1_l[30]), .Y(n6403));
AND2X1 mul_U18860(.A(dpath_mulcore_b3[1]), .B(n11309), .Y(dpath_mulcore_ary1_a0_I1_p0_l[30]));
INVX1 mul_U18861(.A(dpath_mulcore_ary1_a0_I1_p0_l[30]), .Y(n6404));
AND2X1 mul_U18862(.A(dpath_mulcore_b5[1]), .B(n11312), .Y(dpath_mulcore_ary1_a0_I1_p2_l[29]));
INVX1 mul_U18863(.A(dpath_mulcore_ary1_a0_I1_p2_l[29]), .Y(n6405));
AND2X1 mul_U18864(.A(dpath_mulcore_b4[1]), .B(n11315), .Y(dpath_mulcore_ary1_a0_I1_p1_l[29]));
INVX1 mul_U18865(.A(dpath_mulcore_ary1_a0_I1_p1_l[29]), .Y(n6406));
AND2X1 mul_U18866(.A(dpath_mulcore_b3[1]), .B(n11318), .Y(dpath_mulcore_ary1_a0_I1_p0_l[29]));
INVX1 mul_U18867(.A(dpath_mulcore_ary1_a0_I1_p0_l[29]), .Y(n6407));
AND2X1 mul_U18868(.A(dpath_mulcore_b5[1]), .B(n11321), .Y(dpath_mulcore_ary1_a0_I1_p2_l[28]));
INVX1 mul_U18869(.A(dpath_mulcore_ary1_a0_I1_p2_l[28]), .Y(n6408));
AND2X1 mul_U18870(.A(dpath_mulcore_b4[1]), .B(n11324), .Y(dpath_mulcore_ary1_a0_I1_p1_l[28]));
INVX1 mul_U18871(.A(dpath_mulcore_ary1_a0_I1_p1_l[28]), .Y(n6409));
AND2X1 mul_U18872(.A(dpath_mulcore_b3[1]), .B(n11327), .Y(dpath_mulcore_ary1_a0_I1_p0_l[28]));
INVX1 mul_U18873(.A(dpath_mulcore_ary1_a0_I1_p0_l[28]), .Y(n6410));
AND2X1 mul_U18874(.A(dpath_mulcore_b5[1]), .B(n11330), .Y(dpath_mulcore_ary1_a0_I1_p2_l[27]));
INVX1 mul_U18875(.A(dpath_mulcore_ary1_a0_I1_p2_l[27]), .Y(n6411));
AND2X1 mul_U18876(.A(dpath_mulcore_b4[1]), .B(n11333), .Y(dpath_mulcore_ary1_a0_I1_p1_l[27]));
INVX1 mul_U18877(.A(dpath_mulcore_ary1_a0_I1_p1_l[27]), .Y(n6412));
AND2X1 mul_U18878(.A(dpath_mulcore_b3[1]), .B(n11336), .Y(dpath_mulcore_ary1_a0_I1_p0_l[27]));
INVX1 mul_U18879(.A(dpath_mulcore_ary1_a0_I1_p0_l[27]), .Y(n6413));
AND2X1 mul_U18880(.A(dpath_mulcore_b5[1]), .B(n11339), .Y(dpath_mulcore_ary1_a0_I1_p2_l[26]));
INVX1 mul_U18881(.A(dpath_mulcore_ary1_a0_I1_p2_l[26]), .Y(n6414));
AND2X1 mul_U18882(.A(dpath_mulcore_b4[1]), .B(n11342), .Y(dpath_mulcore_ary1_a0_I1_p1_l[26]));
INVX1 mul_U18883(.A(dpath_mulcore_ary1_a0_I1_p1_l[26]), .Y(n6415));
AND2X1 mul_U18884(.A(dpath_mulcore_b3[1]), .B(n11345), .Y(dpath_mulcore_ary1_a0_I1_p0_l[26]));
INVX1 mul_U18885(.A(dpath_mulcore_ary1_a0_I1_p0_l[26]), .Y(n6416));
AND2X1 mul_U18886(.A(dpath_mulcore_b5[1]), .B(n11348), .Y(dpath_mulcore_ary1_a0_I1_p2_l[25]));
INVX1 mul_U18887(.A(dpath_mulcore_ary1_a0_I1_p2_l[25]), .Y(n6417));
AND2X1 mul_U18888(.A(dpath_mulcore_b4[1]), .B(n11351), .Y(dpath_mulcore_ary1_a0_I1_p1_l[25]));
INVX1 mul_U18889(.A(dpath_mulcore_ary1_a0_I1_p1_l[25]), .Y(n6418));
AND2X1 mul_U18890(.A(dpath_mulcore_b3[1]), .B(n11354), .Y(dpath_mulcore_ary1_a0_I1_p0_l[25]));
INVX1 mul_U18891(.A(dpath_mulcore_ary1_a0_I1_p0_l[25]), .Y(n6419));
AND2X1 mul_U18892(.A(dpath_mulcore_b5[1]), .B(n11357), .Y(dpath_mulcore_ary1_a0_I1_p2_l[24]));
INVX1 mul_U18893(.A(dpath_mulcore_ary1_a0_I1_p2_l[24]), .Y(n6420));
AND2X1 mul_U18894(.A(dpath_mulcore_b4[1]), .B(n11360), .Y(dpath_mulcore_ary1_a0_I1_p1_l[24]));
INVX1 mul_U18895(.A(dpath_mulcore_ary1_a0_I1_p1_l[24]), .Y(n6421));
AND2X1 mul_U18896(.A(dpath_mulcore_b3[1]), .B(n11363), .Y(dpath_mulcore_ary1_a0_I1_p0_l[24]));
INVX1 mul_U18897(.A(dpath_mulcore_ary1_a0_I1_p0_l[24]), .Y(n6422));
AND2X1 mul_U18898(.A(dpath_mulcore_b5[1]), .B(n11366), .Y(dpath_mulcore_ary1_a0_I1_p2_l[23]));
INVX1 mul_U18899(.A(dpath_mulcore_ary1_a0_I1_p2_l[23]), .Y(n6423));
AND2X1 mul_U18900(.A(dpath_mulcore_b4[1]), .B(n11369), .Y(dpath_mulcore_ary1_a0_I1_p1_l[23]));
INVX1 mul_U18901(.A(dpath_mulcore_ary1_a0_I1_p1_l[23]), .Y(n6424));
AND2X1 mul_U18902(.A(dpath_mulcore_b3[1]), .B(n11372), .Y(dpath_mulcore_ary1_a0_I1_p0_l[23]));
INVX1 mul_U18903(.A(dpath_mulcore_ary1_a0_I1_p0_l[23]), .Y(n6425));
AND2X1 mul_U18904(.A(dpath_mulcore_b5[1]), .B(n11375), .Y(dpath_mulcore_ary1_a0_I1_p2_l[22]));
INVX1 mul_U18905(.A(dpath_mulcore_ary1_a0_I1_p2_l[22]), .Y(n6426));
AND2X1 mul_U18906(.A(dpath_mulcore_b4[1]), .B(n11378), .Y(dpath_mulcore_ary1_a0_I1_p1_l[22]));
INVX1 mul_U18907(.A(dpath_mulcore_ary1_a0_I1_p1_l[22]), .Y(n6427));
AND2X1 mul_U18908(.A(dpath_mulcore_b3[1]), .B(n11381), .Y(dpath_mulcore_ary1_a0_I1_p0_l[22]));
INVX1 mul_U18909(.A(dpath_mulcore_ary1_a0_I1_p0_l[22]), .Y(n6428));
AND2X1 mul_U18910(.A(dpath_mulcore_b5[1]), .B(n11384), .Y(dpath_mulcore_ary1_a0_I1_p2_l[21]));
INVX1 mul_U18911(.A(dpath_mulcore_ary1_a0_I1_p2_l[21]), .Y(n6429));
AND2X1 mul_U18912(.A(dpath_mulcore_b4[1]), .B(n11387), .Y(dpath_mulcore_ary1_a0_I1_p1_l[21]));
INVX1 mul_U18913(.A(dpath_mulcore_ary1_a0_I1_p1_l[21]), .Y(n6430));
AND2X1 mul_U18914(.A(dpath_mulcore_b3[1]), .B(n11390), .Y(dpath_mulcore_ary1_a0_I1_p0_l[21]));
INVX1 mul_U18915(.A(dpath_mulcore_ary1_a0_I1_p0_l[21]), .Y(n6431));
AND2X1 mul_U18916(.A(dpath_mulcore_b5[1]), .B(n11393), .Y(dpath_mulcore_ary1_a0_I1_p2_l[20]));
INVX1 mul_U18917(.A(dpath_mulcore_ary1_a0_I1_p2_l[20]), .Y(n6432));
AND2X1 mul_U18918(.A(dpath_mulcore_b4[1]), .B(n11396), .Y(dpath_mulcore_ary1_a0_I1_p1_l[20]));
INVX1 mul_U18919(.A(dpath_mulcore_ary1_a0_I1_p1_l[20]), .Y(n6433));
AND2X1 mul_U18920(.A(dpath_mulcore_b3[1]), .B(n11399), .Y(dpath_mulcore_ary1_a0_I1_p0_l[20]));
INVX1 mul_U18921(.A(dpath_mulcore_ary1_a0_I1_p0_l[20]), .Y(n6434));
AND2X1 mul_U18922(.A(dpath_mulcore_b5[1]), .B(n11402), .Y(dpath_mulcore_ary1_a0_I1_p2_l[19]));
INVX1 mul_U18923(.A(dpath_mulcore_ary1_a0_I1_p2_l[19]), .Y(n6435));
AND2X1 mul_U18924(.A(dpath_mulcore_b4[1]), .B(n11405), .Y(dpath_mulcore_ary1_a0_I1_p1_l[19]));
INVX1 mul_U18925(.A(dpath_mulcore_ary1_a0_I1_p1_l[19]), .Y(n6436));
AND2X1 mul_U18926(.A(dpath_mulcore_b3[1]), .B(n11408), .Y(dpath_mulcore_ary1_a0_I1_p0_l[19]));
INVX1 mul_U18927(.A(dpath_mulcore_ary1_a0_I1_p0_l[19]), .Y(n6437));
AND2X1 mul_U18928(.A(dpath_mulcore_b5[1]), .B(n11411), .Y(dpath_mulcore_ary1_a0_I1_p2_l[18]));
INVX1 mul_U18929(.A(dpath_mulcore_ary1_a0_I1_p2_l[18]), .Y(n6438));
AND2X1 mul_U18930(.A(dpath_mulcore_b4[1]), .B(n11414), .Y(dpath_mulcore_ary1_a0_I1_p1_l[18]));
INVX1 mul_U18931(.A(dpath_mulcore_ary1_a0_I1_p1_l[18]), .Y(n6439));
AND2X1 mul_U18932(.A(dpath_mulcore_b3[1]), .B(n11417), .Y(dpath_mulcore_ary1_a0_I1_p0_l[18]));
INVX1 mul_U18933(.A(dpath_mulcore_ary1_a0_I1_p0_l[18]), .Y(n6440));
AND2X1 mul_U18934(.A(dpath_mulcore_b5[1]), .B(n11420), .Y(dpath_mulcore_ary1_a0_I1_p2_l[17]));
INVX1 mul_U18935(.A(dpath_mulcore_ary1_a0_I1_p2_l[17]), .Y(n6441));
AND2X1 mul_U18936(.A(dpath_mulcore_b4[1]), .B(n11423), .Y(dpath_mulcore_ary1_a0_I1_p1_l[17]));
INVX1 mul_U18937(.A(dpath_mulcore_ary1_a0_I1_p1_l[17]), .Y(n6442));
AND2X1 mul_U18938(.A(dpath_mulcore_b3[1]), .B(n11426), .Y(dpath_mulcore_ary1_a0_I1_p0_l[17]));
INVX1 mul_U18939(.A(dpath_mulcore_ary1_a0_I1_p0_l[17]), .Y(n6443));
AND2X1 mul_U18940(.A(dpath_mulcore_b5[1]), .B(n11429), .Y(dpath_mulcore_ary1_a0_I1_p2_l[16]));
INVX1 mul_U18941(.A(dpath_mulcore_ary1_a0_I1_p2_l[16]), .Y(n6444));
AND2X1 mul_U18942(.A(dpath_mulcore_b4[1]), .B(n11432), .Y(dpath_mulcore_ary1_a0_I1_p1_l[16]));
INVX1 mul_U18943(.A(dpath_mulcore_ary1_a0_I1_p1_l[16]), .Y(n6445));
AND2X1 mul_U18944(.A(dpath_mulcore_b3[1]), .B(n11435), .Y(dpath_mulcore_ary1_a0_I1_p0_l[16]));
INVX1 mul_U18945(.A(dpath_mulcore_ary1_a0_I1_p0_l[16]), .Y(n6446));
AND2X1 mul_U18946(.A(dpath_mulcore_b5[1]), .B(n11438), .Y(dpath_mulcore_ary1_a0_I1_p2_l[15]));
INVX1 mul_U18947(.A(dpath_mulcore_ary1_a0_I1_p2_l[15]), .Y(n6447));
AND2X1 mul_U18948(.A(dpath_mulcore_b4[1]), .B(n11441), .Y(dpath_mulcore_ary1_a0_I1_p1_l[15]));
INVX1 mul_U18949(.A(dpath_mulcore_ary1_a0_I1_p1_l[15]), .Y(n6448));
AND2X1 mul_U18950(.A(dpath_mulcore_b3[1]), .B(n11444), .Y(dpath_mulcore_ary1_a0_I1_p0_l[15]));
INVX1 mul_U18951(.A(dpath_mulcore_ary1_a0_I1_p0_l[15]), .Y(n6449));
AND2X1 mul_U18952(.A(dpath_mulcore_b5[1]), .B(n11447), .Y(dpath_mulcore_ary1_a0_I1_p2_l[14]));
INVX1 mul_U18953(.A(dpath_mulcore_ary1_a0_I1_p2_l[14]), .Y(n6450));
AND2X1 mul_U18954(.A(dpath_mulcore_b4[1]), .B(n11450), .Y(dpath_mulcore_ary1_a0_I1_p1_l[14]));
INVX1 mul_U18955(.A(dpath_mulcore_ary1_a0_I1_p1_l[14]), .Y(n6451));
AND2X1 mul_U18956(.A(dpath_mulcore_b3[1]), .B(n11453), .Y(dpath_mulcore_ary1_a0_I1_p0_l[14]));
INVX1 mul_U18957(.A(dpath_mulcore_ary1_a0_I1_p0_l[14]), .Y(n6452));
AND2X1 mul_U18958(.A(dpath_mulcore_b5[1]), .B(n11456), .Y(dpath_mulcore_ary1_a0_I1_p2_l[13]));
INVX1 mul_U18959(.A(dpath_mulcore_ary1_a0_I1_p2_l[13]), .Y(n6453));
AND2X1 mul_U18960(.A(dpath_mulcore_b4[1]), .B(n11459), .Y(dpath_mulcore_ary1_a0_I1_p1_l[13]));
INVX1 mul_U18961(.A(dpath_mulcore_ary1_a0_I1_p1_l[13]), .Y(n6454));
AND2X1 mul_U18962(.A(dpath_mulcore_b3[1]), .B(n11462), .Y(dpath_mulcore_ary1_a0_I1_p0_l[13]));
INVX1 mul_U18963(.A(dpath_mulcore_ary1_a0_I1_p0_l[13]), .Y(n6455));
AND2X1 mul_U18964(.A(dpath_mulcore_b5[1]), .B(n11465), .Y(dpath_mulcore_ary1_a0_I1_p2_l[12]));
INVX1 mul_U18965(.A(dpath_mulcore_ary1_a0_I1_p2_l[12]), .Y(n6456));
AND2X1 mul_U18966(.A(dpath_mulcore_b4[1]), .B(n11468), .Y(dpath_mulcore_ary1_a0_I1_p1_l[12]));
INVX1 mul_U18967(.A(dpath_mulcore_ary1_a0_I1_p1_l[12]), .Y(n6457));
AND2X1 mul_U18968(.A(dpath_mulcore_b3[1]), .B(n11471), .Y(dpath_mulcore_ary1_a0_I1_p0_l[12]));
INVX1 mul_U18969(.A(dpath_mulcore_ary1_a0_I1_p0_l[12]), .Y(n6458));
AND2X1 mul_U18970(.A(dpath_mulcore_b5[1]), .B(n11474), .Y(dpath_mulcore_ary1_a0_I1_p2_l[11]));
INVX1 mul_U18971(.A(dpath_mulcore_ary1_a0_I1_p2_l[11]), .Y(n6459));
AND2X1 mul_U18972(.A(dpath_mulcore_b4[1]), .B(n11477), .Y(dpath_mulcore_ary1_a0_I1_p1_l[11]));
INVX1 mul_U18973(.A(dpath_mulcore_ary1_a0_I1_p1_l[11]), .Y(n6460));
AND2X1 mul_U18974(.A(dpath_mulcore_b3[1]), .B(n11480), .Y(dpath_mulcore_ary1_a0_I1_p0_l[11]));
INVX1 mul_U18975(.A(dpath_mulcore_ary1_a0_I1_p0_l[11]), .Y(n6461));
AND2X1 mul_U18976(.A(dpath_mulcore_b5[1]), .B(n11483), .Y(dpath_mulcore_ary1_a0_I1_p2_l[10]));
INVX1 mul_U18977(.A(dpath_mulcore_ary1_a0_I1_p2_l[10]), .Y(n6462));
AND2X1 mul_U18978(.A(dpath_mulcore_b4[1]), .B(n11486), .Y(dpath_mulcore_ary1_a0_I1_p1_l[10]));
INVX1 mul_U18979(.A(dpath_mulcore_ary1_a0_I1_p1_l[10]), .Y(n6463));
AND2X1 mul_U18980(.A(dpath_mulcore_b3[1]), .B(n11489), .Y(dpath_mulcore_ary1_a0_I1_p0_l[10]));
INVX1 mul_U18981(.A(dpath_mulcore_ary1_a0_I1_p0_l[10]), .Y(n6464));
AND2X1 mul_U18982(.A(dpath_mulcore_b5[1]), .B(n11492), .Y(dpath_mulcore_ary1_a0_I1_p2_l[9]));
INVX1 mul_U18983(.A(dpath_mulcore_ary1_a0_I1_p2_l[9]), .Y(n6465));
AND2X1 mul_U18984(.A(dpath_mulcore_b4[1]), .B(n11495), .Y(dpath_mulcore_ary1_a0_I1_p1_l[9]));
INVX1 mul_U18985(.A(dpath_mulcore_ary1_a0_I1_p1_l[9]), .Y(n6466));
AND2X1 mul_U18986(.A(dpath_mulcore_b3[1]), .B(n11498), .Y(dpath_mulcore_ary1_a0_I1_p0_l[9]));
INVX1 mul_U18987(.A(dpath_mulcore_ary1_a0_I1_p0_l[9]), .Y(n6467));
AND2X1 mul_U18988(.A(dpath_mulcore_b5[1]), .B(n11501), .Y(dpath_mulcore_ary1_a0_I1_p2_l[8]));
INVX1 mul_U18989(.A(dpath_mulcore_ary1_a0_I1_p2_l[8]), .Y(n6468));
AND2X1 mul_U18990(.A(dpath_mulcore_b4[1]), .B(n11504), .Y(dpath_mulcore_ary1_a0_I1_p1_l[8]));
INVX1 mul_U18991(.A(dpath_mulcore_ary1_a0_I1_p1_l[8]), .Y(n6469));
AND2X1 mul_U18992(.A(dpath_mulcore_b3[1]), .B(n11507), .Y(dpath_mulcore_ary1_a0_I1_p0_l[8]));
INVX1 mul_U18993(.A(dpath_mulcore_ary1_a0_I1_p0_l[8]), .Y(n6470));
AND2X1 mul_U18994(.A(dpath_mulcore_b5[1]), .B(n11510), .Y(dpath_mulcore_ary1_a0_I1_p2_l[7]));
INVX1 mul_U18995(.A(dpath_mulcore_ary1_a0_I1_p2_l[7]), .Y(n6471));
AND2X1 mul_U18996(.A(dpath_mulcore_b4[1]), .B(n11513), .Y(dpath_mulcore_ary1_a0_I1_p1_l[7]));
INVX1 mul_U18997(.A(dpath_mulcore_ary1_a0_I1_p1_l[7]), .Y(n6472));
AND2X1 mul_U18998(.A(dpath_mulcore_b3[1]), .B(n11516), .Y(dpath_mulcore_ary1_a0_I1_p0_l[7]));
INVX1 mul_U18999(.A(dpath_mulcore_ary1_a0_I1_p0_l[7]), .Y(n6473));
AND2X1 mul_U19000(.A(dpath_mulcore_b5[1]), .B(n11519), .Y(dpath_mulcore_ary1_a0_I1_p2_l[6]));
INVX1 mul_U19001(.A(dpath_mulcore_ary1_a0_I1_p2_l[6]), .Y(n6474));
AND2X1 mul_U19002(.A(dpath_mulcore_b4[1]), .B(n11522), .Y(dpath_mulcore_ary1_a0_I1_p1_l[6]));
INVX1 mul_U19003(.A(dpath_mulcore_ary1_a0_I1_p1_l[6]), .Y(n6475));
AND2X1 mul_U19004(.A(dpath_mulcore_b3[1]), .B(n11525), .Y(dpath_mulcore_ary1_a0_I1_p0_l[6]));
INVX1 mul_U19005(.A(dpath_mulcore_ary1_a0_I1_p0_l[6]), .Y(n6476));
AND2X1 mul_U19006(.A(dpath_mulcore_b5[1]), .B(n11528), .Y(dpath_mulcore_ary1_a0_I1_p2_l[5]));
INVX1 mul_U19007(.A(dpath_mulcore_ary1_a0_I1_p2_l[5]), .Y(n6477));
AND2X1 mul_U19008(.A(dpath_mulcore_b4[1]), .B(n11531), .Y(dpath_mulcore_ary1_a0_I1_p1_l[5]));
INVX1 mul_U19009(.A(dpath_mulcore_ary1_a0_I1_p1_l[5]), .Y(n6478));
AND2X1 mul_U19010(.A(dpath_mulcore_b3[1]), .B(n11534), .Y(dpath_mulcore_ary1_a0_I1_p0_l[5]));
INVX1 mul_U19011(.A(dpath_mulcore_ary1_a0_I1_p0_l[5]), .Y(n6479));
AND2X1 mul_U19012(.A(dpath_mulcore_b5[1]), .B(n11536), .Y(dpath_mulcore_ary1_a0_I1_p2_l[4]));
INVX1 mul_U19013(.A(dpath_mulcore_ary1_a0_I1_p2_l[4]), .Y(n6480));
AND2X1 mul_U19014(.A(dpath_mulcore_b4[1]), .B(n11539), .Y(dpath_mulcore_ary1_a0_I1_p1_l[4]));
INVX1 mul_U19015(.A(dpath_mulcore_ary1_a0_I1_p1_l[4]), .Y(n6481));
AND2X1 mul_U19016(.A(dpath_mulcore_b3[1]), .B(n11542), .Y(dpath_mulcore_ary1_a0_I1_p0_l[4]));
INVX1 mul_U19017(.A(dpath_mulcore_ary1_a0_I1_p0_l[4]), .Y(n6482));
AND2X1 mul_U19018(.A(dpath_mulcore_b3[1]), .B(n11545), .Y(dpath_mulcore_ary1_a0_I1_p0_l[3]));
INVX1 mul_U19019(.A(dpath_mulcore_ary1_a0_I1_p0_l[3]), .Y(n6483));
AND2X1 mul_U19020(.A(dpath_mulcore_b4[1]), .B(n11548), .Y(dpath_mulcore_ary1_a0_I1_p1_l[3]));
INVX1 mul_U19021(.A(dpath_mulcore_ary1_a0_I1_p1_l[3]), .Y(n6484));
AND2X1 mul_U19022(.A(dpath_mulcore_b3[1]), .B(n11551), .Y(dpath_mulcore_ary1_a0_I1_I0_p0_l_2));
INVX1 mul_U19023(.A(dpath_mulcore_ary1_a0_I1_I0_p0_l_2), .Y(n6485));
AND2X1 mul_U19024(.A(dpath_mulcore_b3[1]), .B(n11554), .Y(dpath_mulcore_ary1_a0_I1_I0_p0_l_1));
INVX1 mul_U19025(.A(dpath_mulcore_ary1_a0_I1_I0_p0_l_1), .Y(n6486));
AND2X1 mul_U19026(.A(dpath_mulcore_b3[1]), .B(n11556), .Y(dpath_mulcore_ary1_a0_I1_I0_p0_l_0));
INVX1 mul_U19027(.A(dpath_mulcore_ary1_a0_I1_I0_p0_l_0), .Y(n6487));
AND2X1 mul_U19028(.A(dpath_mulcore_b4[1]), .B(n11558), .Y(dpath_mulcore_ary1_a0_I1_I0_p1_l_2));
INVX1 mul_U19029(.A(dpath_mulcore_ary1_a0_I1_I0_p1_l_2), .Y(n6488));
AND2X1 mul_U19030(.A(dpath_mulcore_b2[1]), .B(n11561), .Y(dpath_mulcore_ary1_a0_I0_I2_p2_l_67));
INVX1 mul_U19031(.A(dpath_mulcore_ary1_a0_I0_I2_p2_l_67), .Y(n6489));
AND2X1 mul_U19032(.A(dpath_mulcore_b2[1]), .B(n11564), .Y(dpath_mulcore_ary1_a0_I0_I2_p2_l_66));
INVX1 mul_U19033(.A(dpath_mulcore_ary1_a0_I0_I2_p2_l_66), .Y(n6490));
AND2X1 mul_U19034(.A(dpath_mulcore_b2[1]), .B(n11567), .Y(dpath_mulcore_ary1_a0_I0_I2_p2_l_65));
INVX1 mul_U19035(.A(dpath_mulcore_ary1_a0_I0_I2_p2_l_65), .Y(n6491));
AND2X1 mul_U19036(.A(dpath_mulcore_b1[1]), .B(n11570), .Y(dpath_mulcore_ary1_a0_I0_I2_p1_l_65));
INVX1 mul_U19037(.A(dpath_mulcore_ary1_a0_I0_I2_p1_l_65), .Y(n6492));
AND2X1 mul_U19038(.A(dpath_mulcore_b1[1]), .B(n11573), .Y(dpath_mulcore_ary1_a0_I0_I2_p1_l_64));
INVX1 mul_U19039(.A(dpath_mulcore_ary1_a0_I0_I2_p1_l_64), .Y(n6493));
AND2X1 mul_U19040(.A(dpath_mulcore_b2[1]), .B(n11576), .Y(dpath_mulcore_ary1_a0_I0_I2_p2_l_64));
INVX1 mul_U19041(.A(dpath_mulcore_ary1_a0_I0_I2_p2_l_64), .Y(n6494));
AND2X1 mul_U19042(.A(dpath_mulcore_b2[1]), .B(n11579), .Y(dpath_mulcore_ary1_a0_I0_p2_l[63]));
INVX1 mul_U19043(.A(dpath_mulcore_ary1_a0_I0_p2_l[63]), .Y(n6495));
AND2X1 mul_U19044(.A(dpath_mulcore_b1[1]), .B(n11582), .Y(dpath_mulcore_ary1_a0_I0_p1_l[63]));
INVX1 mul_U19045(.A(dpath_mulcore_ary1_a0_I0_p1_l[63]), .Y(n6496));
AND2X1 mul_U19046(.A(dpath_mulcore_b0[1]), .B(n11585), .Y(dpath_mulcore_ary1_a0_I0_p0_l[63]));
INVX1 mul_U19047(.A(dpath_mulcore_ary1_a0_I0_p0_l[63]), .Y(n6497));
AND2X1 mul_U19048(.A(dpath_mulcore_b2[1]), .B(n11588), .Y(dpath_mulcore_ary1_a0_I0_p2_l[62]));
INVX1 mul_U19049(.A(dpath_mulcore_ary1_a0_I0_p2_l[62]), .Y(n6498));
AND2X1 mul_U19050(.A(dpath_mulcore_b1[1]), .B(n11591), .Y(dpath_mulcore_ary1_a0_I0_p1_l[62]));
INVX1 mul_U19051(.A(dpath_mulcore_ary1_a0_I0_p1_l[62]), .Y(n6499));
AND2X1 mul_U19052(.A(dpath_mulcore_b0[1]), .B(n11594), .Y(dpath_mulcore_ary1_a0_I0_p0_l[62]));
INVX1 mul_U19053(.A(dpath_mulcore_ary1_a0_I0_p0_l[62]), .Y(n6500));
AND2X1 mul_U19054(.A(dpath_mulcore_b2[1]), .B(n11597), .Y(dpath_mulcore_ary1_a0_I0_p2_l[61]));
INVX1 mul_U19055(.A(dpath_mulcore_ary1_a0_I0_p2_l[61]), .Y(n6501));
AND2X1 mul_U19056(.A(dpath_mulcore_b1[1]), .B(n11600), .Y(dpath_mulcore_ary1_a0_I0_p1_l[61]));
INVX1 mul_U19057(.A(dpath_mulcore_ary1_a0_I0_p1_l[61]), .Y(n6502));
AND2X1 mul_U19058(.A(dpath_mulcore_b0[1]), .B(n11603), .Y(dpath_mulcore_ary1_a0_I0_p0_l[61]));
INVX1 mul_U19059(.A(dpath_mulcore_ary1_a0_I0_p0_l[61]), .Y(n6503));
AND2X1 mul_U19060(.A(dpath_mulcore_b2[1]), .B(n11606), .Y(dpath_mulcore_ary1_a0_I0_p2_l[60]));
INVX1 mul_U19061(.A(dpath_mulcore_ary1_a0_I0_p2_l[60]), .Y(n6504));
AND2X1 mul_U19062(.A(dpath_mulcore_b1[1]), .B(n11609), .Y(dpath_mulcore_ary1_a0_I0_p1_l[60]));
INVX1 mul_U19063(.A(dpath_mulcore_ary1_a0_I0_p1_l[60]), .Y(n6505));
AND2X1 mul_U19064(.A(dpath_mulcore_b0[1]), .B(n11612), .Y(dpath_mulcore_ary1_a0_I0_p0_l[60]));
INVX1 mul_U19065(.A(dpath_mulcore_ary1_a0_I0_p0_l[60]), .Y(n6506));
AND2X1 mul_U19066(.A(dpath_mulcore_b2[1]), .B(n11615), .Y(dpath_mulcore_ary1_a0_I0_p2_l[59]));
INVX1 mul_U19067(.A(dpath_mulcore_ary1_a0_I0_p2_l[59]), .Y(n6507));
AND2X1 mul_U19068(.A(dpath_mulcore_b1[1]), .B(n11618), .Y(dpath_mulcore_ary1_a0_I0_p1_l[59]));
INVX1 mul_U19069(.A(dpath_mulcore_ary1_a0_I0_p1_l[59]), .Y(n6508));
AND2X1 mul_U19070(.A(dpath_mulcore_b0[1]), .B(n11621), .Y(dpath_mulcore_ary1_a0_I0_p0_l[59]));
INVX1 mul_U19071(.A(dpath_mulcore_ary1_a0_I0_p0_l[59]), .Y(n6509));
AND2X1 mul_U19072(.A(dpath_mulcore_b2[1]), .B(n11624), .Y(dpath_mulcore_ary1_a0_I0_p2_l[58]));
INVX1 mul_U19073(.A(dpath_mulcore_ary1_a0_I0_p2_l[58]), .Y(n6510));
AND2X1 mul_U19074(.A(dpath_mulcore_b1[1]), .B(n11627), .Y(dpath_mulcore_ary1_a0_I0_p1_l[58]));
INVX1 mul_U19075(.A(dpath_mulcore_ary1_a0_I0_p1_l[58]), .Y(n6511));
AND2X1 mul_U19076(.A(dpath_mulcore_b0[1]), .B(n11630), .Y(dpath_mulcore_ary1_a0_I0_p0_l[58]));
INVX1 mul_U19077(.A(dpath_mulcore_ary1_a0_I0_p0_l[58]), .Y(n6512));
AND2X1 mul_U19078(.A(dpath_mulcore_b2[1]), .B(n11633), .Y(dpath_mulcore_ary1_a0_I0_p2_l[57]));
INVX1 mul_U19079(.A(dpath_mulcore_ary1_a0_I0_p2_l[57]), .Y(n6513));
AND2X1 mul_U19080(.A(dpath_mulcore_b1[1]), .B(n11636), .Y(dpath_mulcore_ary1_a0_I0_p1_l[57]));
INVX1 mul_U19081(.A(dpath_mulcore_ary1_a0_I0_p1_l[57]), .Y(n6514));
AND2X1 mul_U19082(.A(dpath_mulcore_b0[1]), .B(n11639), .Y(dpath_mulcore_ary1_a0_I0_p0_l[57]));
INVX1 mul_U19083(.A(dpath_mulcore_ary1_a0_I0_p0_l[57]), .Y(n6515));
AND2X1 mul_U19084(.A(dpath_mulcore_b2[1]), .B(n11642), .Y(dpath_mulcore_ary1_a0_I0_p2_l[56]));
INVX1 mul_U19085(.A(dpath_mulcore_ary1_a0_I0_p2_l[56]), .Y(n6516));
AND2X1 mul_U19086(.A(dpath_mulcore_b1[1]), .B(n11645), .Y(dpath_mulcore_ary1_a0_I0_p1_l[56]));
INVX1 mul_U19087(.A(dpath_mulcore_ary1_a0_I0_p1_l[56]), .Y(n6517));
AND2X1 mul_U19088(.A(dpath_mulcore_b0[1]), .B(n11648), .Y(dpath_mulcore_ary1_a0_I0_p0_l[56]));
INVX1 mul_U19089(.A(dpath_mulcore_ary1_a0_I0_p0_l[56]), .Y(n6518));
AND2X1 mul_U19090(.A(dpath_mulcore_b2[1]), .B(n11651), .Y(dpath_mulcore_ary1_a0_I0_p2_l[55]));
INVX1 mul_U19091(.A(dpath_mulcore_ary1_a0_I0_p2_l[55]), .Y(n6519));
AND2X1 mul_U19092(.A(dpath_mulcore_b1[1]), .B(n11654), .Y(dpath_mulcore_ary1_a0_I0_p1_l[55]));
INVX1 mul_U19093(.A(dpath_mulcore_ary1_a0_I0_p1_l[55]), .Y(n6520));
AND2X1 mul_U19094(.A(dpath_mulcore_b0[1]), .B(n11657), .Y(dpath_mulcore_ary1_a0_I0_p0_l[55]));
INVX1 mul_U19095(.A(dpath_mulcore_ary1_a0_I0_p0_l[55]), .Y(n6521));
AND2X1 mul_U19096(.A(dpath_mulcore_b2[1]), .B(n11660), .Y(dpath_mulcore_ary1_a0_I0_p2_l[54]));
INVX1 mul_U19097(.A(dpath_mulcore_ary1_a0_I0_p2_l[54]), .Y(n6522));
AND2X1 mul_U19098(.A(dpath_mulcore_b1[1]), .B(n11663), .Y(dpath_mulcore_ary1_a0_I0_p1_l[54]));
INVX1 mul_U19099(.A(dpath_mulcore_ary1_a0_I0_p1_l[54]), .Y(n6523));
AND2X1 mul_U19100(.A(dpath_mulcore_b0[1]), .B(n11666), .Y(dpath_mulcore_ary1_a0_I0_p0_l[54]));
INVX1 mul_U19101(.A(dpath_mulcore_ary1_a0_I0_p0_l[54]), .Y(n6524));
AND2X1 mul_U19102(.A(dpath_mulcore_b2[1]), .B(n11669), .Y(dpath_mulcore_ary1_a0_I0_p2_l[53]));
INVX1 mul_U19103(.A(dpath_mulcore_ary1_a0_I0_p2_l[53]), .Y(n6525));
AND2X1 mul_U19104(.A(dpath_mulcore_b1[1]), .B(n11672), .Y(dpath_mulcore_ary1_a0_I0_p1_l[53]));
INVX1 mul_U19105(.A(dpath_mulcore_ary1_a0_I0_p1_l[53]), .Y(n6526));
AND2X1 mul_U19106(.A(dpath_mulcore_b0[1]), .B(n11675), .Y(dpath_mulcore_ary1_a0_I0_p0_l[53]));
INVX1 mul_U19107(.A(dpath_mulcore_ary1_a0_I0_p0_l[53]), .Y(n6527));
AND2X1 mul_U19108(.A(dpath_mulcore_b2[1]), .B(n11678), .Y(dpath_mulcore_ary1_a0_I0_p2_l[52]));
INVX1 mul_U19109(.A(dpath_mulcore_ary1_a0_I0_p2_l[52]), .Y(n6528));
AND2X1 mul_U19110(.A(dpath_mulcore_b1[1]), .B(n11681), .Y(dpath_mulcore_ary1_a0_I0_p1_l[52]));
INVX1 mul_U19111(.A(dpath_mulcore_ary1_a0_I0_p1_l[52]), .Y(n6529));
AND2X1 mul_U19112(.A(dpath_mulcore_b0[1]), .B(n11684), .Y(dpath_mulcore_ary1_a0_I0_p0_l[52]));
INVX1 mul_U19113(.A(dpath_mulcore_ary1_a0_I0_p0_l[52]), .Y(n6530));
AND2X1 mul_U19114(.A(dpath_mulcore_b2[1]), .B(n11687), .Y(dpath_mulcore_ary1_a0_I0_p2_l[51]));
INVX1 mul_U19115(.A(dpath_mulcore_ary1_a0_I0_p2_l[51]), .Y(n6531));
AND2X1 mul_U19116(.A(dpath_mulcore_b1[1]), .B(n11690), .Y(dpath_mulcore_ary1_a0_I0_p1_l[51]));
INVX1 mul_U19117(.A(dpath_mulcore_ary1_a0_I0_p1_l[51]), .Y(n6532));
AND2X1 mul_U19118(.A(dpath_mulcore_b0[1]), .B(n11693), .Y(dpath_mulcore_ary1_a0_I0_p0_l[51]));
INVX1 mul_U19119(.A(dpath_mulcore_ary1_a0_I0_p0_l[51]), .Y(n6533));
AND2X1 mul_U19120(.A(dpath_mulcore_b2[1]), .B(n11696), .Y(dpath_mulcore_ary1_a0_I0_p2_l[50]));
INVX1 mul_U19121(.A(dpath_mulcore_ary1_a0_I0_p2_l[50]), .Y(n6534));
AND2X1 mul_U19122(.A(dpath_mulcore_b1[1]), .B(n11699), .Y(dpath_mulcore_ary1_a0_I0_p1_l[50]));
INVX1 mul_U19123(.A(dpath_mulcore_ary1_a0_I0_p1_l[50]), .Y(n6535));
AND2X1 mul_U19124(.A(dpath_mulcore_b0[1]), .B(n11702), .Y(dpath_mulcore_ary1_a0_I0_p0_l[50]));
INVX1 mul_U19125(.A(dpath_mulcore_ary1_a0_I0_p0_l[50]), .Y(n6536));
AND2X1 mul_U19126(.A(dpath_mulcore_b2[1]), .B(n11705), .Y(dpath_mulcore_ary1_a0_I0_p2_l[49]));
INVX1 mul_U19127(.A(dpath_mulcore_ary1_a0_I0_p2_l[49]), .Y(n6537));
AND2X1 mul_U19128(.A(dpath_mulcore_b1[1]), .B(n11708), .Y(dpath_mulcore_ary1_a0_I0_p1_l[49]));
INVX1 mul_U19129(.A(dpath_mulcore_ary1_a0_I0_p1_l[49]), .Y(n6538));
AND2X1 mul_U19130(.A(dpath_mulcore_b0[1]), .B(n11711), .Y(dpath_mulcore_ary1_a0_I0_p0_l[49]));
INVX1 mul_U19131(.A(dpath_mulcore_ary1_a0_I0_p0_l[49]), .Y(n6539));
AND2X1 mul_U19132(.A(dpath_mulcore_b2[1]), .B(n11714), .Y(dpath_mulcore_ary1_a0_I0_p2_l[48]));
INVX1 mul_U19133(.A(dpath_mulcore_ary1_a0_I0_p2_l[48]), .Y(n6540));
AND2X1 mul_U19134(.A(dpath_mulcore_b1[1]), .B(n11717), .Y(dpath_mulcore_ary1_a0_I0_p1_l[48]));
INVX1 mul_U19135(.A(dpath_mulcore_ary1_a0_I0_p1_l[48]), .Y(n6541));
AND2X1 mul_U19136(.A(dpath_mulcore_b0[1]), .B(n11720), .Y(dpath_mulcore_ary1_a0_I0_p0_l[48]));
INVX1 mul_U19137(.A(dpath_mulcore_ary1_a0_I0_p0_l[48]), .Y(n6542));
AND2X1 mul_U19138(.A(dpath_mulcore_b2[1]), .B(n11723), .Y(dpath_mulcore_ary1_a0_I0_p2_l[47]));
INVX1 mul_U19139(.A(dpath_mulcore_ary1_a0_I0_p2_l[47]), .Y(n6543));
AND2X1 mul_U19140(.A(dpath_mulcore_b1[1]), .B(n11726), .Y(dpath_mulcore_ary1_a0_I0_p1_l[47]));
INVX1 mul_U19141(.A(dpath_mulcore_ary1_a0_I0_p1_l[47]), .Y(n6544));
AND2X1 mul_U19142(.A(dpath_mulcore_b0[1]), .B(n11729), .Y(dpath_mulcore_ary1_a0_I0_p0_l[47]));
INVX1 mul_U19143(.A(dpath_mulcore_ary1_a0_I0_p0_l[47]), .Y(n6545));
AND2X1 mul_U19144(.A(dpath_mulcore_b2[1]), .B(n11732), .Y(dpath_mulcore_ary1_a0_I0_p2_l[46]));
INVX1 mul_U19145(.A(dpath_mulcore_ary1_a0_I0_p2_l[46]), .Y(n6546));
AND2X1 mul_U19146(.A(dpath_mulcore_b1[1]), .B(n11735), .Y(dpath_mulcore_ary1_a0_I0_p1_l[46]));
INVX1 mul_U19147(.A(dpath_mulcore_ary1_a0_I0_p1_l[46]), .Y(n6547));
AND2X1 mul_U19148(.A(dpath_mulcore_b0[1]), .B(n11738), .Y(dpath_mulcore_ary1_a0_I0_p0_l[46]));
INVX1 mul_U19149(.A(dpath_mulcore_ary1_a0_I0_p0_l[46]), .Y(n6548));
AND2X1 mul_U19150(.A(dpath_mulcore_b2[1]), .B(n11741), .Y(dpath_mulcore_ary1_a0_I0_p2_l[45]));
INVX1 mul_U19151(.A(dpath_mulcore_ary1_a0_I0_p2_l[45]), .Y(n6549));
AND2X1 mul_U19152(.A(dpath_mulcore_b1[1]), .B(n11744), .Y(dpath_mulcore_ary1_a0_I0_p1_l[45]));
INVX1 mul_U19153(.A(dpath_mulcore_ary1_a0_I0_p1_l[45]), .Y(n6550));
AND2X1 mul_U19154(.A(dpath_mulcore_b0[1]), .B(n11747), .Y(dpath_mulcore_ary1_a0_I0_p0_l[45]));
INVX1 mul_U19155(.A(dpath_mulcore_ary1_a0_I0_p0_l[45]), .Y(n6551));
AND2X1 mul_U19156(.A(dpath_mulcore_b2[1]), .B(n11750), .Y(dpath_mulcore_ary1_a0_I0_p2_l[44]));
INVX1 mul_U19157(.A(dpath_mulcore_ary1_a0_I0_p2_l[44]), .Y(n6552));
AND2X1 mul_U19158(.A(dpath_mulcore_b1[1]), .B(n11753), .Y(dpath_mulcore_ary1_a0_I0_p1_l[44]));
INVX1 mul_U19159(.A(dpath_mulcore_ary1_a0_I0_p1_l[44]), .Y(n6553));
AND2X1 mul_U19160(.A(dpath_mulcore_b0[1]), .B(n11756), .Y(dpath_mulcore_ary1_a0_I0_p0_l[44]));
INVX1 mul_U19161(.A(dpath_mulcore_ary1_a0_I0_p0_l[44]), .Y(n6554));
AND2X1 mul_U19162(.A(dpath_mulcore_b2[1]), .B(n11759), .Y(dpath_mulcore_ary1_a0_I0_p2_l[43]));
INVX1 mul_U19163(.A(dpath_mulcore_ary1_a0_I0_p2_l[43]), .Y(n6555));
AND2X1 mul_U19164(.A(dpath_mulcore_b1[1]), .B(n11762), .Y(dpath_mulcore_ary1_a0_I0_p1_l[43]));
INVX1 mul_U19165(.A(dpath_mulcore_ary1_a0_I0_p1_l[43]), .Y(n6556));
AND2X1 mul_U19166(.A(dpath_mulcore_b0[1]), .B(n11765), .Y(dpath_mulcore_ary1_a0_I0_p0_l[43]));
INVX1 mul_U19167(.A(dpath_mulcore_ary1_a0_I0_p0_l[43]), .Y(n6557));
AND2X1 mul_U19168(.A(dpath_mulcore_b2[1]), .B(n11768), .Y(dpath_mulcore_ary1_a0_I0_p2_l[42]));
INVX1 mul_U19169(.A(dpath_mulcore_ary1_a0_I0_p2_l[42]), .Y(n6558));
AND2X1 mul_U19170(.A(dpath_mulcore_b1[1]), .B(n11771), .Y(dpath_mulcore_ary1_a0_I0_p1_l[42]));
INVX1 mul_U19171(.A(dpath_mulcore_ary1_a0_I0_p1_l[42]), .Y(n6559));
AND2X1 mul_U19172(.A(dpath_mulcore_b0[1]), .B(n11774), .Y(dpath_mulcore_ary1_a0_I0_p0_l[42]));
INVX1 mul_U19173(.A(dpath_mulcore_ary1_a0_I0_p0_l[42]), .Y(n6560));
AND2X1 mul_U19174(.A(dpath_mulcore_b2[1]), .B(n11777), .Y(dpath_mulcore_ary1_a0_I0_p2_l[41]));
INVX1 mul_U19175(.A(dpath_mulcore_ary1_a0_I0_p2_l[41]), .Y(n6561));
AND2X1 mul_U19176(.A(dpath_mulcore_b1[1]), .B(n11780), .Y(dpath_mulcore_ary1_a0_I0_p1_l[41]));
INVX1 mul_U19177(.A(dpath_mulcore_ary1_a0_I0_p1_l[41]), .Y(n6562));
AND2X1 mul_U19178(.A(dpath_mulcore_b0[1]), .B(n11783), .Y(dpath_mulcore_ary1_a0_I0_p0_l[41]));
INVX1 mul_U19179(.A(dpath_mulcore_ary1_a0_I0_p0_l[41]), .Y(n6563));
AND2X1 mul_U19180(.A(dpath_mulcore_b2[1]), .B(n11786), .Y(dpath_mulcore_ary1_a0_I0_p2_l[40]));
INVX1 mul_U19181(.A(dpath_mulcore_ary1_a0_I0_p2_l[40]), .Y(n6564));
AND2X1 mul_U19182(.A(dpath_mulcore_b1[1]), .B(n11789), .Y(dpath_mulcore_ary1_a0_I0_p1_l[40]));
INVX1 mul_U19183(.A(dpath_mulcore_ary1_a0_I0_p1_l[40]), .Y(n6565));
AND2X1 mul_U19184(.A(dpath_mulcore_b0[1]), .B(n11792), .Y(dpath_mulcore_ary1_a0_I0_p0_l[40]));
INVX1 mul_U19185(.A(dpath_mulcore_ary1_a0_I0_p0_l[40]), .Y(n6566));
AND2X1 mul_U19186(.A(dpath_mulcore_b2[1]), .B(n11795), .Y(dpath_mulcore_ary1_a0_I0_p2_l[39]));
INVX1 mul_U19187(.A(dpath_mulcore_ary1_a0_I0_p2_l[39]), .Y(n6567));
AND2X1 mul_U19188(.A(dpath_mulcore_b1[1]), .B(n11798), .Y(dpath_mulcore_ary1_a0_I0_p1_l[39]));
INVX1 mul_U19189(.A(dpath_mulcore_ary1_a0_I0_p1_l[39]), .Y(n6568));
AND2X1 mul_U19190(.A(dpath_mulcore_b0[1]), .B(n11801), .Y(dpath_mulcore_ary1_a0_I0_p0_l[39]));
INVX1 mul_U19191(.A(dpath_mulcore_ary1_a0_I0_p0_l[39]), .Y(n6569));
AND2X1 mul_U19192(.A(dpath_mulcore_b2[1]), .B(n11804), .Y(dpath_mulcore_ary1_a0_I0_p2_l[38]));
INVX1 mul_U19193(.A(dpath_mulcore_ary1_a0_I0_p2_l[38]), .Y(n6570));
AND2X1 mul_U19194(.A(dpath_mulcore_b1[1]), .B(n11807), .Y(dpath_mulcore_ary1_a0_I0_p1_l[38]));
INVX1 mul_U19195(.A(dpath_mulcore_ary1_a0_I0_p1_l[38]), .Y(n6571));
AND2X1 mul_U19196(.A(dpath_mulcore_b0[1]), .B(n11810), .Y(dpath_mulcore_ary1_a0_I0_p0_l[38]));
INVX1 mul_U19197(.A(dpath_mulcore_ary1_a0_I0_p0_l[38]), .Y(n6572));
AND2X1 mul_U19198(.A(dpath_mulcore_b2[1]), .B(n11813), .Y(dpath_mulcore_ary1_a0_I0_p2_l[37]));
INVX1 mul_U19199(.A(dpath_mulcore_ary1_a0_I0_p2_l[37]), .Y(n6573));
AND2X1 mul_U19200(.A(dpath_mulcore_b1[1]), .B(n11816), .Y(dpath_mulcore_ary1_a0_I0_p1_l[37]));
INVX1 mul_U19201(.A(dpath_mulcore_ary1_a0_I0_p1_l[37]), .Y(n6574));
AND2X1 mul_U19202(.A(dpath_mulcore_b0[1]), .B(n11819), .Y(dpath_mulcore_ary1_a0_I0_p0_l[37]));
INVX1 mul_U19203(.A(dpath_mulcore_ary1_a0_I0_p0_l[37]), .Y(n6575));
AND2X1 mul_U19204(.A(dpath_mulcore_b2[1]), .B(n11822), .Y(dpath_mulcore_ary1_a0_I0_p2_l[36]));
INVX1 mul_U19205(.A(dpath_mulcore_ary1_a0_I0_p2_l[36]), .Y(n6576));
AND2X1 mul_U19206(.A(dpath_mulcore_b1[1]), .B(n11825), .Y(dpath_mulcore_ary1_a0_I0_p1_l[36]));
INVX1 mul_U19207(.A(dpath_mulcore_ary1_a0_I0_p1_l[36]), .Y(n6577));
AND2X1 mul_U19208(.A(dpath_mulcore_b0[1]), .B(n11828), .Y(dpath_mulcore_ary1_a0_I0_p0_l[36]));
INVX1 mul_U19209(.A(dpath_mulcore_ary1_a0_I0_p0_l[36]), .Y(n6578));
AND2X1 mul_U19210(.A(dpath_mulcore_b2[1]), .B(n11831), .Y(dpath_mulcore_ary1_a0_I0_p2_l[35]));
INVX1 mul_U19211(.A(dpath_mulcore_ary1_a0_I0_p2_l[35]), .Y(n6579));
AND2X1 mul_U19212(.A(dpath_mulcore_b1[1]), .B(n11834), .Y(dpath_mulcore_ary1_a0_I0_p1_l[35]));
INVX1 mul_U19213(.A(dpath_mulcore_ary1_a0_I0_p1_l[35]), .Y(n6580));
AND2X1 mul_U19214(.A(dpath_mulcore_b0[1]), .B(n11837), .Y(dpath_mulcore_ary1_a0_I0_p0_l[35]));
INVX1 mul_U19215(.A(dpath_mulcore_ary1_a0_I0_p0_l[35]), .Y(n6581));
AND2X1 mul_U19216(.A(dpath_mulcore_b2[1]), .B(n11840), .Y(dpath_mulcore_ary1_a0_I0_p2_l[34]));
INVX1 mul_U19217(.A(dpath_mulcore_ary1_a0_I0_p2_l[34]), .Y(n6582));
AND2X1 mul_U19218(.A(dpath_mulcore_b1[1]), .B(n11843), .Y(dpath_mulcore_ary1_a0_I0_p1_l[34]));
INVX1 mul_U19219(.A(dpath_mulcore_ary1_a0_I0_p1_l[34]), .Y(n6583));
AND2X1 mul_U19220(.A(dpath_mulcore_b0[1]), .B(n11846), .Y(dpath_mulcore_ary1_a0_I0_p0_l[34]));
INVX1 mul_U19221(.A(dpath_mulcore_ary1_a0_I0_p0_l[34]), .Y(n6584));
AND2X1 mul_U19222(.A(dpath_mulcore_b2[1]), .B(n11849), .Y(dpath_mulcore_ary1_a0_I0_p2_l[33]));
INVX1 mul_U19223(.A(dpath_mulcore_ary1_a0_I0_p2_l[33]), .Y(n6585));
AND2X1 mul_U19224(.A(dpath_mulcore_b1[1]), .B(n11852), .Y(dpath_mulcore_ary1_a0_I0_p1_l[33]));
INVX1 mul_U19225(.A(dpath_mulcore_ary1_a0_I0_p1_l[33]), .Y(n6586));
AND2X1 mul_U19226(.A(dpath_mulcore_b0[1]), .B(n11855), .Y(dpath_mulcore_ary1_a0_I0_p0_l[33]));
INVX1 mul_U19227(.A(dpath_mulcore_ary1_a0_I0_p0_l[33]), .Y(n6587));
AND2X1 mul_U19228(.A(dpath_mulcore_b2[1]), .B(n11858), .Y(dpath_mulcore_ary1_a0_I0_p2_l[32]));
INVX1 mul_U19229(.A(dpath_mulcore_ary1_a0_I0_p2_l[32]), .Y(n6588));
AND2X1 mul_U19230(.A(dpath_mulcore_b1[1]), .B(n11861), .Y(dpath_mulcore_ary1_a0_I0_p1_l[32]));
INVX1 mul_U19231(.A(dpath_mulcore_ary1_a0_I0_p1_l[32]), .Y(n6589));
AND2X1 mul_U19232(.A(dpath_mulcore_b0[1]), .B(n11864), .Y(dpath_mulcore_ary1_a0_I0_p0_l[32]));
INVX1 mul_U19233(.A(dpath_mulcore_ary1_a0_I0_p0_l[32]), .Y(n6590));
AND2X1 mul_U19234(.A(dpath_mulcore_b2[1]), .B(n11867), .Y(dpath_mulcore_ary1_a0_I0_p2_l[31]));
INVX1 mul_U19235(.A(dpath_mulcore_ary1_a0_I0_p2_l[31]), .Y(n6591));
AND2X1 mul_U19236(.A(dpath_mulcore_b1[1]), .B(n11870), .Y(dpath_mulcore_ary1_a0_I0_p1_l[31]));
INVX1 mul_U19237(.A(dpath_mulcore_ary1_a0_I0_p1_l[31]), .Y(n6592));
AND2X1 mul_U19238(.A(dpath_mulcore_b0[1]), .B(n11873), .Y(dpath_mulcore_ary1_a0_I0_p0_l[31]));
INVX1 mul_U19239(.A(dpath_mulcore_ary1_a0_I0_p0_l[31]), .Y(n6593));
AND2X1 mul_U19240(.A(dpath_mulcore_b2[1]), .B(n11876), .Y(dpath_mulcore_ary1_a0_I0_p2_l[30]));
INVX1 mul_U19241(.A(dpath_mulcore_ary1_a0_I0_p2_l[30]), .Y(n6594));
AND2X1 mul_U19242(.A(dpath_mulcore_b1[1]), .B(n11879), .Y(dpath_mulcore_ary1_a0_I0_p1_l[30]));
INVX1 mul_U19243(.A(dpath_mulcore_ary1_a0_I0_p1_l[30]), .Y(n6595));
AND2X1 mul_U19244(.A(dpath_mulcore_b0[1]), .B(n11882), .Y(dpath_mulcore_ary1_a0_I0_p0_l[30]));
INVX1 mul_U19245(.A(dpath_mulcore_ary1_a0_I0_p0_l[30]), .Y(n6596));
AND2X1 mul_U19246(.A(dpath_mulcore_b2[1]), .B(n11885), .Y(dpath_mulcore_ary1_a0_I0_p2_l[29]));
INVX1 mul_U19247(.A(dpath_mulcore_ary1_a0_I0_p2_l[29]), .Y(n6597));
AND2X1 mul_U19248(.A(dpath_mulcore_b1[1]), .B(n11888), .Y(dpath_mulcore_ary1_a0_I0_p1_l[29]));
INVX1 mul_U19249(.A(dpath_mulcore_ary1_a0_I0_p1_l[29]), .Y(n6598));
AND2X1 mul_U19250(.A(dpath_mulcore_b0[1]), .B(n11891), .Y(dpath_mulcore_ary1_a0_I0_p0_l[29]));
INVX1 mul_U19251(.A(dpath_mulcore_ary1_a0_I0_p0_l[29]), .Y(n6599));
AND2X1 mul_U19252(.A(dpath_mulcore_b2[1]), .B(n11894), .Y(dpath_mulcore_ary1_a0_I0_p2_l[28]));
INVX1 mul_U19253(.A(dpath_mulcore_ary1_a0_I0_p2_l[28]), .Y(n6600));
AND2X1 mul_U19254(.A(dpath_mulcore_b1[1]), .B(n11897), .Y(dpath_mulcore_ary1_a0_I0_p1_l[28]));
INVX1 mul_U19255(.A(dpath_mulcore_ary1_a0_I0_p1_l[28]), .Y(n6601));
AND2X1 mul_U19256(.A(dpath_mulcore_b0[1]), .B(n11900), .Y(dpath_mulcore_ary1_a0_I0_p0_l[28]));
INVX1 mul_U19257(.A(dpath_mulcore_ary1_a0_I0_p0_l[28]), .Y(n6602));
AND2X1 mul_U19258(.A(dpath_mulcore_b2[1]), .B(n11903), .Y(dpath_mulcore_ary1_a0_I0_p2_l[27]));
INVX1 mul_U19259(.A(dpath_mulcore_ary1_a0_I0_p2_l[27]), .Y(n6603));
AND2X1 mul_U19260(.A(dpath_mulcore_b1[1]), .B(n11906), .Y(dpath_mulcore_ary1_a0_I0_p1_l[27]));
INVX1 mul_U19261(.A(dpath_mulcore_ary1_a0_I0_p1_l[27]), .Y(n6604));
AND2X1 mul_U19262(.A(dpath_mulcore_b0[1]), .B(n11909), .Y(dpath_mulcore_ary1_a0_I0_p0_l[27]));
INVX1 mul_U19263(.A(dpath_mulcore_ary1_a0_I0_p0_l[27]), .Y(n6605));
AND2X1 mul_U19264(.A(dpath_mulcore_b2[1]), .B(n11912), .Y(dpath_mulcore_ary1_a0_I0_p2_l[26]));
INVX1 mul_U19265(.A(dpath_mulcore_ary1_a0_I0_p2_l[26]), .Y(n6606));
AND2X1 mul_U19266(.A(dpath_mulcore_b1[1]), .B(n11915), .Y(dpath_mulcore_ary1_a0_I0_p1_l[26]));
INVX1 mul_U19267(.A(dpath_mulcore_ary1_a0_I0_p1_l[26]), .Y(n6607));
AND2X1 mul_U19268(.A(dpath_mulcore_b0[1]), .B(n11918), .Y(dpath_mulcore_ary1_a0_I0_p0_l[26]));
INVX1 mul_U19269(.A(dpath_mulcore_ary1_a0_I0_p0_l[26]), .Y(n6608));
AND2X1 mul_U19270(.A(dpath_mulcore_b2[1]), .B(n11921), .Y(dpath_mulcore_ary1_a0_I0_p2_l[25]));
INVX1 mul_U19271(.A(dpath_mulcore_ary1_a0_I0_p2_l[25]), .Y(n6609));
AND2X1 mul_U19272(.A(dpath_mulcore_b1[1]), .B(n11924), .Y(dpath_mulcore_ary1_a0_I0_p1_l[25]));
INVX1 mul_U19273(.A(dpath_mulcore_ary1_a0_I0_p1_l[25]), .Y(n6610));
AND2X1 mul_U19274(.A(dpath_mulcore_b0[1]), .B(n11927), .Y(dpath_mulcore_ary1_a0_I0_p0_l[25]));
INVX1 mul_U19275(.A(dpath_mulcore_ary1_a0_I0_p0_l[25]), .Y(n6611));
AND2X1 mul_U19276(.A(dpath_mulcore_b2[1]), .B(n11930), .Y(dpath_mulcore_ary1_a0_I0_p2_l[24]));
INVX1 mul_U19277(.A(dpath_mulcore_ary1_a0_I0_p2_l[24]), .Y(n6612));
AND2X1 mul_U19278(.A(dpath_mulcore_b1[1]), .B(n11933), .Y(dpath_mulcore_ary1_a0_I0_p1_l[24]));
INVX1 mul_U19279(.A(dpath_mulcore_ary1_a0_I0_p1_l[24]), .Y(n6613));
AND2X1 mul_U19280(.A(dpath_mulcore_b0[1]), .B(n11936), .Y(dpath_mulcore_ary1_a0_I0_p0_l[24]));
INVX1 mul_U19281(.A(dpath_mulcore_ary1_a0_I0_p0_l[24]), .Y(n6614));
AND2X1 mul_U19282(.A(dpath_mulcore_b2[1]), .B(n11939), .Y(dpath_mulcore_ary1_a0_I0_p2_l[23]));
INVX1 mul_U19283(.A(dpath_mulcore_ary1_a0_I0_p2_l[23]), .Y(n6615));
AND2X1 mul_U19284(.A(dpath_mulcore_b1[1]), .B(n11942), .Y(dpath_mulcore_ary1_a0_I0_p1_l[23]));
INVX1 mul_U19285(.A(dpath_mulcore_ary1_a0_I0_p1_l[23]), .Y(n6616));
AND2X1 mul_U19286(.A(dpath_mulcore_b0[1]), .B(n11945), .Y(dpath_mulcore_ary1_a0_I0_p0_l[23]));
INVX1 mul_U19287(.A(dpath_mulcore_ary1_a0_I0_p0_l[23]), .Y(n6617));
AND2X1 mul_U19288(.A(dpath_mulcore_b2[1]), .B(n11948), .Y(dpath_mulcore_ary1_a0_I0_p2_l[22]));
INVX1 mul_U19289(.A(dpath_mulcore_ary1_a0_I0_p2_l[22]), .Y(n6618));
AND2X1 mul_U19290(.A(dpath_mulcore_b1[1]), .B(n11951), .Y(dpath_mulcore_ary1_a0_I0_p1_l[22]));
INVX1 mul_U19291(.A(dpath_mulcore_ary1_a0_I0_p1_l[22]), .Y(n6619));
AND2X1 mul_U19292(.A(dpath_mulcore_b0[1]), .B(n11954), .Y(dpath_mulcore_ary1_a0_I0_p0_l[22]));
INVX1 mul_U19293(.A(dpath_mulcore_ary1_a0_I0_p0_l[22]), .Y(n6620));
AND2X1 mul_U19294(.A(dpath_mulcore_b2[1]), .B(n11957), .Y(dpath_mulcore_ary1_a0_I0_p2_l[21]));
INVX1 mul_U19295(.A(dpath_mulcore_ary1_a0_I0_p2_l[21]), .Y(n6621));
AND2X1 mul_U19296(.A(dpath_mulcore_b1[1]), .B(n11960), .Y(dpath_mulcore_ary1_a0_I0_p1_l[21]));
INVX1 mul_U19297(.A(dpath_mulcore_ary1_a0_I0_p1_l[21]), .Y(n6622));
AND2X1 mul_U19298(.A(dpath_mulcore_b0[1]), .B(n11963), .Y(dpath_mulcore_ary1_a0_I0_p0_l[21]));
INVX1 mul_U19299(.A(dpath_mulcore_ary1_a0_I0_p0_l[21]), .Y(n6623));
AND2X1 mul_U19300(.A(dpath_mulcore_b2[1]), .B(n11966), .Y(dpath_mulcore_ary1_a0_I0_p2_l[20]));
INVX1 mul_U19301(.A(dpath_mulcore_ary1_a0_I0_p2_l[20]), .Y(n6624));
AND2X1 mul_U19302(.A(dpath_mulcore_b1[1]), .B(n11969), .Y(dpath_mulcore_ary1_a0_I0_p1_l[20]));
INVX1 mul_U19303(.A(dpath_mulcore_ary1_a0_I0_p1_l[20]), .Y(n6625));
AND2X1 mul_U19304(.A(dpath_mulcore_b0[1]), .B(n11972), .Y(dpath_mulcore_ary1_a0_I0_p0_l[20]));
INVX1 mul_U19305(.A(dpath_mulcore_ary1_a0_I0_p0_l[20]), .Y(n6626));
AND2X1 mul_U19306(.A(dpath_mulcore_b2[1]), .B(n11975), .Y(dpath_mulcore_ary1_a0_I0_p2_l[19]));
INVX1 mul_U19307(.A(dpath_mulcore_ary1_a0_I0_p2_l[19]), .Y(n6627));
AND2X1 mul_U19308(.A(dpath_mulcore_b1[1]), .B(n11978), .Y(dpath_mulcore_ary1_a0_I0_p1_l[19]));
INVX1 mul_U19309(.A(dpath_mulcore_ary1_a0_I0_p1_l[19]), .Y(n6628));
AND2X1 mul_U19310(.A(dpath_mulcore_b0[1]), .B(n11981), .Y(dpath_mulcore_ary1_a0_I0_p0_l[19]));
INVX1 mul_U19311(.A(dpath_mulcore_ary1_a0_I0_p0_l[19]), .Y(n6629));
AND2X1 mul_U19312(.A(dpath_mulcore_b2[1]), .B(n11984), .Y(dpath_mulcore_ary1_a0_I0_p2_l[18]));
INVX1 mul_U19313(.A(dpath_mulcore_ary1_a0_I0_p2_l[18]), .Y(n6630));
AND2X1 mul_U19314(.A(dpath_mulcore_b1[1]), .B(n11987), .Y(dpath_mulcore_ary1_a0_I0_p1_l[18]));
INVX1 mul_U19315(.A(dpath_mulcore_ary1_a0_I0_p1_l[18]), .Y(n6631));
AND2X1 mul_U19316(.A(dpath_mulcore_b0[1]), .B(n11990), .Y(dpath_mulcore_ary1_a0_I0_p0_l[18]));
INVX1 mul_U19317(.A(dpath_mulcore_ary1_a0_I0_p0_l[18]), .Y(n6632));
AND2X1 mul_U19318(.A(dpath_mulcore_b2[1]), .B(n11993), .Y(dpath_mulcore_ary1_a0_I0_p2_l[17]));
INVX1 mul_U19319(.A(dpath_mulcore_ary1_a0_I0_p2_l[17]), .Y(n6633));
AND2X1 mul_U19320(.A(dpath_mulcore_b1[1]), .B(n11996), .Y(dpath_mulcore_ary1_a0_I0_p1_l[17]));
INVX1 mul_U19321(.A(dpath_mulcore_ary1_a0_I0_p1_l[17]), .Y(n6634));
AND2X1 mul_U19322(.A(dpath_mulcore_b0[1]), .B(n11999), .Y(dpath_mulcore_ary1_a0_I0_p0_l[17]));
INVX1 mul_U19323(.A(dpath_mulcore_ary1_a0_I0_p0_l[17]), .Y(n6635));
AND2X1 mul_U19324(.A(dpath_mulcore_b2[1]), .B(n12002), .Y(dpath_mulcore_ary1_a0_I0_p2_l[16]));
INVX1 mul_U19325(.A(dpath_mulcore_ary1_a0_I0_p2_l[16]), .Y(n6636));
AND2X1 mul_U19326(.A(dpath_mulcore_b1[1]), .B(n12005), .Y(dpath_mulcore_ary1_a0_I0_p1_l[16]));
INVX1 mul_U19327(.A(dpath_mulcore_ary1_a0_I0_p1_l[16]), .Y(n6637));
AND2X1 mul_U19328(.A(dpath_mulcore_b0[1]), .B(n12008), .Y(dpath_mulcore_ary1_a0_I0_p0_l[16]));
INVX1 mul_U19329(.A(dpath_mulcore_ary1_a0_I0_p0_l[16]), .Y(n6638));
AND2X1 mul_U19330(.A(dpath_mulcore_b2[1]), .B(n12011), .Y(dpath_mulcore_ary1_a0_I0_p2_l[15]));
INVX1 mul_U19331(.A(dpath_mulcore_ary1_a0_I0_p2_l[15]), .Y(n6639));
AND2X1 mul_U19332(.A(dpath_mulcore_b1[1]), .B(n12014), .Y(dpath_mulcore_ary1_a0_I0_p1_l[15]));
INVX1 mul_U19333(.A(dpath_mulcore_ary1_a0_I0_p1_l[15]), .Y(n6640));
AND2X1 mul_U19334(.A(dpath_mulcore_b0[1]), .B(n12017), .Y(dpath_mulcore_ary1_a0_I0_p0_l[15]));
INVX1 mul_U19335(.A(dpath_mulcore_ary1_a0_I0_p0_l[15]), .Y(n6641));
AND2X1 mul_U19336(.A(dpath_mulcore_b2[1]), .B(n12020), .Y(dpath_mulcore_ary1_a0_I0_p2_l[14]));
INVX1 mul_U19337(.A(dpath_mulcore_ary1_a0_I0_p2_l[14]), .Y(n6642));
AND2X1 mul_U19338(.A(dpath_mulcore_b1[1]), .B(n12023), .Y(dpath_mulcore_ary1_a0_I0_p1_l[14]));
INVX1 mul_U19339(.A(dpath_mulcore_ary1_a0_I0_p1_l[14]), .Y(n6643));
AND2X1 mul_U19340(.A(dpath_mulcore_b0[1]), .B(n12026), .Y(dpath_mulcore_ary1_a0_I0_p0_l[14]));
INVX1 mul_U19341(.A(dpath_mulcore_ary1_a0_I0_p0_l[14]), .Y(n6644));
AND2X1 mul_U19342(.A(dpath_mulcore_b2[1]), .B(n12029), .Y(dpath_mulcore_ary1_a0_I0_p2_l[13]));
INVX1 mul_U19343(.A(dpath_mulcore_ary1_a0_I0_p2_l[13]), .Y(n6645));
AND2X1 mul_U19344(.A(dpath_mulcore_b1[1]), .B(n12032), .Y(dpath_mulcore_ary1_a0_I0_p1_l[13]));
INVX1 mul_U19345(.A(dpath_mulcore_ary1_a0_I0_p1_l[13]), .Y(n6646));
AND2X1 mul_U19346(.A(dpath_mulcore_b0[1]), .B(n12035), .Y(dpath_mulcore_ary1_a0_I0_p0_l[13]));
INVX1 mul_U19347(.A(dpath_mulcore_ary1_a0_I0_p0_l[13]), .Y(n6647));
AND2X1 mul_U19348(.A(dpath_mulcore_b2[1]), .B(n12038), .Y(dpath_mulcore_ary1_a0_I0_p2_l[12]));
INVX1 mul_U19349(.A(dpath_mulcore_ary1_a0_I0_p2_l[12]), .Y(n6648));
AND2X1 mul_U19350(.A(dpath_mulcore_b1[1]), .B(n12041), .Y(dpath_mulcore_ary1_a0_I0_p1_l[12]));
INVX1 mul_U19351(.A(dpath_mulcore_ary1_a0_I0_p1_l[12]), .Y(n6649));
AND2X1 mul_U19352(.A(dpath_mulcore_b0[1]), .B(n12044), .Y(dpath_mulcore_ary1_a0_I0_p0_l[12]));
INVX1 mul_U19353(.A(dpath_mulcore_ary1_a0_I0_p0_l[12]), .Y(n6650));
AND2X1 mul_U19354(.A(dpath_mulcore_b2[1]), .B(n12047), .Y(dpath_mulcore_ary1_a0_I0_p2_l[11]));
INVX1 mul_U19355(.A(dpath_mulcore_ary1_a0_I0_p2_l[11]), .Y(n6651));
AND2X1 mul_U19356(.A(dpath_mulcore_b1[1]), .B(n12050), .Y(dpath_mulcore_ary1_a0_I0_p1_l[11]));
INVX1 mul_U19357(.A(dpath_mulcore_ary1_a0_I0_p1_l[11]), .Y(n6652));
AND2X1 mul_U19358(.A(dpath_mulcore_b0[1]), .B(n12053), .Y(dpath_mulcore_ary1_a0_I0_p0_l[11]));
INVX1 mul_U19359(.A(dpath_mulcore_ary1_a0_I0_p0_l[11]), .Y(n6653));
AND2X1 mul_U19360(.A(dpath_mulcore_b2[1]), .B(n12056), .Y(dpath_mulcore_ary1_a0_I0_p2_l[10]));
INVX1 mul_U19361(.A(dpath_mulcore_ary1_a0_I0_p2_l[10]), .Y(n6654));
AND2X1 mul_U19362(.A(dpath_mulcore_b1[1]), .B(n12059), .Y(dpath_mulcore_ary1_a0_I0_p1_l[10]));
INVX1 mul_U19363(.A(dpath_mulcore_ary1_a0_I0_p1_l[10]), .Y(n6655));
AND2X1 mul_U19364(.A(dpath_mulcore_b0[1]), .B(n12062), .Y(dpath_mulcore_ary1_a0_I0_p0_l[10]));
INVX1 mul_U19365(.A(dpath_mulcore_ary1_a0_I0_p0_l[10]), .Y(n6656));
AND2X1 mul_U19366(.A(dpath_mulcore_b2[1]), .B(n12065), .Y(dpath_mulcore_ary1_a0_I0_p2_l[9]));
INVX1 mul_U19367(.A(dpath_mulcore_ary1_a0_I0_p2_l[9]), .Y(n6657));
AND2X1 mul_U19368(.A(dpath_mulcore_b1[1]), .B(n12068), .Y(dpath_mulcore_ary1_a0_I0_p1_l[9]));
INVX1 mul_U19369(.A(dpath_mulcore_ary1_a0_I0_p1_l[9]), .Y(n6658));
AND2X1 mul_U19370(.A(dpath_mulcore_b0[1]), .B(n12071), .Y(dpath_mulcore_ary1_a0_I0_p0_l[9]));
INVX1 mul_U19371(.A(dpath_mulcore_ary1_a0_I0_p0_l[9]), .Y(n6659));
AND2X1 mul_U19372(.A(dpath_mulcore_b2[1]), .B(n12074), .Y(dpath_mulcore_ary1_a0_I0_p2_l[8]));
INVX1 mul_U19373(.A(dpath_mulcore_ary1_a0_I0_p2_l[8]), .Y(n6660));
AND2X1 mul_U19374(.A(dpath_mulcore_b1[1]), .B(n12077), .Y(dpath_mulcore_ary1_a0_I0_p1_l[8]));
INVX1 mul_U19375(.A(dpath_mulcore_ary1_a0_I0_p1_l[8]), .Y(n6661));
AND2X1 mul_U19376(.A(dpath_mulcore_b0[1]), .B(n12080), .Y(dpath_mulcore_ary1_a0_I0_p0_l[8]));
INVX1 mul_U19377(.A(dpath_mulcore_ary1_a0_I0_p0_l[8]), .Y(n6662));
AND2X1 mul_U19378(.A(dpath_mulcore_b2[1]), .B(n12083), .Y(dpath_mulcore_ary1_a0_I0_p2_l[7]));
INVX1 mul_U19379(.A(dpath_mulcore_ary1_a0_I0_p2_l[7]), .Y(n6663));
AND2X1 mul_U19380(.A(dpath_mulcore_b1[1]), .B(n12086), .Y(dpath_mulcore_ary1_a0_I0_p1_l[7]));
INVX1 mul_U19381(.A(dpath_mulcore_ary1_a0_I0_p1_l[7]), .Y(n6664));
AND2X1 mul_U19382(.A(dpath_mulcore_b0[1]), .B(n12089), .Y(dpath_mulcore_ary1_a0_I0_p0_l[7]));
INVX1 mul_U19383(.A(dpath_mulcore_ary1_a0_I0_p0_l[7]), .Y(n6665));
AND2X1 mul_U19384(.A(dpath_mulcore_b2[1]), .B(n12092), .Y(dpath_mulcore_ary1_a0_I0_p2_l[6]));
INVX1 mul_U19385(.A(dpath_mulcore_ary1_a0_I0_p2_l[6]), .Y(n6666));
AND2X1 mul_U19386(.A(dpath_mulcore_b1[1]), .B(n12095), .Y(dpath_mulcore_ary1_a0_I0_p1_l[6]));
INVX1 mul_U19387(.A(dpath_mulcore_ary1_a0_I0_p1_l[6]), .Y(n6667));
AND2X1 mul_U19388(.A(dpath_mulcore_b0[1]), .B(n12098), .Y(dpath_mulcore_ary1_a0_I0_p0_l[6]));
INVX1 mul_U19389(.A(dpath_mulcore_ary1_a0_I0_p0_l[6]), .Y(n6668));
AND2X1 mul_U19390(.A(dpath_mulcore_b2[1]), .B(n12101), .Y(dpath_mulcore_ary1_a0_I0_p2_l[5]));
INVX1 mul_U19391(.A(dpath_mulcore_ary1_a0_I0_p2_l[5]), .Y(n6669));
AND2X1 mul_U19392(.A(dpath_mulcore_b1[1]), .B(n12104), .Y(dpath_mulcore_ary1_a0_I0_p1_l[5]));
INVX1 mul_U19393(.A(dpath_mulcore_ary1_a0_I0_p1_l[5]), .Y(n6670));
AND2X1 mul_U19394(.A(dpath_mulcore_b0[1]), .B(n12107), .Y(dpath_mulcore_ary1_a0_I0_p0_l[5]));
INVX1 mul_U19395(.A(dpath_mulcore_ary1_a0_I0_p0_l[5]), .Y(n6671));
AND2X1 mul_U19396(.A(dpath_mulcore_b2[1]), .B(n12109), .Y(dpath_mulcore_ary1_a0_I0_p2_l[4]));
INVX1 mul_U19397(.A(dpath_mulcore_ary1_a0_I0_p2_l[4]), .Y(n6672));
AND2X1 mul_U19398(.A(dpath_mulcore_b1[1]), .B(n12112), .Y(dpath_mulcore_ary1_a0_I0_p1_l[4]));
INVX1 mul_U19399(.A(dpath_mulcore_ary1_a0_I0_p1_l[4]), .Y(n6673));
AND2X1 mul_U19400(.A(dpath_mulcore_b0[1]), .B(n12115), .Y(dpath_mulcore_ary1_a0_I0_p0_l[4]));
INVX1 mul_U19401(.A(dpath_mulcore_ary1_a0_I0_p0_l[4]), .Y(n6674));
AND2X1 mul_U19402(.A(dpath_mulcore_b0[1]), .B(n12118), .Y(dpath_mulcore_ary1_a0_I0_p0_l[3]));
INVX1 mul_U19403(.A(dpath_mulcore_ary1_a0_I0_p0_l[3]), .Y(n6675));
AND2X1 mul_U19404(.A(dpath_mulcore_b1[1]), .B(n12121), .Y(dpath_mulcore_ary1_a0_I0_p1_l[3]));
INVX1 mul_U19405(.A(dpath_mulcore_ary1_a0_I0_p1_l[3]), .Y(n6676));
AND2X1 mul_U19406(.A(dpath_mulcore_b0[1]), .B(n12124), .Y(dpath_mulcore_ary1_a0_I0_I0_p0_l_2));
INVX1 mul_U19407(.A(dpath_mulcore_ary1_a0_I0_I0_p0_l_2), .Y(n6677));
AND2X1 mul_U19408(.A(dpath_mulcore_b0[1]), .B(n12127), .Y(dpath_mulcore_ary1_a0_I0_I0_p0_l_1));
INVX1 mul_U19409(.A(dpath_mulcore_ary1_a0_I0_I0_p0_l_1), .Y(n6678));
AND2X1 mul_U19410(.A(dpath_mulcore_b0[1]), .B(n12129), .Y(dpath_mulcore_ary1_a0_I0_I0_p0_l_0));
INVX1 mul_U19411(.A(dpath_mulcore_ary1_a0_I0_I0_p0_l_0), .Y(n6679));
AND2X1 mul_U19412(.A(dpath_mulcore_b1[1]), .B(n12131), .Y(dpath_mulcore_ary1_a0_I0_I0_p1_l_2));
INVX1 mul_U19413(.A(dpath_mulcore_ary1_a0_I0_I0_p1_l_2), .Y(n6680));
AND2X1 mul_U19414(.A(dpath_mulcore_b15[1]), .B(n12134), .Y(dpath_mulcore_ary1_a1_I2_I2_p1_l_65));
INVX1 mul_U19415(.A(dpath_mulcore_ary1_a1_I2_I2_p1_l_65), .Y(n6681));
AND2X1 mul_U19416(.A(dpath_mulcore_b15[1]), .B(n12137), .Y(dpath_mulcore_ary1_a1_I2_I2_p1_l_64));
INVX1 mul_U19417(.A(dpath_mulcore_ary1_a1_I2_I2_p1_l_64), .Y(n6682));
AND2X1 mul_U19418(.A(dpath_mulcore_b15[1]), .B(n12140), .Y(dpath_mulcore_ary1_a1_I2_p1_l[63]));
INVX1 mul_U19419(.A(dpath_mulcore_ary1_a1_I2_p1_l[63]), .Y(n6683));
AND2X1 mul_U19420(.A(dpath_mulcore_b14[1]), .B(n12143), .Y(dpath_mulcore_ary1_a1_I2_p0_l[63]));
INVX1 mul_U19421(.A(dpath_mulcore_ary1_a1_I2_p0_l[63]), .Y(n6684));
AND2X1 mul_U19422(.A(dpath_mulcore_b15[1]), .B(n12146), .Y(dpath_mulcore_ary1_a1_I2_p1_l[62]));
INVX1 mul_U19423(.A(dpath_mulcore_ary1_a1_I2_p1_l[62]), .Y(n6685));
AND2X1 mul_U19424(.A(dpath_mulcore_b14[1]), .B(n12149), .Y(dpath_mulcore_ary1_a1_I2_p0_l[62]));
INVX1 mul_U19425(.A(dpath_mulcore_ary1_a1_I2_p0_l[62]), .Y(n6686));
AND2X1 mul_U19426(.A(dpath_mulcore_b15[1]), .B(n12152), .Y(dpath_mulcore_ary1_a1_I2_p1_l[61]));
INVX1 mul_U19427(.A(dpath_mulcore_ary1_a1_I2_p1_l[61]), .Y(n6687));
AND2X1 mul_U19428(.A(dpath_mulcore_b14[1]), .B(n12155), .Y(dpath_mulcore_ary1_a1_I2_p0_l[61]));
INVX1 mul_U19429(.A(dpath_mulcore_ary1_a1_I2_p0_l[61]), .Y(n6688));
AND2X1 mul_U19430(.A(dpath_mulcore_b15[1]), .B(n12158), .Y(dpath_mulcore_ary1_a1_I2_p1_l[60]));
INVX1 mul_U19431(.A(dpath_mulcore_ary1_a1_I2_p1_l[60]), .Y(n6689));
AND2X1 mul_U19432(.A(dpath_mulcore_b14[1]), .B(n12161), .Y(dpath_mulcore_ary1_a1_I2_p0_l[60]));
INVX1 mul_U19433(.A(dpath_mulcore_ary1_a1_I2_p0_l[60]), .Y(n6690));
AND2X1 mul_U19434(.A(dpath_mulcore_b15[1]), .B(n12164), .Y(dpath_mulcore_ary1_a1_I2_p1_l[59]));
INVX1 mul_U19435(.A(dpath_mulcore_ary1_a1_I2_p1_l[59]), .Y(n6691));
AND2X1 mul_U19436(.A(dpath_mulcore_b14[1]), .B(n12167), .Y(dpath_mulcore_ary1_a1_I2_p0_l[59]));
INVX1 mul_U19437(.A(dpath_mulcore_ary1_a1_I2_p0_l[59]), .Y(n6692));
AND2X1 mul_U19438(.A(dpath_mulcore_b15[1]), .B(n12170), .Y(dpath_mulcore_ary1_a1_I2_p1_l[58]));
INVX1 mul_U19439(.A(dpath_mulcore_ary1_a1_I2_p1_l[58]), .Y(n6693));
AND2X1 mul_U19440(.A(dpath_mulcore_b14[1]), .B(n12173), .Y(dpath_mulcore_ary1_a1_I2_p0_l[58]));
INVX1 mul_U19441(.A(dpath_mulcore_ary1_a1_I2_p0_l[58]), .Y(n6694));
AND2X1 mul_U19442(.A(dpath_mulcore_b15[1]), .B(n12176), .Y(dpath_mulcore_ary1_a1_I2_p1_l[57]));
INVX1 mul_U19443(.A(dpath_mulcore_ary1_a1_I2_p1_l[57]), .Y(n6695));
AND2X1 mul_U19444(.A(dpath_mulcore_b14[1]), .B(n12179), .Y(dpath_mulcore_ary1_a1_I2_p0_l[57]));
INVX1 mul_U19445(.A(dpath_mulcore_ary1_a1_I2_p0_l[57]), .Y(n6696));
AND2X1 mul_U19446(.A(dpath_mulcore_b15[1]), .B(n12182), .Y(dpath_mulcore_ary1_a1_I2_p1_l[56]));
INVX1 mul_U19447(.A(dpath_mulcore_ary1_a1_I2_p1_l[56]), .Y(n6697));
AND2X1 mul_U19448(.A(dpath_mulcore_b14[1]), .B(n12185), .Y(dpath_mulcore_ary1_a1_I2_p0_l[56]));
INVX1 mul_U19449(.A(dpath_mulcore_ary1_a1_I2_p0_l[56]), .Y(n6698));
AND2X1 mul_U19450(.A(dpath_mulcore_b15[1]), .B(n12188), .Y(dpath_mulcore_ary1_a1_I2_p1_l[55]));
INVX1 mul_U19451(.A(dpath_mulcore_ary1_a1_I2_p1_l[55]), .Y(n6699));
AND2X1 mul_U19452(.A(dpath_mulcore_b14[1]), .B(n12191), .Y(dpath_mulcore_ary1_a1_I2_p0_l[55]));
INVX1 mul_U19453(.A(dpath_mulcore_ary1_a1_I2_p0_l[55]), .Y(n6700));
AND2X1 mul_U19454(.A(dpath_mulcore_b15[1]), .B(n12194), .Y(dpath_mulcore_ary1_a1_I2_p1_l[54]));
INVX1 mul_U19455(.A(dpath_mulcore_ary1_a1_I2_p1_l[54]), .Y(n6701));
AND2X1 mul_U19456(.A(dpath_mulcore_b14[1]), .B(n12197), .Y(dpath_mulcore_ary1_a1_I2_p0_l[54]));
INVX1 mul_U19457(.A(dpath_mulcore_ary1_a1_I2_p0_l[54]), .Y(n6702));
AND2X1 mul_U19458(.A(dpath_mulcore_b15[1]), .B(n12200), .Y(dpath_mulcore_ary1_a1_I2_p1_l[53]));
INVX1 mul_U19459(.A(dpath_mulcore_ary1_a1_I2_p1_l[53]), .Y(n6703));
AND2X1 mul_U19460(.A(dpath_mulcore_b14[1]), .B(n12203), .Y(dpath_mulcore_ary1_a1_I2_p0_l[53]));
INVX1 mul_U19461(.A(dpath_mulcore_ary1_a1_I2_p0_l[53]), .Y(n6704));
AND2X1 mul_U19462(.A(dpath_mulcore_b15[1]), .B(n12206), .Y(dpath_mulcore_ary1_a1_I2_p1_l[52]));
INVX1 mul_U19463(.A(dpath_mulcore_ary1_a1_I2_p1_l[52]), .Y(n6705));
AND2X1 mul_U19464(.A(dpath_mulcore_b14[1]), .B(n12209), .Y(dpath_mulcore_ary1_a1_I2_p0_l[52]));
INVX1 mul_U19465(.A(dpath_mulcore_ary1_a1_I2_p0_l[52]), .Y(n6706));
AND2X1 mul_U19466(.A(dpath_mulcore_b15[1]), .B(n12212), .Y(dpath_mulcore_ary1_a1_I2_p1_l[51]));
INVX1 mul_U19467(.A(dpath_mulcore_ary1_a1_I2_p1_l[51]), .Y(n6707));
AND2X1 mul_U19468(.A(dpath_mulcore_b14[1]), .B(n12215), .Y(dpath_mulcore_ary1_a1_I2_p0_l[51]));
INVX1 mul_U19469(.A(dpath_mulcore_ary1_a1_I2_p0_l[51]), .Y(n6708));
AND2X1 mul_U19470(.A(dpath_mulcore_b15[1]), .B(n12218), .Y(dpath_mulcore_ary1_a1_I2_p1_l[50]));
INVX1 mul_U19471(.A(dpath_mulcore_ary1_a1_I2_p1_l[50]), .Y(n6709));
AND2X1 mul_U19472(.A(dpath_mulcore_b14[1]), .B(n12221), .Y(dpath_mulcore_ary1_a1_I2_p0_l[50]));
INVX1 mul_U19473(.A(dpath_mulcore_ary1_a1_I2_p0_l[50]), .Y(n6710));
AND2X1 mul_U19474(.A(dpath_mulcore_b15[1]), .B(n12224), .Y(dpath_mulcore_ary1_a1_I2_p1_l[49]));
INVX1 mul_U19475(.A(dpath_mulcore_ary1_a1_I2_p1_l[49]), .Y(n6711));
AND2X1 mul_U19476(.A(dpath_mulcore_b14[1]), .B(n12227), .Y(dpath_mulcore_ary1_a1_I2_p0_l[49]));
INVX1 mul_U19477(.A(dpath_mulcore_ary1_a1_I2_p0_l[49]), .Y(n6712));
AND2X1 mul_U19478(.A(dpath_mulcore_b15[1]), .B(n12230), .Y(dpath_mulcore_ary1_a1_I2_p1_l[48]));
INVX1 mul_U19479(.A(dpath_mulcore_ary1_a1_I2_p1_l[48]), .Y(n6713));
AND2X1 mul_U19480(.A(dpath_mulcore_b14[1]), .B(n12233), .Y(dpath_mulcore_ary1_a1_I2_p0_l[48]));
INVX1 mul_U19481(.A(dpath_mulcore_ary1_a1_I2_p0_l[48]), .Y(n6714));
AND2X1 mul_U19482(.A(dpath_mulcore_b15[1]), .B(n12236), .Y(dpath_mulcore_ary1_a1_I2_p1_l[47]));
INVX1 mul_U19483(.A(dpath_mulcore_ary1_a1_I2_p1_l[47]), .Y(n6715));
AND2X1 mul_U19484(.A(dpath_mulcore_b14[1]), .B(n12239), .Y(dpath_mulcore_ary1_a1_I2_p0_l[47]));
INVX1 mul_U19485(.A(dpath_mulcore_ary1_a1_I2_p0_l[47]), .Y(n6716));
AND2X1 mul_U19486(.A(dpath_mulcore_b15[1]), .B(n12242), .Y(dpath_mulcore_ary1_a1_I2_p1_l[46]));
INVX1 mul_U19487(.A(dpath_mulcore_ary1_a1_I2_p1_l[46]), .Y(n6717));
AND2X1 mul_U19488(.A(dpath_mulcore_b14[1]), .B(n12245), .Y(dpath_mulcore_ary1_a1_I2_p0_l[46]));
INVX1 mul_U19489(.A(dpath_mulcore_ary1_a1_I2_p0_l[46]), .Y(n6718));
AND2X1 mul_U19490(.A(dpath_mulcore_b15[1]), .B(n12248), .Y(dpath_mulcore_ary1_a1_I2_p1_l[45]));
INVX1 mul_U19491(.A(dpath_mulcore_ary1_a1_I2_p1_l[45]), .Y(n6719));
AND2X1 mul_U19492(.A(dpath_mulcore_b14[1]), .B(n12251), .Y(dpath_mulcore_ary1_a1_I2_p0_l[45]));
INVX1 mul_U19493(.A(dpath_mulcore_ary1_a1_I2_p0_l[45]), .Y(n6720));
AND2X1 mul_U19494(.A(dpath_mulcore_b15[1]), .B(n12254), .Y(dpath_mulcore_ary1_a1_I2_p1_l[44]));
INVX1 mul_U19495(.A(dpath_mulcore_ary1_a1_I2_p1_l[44]), .Y(n6721));
AND2X1 mul_U19496(.A(dpath_mulcore_b14[1]), .B(n12257), .Y(dpath_mulcore_ary1_a1_I2_p0_l[44]));
INVX1 mul_U19497(.A(dpath_mulcore_ary1_a1_I2_p0_l[44]), .Y(n6722));
AND2X1 mul_U19498(.A(dpath_mulcore_b15[1]), .B(n12260), .Y(dpath_mulcore_ary1_a1_I2_p1_l[43]));
INVX1 mul_U19499(.A(dpath_mulcore_ary1_a1_I2_p1_l[43]), .Y(n6723));
AND2X1 mul_U19500(.A(dpath_mulcore_b14[1]), .B(n12263), .Y(dpath_mulcore_ary1_a1_I2_p0_l[43]));
INVX1 mul_U19501(.A(dpath_mulcore_ary1_a1_I2_p0_l[43]), .Y(n6724));
AND2X1 mul_U19502(.A(dpath_mulcore_b15[1]), .B(n12266), .Y(dpath_mulcore_ary1_a1_I2_p1_l[42]));
INVX1 mul_U19503(.A(dpath_mulcore_ary1_a1_I2_p1_l[42]), .Y(n6725));
AND2X1 mul_U19504(.A(dpath_mulcore_b14[1]), .B(n12269), .Y(dpath_mulcore_ary1_a1_I2_p0_l[42]));
INVX1 mul_U19505(.A(dpath_mulcore_ary1_a1_I2_p0_l[42]), .Y(n6726));
AND2X1 mul_U19506(.A(dpath_mulcore_b15[1]), .B(n12272), .Y(dpath_mulcore_ary1_a1_I2_p1_l[41]));
INVX1 mul_U19507(.A(dpath_mulcore_ary1_a1_I2_p1_l[41]), .Y(n6727));
AND2X1 mul_U19508(.A(dpath_mulcore_b14[1]), .B(n12275), .Y(dpath_mulcore_ary1_a1_I2_p0_l[41]));
INVX1 mul_U19509(.A(dpath_mulcore_ary1_a1_I2_p0_l[41]), .Y(n6728));
AND2X1 mul_U19510(.A(dpath_mulcore_b15[1]), .B(n12278), .Y(dpath_mulcore_ary1_a1_I2_p1_l[40]));
INVX1 mul_U19511(.A(dpath_mulcore_ary1_a1_I2_p1_l[40]), .Y(n6729));
AND2X1 mul_U19512(.A(dpath_mulcore_b14[1]), .B(n12281), .Y(dpath_mulcore_ary1_a1_I2_p0_l[40]));
INVX1 mul_U19513(.A(dpath_mulcore_ary1_a1_I2_p0_l[40]), .Y(n6730));
AND2X1 mul_U19514(.A(dpath_mulcore_b15[1]), .B(n12284), .Y(dpath_mulcore_ary1_a1_I2_p1_l[39]));
INVX1 mul_U19515(.A(dpath_mulcore_ary1_a1_I2_p1_l[39]), .Y(n6731));
AND2X1 mul_U19516(.A(dpath_mulcore_b14[1]), .B(n12287), .Y(dpath_mulcore_ary1_a1_I2_p0_l[39]));
INVX1 mul_U19517(.A(dpath_mulcore_ary1_a1_I2_p0_l[39]), .Y(n6732));
AND2X1 mul_U19518(.A(dpath_mulcore_b15[1]), .B(n12290), .Y(dpath_mulcore_ary1_a1_I2_p1_l[38]));
INVX1 mul_U19519(.A(dpath_mulcore_ary1_a1_I2_p1_l[38]), .Y(n6733));
AND2X1 mul_U19520(.A(dpath_mulcore_b14[1]), .B(n12293), .Y(dpath_mulcore_ary1_a1_I2_p0_l[38]));
INVX1 mul_U19521(.A(dpath_mulcore_ary1_a1_I2_p0_l[38]), .Y(n6734));
AND2X1 mul_U19522(.A(dpath_mulcore_b15[1]), .B(n12296), .Y(dpath_mulcore_ary1_a1_I2_p1_l[37]));
INVX1 mul_U19523(.A(dpath_mulcore_ary1_a1_I2_p1_l[37]), .Y(n6735));
AND2X1 mul_U19524(.A(dpath_mulcore_b14[1]), .B(n12299), .Y(dpath_mulcore_ary1_a1_I2_p0_l[37]));
INVX1 mul_U19525(.A(dpath_mulcore_ary1_a1_I2_p0_l[37]), .Y(n6736));
AND2X1 mul_U19526(.A(dpath_mulcore_b15[1]), .B(n12302), .Y(dpath_mulcore_ary1_a1_I2_p1_l[36]));
INVX1 mul_U19527(.A(dpath_mulcore_ary1_a1_I2_p1_l[36]), .Y(n6737));
AND2X1 mul_U19528(.A(dpath_mulcore_b14[1]), .B(n12305), .Y(dpath_mulcore_ary1_a1_I2_p0_l[36]));
INVX1 mul_U19529(.A(dpath_mulcore_ary1_a1_I2_p0_l[36]), .Y(n6738));
AND2X1 mul_U19530(.A(dpath_mulcore_b15[1]), .B(n12308), .Y(dpath_mulcore_ary1_a1_I2_p1_l[35]));
INVX1 mul_U19531(.A(dpath_mulcore_ary1_a1_I2_p1_l[35]), .Y(n6739));
AND2X1 mul_U19532(.A(dpath_mulcore_b14[1]), .B(n12311), .Y(dpath_mulcore_ary1_a1_I2_p0_l[35]));
INVX1 mul_U19533(.A(dpath_mulcore_ary1_a1_I2_p0_l[35]), .Y(n6740));
AND2X1 mul_U19534(.A(dpath_mulcore_b15[1]), .B(n12314), .Y(dpath_mulcore_ary1_a1_I2_p1_l[34]));
INVX1 mul_U19535(.A(dpath_mulcore_ary1_a1_I2_p1_l[34]), .Y(n6741));
AND2X1 mul_U19536(.A(dpath_mulcore_b14[1]), .B(n12317), .Y(dpath_mulcore_ary1_a1_I2_p0_l[34]));
INVX1 mul_U19537(.A(dpath_mulcore_ary1_a1_I2_p0_l[34]), .Y(n6742));
AND2X1 mul_U19538(.A(dpath_mulcore_b15[1]), .B(n12320), .Y(dpath_mulcore_ary1_a1_I2_p1_l[33]));
INVX1 mul_U19539(.A(dpath_mulcore_ary1_a1_I2_p1_l[33]), .Y(n6743));
AND2X1 mul_U19540(.A(dpath_mulcore_b14[1]), .B(n12323), .Y(dpath_mulcore_ary1_a1_I2_p0_l[33]));
INVX1 mul_U19541(.A(dpath_mulcore_ary1_a1_I2_p0_l[33]), .Y(n6744));
AND2X1 mul_U19542(.A(dpath_mulcore_b15[1]), .B(n12326), .Y(dpath_mulcore_ary1_a1_I2_p1_l[32]));
INVX1 mul_U19543(.A(dpath_mulcore_ary1_a1_I2_p1_l[32]), .Y(n6745));
AND2X1 mul_U19544(.A(dpath_mulcore_b14[1]), .B(n12329), .Y(dpath_mulcore_ary1_a1_I2_p0_l[32]));
INVX1 mul_U19545(.A(dpath_mulcore_ary1_a1_I2_p0_l[32]), .Y(n6746));
AND2X1 mul_U19546(.A(dpath_mulcore_b15[1]), .B(n12332), .Y(dpath_mulcore_ary1_a1_I2_p1_l[31]));
INVX1 mul_U19547(.A(dpath_mulcore_ary1_a1_I2_p1_l[31]), .Y(n6747));
AND2X1 mul_U19548(.A(dpath_mulcore_b14[1]), .B(n12335), .Y(dpath_mulcore_ary1_a1_I2_p0_l[31]));
INVX1 mul_U19549(.A(dpath_mulcore_ary1_a1_I2_p0_l[31]), .Y(n6748));
AND2X1 mul_U19550(.A(dpath_mulcore_b15[1]), .B(n12338), .Y(dpath_mulcore_ary1_a1_I2_p1_l[30]));
INVX1 mul_U19551(.A(dpath_mulcore_ary1_a1_I2_p1_l[30]), .Y(n6749));
AND2X1 mul_U19552(.A(dpath_mulcore_b14[1]), .B(n12341), .Y(dpath_mulcore_ary1_a1_I2_p0_l[30]));
INVX1 mul_U19553(.A(dpath_mulcore_ary1_a1_I2_p0_l[30]), .Y(n6750));
AND2X1 mul_U19554(.A(dpath_mulcore_b15[1]), .B(n12344), .Y(dpath_mulcore_ary1_a1_I2_p1_l[29]));
INVX1 mul_U19555(.A(dpath_mulcore_ary1_a1_I2_p1_l[29]), .Y(n6751));
AND2X1 mul_U19556(.A(dpath_mulcore_b14[1]), .B(n12347), .Y(dpath_mulcore_ary1_a1_I2_p0_l[29]));
INVX1 mul_U19557(.A(dpath_mulcore_ary1_a1_I2_p0_l[29]), .Y(n6752));
AND2X1 mul_U19558(.A(dpath_mulcore_b15[1]), .B(n12350), .Y(dpath_mulcore_ary1_a1_I2_p1_l[28]));
INVX1 mul_U19559(.A(dpath_mulcore_ary1_a1_I2_p1_l[28]), .Y(n6753));
AND2X1 mul_U19560(.A(dpath_mulcore_b14[1]), .B(n12353), .Y(dpath_mulcore_ary1_a1_I2_p0_l[28]));
INVX1 mul_U19561(.A(dpath_mulcore_ary1_a1_I2_p0_l[28]), .Y(n6754));
AND2X1 mul_U19562(.A(dpath_mulcore_b15[1]), .B(n12356), .Y(dpath_mulcore_ary1_a1_I2_p1_l[27]));
INVX1 mul_U19563(.A(dpath_mulcore_ary1_a1_I2_p1_l[27]), .Y(n6755));
AND2X1 mul_U19564(.A(dpath_mulcore_b14[1]), .B(n12359), .Y(dpath_mulcore_ary1_a1_I2_p0_l[27]));
INVX1 mul_U19565(.A(dpath_mulcore_ary1_a1_I2_p0_l[27]), .Y(n6756));
AND2X1 mul_U19566(.A(dpath_mulcore_b15[1]), .B(n12362), .Y(dpath_mulcore_ary1_a1_I2_p1_l[26]));
INVX1 mul_U19567(.A(dpath_mulcore_ary1_a1_I2_p1_l[26]), .Y(n6757));
AND2X1 mul_U19568(.A(dpath_mulcore_b14[1]), .B(n12365), .Y(dpath_mulcore_ary1_a1_I2_p0_l[26]));
INVX1 mul_U19569(.A(dpath_mulcore_ary1_a1_I2_p0_l[26]), .Y(n6758));
AND2X1 mul_U19570(.A(dpath_mulcore_b15[1]), .B(n12368), .Y(dpath_mulcore_ary1_a1_I2_p1_l[25]));
INVX1 mul_U19571(.A(dpath_mulcore_ary1_a1_I2_p1_l[25]), .Y(n6759));
AND2X1 mul_U19572(.A(dpath_mulcore_b14[1]), .B(n12371), .Y(dpath_mulcore_ary1_a1_I2_p0_l[25]));
INVX1 mul_U19573(.A(dpath_mulcore_ary1_a1_I2_p0_l[25]), .Y(n6760));
AND2X1 mul_U19574(.A(dpath_mulcore_b15[1]), .B(n12374), .Y(dpath_mulcore_ary1_a1_I2_p1_l[24]));
INVX1 mul_U19575(.A(dpath_mulcore_ary1_a1_I2_p1_l[24]), .Y(n6761));
AND2X1 mul_U19576(.A(dpath_mulcore_b14[1]), .B(n12377), .Y(dpath_mulcore_ary1_a1_I2_p0_l[24]));
INVX1 mul_U19577(.A(dpath_mulcore_ary1_a1_I2_p0_l[24]), .Y(n6762));
AND2X1 mul_U19578(.A(dpath_mulcore_b15[1]), .B(n12380), .Y(dpath_mulcore_ary1_a1_I2_p1_l[23]));
INVX1 mul_U19579(.A(dpath_mulcore_ary1_a1_I2_p1_l[23]), .Y(n6763));
AND2X1 mul_U19580(.A(dpath_mulcore_b14[1]), .B(n12383), .Y(dpath_mulcore_ary1_a1_I2_p0_l[23]));
INVX1 mul_U19581(.A(dpath_mulcore_ary1_a1_I2_p0_l[23]), .Y(n6764));
AND2X1 mul_U19582(.A(dpath_mulcore_b15[1]), .B(n12386), .Y(dpath_mulcore_ary1_a1_I2_p1_l[22]));
INVX1 mul_U19583(.A(dpath_mulcore_ary1_a1_I2_p1_l[22]), .Y(n6765));
AND2X1 mul_U19584(.A(dpath_mulcore_b14[1]), .B(n12389), .Y(dpath_mulcore_ary1_a1_I2_p0_l[22]));
INVX1 mul_U19585(.A(dpath_mulcore_ary1_a1_I2_p0_l[22]), .Y(n6766));
AND2X1 mul_U19586(.A(dpath_mulcore_b15[1]), .B(n12392), .Y(dpath_mulcore_ary1_a1_I2_p1_l[21]));
INVX1 mul_U19587(.A(dpath_mulcore_ary1_a1_I2_p1_l[21]), .Y(n6767));
AND2X1 mul_U19588(.A(dpath_mulcore_b14[1]), .B(n12395), .Y(dpath_mulcore_ary1_a1_I2_p0_l[21]));
INVX1 mul_U19589(.A(dpath_mulcore_ary1_a1_I2_p0_l[21]), .Y(n6768));
AND2X1 mul_U19590(.A(dpath_mulcore_b15[1]), .B(n12398), .Y(dpath_mulcore_ary1_a1_I2_p1_l[20]));
INVX1 mul_U19591(.A(dpath_mulcore_ary1_a1_I2_p1_l[20]), .Y(n6769));
AND2X1 mul_U19592(.A(dpath_mulcore_b14[1]), .B(n12401), .Y(dpath_mulcore_ary1_a1_I2_p0_l[20]));
INVX1 mul_U19593(.A(dpath_mulcore_ary1_a1_I2_p0_l[20]), .Y(n6770));
AND2X1 mul_U19594(.A(dpath_mulcore_b15[1]), .B(n12404), .Y(dpath_mulcore_ary1_a1_I2_p1_l[19]));
INVX1 mul_U19595(.A(dpath_mulcore_ary1_a1_I2_p1_l[19]), .Y(n6771));
AND2X1 mul_U19596(.A(dpath_mulcore_b14[1]), .B(n12407), .Y(dpath_mulcore_ary1_a1_I2_p0_l[19]));
INVX1 mul_U19597(.A(dpath_mulcore_ary1_a1_I2_p0_l[19]), .Y(n6772));
AND2X1 mul_U19598(.A(dpath_mulcore_b15[1]), .B(n12410), .Y(dpath_mulcore_ary1_a1_I2_p1_l[18]));
INVX1 mul_U19599(.A(dpath_mulcore_ary1_a1_I2_p1_l[18]), .Y(n6773));
AND2X1 mul_U19600(.A(dpath_mulcore_b14[1]), .B(n12413), .Y(dpath_mulcore_ary1_a1_I2_p0_l[18]));
INVX1 mul_U19601(.A(dpath_mulcore_ary1_a1_I2_p0_l[18]), .Y(n6774));
AND2X1 mul_U19602(.A(dpath_mulcore_b15[1]), .B(n12416), .Y(dpath_mulcore_ary1_a1_I2_p1_l[17]));
INVX1 mul_U19603(.A(dpath_mulcore_ary1_a1_I2_p1_l[17]), .Y(n6775));
AND2X1 mul_U19604(.A(dpath_mulcore_b14[1]), .B(n12419), .Y(dpath_mulcore_ary1_a1_I2_p0_l[17]));
INVX1 mul_U19605(.A(dpath_mulcore_ary1_a1_I2_p0_l[17]), .Y(n6776));
AND2X1 mul_U19606(.A(dpath_mulcore_b15[1]), .B(n12422), .Y(dpath_mulcore_ary1_a1_I2_p1_l[16]));
INVX1 mul_U19607(.A(dpath_mulcore_ary1_a1_I2_p1_l[16]), .Y(n6777));
AND2X1 mul_U19608(.A(dpath_mulcore_b14[1]), .B(n12425), .Y(dpath_mulcore_ary1_a1_I2_p0_l[16]));
INVX1 mul_U19609(.A(dpath_mulcore_ary1_a1_I2_p0_l[16]), .Y(n6778));
AND2X1 mul_U19610(.A(dpath_mulcore_b15[1]), .B(n12428), .Y(dpath_mulcore_ary1_a1_I2_p1_l[15]));
INVX1 mul_U19611(.A(dpath_mulcore_ary1_a1_I2_p1_l[15]), .Y(n6779));
AND2X1 mul_U19612(.A(dpath_mulcore_b14[1]), .B(n12431), .Y(dpath_mulcore_ary1_a1_I2_p0_l[15]));
INVX1 mul_U19613(.A(dpath_mulcore_ary1_a1_I2_p0_l[15]), .Y(n6780));
AND2X1 mul_U19614(.A(dpath_mulcore_b15[1]), .B(n12434), .Y(dpath_mulcore_ary1_a1_I2_p1_l[14]));
INVX1 mul_U19615(.A(dpath_mulcore_ary1_a1_I2_p1_l[14]), .Y(n6781));
AND2X1 mul_U19616(.A(dpath_mulcore_b14[1]), .B(n12437), .Y(dpath_mulcore_ary1_a1_I2_p0_l[14]));
INVX1 mul_U19617(.A(dpath_mulcore_ary1_a1_I2_p0_l[14]), .Y(n6782));
AND2X1 mul_U19618(.A(dpath_mulcore_b15[1]), .B(n12440), .Y(dpath_mulcore_ary1_a1_I2_p1_l[13]));
INVX1 mul_U19619(.A(dpath_mulcore_ary1_a1_I2_p1_l[13]), .Y(n6783));
AND2X1 mul_U19620(.A(dpath_mulcore_b14[1]), .B(n12443), .Y(dpath_mulcore_ary1_a1_I2_p0_l[13]));
INVX1 mul_U19621(.A(dpath_mulcore_ary1_a1_I2_p0_l[13]), .Y(n6784));
AND2X1 mul_U19622(.A(dpath_mulcore_b15[1]), .B(n12446), .Y(dpath_mulcore_ary1_a1_I2_p1_l[12]));
INVX1 mul_U19623(.A(dpath_mulcore_ary1_a1_I2_p1_l[12]), .Y(n6785));
AND2X1 mul_U19624(.A(dpath_mulcore_b14[1]), .B(n12449), .Y(dpath_mulcore_ary1_a1_I2_p0_l[12]));
INVX1 mul_U19625(.A(dpath_mulcore_ary1_a1_I2_p0_l[12]), .Y(n6786));
AND2X1 mul_U19626(.A(dpath_mulcore_b15[1]), .B(n12452), .Y(dpath_mulcore_ary1_a1_I2_p1_l[11]));
INVX1 mul_U19627(.A(dpath_mulcore_ary1_a1_I2_p1_l[11]), .Y(n6787));
AND2X1 mul_U19628(.A(dpath_mulcore_b14[1]), .B(n12455), .Y(dpath_mulcore_ary1_a1_I2_p0_l[11]));
INVX1 mul_U19629(.A(dpath_mulcore_ary1_a1_I2_p0_l[11]), .Y(n6788));
AND2X1 mul_U19630(.A(dpath_mulcore_b15[1]), .B(n12458), .Y(dpath_mulcore_ary1_a1_I2_p1_l[10]));
INVX1 mul_U19631(.A(dpath_mulcore_ary1_a1_I2_p1_l[10]), .Y(n6789));
AND2X1 mul_U19632(.A(dpath_mulcore_b14[1]), .B(n12461), .Y(dpath_mulcore_ary1_a1_I2_p0_l[10]));
INVX1 mul_U19633(.A(dpath_mulcore_ary1_a1_I2_p0_l[10]), .Y(n6790));
AND2X1 mul_U19634(.A(dpath_mulcore_b15[1]), .B(n12464), .Y(dpath_mulcore_ary1_a1_I2_p1_l[9]));
INVX1 mul_U19635(.A(dpath_mulcore_ary1_a1_I2_p1_l[9]), .Y(n6791));
AND2X1 mul_U19636(.A(dpath_mulcore_b14[1]), .B(n12467), .Y(dpath_mulcore_ary1_a1_I2_p0_l[9]));
INVX1 mul_U19637(.A(dpath_mulcore_ary1_a1_I2_p0_l[9]), .Y(n6792));
AND2X1 mul_U19638(.A(dpath_mulcore_b15[1]), .B(n12470), .Y(dpath_mulcore_ary1_a1_I2_p1_l[8]));
INVX1 mul_U19639(.A(dpath_mulcore_ary1_a1_I2_p1_l[8]), .Y(n6793));
AND2X1 mul_U19640(.A(dpath_mulcore_b14[1]), .B(n12473), .Y(dpath_mulcore_ary1_a1_I2_p0_l[8]));
INVX1 mul_U19641(.A(dpath_mulcore_ary1_a1_I2_p0_l[8]), .Y(n6794));
AND2X1 mul_U19642(.A(dpath_mulcore_b15[1]), .B(n12476), .Y(dpath_mulcore_ary1_a1_I2_p1_l[7]));
INVX1 mul_U19643(.A(dpath_mulcore_ary1_a1_I2_p1_l[7]), .Y(n6795));
AND2X1 mul_U19644(.A(dpath_mulcore_b14[1]), .B(n12479), .Y(dpath_mulcore_ary1_a1_I2_p0_l[7]));
INVX1 mul_U19645(.A(dpath_mulcore_ary1_a1_I2_p0_l[7]), .Y(n6796));
AND2X1 mul_U19646(.A(dpath_mulcore_b15[1]), .B(n12482), .Y(dpath_mulcore_ary1_a1_I2_p1_l[6]));
INVX1 mul_U19647(.A(dpath_mulcore_ary1_a1_I2_p1_l[6]), .Y(n6797));
AND2X1 mul_U19648(.A(dpath_mulcore_b14[1]), .B(n12485), .Y(dpath_mulcore_ary1_a1_I2_p0_l[6]));
INVX1 mul_U19649(.A(dpath_mulcore_ary1_a1_I2_p0_l[6]), .Y(n6798));
AND2X1 mul_U19650(.A(dpath_mulcore_b15[1]), .B(n12488), .Y(dpath_mulcore_ary1_a1_I2_p1_l[5]));
INVX1 mul_U19651(.A(dpath_mulcore_ary1_a1_I2_p1_l[5]), .Y(n6799));
AND2X1 mul_U19652(.A(dpath_mulcore_b14[1]), .B(n12491), .Y(dpath_mulcore_ary1_a1_I2_p0_l[5]));
INVX1 mul_U19653(.A(dpath_mulcore_ary1_a1_I2_p0_l[5]), .Y(n6800));
AND2X1 mul_U19654(.A(dpath_mulcore_b15[1]), .B(n12494), .Y(dpath_mulcore_ary1_a1_I2_p1_l[4]));
INVX1 mul_U19655(.A(dpath_mulcore_ary1_a1_I2_p1_l[4]), .Y(n6801));
AND2X1 mul_U19656(.A(dpath_mulcore_b14[1]), .B(n12497), .Y(dpath_mulcore_ary1_a1_I2_p0_l[4]));
INVX1 mul_U19657(.A(dpath_mulcore_ary1_a1_I2_p0_l[4]), .Y(n6802));
AND2X1 mul_U19658(.A(dpath_mulcore_b14[1]), .B(n12500), .Y(dpath_mulcore_ary1_a1_I2_p0_l[3]));
INVX1 mul_U19659(.A(dpath_mulcore_ary1_a1_I2_p0_l[3]), .Y(n6803));
AND2X1 mul_U19660(.A(dpath_mulcore_b15[1]), .B(n12503), .Y(dpath_mulcore_ary1_a1_I2_p1_l[3]));
INVX1 mul_U19661(.A(dpath_mulcore_ary1_a1_I2_p1_l[3]), .Y(n6804));
AND2X1 mul_U19662(.A(dpath_mulcore_b14[1]), .B(n12506), .Y(dpath_mulcore_ary1_a1_I2_I0_p0_l_2));
INVX1 mul_U19663(.A(dpath_mulcore_ary1_a1_I2_I0_p0_l_2), .Y(n6805));
AND2X1 mul_U19664(.A(dpath_mulcore_b14[1]), .B(n12509), .Y(dpath_mulcore_ary1_a1_I2_I0_p0_l_1));
INVX1 mul_U19665(.A(dpath_mulcore_ary1_a1_I2_I0_p0_l_1), .Y(n6806));
AND2X1 mul_U19666(.A(dpath_mulcore_b14[1]), .B(n12511), .Y(dpath_mulcore_ary1_a1_I2_I0_p0_l_0));
INVX1 mul_U19667(.A(dpath_mulcore_ary1_a1_I2_I0_p0_l_0), .Y(n6807));
AND2X1 mul_U19668(.A(dpath_mulcore_b15[1]), .B(n12513), .Y(dpath_mulcore_ary1_a1_I2_I0_p1_l_2));
INVX1 mul_U19669(.A(dpath_mulcore_ary1_a1_I2_I0_p1_l_2), .Y(n6808));
AND2X1 mul_U19670(.A(dpath_mulcore_b13[1]), .B(n12516), .Y(dpath_mulcore_ary1_a1_I1_I2_p2_l_67));
INVX1 mul_U19671(.A(dpath_mulcore_ary1_a1_I1_I2_p2_l_67), .Y(n6809));
AND2X1 mul_U19672(.A(dpath_mulcore_b13[1]), .B(n12519), .Y(dpath_mulcore_ary1_a1_I1_I2_p2_l_66));
INVX1 mul_U19673(.A(dpath_mulcore_ary1_a1_I1_I2_p2_l_66), .Y(n6810));
AND2X1 mul_U19674(.A(dpath_mulcore_b13[1]), .B(n12522), .Y(dpath_mulcore_ary1_a1_I1_I2_p2_l_65));
INVX1 mul_U19675(.A(dpath_mulcore_ary1_a1_I1_I2_p2_l_65), .Y(n6811));
AND2X1 mul_U19676(.A(dpath_mulcore_b12[1]), .B(n12525), .Y(dpath_mulcore_ary1_a1_I1_I2_p1_l_65));
INVX1 mul_U19677(.A(dpath_mulcore_ary1_a1_I1_I2_p1_l_65), .Y(n6812));
AND2X1 mul_U19678(.A(dpath_mulcore_b12[1]), .B(n12528), .Y(dpath_mulcore_ary1_a1_I1_I2_p1_l_64));
INVX1 mul_U19679(.A(dpath_mulcore_ary1_a1_I1_I2_p1_l_64), .Y(n6813));
AND2X1 mul_U19680(.A(dpath_mulcore_b13[1]), .B(n12531), .Y(dpath_mulcore_ary1_a1_I1_I2_p2_l_64));
INVX1 mul_U19681(.A(dpath_mulcore_ary1_a1_I1_I2_p2_l_64), .Y(n6814));
AND2X1 mul_U19682(.A(dpath_mulcore_b13[1]), .B(n12534), .Y(dpath_mulcore_ary1_a1_I1_p2_l[63]));
INVX1 mul_U19683(.A(dpath_mulcore_ary1_a1_I1_p2_l[63]), .Y(n6815));
AND2X1 mul_U19684(.A(dpath_mulcore_b12[1]), .B(n12537), .Y(dpath_mulcore_ary1_a1_I1_p1_l[63]));
INVX1 mul_U19685(.A(dpath_mulcore_ary1_a1_I1_p1_l[63]), .Y(n6816));
AND2X1 mul_U19686(.A(dpath_mulcore_b11[1]), .B(n12540), .Y(dpath_mulcore_ary1_a1_I1_p0_l[63]));
INVX1 mul_U19687(.A(dpath_mulcore_ary1_a1_I1_p0_l[63]), .Y(n6817));
AND2X1 mul_U19688(.A(dpath_mulcore_b13[1]), .B(n12543), .Y(dpath_mulcore_ary1_a1_I1_p2_l[62]));
INVX1 mul_U19689(.A(dpath_mulcore_ary1_a1_I1_p2_l[62]), .Y(n6818));
AND2X1 mul_U19690(.A(dpath_mulcore_b12[1]), .B(n12546), .Y(dpath_mulcore_ary1_a1_I1_p1_l[62]));
INVX1 mul_U19691(.A(dpath_mulcore_ary1_a1_I1_p1_l[62]), .Y(n6819));
AND2X1 mul_U19692(.A(dpath_mulcore_b11[1]), .B(n12549), .Y(dpath_mulcore_ary1_a1_I1_p0_l[62]));
INVX1 mul_U19693(.A(dpath_mulcore_ary1_a1_I1_p0_l[62]), .Y(n6820));
AND2X1 mul_U19694(.A(dpath_mulcore_b13[1]), .B(n12552), .Y(dpath_mulcore_ary1_a1_I1_p2_l[61]));
INVX1 mul_U19695(.A(dpath_mulcore_ary1_a1_I1_p2_l[61]), .Y(n6821));
AND2X1 mul_U19696(.A(dpath_mulcore_b12[1]), .B(n12555), .Y(dpath_mulcore_ary1_a1_I1_p1_l[61]));
INVX1 mul_U19697(.A(dpath_mulcore_ary1_a1_I1_p1_l[61]), .Y(n6822));
AND2X1 mul_U19698(.A(dpath_mulcore_b11[1]), .B(n12558), .Y(dpath_mulcore_ary1_a1_I1_p0_l[61]));
INVX1 mul_U19699(.A(dpath_mulcore_ary1_a1_I1_p0_l[61]), .Y(n6823));
AND2X1 mul_U19700(.A(dpath_mulcore_b13[1]), .B(n12561), .Y(dpath_mulcore_ary1_a1_I1_p2_l[60]));
INVX1 mul_U19701(.A(dpath_mulcore_ary1_a1_I1_p2_l[60]), .Y(n6824));
AND2X1 mul_U19702(.A(dpath_mulcore_b12[1]), .B(n12564), .Y(dpath_mulcore_ary1_a1_I1_p1_l[60]));
INVX1 mul_U19703(.A(dpath_mulcore_ary1_a1_I1_p1_l[60]), .Y(n6825));
AND2X1 mul_U19704(.A(dpath_mulcore_b11[1]), .B(n12567), .Y(dpath_mulcore_ary1_a1_I1_p0_l[60]));
INVX1 mul_U19705(.A(dpath_mulcore_ary1_a1_I1_p0_l[60]), .Y(n6826));
AND2X1 mul_U19706(.A(dpath_mulcore_b13[1]), .B(n12570), .Y(dpath_mulcore_ary1_a1_I1_p2_l[59]));
INVX1 mul_U19707(.A(dpath_mulcore_ary1_a1_I1_p2_l[59]), .Y(n6827));
AND2X1 mul_U19708(.A(dpath_mulcore_b12[1]), .B(n12573), .Y(dpath_mulcore_ary1_a1_I1_p1_l[59]));
INVX1 mul_U19709(.A(dpath_mulcore_ary1_a1_I1_p1_l[59]), .Y(n6828));
AND2X1 mul_U19710(.A(dpath_mulcore_b11[1]), .B(n12576), .Y(dpath_mulcore_ary1_a1_I1_p0_l[59]));
INVX1 mul_U19711(.A(dpath_mulcore_ary1_a1_I1_p0_l[59]), .Y(n6829));
AND2X1 mul_U19712(.A(dpath_mulcore_b13[1]), .B(n12579), .Y(dpath_mulcore_ary1_a1_I1_p2_l[58]));
INVX1 mul_U19713(.A(dpath_mulcore_ary1_a1_I1_p2_l[58]), .Y(n6830));
AND2X1 mul_U19714(.A(dpath_mulcore_b12[1]), .B(n12582), .Y(dpath_mulcore_ary1_a1_I1_p1_l[58]));
INVX1 mul_U19715(.A(dpath_mulcore_ary1_a1_I1_p1_l[58]), .Y(n6831));
AND2X1 mul_U19716(.A(dpath_mulcore_b11[1]), .B(n12585), .Y(dpath_mulcore_ary1_a1_I1_p0_l[58]));
INVX1 mul_U19717(.A(dpath_mulcore_ary1_a1_I1_p0_l[58]), .Y(n6832));
AND2X1 mul_U19718(.A(dpath_mulcore_b13[1]), .B(n12588), .Y(dpath_mulcore_ary1_a1_I1_p2_l[57]));
INVX1 mul_U19719(.A(dpath_mulcore_ary1_a1_I1_p2_l[57]), .Y(n6833));
AND2X1 mul_U19720(.A(dpath_mulcore_b12[1]), .B(n12591), .Y(dpath_mulcore_ary1_a1_I1_p1_l[57]));
INVX1 mul_U19721(.A(dpath_mulcore_ary1_a1_I1_p1_l[57]), .Y(n6834));
AND2X1 mul_U19722(.A(dpath_mulcore_b11[1]), .B(n12594), .Y(dpath_mulcore_ary1_a1_I1_p0_l[57]));
INVX1 mul_U19723(.A(dpath_mulcore_ary1_a1_I1_p0_l[57]), .Y(n6835));
AND2X1 mul_U19724(.A(dpath_mulcore_b13[1]), .B(n12597), .Y(dpath_mulcore_ary1_a1_I1_p2_l[56]));
INVX1 mul_U19725(.A(dpath_mulcore_ary1_a1_I1_p2_l[56]), .Y(n6836));
AND2X1 mul_U19726(.A(dpath_mulcore_b12[1]), .B(n12600), .Y(dpath_mulcore_ary1_a1_I1_p1_l[56]));
INVX1 mul_U19727(.A(dpath_mulcore_ary1_a1_I1_p1_l[56]), .Y(n6837));
AND2X1 mul_U19728(.A(dpath_mulcore_b11[1]), .B(n12603), .Y(dpath_mulcore_ary1_a1_I1_p0_l[56]));
INVX1 mul_U19729(.A(dpath_mulcore_ary1_a1_I1_p0_l[56]), .Y(n6838));
AND2X1 mul_U19730(.A(dpath_mulcore_b13[1]), .B(n12606), .Y(dpath_mulcore_ary1_a1_I1_p2_l[55]));
INVX1 mul_U19731(.A(dpath_mulcore_ary1_a1_I1_p2_l[55]), .Y(n6839));
AND2X1 mul_U19732(.A(dpath_mulcore_b12[1]), .B(n12609), .Y(dpath_mulcore_ary1_a1_I1_p1_l[55]));
INVX1 mul_U19733(.A(dpath_mulcore_ary1_a1_I1_p1_l[55]), .Y(n6840));
AND2X1 mul_U19734(.A(dpath_mulcore_b11[1]), .B(n12612), .Y(dpath_mulcore_ary1_a1_I1_p0_l[55]));
INVX1 mul_U19735(.A(dpath_mulcore_ary1_a1_I1_p0_l[55]), .Y(n6841));
AND2X1 mul_U19736(.A(dpath_mulcore_b13[1]), .B(n12615), .Y(dpath_mulcore_ary1_a1_I1_p2_l[54]));
INVX1 mul_U19737(.A(dpath_mulcore_ary1_a1_I1_p2_l[54]), .Y(n6842));
AND2X1 mul_U19738(.A(dpath_mulcore_b12[1]), .B(n12618), .Y(dpath_mulcore_ary1_a1_I1_p1_l[54]));
INVX1 mul_U19739(.A(dpath_mulcore_ary1_a1_I1_p1_l[54]), .Y(n6843));
AND2X1 mul_U19740(.A(dpath_mulcore_b11[1]), .B(n12621), .Y(dpath_mulcore_ary1_a1_I1_p0_l[54]));
INVX1 mul_U19741(.A(dpath_mulcore_ary1_a1_I1_p0_l[54]), .Y(n6844));
AND2X1 mul_U19742(.A(dpath_mulcore_b13[1]), .B(n12624), .Y(dpath_mulcore_ary1_a1_I1_p2_l[53]));
INVX1 mul_U19743(.A(dpath_mulcore_ary1_a1_I1_p2_l[53]), .Y(n6845));
AND2X1 mul_U19744(.A(dpath_mulcore_b12[1]), .B(n12627), .Y(dpath_mulcore_ary1_a1_I1_p1_l[53]));
INVX1 mul_U19745(.A(dpath_mulcore_ary1_a1_I1_p1_l[53]), .Y(n6846));
AND2X1 mul_U19746(.A(dpath_mulcore_b11[1]), .B(n12630), .Y(dpath_mulcore_ary1_a1_I1_p0_l[53]));
INVX1 mul_U19747(.A(dpath_mulcore_ary1_a1_I1_p0_l[53]), .Y(n6847));
AND2X1 mul_U19748(.A(dpath_mulcore_b13[1]), .B(n12633), .Y(dpath_mulcore_ary1_a1_I1_p2_l[52]));
INVX1 mul_U19749(.A(dpath_mulcore_ary1_a1_I1_p2_l[52]), .Y(n6848));
AND2X1 mul_U19750(.A(dpath_mulcore_b12[1]), .B(n12636), .Y(dpath_mulcore_ary1_a1_I1_p1_l[52]));
INVX1 mul_U19751(.A(dpath_mulcore_ary1_a1_I1_p1_l[52]), .Y(n6849));
AND2X1 mul_U19752(.A(dpath_mulcore_b11[1]), .B(n12639), .Y(dpath_mulcore_ary1_a1_I1_p0_l[52]));
INVX1 mul_U19753(.A(dpath_mulcore_ary1_a1_I1_p0_l[52]), .Y(n6850));
AND2X1 mul_U19754(.A(dpath_mulcore_b13[1]), .B(n12642), .Y(dpath_mulcore_ary1_a1_I1_p2_l[51]));
INVX1 mul_U19755(.A(dpath_mulcore_ary1_a1_I1_p2_l[51]), .Y(n6851));
AND2X1 mul_U19756(.A(dpath_mulcore_b12[1]), .B(n12645), .Y(dpath_mulcore_ary1_a1_I1_p1_l[51]));
INVX1 mul_U19757(.A(dpath_mulcore_ary1_a1_I1_p1_l[51]), .Y(n6852));
AND2X1 mul_U19758(.A(dpath_mulcore_b11[1]), .B(n12648), .Y(dpath_mulcore_ary1_a1_I1_p0_l[51]));
INVX1 mul_U19759(.A(dpath_mulcore_ary1_a1_I1_p0_l[51]), .Y(n6853));
AND2X1 mul_U19760(.A(dpath_mulcore_b13[1]), .B(n12651), .Y(dpath_mulcore_ary1_a1_I1_p2_l[50]));
INVX1 mul_U19761(.A(dpath_mulcore_ary1_a1_I1_p2_l[50]), .Y(n6854));
AND2X1 mul_U19762(.A(dpath_mulcore_b12[1]), .B(n12654), .Y(dpath_mulcore_ary1_a1_I1_p1_l[50]));
INVX1 mul_U19763(.A(dpath_mulcore_ary1_a1_I1_p1_l[50]), .Y(n6855));
AND2X1 mul_U19764(.A(dpath_mulcore_b11[1]), .B(n12657), .Y(dpath_mulcore_ary1_a1_I1_p0_l[50]));
INVX1 mul_U19765(.A(dpath_mulcore_ary1_a1_I1_p0_l[50]), .Y(n6856));
AND2X1 mul_U19766(.A(dpath_mulcore_b13[1]), .B(n12660), .Y(dpath_mulcore_ary1_a1_I1_p2_l[49]));
INVX1 mul_U19767(.A(dpath_mulcore_ary1_a1_I1_p2_l[49]), .Y(n6857));
AND2X1 mul_U19768(.A(dpath_mulcore_b12[1]), .B(n12663), .Y(dpath_mulcore_ary1_a1_I1_p1_l[49]));
INVX1 mul_U19769(.A(dpath_mulcore_ary1_a1_I1_p1_l[49]), .Y(n6858));
AND2X1 mul_U19770(.A(dpath_mulcore_b11[1]), .B(n12666), .Y(dpath_mulcore_ary1_a1_I1_p0_l[49]));
INVX1 mul_U19771(.A(dpath_mulcore_ary1_a1_I1_p0_l[49]), .Y(n6859));
AND2X1 mul_U19772(.A(dpath_mulcore_b13[1]), .B(n12669), .Y(dpath_mulcore_ary1_a1_I1_p2_l[48]));
INVX1 mul_U19773(.A(dpath_mulcore_ary1_a1_I1_p2_l[48]), .Y(n6860));
AND2X1 mul_U19774(.A(dpath_mulcore_b12[1]), .B(n12672), .Y(dpath_mulcore_ary1_a1_I1_p1_l[48]));
INVX1 mul_U19775(.A(dpath_mulcore_ary1_a1_I1_p1_l[48]), .Y(n6861));
AND2X1 mul_U19776(.A(dpath_mulcore_b11[1]), .B(n12675), .Y(dpath_mulcore_ary1_a1_I1_p0_l[48]));
INVX1 mul_U19777(.A(dpath_mulcore_ary1_a1_I1_p0_l[48]), .Y(n6862));
AND2X1 mul_U19778(.A(dpath_mulcore_b13[1]), .B(n12678), .Y(dpath_mulcore_ary1_a1_I1_p2_l[47]));
INVX1 mul_U19779(.A(dpath_mulcore_ary1_a1_I1_p2_l[47]), .Y(n6863));
AND2X1 mul_U19780(.A(dpath_mulcore_b12[1]), .B(n12681), .Y(dpath_mulcore_ary1_a1_I1_p1_l[47]));
INVX1 mul_U19781(.A(dpath_mulcore_ary1_a1_I1_p1_l[47]), .Y(n6864));
AND2X1 mul_U19782(.A(dpath_mulcore_b11[1]), .B(n12684), .Y(dpath_mulcore_ary1_a1_I1_p0_l[47]));
INVX1 mul_U19783(.A(dpath_mulcore_ary1_a1_I1_p0_l[47]), .Y(n6865));
AND2X1 mul_U19784(.A(dpath_mulcore_b13[1]), .B(n12687), .Y(dpath_mulcore_ary1_a1_I1_p2_l[46]));
INVX1 mul_U19785(.A(dpath_mulcore_ary1_a1_I1_p2_l[46]), .Y(n6866));
AND2X1 mul_U19786(.A(dpath_mulcore_b12[1]), .B(n12690), .Y(dpath_mulcore_ary1_a1_I1_p1_l[46]));
INVX1 mul_U19787(.A(dpath_mulcore_ary1_a1_I1_p1_l[46]), .Y(n6867));
AND2X1 mul_U19788(.A(dpath_mulcore_b11[1]), .B(n12693), .Y(dpath_mulcore_ary1_a1_I1_p0_l[46]));
INVX1 mul_U19789(.A(dpath_mulcore_ary1_a1_I1_p0_l[46]), .Y(n6868));
AND2X1 mul_U19790(.A(dpath_mulcore_b13[1]), .B(n12696), .Y(dpath_mulcore_ary1_a1_I1_p2_l[45]));
INVX1 mul_U19791(.A(dpath_mulcore_ary1_a1_I1_p2_l[45]), .Y(n6869));
AND2X1 mul_U19792(.A(dpath_mulcore_b12[1]), .B(n12699), .Y(dpath_mulcore_ary1_a1_I1_p1_l[45]));
INVX1 mul_U19793(.A(dpath_mulcore_ary1_a1_I1_p1_l[45]), .Y(n6870));
AND2X1 mul_U19794(.A(dpath_mulcore_b11[1]), .B(n12702), .Y(dpath_mulcore_ary1_a1_I1_p0_l[45]));
INVX1 mul_U19795(.A(dpath_mulcore_ary1_a1_I1_p0_l[45]), .Y(n6871));
AND2X1 mul_U19796(.A(dpath_mulcore_b13[1]), .B(n12705), .Y(dpath_mulcore_ary1_a1_I1_p2_l[44]));
INVX1 mul_U19797(.A(dpath_mulcore_ary1_a1_I1_p2_l[44]), .Y(n6872));
AND2X1 mul_U19798(.A(dpath_mulcore_b12[1]), .B(n12708), .Y(dpath_mulcore_ary1_a1_I1_p1_l[44]));
INVX1 mul_U19799(.A(dpath_mulcore_ary1_a1_I1_p1_l[44]), .Y(n6873));
AND2X1 mul_U19800(.A(dpath_mulcore_b11[1]), .B(n12711), .Y(dpath_mulcore_ary1_a1_I1_p0_l[44]));
INVX1 mul_U19801(.A(dpath_mulcore_ary1_a1_I1_p0_l[44]), .Y(n6874));
AND2X1 mul_U19802(.A(dpath_mulcore_b13[1]), .B(n12714), .Y(dpath_mulcore_ary1_a1_I1_p2_l[43]));
INVX1 mul_U19803(.A(dpath_mulcore_ary1_a1_I1_p2_l[43]), .Y(n6875));
AND2X1 mul_U19804(.A(dpath_mulcore_b12[1]), .B(n12717), .Y(dpath_mulcore_ary1_a1_I1_p1_l[43]));
INVX1 mul_U19805(.A(dpath_mulcore_ary1_a1_I1_p1_l[43]), .Y(n6876));
AND2X1 mul_U19806(.A(dpath_mulcore_b11[1]), .B(n12720), .Y(dpath_mulcore_ary1_a1_I1_p0_l[43]));
INVX1 mul_U19807(.A(dpath_mulcore_ary1_a1_I1_p0_l[43]), .Y(n6877));
AND2X1 mul_U19808(.A(dpath_mulcore_b13[1]), .B(n12723), .Y(dpath_mulcore_ary1_a1_I1_p2_l[42]));
INVX1 mul_U19809(.A(dpath_mulcore_ary1_a1_I1_p2_l[42]), .Y(n6878));
AND2X1 mul_U19810(.A(dpath_mulcore_b12[1]), .B(n12726), .Y(dpath_mulcore_ary1_a1_I1_p1_l[42]));
INVX1 mul_U19811(.A(dpath_mulcore_ary1_a1_I1_p1_l[42]), .Y(n6879));
AND2X1 mul_U19812(.A(dpath_mulcore_b11[1]), .B(n12729), .Y(dpath_mulcore_ary1_a1_I1_p0_l[42]));
INVX1 mul_U19813(.A(dpath_mulcore_ary1_a1_I1_p0_l[42]), .Y(n6880));
AND2X1 mul_U19814(.A(dpath_mulcore_b13[1]), .B(n12732), .Y(dpath_mulcore_ary1_a1_I1_p2_l[41]));
INVX1 mul_U19815(.A(dpath_mulcore_ary1_a1_I1_p2_l[41]), .Y(n6881));
AND2X1 mul_U19816(.A(dpath_mulcore_b12[1]), .B(n12735), .Y(dpath_mulcore_ary1_a1_I1_p1_l[41]));
INVX1 mul_U19817(.A(dpath_mulcore_ary1_a1_I1_p1_l[41]), .Y(n6882));
AND2X1 mul_U19818(.A(dpath_mulcore_b11[1]), .B(n12738), .Y(dpath_mulcore_ary1_a1_I1_p0_l[41]));
INVX1 mul_U19819(.A(dpath_mulcore_ary1_a1_I1_p0_l[41]), .Y(n6883));
AND2X1 mul_U19820(.A(dpath_mulcore_b13[1]), .B(n12741), .Y(dpath_mulcore_ary1_a1_I1_p2_l[40]));
INVX1 mul_U19821(.A(dpath_mulcore_ary1_a1_I1_p2_l[40]), .Y(n6884));
AND2X1 mul_U19822(.A(dpath_mulcore_b12[1]), .B(n12744), .Y(dpath_mulcore_ary1_a1_I1_p1_l[40]));
INVX1 mul_U19823(.A(dpath_mulcore_ary1_a1_I1_p1_l[40]), .Y(n6885));
AND2X1 mul_U19824(.A(dpath_mulcore_b11[1]), .B(n12747), .Y(dpath_mulcore_ary1_a1_I1_p0_l[40]));
INVX1 mul_U19825(.A(dpath_mulcore_ary1_a1_I1_p0_l[40]), .Y(n6886));
AND2X1 mul_U19826(.A(dpath_mulcore_b13[1]), .B(n12750), .Y(dpath_mulcore_ary1_a1_I1_p2_l[39]));
INVX1 mul_U19827(.A(dpath_mulcore_ary1_a1_I1_p2_l[39]), .Y(n6887));
AND2X1 mul_U19828(.A(dpath_mulcore_b12[1]), .B(n12753), .Y(dpath_mulcore_ary1_a1_I1_p1_l[39]));
INVX1 mul_U19829(.A(dpath_mulcore_ary1_a1_I1_p1_l[39]), .Y(n6888));
AND2X1 mul_U19830(.A(dpath_mulcore_b11[1]), .B(n12756), .Y(dpath_mulcore_ary1_a1_I1_p0_l[39]));
INVX1 mul_U19831(.A(dpath_mulcore_ary1_a1_I1_p0_l[39]), .Y(n6889));
AND2X1 mul_U19832(.A(dpath_mulcore_b13[1]), .B(n12759), .Y(dpath_mulcore_ary1_a1_I1_p2_l[38]));
INVX1 mul_U19833(.A(dpath_mulcore_ary1_a1_I1_p2_l[38]), .Y(n6890));
AND2X1 mul_U19834(.A(dpath_mulcore_b12[1]), .B(n12762), .Y(dpath_mulcore_ary1_a1_I1_p1_l[38]));
INVX1 mul_U19835(.A(dpath_mulcore_ary1_a1_I1_p1_l[38]), .Y(n6891));
AND2X1 mul_U19836(.A(dpath_mulcore_b11[1]), .B(n12765), .Y(dpath_mulcore_ary1_a1_I1_p0_l[38]));
INVX1 mul_U19837(.A(dpath_mulcore_ary1_a1_I1_p0_l[38]), .Y(n6892));
AND2X1 mul_U19838(.A(dpath_mulcore_b13[1]), .B(n12768), .Y(dpath_mulcore_ary1_a1_I1_p2_l[37]));
INVX1 mul_U19839(.A(dpath_mulcore_ary1_a1_I1_p2_l[37]), .Y(n6893));
AND2X1 mul_U19840(.A(dpath_mulcore_b12[1]), .B(n12771), .Y(dpath_mulcore_ary1_a1_I1_p1_l[37]));
INVX1 mul_U19841(.A(dpath_mulcore_ary1_a1_I1_p1_l[37]), .Y(n6894));
AND2X1 mul_U19842(.A(dpath_mulcore_b11[1]), .B(n12774), .Y(dpath_mulcore_ary1_a1_I1_p0_l[37]));
INVX1 mul_U19843(.A(dpath_mulcore_ary1_a1_I1_p0_l[37]), .Y(n6895));
AND2X1 mul_U19844(.A(dpath_mulcore_b13[1]), .B(n12777), .Y(dpath_mulcore_ary1_a1_I1_p2_l[36]));
INVX1 mul_U19845(.A(dpath_mulcore_ary1_a1_I1_p2_l[36]), .Y(n6896));
AND2X1 mul_U19846(.A(dpath_mulcore_b12[1]), .B(n12780), .Y(dpath_mulcore_ary1_a1_I1_p1_l[36]));
INVX1 mul_U19847(.A(dpath_mulcore_ary1_a1_I1_p1_l[36]), .Y(n6897));
AND2X1 mul_U19848(.A(dpath_mulcore_b11[1]), .B(n12783), .Y(dpath_mulcore_ary1_a1_I1_p0_l[36]));
INVX1 mul_U19849(.A(dpath_mulcore_ary1_a1_I1_p0_l[36]), .Y(n6898));
AND2X1 mul_U19850(.A(dpath_mulcore_b13[1]), .B(n12786), .Y(dpath_mulcore_ary1_a1_I1_p2_l[35]));
INVX1 mul_U19851(.A(dpath_mulcore_ary1_a1_I1_p2_l[35]), .Y(n6899));
AND2X1 mul_U19852(.A(dpath_mulcore_b12[1]), .B(n12789), .Y(dpath_mulcore_ary1_a1_I1_p1_l[35]));
INVX1 mul_U19853(.A(dpath_mulcore_ary1_a1_I1_p1_l[35]), .Y(n6900));
AND2X1 mul_U19854(.A(dpath_mulcore_b11[1]), .B(n12792), .Y(dpath_mulcore_ary1_a1_I1_p0_l[35]));
INVX1 mul_U19855(.A(dpath_mulcore_ary1_a1_I1_p0_l[35]), .Y(n6901));
AND2X1 mul_U19856(.A(dpath_mulcore_b13[1]), .B(n12795), .Y(dpath_mulcore_ary1_a1_I1_p2_l[34]));
INVX1 mul_U19857(.A(dpath_mulcore_ary1_a1_I1_p2_l[34]), .Y(n6902));
AND2X1 mul_U19858(.A(dpath_mulcore_b12[1]), .B(n12798), .Y(dpath_mulcore_ary1_a1_I1_p1_l[34]));
INVX1 mul_U19859(.A(dpath_mulcore_ary1_a1_I1_p1_l[34]), .Y(n6903));
AND2X1 mul_U19860(.A(dpath_mulcore_b11[1]), .B(n12801), .Y(dpath_mulcore_ary1_a1_I1_p0_l[34]));
INVX1 mul_U19861(.A(dpath_mulcore_ary1_a1_I1_p0_l[34]), .Y(n6904));
AND2X1 mul_U19862(.A(dpath_mulcore_b13[1]), .B(n12804), .Y(dpath_mulcore_ary1_a1_I1_p2_l[33]));
INVX1 mul_U19863(.A(dpath_mulcore_ary1_a1_I1_p2_l[33]), .Y(n6905));
AND2X1 mul_U19864(.A(dpath_mulcore_b12[1]), .B(n12807), .Y(dpath_mulcore_ary1_a1_I1_p1_l[33]));
INVX1 mul_U19865(.A(dpath_mulcore_ary1_a1_I1_p1_l[33]), .Y(n6906));
AND2X1 mul_U19866(.A(dpath_mulcore_b11[1]), .B(n12810), .Y(dpath_mulcore_ary1_a1_I1_p0_l[33]));
INVX1 mul_U19867(.A(dpath_mulcore_ary1_a1_I1_p0_l[33]), .Y(n6907));
AND2X1 mul_U19868(.A(dpath_mulcore_b13[1]), .B(n12813), .Y(dpath_mulcore_ary1_a1_I1_p2_l[32]));
INVX1 mul_U19869(.A(dpath_mulcore_ary1_a1_I1_p2_l[32]), .Y(n6908));
AND2X1 mul_U19870(.A(dpath_mulcore_b12[1]), .B(n12816), .Y(dpath_mulcore_ary1_a1_I1_p1_l[32]));
INVX1 mul_U19871(.A(dpath_mulcore_ary1_a1_I1_p1_l[32]), .Y(n6909));
AND2X1 mul_U19872(.A(dpath_mulcore_b11[1]), .B(n12819), .Y(dpath_mulcore_ary1_a1_I1_p0_l[32]));
INVX1 mul_U19873(.A(dpath_mulcore_ary1_a1_I1_p0_l[32]), .Y(n6910));
AND2X1 mul_U19874(.A(dpath_mulcore_b13[1]), .B(n12822), .Y(dpath_mulcore_ary1_a1_I1_p2_l[31]));
INVX1 mul_U19875(.A(dpath_mulcore_ary1_a1_I1_p2_l[31]), .Y(n6911));
AND2X1 mul_U19876(.A(dpath_mulcore_b12[1]), .B(n12825), .Y(dpath_mulcore_ary1_a1_I1_p1_l[31]));
INVX1 mul_U19877(.A(dpath_mulcore_ary1_a1_I1_p1_l[31]), .Y(n6912));
AND2X1 mul_U19878(.A(dpath_mulcore_b11[1]), .B(n12828), .Y(dpath_mulcore_ary1_a1_I1_p0_l[31]));
INVX1 mul_U19879(.A(dpath_mulcore_ary1_a1_I1_p0_l[31]), .Y(n6913));
AND2X1 mul_U19880(.A(dpath_mulcore_b13[1]), .B(n12831), .Y(dpath_mulcore_ary1_a1_I1_p2_l[30]));
INVX1 mul_U19881(.A(dpath_mulcore_ary1_a1_I1_p2_l[30]), .Y(n6914));
AND2X1 mul_U19882(.A(dpath_mulcore_b12[1]), .B(n12834), .Y(dpath_mulcore_ary1_a1_I1_p1_l[30]));
INVX1 mul_U19883(.A(dpath_mulcore_ary1_a1_I1_p1_l[30]), .Y(n6915));
AND2X1 mul_U19884(.A(dpath_mulcore_b11[1]), .B(n12837), .Y(dpath_mulcore_ary1_a1_I1_p0_l[30]));
INVX1 mul_U19885(.A(dpath_mulcore_ary1_a1_I1_p0_l[30]), .Y(n6916));
AND2X1 mul_U19886(.A(dpath_mulcore_b13[1]), .B(n12840), .Y(dpath_mulcore_ary1_a1_I1_p2_l[29]));
INVX1 mul_U19887(.A(dpath_mulcore_ary1_a1_I1_p2_l[29]), .Y(n6917));
AND2X1 mul_U19888(.A(dpath_mulcore_b12[1]), .B(n12843), .Y(dpath_mulcore_ary1_a1_I1_p1_l[29]));
INVX1 mul_U19889(.A(dpath_mulcore_ary1_a1_I1_p1_l[29]), .Y(n6918));
AND2X1 mul_U19890(.A(dpath_mulcore_b11[1]), .B(n12846), .Y(dpath_mulcore_ary1_a1_I1_p0_l[29]));
INVX1 mul_U19891(.A(dpath_mulcore_ary1_a1_I1_p0_l[29]), .Y(n6919));
AND2X1 mul_U19892(.A(dpath_mulcore_b13[1]), .B(n12849), .Y(dpath_mulcore_ary1_a1_I1_p2_l[28]));
INVX1 mul_U19893(.A(dpath_mulcore_ary1_a1_I1_p2_l[28]), .Y(n6920));
AND2X1 mul_U19894(.A(dpath_mulcore_b12[1]), .B(n12852), .Y(dpath_mulcore_ary1_a1_I1_p1_l[28]));
INVX1 mul_U19895(.A(dpath_mulcore_ary1_a1_I1_p1_l[28]), .Y(n6921));
AND2X1 mul_U19896(.A(dpath_mulcore_b11[1]), .B(n12855), .Y(dpath_mulcore_ary1_a1_I1_p0_l[28]));
INVX1 mul_U19897(.A(dpath_mulcore_ary1_a1_I1_p0_l[28]), .Y(n6922));
AND2X1 mul_U19898(.A(dpath_mulcore_b13[1]), .B(n12858), .Y(dpath_mulcore_ary1_a1_I1_p2_l[27]));
INVX1 mul_U19899(.A(dpath_mulcore_ary1_a1_I1_p2_l[27]), .Y(n6923));
AND2X1 mul_U19900(.A(dpath_mulcore_b12[1]), .B(n12861), .Y(dpath_mulcore_ary1_a1_I1_p1_l[27]));
INVX1 mul_U19901(.A(dpath_mulcore_ary1_a1_I1_p1_l[27]), .Y(n6924));
AND2X1 mul_U19902(.A(dpath_mulcore_b11[1]), .B(n12864), .Y(dpath_mulcore_ary1_a1_I1_p0_l[27]));
INVX1 mul_U19903(.A(dpath_mulcore_ary1_a1_I1_p0_l[27]), .Y(n6925));
AND2X1 mul_U19904(.A(dpath_mulcore_b13[1]), .B(n12867), .Y(dpath_mulcore_ary1_a1_I1_p2_l[26]));
INVX1 mul_U19905(.A(dpath_mulcore_ary1_a1_I1_p2_l[26]), .Y(n6926));
AND2X1 mul_U19906(.A(dpath_mulcore_b12[1]), .B(n12870), .Y(dpath_mulcore_ary1_a1_I1_p1_l[26]));
INVX1 mul_U19907(.A(dpath_mulcore_ary1_a1_I1_p1_l[26]), .Y(n6927));
AND2X1 mul_U19908(.A(dpath_mulcore_b11[1]), .B(n12873), .Y(dpath_mulcore_ary1_a1_I1_p0_l[26]));
INVX1 mul_U19909(.A(dpath_mulcore_ary1_a1_I1_p0_l[26]), .Y(n6928));
AND2X1 mul_U19910(.A(dpath_mulcore_b13[1]), .B(n12876), .Y(dpath_mulcore_ary1_a1_I1_p2_l[25]));
INVX1 mul_U19911(.A(dpath_mulcore_ary1_a1_I1_p2_l[25]), .Y(n6929));
AND2X1 mul_U19912(.A(dpath_mulcore_b12[1]), .B(n12879), .Y(dpath_mulcore_ary1_a1_I1_p1_l[25]));
INVX1 mul_U19913(.A(dpath_mulcore_ary1_a1_I1_p1_l[25]), .Y(n6930));
AND2X1 mul_U19914(.A(dpath_mulcore_b11[1]), .B(n12882), .Y(dpath_mulcore_ary1_a1_I1_p0_l[25]));
INVX1 mul_U19915(.A(dpath_mulcore_ary1_a1_I1_p0_l[25]), .Y(n6931));
AND2X1 mul_U19916(.A(dpath_mulcore_b13[1]), .B(n12885), .Y(dpath_mulcore_ary1_a1_I1_p2_l[24]));
INVX1 mul_U19917(.A(dpath_mulcore_ary1_a1_I1_p2_l[24]), .Y(n6932));
AND2X1 mul_U19918(.A(dpath_mulcore_b12[1]), .B(n12888), .Y(dpath_mulcore_ary1_a1_I1_p1_l[24]));
INVX1 mul_U19919(.A(dpath_mulcore_ary1_a1_I1_p1_l[24]), .Y(n6933));
AND2X1 mul_U19920(.A(dpath_mulcore_b11[1]), .B(n12891), .Y(dpath_mulcore_ary1_a1_I1_p0_l[24]));
INVX1 mul_U19921(.A(dpath_mulcore_ary1_a1_I1_p0_l[24]), .Y(n6934));
AND2X1 mul_U19922(.A(dpath_mulcore_b13[1]), .B(n12894), .Y(dpath_mulcore_ary1_a1_I1_p2_l[23]));
INVX1 mul_U19923(.A(dpath_mulcore_ary1_a1_I1_p2_l[23]), .Y(n6935));
AND2X1 mul_U19924(.A(dpath_mulcore_b12[1]), .B(n12897), .Y(dpath_mulcore_ary1_a1_I1_p1_l[23]));
INVX1 mul_U19925(.A(dpath_mulcore_ary1_a1_I1_p1_l[23]), .Y(n6936));
AND2X1 mul_U19926(.A(dpath_mulcore_b11[1]), .B(n12900), .Y(dpath_mulcore_ary1_a1_I1_p0_l[23]));
INVX1 mul_U19927(.A(dpath_mulcore_ary1_a1_I1_p0_l[23]), .Y(n6937));
AND2X1 mul_U19928(.A(dpath_mulcore_b13[1]), .B(n12903), .Y(dpath_mulcore_ary1_a1_I1_p2_l[22]));
INVX1 mul_U19929(.A(dpath_mulcore_ary1_a1_I1_p2_l[22]), .Y(n6938));
AND2X1 mul_U19930(.A(dpath_mulcore_b12[1]), .B(n12906), .Y(dpath_mulcore_ary1_a1_I1_p1_l[22]));
INVX1 mul_U19931(.A(dpath_mulcore_ary1_a1_I1_p1_l[22]), .Y(n6939));
AND2X1 mul_U19932(.A(dpath_mulcore_b11[1]), .B(n12909), .Y(dpath_mulcore_ary1_a1_I1_p0_l[22]));
INVX1 mul_U19933(.A(dpath_mulcore_ary1_a1_I1_p0_l[22]), .Y(n6940));
AND2X1 mul_U19934(.A(dpath_mulcore_b13[1]), .B(n12912), .Y(dpath_mulcore_ary1_a1_I1_p2_l[21]));
INVX1 mul_U19935(.A(dpath_mulcore_ary1_a1_I1_p2_l[21]), .Y(n6941));
AND2X1 mul_U19936(.A(dpath_mulcore_b12[1]), .B(n12915), .Y(dpath_mulcore_ary1_a1_I1_p1_l[21]));
INVX1 mul_U19937(.A(dpath_mulcore_ary1_a1_I1_p1_l[21]), .Y(n6942));
AND2X1 mul_U19938(.A(dpath_mulcore_b11[1]), .B(n12918), .Y(dpath_mulcore_ary1_a1_I1_p0_l[21]));
INVX1 mul_U19939(.A(dpath_mulcore_ary1_a1_I1_p0_l[21]), .Y(n6943));
AND2X1 mul_U19940(.A(dpath_mulcore_b13[1]), .B(n12921), .Y(dpath_mulcore_ary1_a1_I1_p2_l[20]));
INVX1 mul_U19941(.A(dpath_mulcore_ary1_a1_I1_p2_l[20]), .Y(n6944));
AND2X1 mul_U19942(.A(dpath_mulcore_b12[1]), .B(n12924), .Y(dpath_mulcore_ary1_a1_I1_p1_l[20]));
INVX1 mul_U19943(.A(dpath_mulcore_ary1_a1_I1_p1_l[20]), .Y(n6945));
AND2X1 mul_U19944(.A(dpath_mulcore_b11[1]), .B(n12927), .Y(dpath_mulcore_ary1_a1_I1_p0_l[20]));
INVX1 mul_U19945(.A(dpath_mulcore_ary1_a1_I1_p0_l[20]), .Y(n6946));
AND2X1 mul_U19946(.A(dpath_mulcore_b13[1]), .B(n12930), .Y(dpath_mulcore_ary1_a1_I1_p2_l[19]));
INVX1 mul_U19947(.A(dpath_mulcore_ary1_a1_I1_p2_l[19]), .Y(n6947));
AND2X1 mul_U19948(.A(dpath_mulcore_b12[1]), .B(n12933), .Y(dpath_mulcore_ary1_a1_I1_p1_l[19]));
INVX1 mul_U19949(.A(dpath_mulcore_ary1_a1_I1_p1_l[19]), .Y(n6948));
AND2X1 mul_U19950(.A(dpath_mulcore_b11[1]), .B(n12936), .Y(dpath_mulcore_ary1_a1_I1_p0_l[19]));
INVX1 mul_U19951(.A(dpath_mulcore_ary1_a1_I1_p0_l[19]), .Y(n6949));
AND2X1 mul_U19952(.A(dpath_mulcore_b13[1]), .B(n12939), .Y(dpath_mulcore_ary1_a1_I1_p2_l[18]));
INVX1 mul_U19953(.A(dpath_mulcore_ary1_a1_I1_p2_l[18]), .Y(n6950));
AND2X1 mul_U19954(.A(dpath_mulcore_b12[1]), .B(n12942), .Y(dpath_mulcore_ary1_a1_I1_p1_l[18]));
INVX1 mul_U19955(.A(dpath_mulcore_ary1_a1_I1_p1_l[18]), .Y(n6951));
AND2X1 mul_U19956(.A(dpath_mulcore_b11[1]), .B(n12945), .Y(dpath_mulcore_ary1_a1_I1_p0_l[18]));
INVX1 mul_U19957(.A(dpath_mulcore_ary1_a1_I1_p0_l[18]), .Y(n6952));
AND2X1 mul_U19958(.A(dpath_mulcore_b13[1]), .B(n12948), .Y(dpath_mulcore_ary1_a1_I1_p2_l[17]));
INVX1 mul_U19959(.A(dpath_mulcore_ary1_a1_I1_p2_l[17]), .Y(n6953));
AND2X1 mul_U19960(.A(dpath_mulcore_b12[1]), .B(n12951), .Y(dpath_mulcore_ary1_a1_I1_p1_l[17]));
INVX1 mul_U19961(.A(dpath_mulcore_ary1_a1_I1_p1_l[17]), .Y(n6954));
AND2X1 mul_U19962(.A(dpath_mulcore_b11[1]), .B(n12954), .Y(dpath_mulcore_ary1_a1_I1_p0_l[17]));
INVX1 mul_U19963(.A(dpath_mulcore_ary1_a1_I1_p0_l[17]), .Y(n6955));
AND2X1 mul_U19964(.A(dpath_mulcore_b13[1]), .B(n12957), .Y(dpath_mulcore_ary1_a1_I1_p2_l[16]));
INVX1 mul_U19965(.A(dpath_mulcore_ary1_a1_I1_p2_l[16]), .Y(n6956));
AND2X1 mul_U19966(.A(dpath_mulcore_b12[1]), .B(n12960), .Y(dpath_mulcore_ary1_a1_I1_p1_l[16]));
INVX1 mul_U19967(.A(dpath_mulcore_ary1_a1_I1_p1_l[16]), .Y(n6957));
AND2X1 mul_U19968(.A(dpath_mulcore_b11[1]), .B(n12963), .Y(dpath_mulcore_ary1_a1_I1_p0_l[16]));
INVX1 mul_U19969(.A(dpath_mulcore_ary1_a1_I1_p0_l[16]), .Y(n6958));
AND2X1 mul_U19970(.A(dpath_mulcore_b13[1]), .B(n12966), .Y(dpath_mulcore_ary1_a1_I1_p2_l[15]));
INVX1 mul_U19971(.A(dpath_mulcore_ary1_a1_I1_p2_l[15]), .Y(n6959));
AND2X1 mul_U19972(.A(dpath_mulcore_b12[1]), .B(n12969), .Y(dpath_mulcore_ary1_a1_I1_p1_l[15]));
INVX1 mul_U19973(.A(dpath_mulcore_ary1_a1_I1_p1_l[15]), .Y(n6960));
AND2X1 mul_U19974(.A(dpath_mulcore_b11[1]), .B(n12972), .Y(dpath_mulcore_ary1_a1_I1_p0_l[15]));
INVX1 mul_U19975(.A(dpath_mulcore_ary1_a1_I1_p0_l[15]), .Y(n6961));
AND2X1 mul_U19976(.A(dpath_mulcore_b13[1]), .B(n12975), .Y(dpath_mulcore_ary1_a1_I1_p2_l[14]));
INVX1 mul_U19977(.A(dpath_mulcore_ary1_a1_I1_p2_l[14]), .Y(n6962));
AND2X1 mul_U19978(.A(dpath_mulcore_b12[1]), .B(n12978), .Y(dpath_mulcore_ary1_a1_I1_p1_l[14]));
INVX1 mul_U19979(.A(dpath_mulcore_ary1_a1_I1_p1_l[14]), .Y(n6963));
AND2X1 mul_U19980(.A(dpath_mulcore_b11[1]), .B(n12981), .Y(dpath_mulcore_ary1_a1_I1_p0_l[14]));
INVX1 mul_U19981(.A(dpath_mulcore_ary1_a1_I1_p0_l[14]), .Y(n6964));
AND2X1 mul_U19982(.A(dpath_mulcore_b13[1]), .B(n12984), .Y(dpath_mulcore_ary1_a1_I1_p2_l[13]));
INVX1 mul_U19983(.A(dpath_mulcore_ary1_a1_I1_p2_l[13]), .Y(n6965));
AND2X1 mul_U19984(.A(dpath_mulcore_b12[1]), .B(n12987), .Y(dpath_mulcore_ary1_a1_I1_p1_l[13]));
INVX1 mul_U19985(.A(dpath_mulcore_ary1_a1_I1_p1_l[13]), .Y(n6966));
AND2X1 mul_U19986(.A(dpath_mulcore_b11[1]), .B(n12990), .Y(dpath_mulcore_ary1_a1_I1_p0_l[13]));
INVX1 mul_U19987(.A(dpath_mulcore_ary1_a1_I1_p0_l[13]), .Y(n6967));
AND2X1 mul_U19988(.A(dpath_mulcore_b13[1]), .B(n12993), .Y(dpath_mulcore_ary1_a1_I1_p2_l[12]));
INVX1 mul_U19989(.A(dpath_mulcore_ary1_a1_I1_p2_l[12]), .Y(n6968));
AND2X1 mul_U19990(.A(dpath_mulcore_b12[1]), .B(n12996), .Y(dpath_mulcore_ary1_a1_I1_p1_l[12]));
INVX1 mul_U19991(.A(dpath_mulcore_ary1_a1_I1_p1_l[12]), .Y(n6969));
AND2X1 mul_U19992(.A(dpath_mulcore_b11[1]), .B(n12999), .Y(dpath_mulcore_ary1_a1_I1_p0_l[12]));
INVX1 mul_U19993(.A(dpath_mulcore_ary1_a1_I1_p0_l[12]), .Y(n6970));
AND2X1 mul_U19994(.A(dpath_mulcore_b13[1]), .B(n13002), .Y(dpath_mulcore_ary1_a1_I1_p2_l[11]));
INVX1 mul_U19995(.A(dpath_mulcore_ary1_a1_I1_p2_l[11]), .Y(n6971));
AND2X1 mul_U19996(.A(dpath_mulcore_b12[1]), .B(n13005), .Y(dpath_mulcore_ary1_a1_I1_p1_l[11]));
INVX1 mul_U19997(.A(dpath_mulcore_ary1_a1_I1_p1_l[11]), .Y(n6972));
AND2X1 mul_U19998(.A(dpath_mulcore_b11[1]), .B(n13008), .Y(dpath_mulcore_ary1_a1_I1_p0_l[11]));
INVX1 mul_U19999(.A(dpath_mulcore_ary1_a1_I1_p0_l[11]), .Y(n6973));
AND2X1 mul_U20000(.A(dpath_mulcore_b13[1]), .B(n13011), .Y(dpath_mulcore_ary1_a1_I1_p2_l[10]));
INVX1 mul_U20001(.A(dpath_mulcore_ary1_a1_I1_p2_l[10]), .Y(n6974));
AND2X1 mul_U20002(.A(dpath_mulcore_b12[1]), .B(n13014), .Y(dpath_mulcore_ary1_a1_I1_p1_l[10]));
INVX1 mul_U20003(.A(dpath_mulcore_ary1_a1_I1_p1_l[10]), .Y(n6975));
AND2X1 mul_U20004(.A(dpath_mulcore_b11[1]), .B(n13017), .Y(dpath_mulcore_ary1_a1_I1_p0_l[10]));
INVX1 mul_U20005(.A(dpath_mulcore_ary1_a1_I1_p0_l[10]), .Y(n6976));
AND2X1 mul_U20006(.A(dpath_mulcore_b13[1]), .B(n13020), .Y(dpath_mulcore_ary1_a1_I1_p2_l[9]));
INVX1 mul_U20007(.A(dpath_mulcore_ary1_a1_I1_p2_l[9]), .Y(n6977));
AND2X1 mul_U20008(.A(dpath_mulcore_b12[1]), .B(n13023), .Y(dpath_mulcore_ary1_a1_I1_p1_l[9]));
INVX1 mul_U20009(.A(dpath_mulcore_ary1_a1_I1_p1_l[9]), .Y(n6978));
AND2X1 mul_U20010(.A(dpath_mulcore_b11[1]), .B(n13026), .Y(dpath_mulcore_ary1_a1_I1_p0_l[9]));
INVX1 mul_U20011(.A(dpath_mulcore_ary1_a1_I1_p0_l[9]), .Y(n6979));
AND2X1 mul_U20012(.A(dpath_mulcore_b13[1]), .B(n13029), .Y(dpath_mulcore_ary1_a1_I1_p2_l[8]));
INVX1 mul_U20013(.A(dpath_mulcore_ary1_a1_I1_p2_l[8]), .Y(n6980));
AND2X1 mul_U20014(.A(dpath_mulcore_b12[1]), .B(n13032), .Y(dpath_mulcore_ary1_a1_I1_p1_l[8]));
INVX1 mul_U20015(.A(dpath_mulcore_ary1_a1_I1_p1_l[8]), .Y(n6981));
AND2X1 mul_U20016(.A(dpath_mulcore_b11[1]), .B(n13035), .Y(dpath_mulcore_ary1_a1_I1_p0_l[8]));
INVX1 mul_U20017(.A(dpath_mulcore_ary1_a1_I1_p0_l[8]), .Y(n6982));
AND2X1 mul_U20018(.A(dpath_mulcore_b13[1]), .B(n13038), .Y(dpath_mulcore_ary1_a1_I1_p2_l[7]));
INVX1 mul_U20019(.A(dpath_mulcore_ary1_a1_I1_p2_l[7]), .Y(n6983));
AND2X1 mul_U20020(.A(dpath_mulcore_b12[1]), .B(n13041), .Y(dpath_mulcore_ary1_a1_I1_p1_l[7]));
INVX1 mul_U20021(.A(dpath_mulcore_ary1_a1_I1_p1_l[7]), .Y(n6984));
AND2X1 mul_U20022(.A(dpath_mulcore_b11[1]), .B(n13044), .Y(dpath_mulcore_ary1_a1_I1_p0_l[7]));
INVX1 mul_U20023(.A(dpath_mulcore_ary1_a1_I1_p0_l[7]), .Y(n6985));
AND2X1 mul_U20024(.A(dpath_mulcore_b13[1]), .B(n13047), .Y(dpath_mulcore_ary1_a1_I1_p2_l[6]));
INVX1 mul_U20025(.A(dpath_mulcore_ary1_a1_I1_p2_l[6]), .Y(n6986));
AND2X1 mul_U20026(.A(dpath_mulcore_b12[1]), .B(n13050), .Y(dpath_mulcore_ary1_a1_I1_p1_l[6]));
INVX1 mul_U20027(.A(dpath_mulcore_ary1_a1_I1_p1_l[6]), .Y(n6987));
AND2X1 mul_U20028(.A(dpath_mulcore_b11[1]), .B(n13053), .Y(dpath_mulcore_ary1_a1_I1_p0_l[6]));
INVX1 mul_U20029(.A(dpath_mulcore_ary1_a1_I1_p0_l[6]), .Y(n6988));
AND2X1 mul_U20030(.A(dpath_mulcore_b13[1]), .B(n13056), .Y(dpath_mulcore_ary1_a1_I1_p2_l[5]));
INVX1 mul_U20031(.A(dpath_mulcore_ary1_a1_I1_p2_l[5]), .Y(n6989));
AND2X1 mul_U20032(.A(dpath_mulcore_b12[1]), .B(n13059), .Y(dpath_mulcore_ary1_a1_I1_p1_l[5]));
INVX1 mul_U20033(.A(dpath_mulcore_ary1_a1_I1_p1_l[5]), .Y(n6990));
AND2X1 mul_U20034(.A(dpath_mulcore_b11[1]), .B(n13062), .Y(dpath_mulcore_ary1_a1_I1_p0_l[5]));
INVX1 mul_U20035(.A(dpath_mulcore_ary1_a1_I1_p0_l[5]), .Y(n6991));
AND2X1 mul_U20036(.A(dpath_mulcore_b13[1]), .B(n13064), .Y(dpath_mulcore_ary1_a1_I1_p2_l[4]));
INVX1 mul_U20037(.A(dpath_mulcore_ary1_a1_I1_p2_l[4]), .Y(n6992));
AND2X1 mul_U20038(.A(dpath_mulcore_b12[1]), .B(n13067), .Y(dpath_mulcore_ary1_a1_I1_p1_l[4]));
INVX1 mul_U20039(.A(dpath_mulcore_ary1_a1_I1_p1_l[4]), .Y(n6993));
AND2X1 mul_U20040(.A(dpath_mulcore_b11[1]), .B(n13070), .Y(dpath_mulcore_ary1_a1_I1_p0_l[4]));
INVX1 mul_U20041(.A(dpath_mulcore_ary1_a1_I1_p0_l[4]), .Y(n6994));
AND2X1 mul_U20042(.A(dpath_mulcore_b11[1]), .B(n13073), .Y(dpath_mulcore_ary1_a1_I1_p0_l[3]));
INVX1 mul_U20043(.A(dpath_mulcore_ary1_a1_I1_p0_l[3]), .Y(n6995));
AND2X1 mul_U20044(.A(dpath_mulcore_b12[1]), .B(n13076), .Y(dpath_mulcore_ary1_a1_I1_p1_l[3]));
INVX1 mul_U20045(.A(dpath_mulcore_ary1_a1_I1_p1_l[3]), .Y(n6996));
AND2X1 mul_U20046(.A(dpath_mulcore_b11[1]), .B(n13079), .Y(dpath_mulcore_ary1_a1_I1_I0_p0_l_2));
INVX1 mul_U20047(.A(dpath_mulcore_ary1_a1_I1_I0_p0_l_2), .Y(n6997));
AND2X1 mul_U20048(.A(dpath_mulcore_b11[1]), .B(n13082), .Y(dpath_mulcore_ary1_a1_I1_I0_p0_l_1));
INVX1 mul_U20049(.A(dpath_mulcore_ary1_a1_I1_I0_p0_l_1), .Y(n6998));
AND2X1 mul_U20050(.A(dpath_mulcore_b11[1]), .B(n13084), .Y(dpath_mulcore_ary1_a1_I1_I0_p0_l_0));
INVX1 mul_U20051(.A(dpath_mulcore_ary1_a1_I1_I0_p0_l_0), .Y(n6999));
AND2X1 mul_U20052(.A(dpath_mulcore_b12[1]), .B(n13086), .Y(dpath_mulcore_ary1_a1_I1_I0_p1_l_2));
INVX1 mul_U20053(.A(dpath_mulcore_ary1_a1_I1_I0_p1_l_2), .Y(n7000));
AND2X1 mul_U20054(.A(dpath_mulcore_b10[1]), .B(n13089), .Y(dpath_mulcore_ary1_a1_I0_I2_p2_l_67));
INVX1 mul_U20055(.A(dpath_mulcore_ary1_a1_I0_I2_p2_l_67), .Y(n7001));
AND2X1 mul_U20056(.A(dpath_mulcore_b10[1]), .B(n13092), .Y(dpath_mulcore_ary1_a1_I0_I2_p2_l_66));
INVX1 mul_U20057(.A(dpath_mulcore_ary1_a1_I0_I2_p2_l_66), .Y(n7002));
AND2X1 mul_U20058(.A(dpath_mulcore_b10[1]), .B(n13095), .Y(dpath_mulcore_ary1_a1_I0_I2_p2_l_65));
INVX1 mul_U20059(.A(dpath_mulcore_ary1_a1_I0_I2_p2_l_65), .Y(n7003));
AND2X1 mul_U20060(.A(dpath_mulcore_b9[1]), .B(n13098), .Y(dpath_mulcore_ary1_a1_I0_I2_p1_l_65));
INVX1 mul_U20061(.A(dpath_mulcore_ary1_a1_I0_I2_p1_l_65), .Y(n7004));
AND2X1 mul_U20062(.A(dpath_mulcore_b9[1]), .B(n13101), .Y(dpath_mulcore_ary1_a1_I0_I2_p1_l_64));
INVX1 mul_U20063(.A(dpath_mulcore_ary1_a1_I0_I2_p1_l_64), .Y(n7005));
AND2X1 mul_U20064(.A(dpath_mulcore_b10[1]), .B(n13104), .Y(dpath_mulcore_ary1_a1_I0_I2_p2_l_64));
INVX1 mul_U20065(.A(dpath_mulcore_ary1_a1_I0_I2_p2_l_64), .Y(n7006));
AND2X1 mul_U20066(.A(dpath_mulcore_b10[1]), .B(n13107), .Y(dpath_mulcore_ary1_a1_I0_p2_l[63]));
INVX1 mul_U20067(.A(dpath_mulcore_ary1_a1_I0_p2_l[63]), .Y(n7007));
AND2X1 mul_U20068(.A(dpath_mulcore_b9[1]), .B(n13110), .Y(dpath_mulcore_ary1_a1_I0_p1_l[63]));
INVX1 mul_U20069(.A(dpath_mulcore_ary1_a1_I0_p1_l[63]), .Y(n7008));
AND2X1 mul_U20070(.A(dpath_mulcore_b8[1]), .B(n13113), .Y(dpath_mulcore_ary1_a1_I0_p0_l[63]));
INVX1 mul_U20071(.A(dpath_mulcore_ary1_a1_I0_p0_l[63]), .Y(n7009));
AND2X1 mul_U20072(.A(dpath_mulcore_b10[1]), .B(n13116), .Y(dpath_mulcore_ary1_a1_I0_p2_l[62]));
INVX1 mul_U20073(.A(dpath_mulcore_ary1_a1_I0_p2_l[62]), .Y(n7010));
AND2X1 mul_U20074(.A(dpath_mulcore_b9[1]), .B(n13119), .Y(dpath_mulcore_ary1_a1_I0_p1_l[62]));
INVX1 mul_U20075(.A(dpath_mulcore_ary1_a1_I0_p1_l[62]), .Y(n7011));
AND2X1 mul_U20076(.A(dpath_mulcore_b8[1]), .B(n13122), .Y(dpath_mulcore_ary1_a1_I0_p0_l[62]));
INVX1 mul_U20077(.A(dpath_mulcore_ary1_a1_I0_p0_l[62]), .Y(n7012));
AND2X1 mul_U20078(.A(dpath_mulcore_b10[1]), .B(n13125), .Y(dpath_mulcore_ary1_a1_I0_p2_l[61]));
INVX1 mul_U20079(.A(dpath_mulcore_ary1_a1_I0_p2_l[61]), .Y(n7013));
AND2X1 mul_U20080(.A(dpath_mulcore_b9[1]), .B(n13128), .Y(dpath_mulcore_ary1_a1_I0_p1_l[61]));
INVX1 mul_U20081(.A(dpath_mulcore_ary1_a1_I0_p1_l[61]), .Y(n7014));
AND2X1 mul_U20082(.A(dpath_mulcore_b8[1]), .B(n13131), .Y(dpath_mulcore_ary1_a1_I0_p0_l[61]));
INVX1 mul_U20083(.A(dpath_mulcore_ary1_a1_I0_p0_l[61]), .Y(n7015));
AND2X1 mul_U20084(.A(dpath_mulcore_b10[1]), .B(n13134), .Y(dpath_mulcore_ary1_a1_I0_p2_l[60]));
INVX1 mul_U20085(.A(dpath_mulcore_ary1_a1_I0_p2_l[60]), .Y(n7016));
AND2X1 mul_U20086(.A(dpath_mulcore_b9[1]), .B(n13137), .Y(dpath_mulcore_ary1_a1_I0_p1_l[60]));
INVX1 mul_U20087(.A(dpath_mulcore_ary1_a1_I0_p1_l[60]), .Y(n7017));
AND2X1 mul_U20088(.A(dpath_mulcore_b8[1]), .B(n13140), .Y(dpath_mulcore_ary1_a1_I0_p0_l[60]));
INVX1 mul_U20089(.A(dpath_mulcore_ary1_a1_I0_p0_l[60]), .Y(n7018));
AND2X1 mul_U20090(.A(dpath_mulcore_b10[1]), .B(n13143), .Y(dpath_mulcore_ary1_a1_I0_p2_l[59]));
INVX1 mul_U20091(.A(dpath_mulcore_ary1_a1_I0_p2_l[59]), .Y(n7019));
AND2X1 mul_U20092(.A(dpath_mulcore_b9[1]), .B(n13146), .Y(dpath_mulcore_ary1_a1_I0_p1_l[59]));
INVX1 mul_U20093(.A(dpath_mulcore_ary1_a1_I0_p1_l[59]), .Y(n7020));
AND2X1 mul_U20094(.A(dpath_mulcore_b8[1]), .B(n13149), .Y(dpath_mulcore_ary1_a1_I0_p0_l[59]));
INVX1 mul_U20095(.A(dpath_mulcore_ary1_a1_I0_p0_l[59]), .Y(n7021));
AND2X1 mul_U20096(.A(dpath_mulcore_b10[1]), .B(n13152), .Y(dpath_mulcore_ary1_a1_I0_p2_l[58]));
INVX1 mul_U20097(.A(dpath_mulcore_ary1_a1_I0_p2_l[58]), .Y(n7022));
AND2X1 mul_U20098(.A(dpath_mulcore_b9[1]), .B(n13155), .Y(dpath_mulcore_ary1_a1_I0_p1_l[58]));
INVX1 mul_U20099(.A(dpath_mulcore_ary1_a1_I0_p1_l[58]), .Y(n7023));
AND2X1 mul_U20100(.A(dpath_mulcore_b8[1]), .B(n13158), .Y(dpath_mulcore_ary1_a1_I0_p0_l[58]));
INVX1 mul_U20101(.A(dpath_mulcore_ary1_a1_I0_p0_l[58]), .Y(n7024));
AND2X1 mul_U20102(.A(dpath_mulcore_b10[1]), .B(n13161), .Y(dpath_mulcore_ary1_a1_I0_p2_l[57]));
INVX1 mul_U20103(.A(dpath_mulcore_ary1_a1_I0_p2_l[57]), .Y(n7025));
AND2X1 mul_U20104(.A(dpath_mulcore_b9[1]), .B(n13164), .Y(dpath_mulcore_ary1_a1_I0_p1_l[57]));
INVX1 mul_U20105(.A(dpath_mulcore_ary1_a1_I0_p1_l[57]), .Y(n7026));
AND2X1 mul_U20106(.A(dpath_mulcore_b8[1]), .B(n13167), .Y(dpath_mulcore_ary1_a1_I0_p0_l[57]));
INVX1 mul_U20107(.A(dpath_mulcore_ary1_a1_I0_p0_l[57]), .Y(n7027));
AND2X1 mul_U20108(.A(dpath_mulcore_b10[1]), .B(n13170), .Y(dpath_mulcore_ary1_a1_I0_p2_l[56]));
INVX1 mul_U20109(.A(dpath_mulcore_ary1_a1_I0_p2_l[56]), .Y(n7028));
AND2X1 mul_U20110(.A(dpath_mulcore_b9[1]), .B(n13173), .Y(dpath_mulcore_ary1_a1_I0_p1_l[56]));
INVX1 mul_U20111(.A(dpath_mulcore_ary1_a1_I0_p1_l[56]), .Y(n7029));
AND2X1 mul_U20112(.A(dpath_mulcore_b8[1]), .B(n13176), .Y(dpath_mulcore_ary1_a1_I0_p0_l[56]));
INVX1 mul_U20113(.A(dpath_mulcore_ary1_a1_I0_p0_l[56]), .Y(n7030));
AND2X1 mul_U20114(.A(dpath_mulcore_b10[1]), .B(n13179), .Y(dpath_mulcore_ary1_a1_I0_p2_l[55]));
INVX1 mul_U20115(.A(dpath_mulcore_ary1_a1_I0_p2_l[55]), .Y(n7031));
AND2X1 mul_U20116(.A(dpath_mulcore_b9[1]), .B(n13182), .Y(dpath_mulcore_ary1_a1_I0_p1_l[55]));
INVX1 mul_U20117(.A(dpath_mulcore_ary1_a1_I0_p1_l[55]), .Y(n7032));
AND2X1 mul_U20118(.A(dpath_mulcore_b8[1]), .B(n13185), .Y(dpath_mulcore_ary1_a1_I0_p0_l[55]));
INVX1 mul_U20119(.A(dpath_mulcore_ary1_a1_I0_p0_l[55]), .Y(n7033));
AND2X1 mul_U20120(.A(dpath_mulcore_b10[1]), .B(n13188), .Y(dpath_mulcore_ary1_a1_I0_p2_l[54]));
INVX1 mul_U20121(.A(dpath_mulcore_ary1_a1_I0_p2_l[54]), .Y(n7034));
AND2X1 mul_U20122(.A(dpath_mulcore_b9[1]), .B(n13191), .Y(dpath_mulcore_ary1_a1_I0_p1_l[54]));
INVX1 mul_U20123(.A(dpath_mulcore_ary1_a1_I0_p1_l[54]), .Y(n7035));
AND2X1 mul_U20124(.A(dpath_mulcore_b8[1]), .B(n13194), .Y(dpath_mulcore_ary1_a1_I0_p0_l[54]));
INVX1 mul_U20125(.A(dpath_mulcore_ary1_a1_I0_p0_l[54]), .Y(n7036));
AND2X1 mul_U20126(.A(dpath_mulcore_b10[1]), .B(n13197), .Y(dpath_mulcore_ary1_a1_I0_p2_l[53]));
INVX1 mul_U20127(.A(dpath_mulcore_ary1_a1_I0_p2_l[53]), .Y(n7037));
AND2X1 mul_U20128(.A(dpath_mulcore_b9[1]), .B(n13200), .Y(dpath_mulcore_ary1_a1_I0_p1_l[53]));
INVX1 mul_U20129(.A(dpath_mulcore_ary1_a1_I0_p1_l[53]), .Y(n7038));
AND2X1 mul_U20130(.A(dpath_mulcore_b8[1]), .B(n13203), .Y(dpath_mulcore_ary1_a1_I0_p0_l[53]));
INVX1 mul_U20131(.A(dpath_mulcore_ary1_a1_I0_p0_l[53]), .Y(n7039));
AND2X1 mul_U20132(.A(dpath_mulcore_b10[1]), .B(n13206), .Y(dpath_mulcore_ary1_a1_I0_p2_l[52]));
INVX1 mul_U20133(.A(dpath_mulcore_ary1_a1_I0_p2_l[52]), .Y(n7040));
AND2X1 mul_U20134(.A(dpath_mulcore_b9[1]), .B(n13209), .Y(dpath_mulcore_ary1_a1_I0_p1_l[52]));
INVX1 mul_U20135(.A(dpath_mulcore_ary1_a1_I0_p1_l[52]), .Y(n7041));
AND2X1 mul_U20136(.A(dpath_mulcore_b8[1]), .B(n13212), .Y(dpath_mulcore_ary1_a1_I0_p0_l[52]));
INVX1 mul_U20137(.A(dpath_mulcore_ary1_a1_I0_p0_l[52]), .Y(n7042));
AND2X1 mul_U20138(.A(dpath_mulcore_b10[1]), .B(n13215), .Y(dpath_mulcore_ary1_a1_I0_p2_l[51]));
INVX1 mul_U20139(.A(dpath_mulcore_ary1_a1_I0_p2_l[51]), .Y(n7043));
AND2X1 mul_U20140(.A(dpath_mulcore_b9[1]), .B(n13218), .Y(dpath_mulcore_ary1_a1_I0_p1_l[51]));
INVX1 mul_U20141(.A(dpath_mulcore_ary1_a1_I0_p1_l[51]), .Y(n7044));
AND2X1 mul_U20142(.A(dpath_mulcore_b8[1]), .B(n13221), .Y(dpath_mulcore_ary1_a1_I0_p0_l[51]));
INVX1 mul_U20143(.A(dpath_mulcore_ary1_a1_I0_p0_l[51]), .Y(n7045));
AND2X1 mul_U20144(.A(dpath_mulcore_b10[1]), .B(n13224), .Y(dpath_mulcore_ary1_a1_I0_p2_l[50]));
INVX1 mul_U20145(.A(dpath_mulcore_ary1_a1_I0_p2_l[50]), .Y(n7046));
AND2X1 mul_U20146(.A(dpath_mulcore_b9[1]), .B(n13227), .Y(dpath_mulcore_ary1_a1_I0_p1_l[50]));
INVX1 mul_U20147(.A(dpath_mulcore_ary1_a1_I0_p1_l[50]), .Y(n7047));
AND2X1 mul_U20148(.A(dpath_mulcore_b8[1]), .B(n13230), .Y(dpath_mulcore_ary1_a1_I0_p0_l[50]));
INVX1 mul_U20149(.A(dpath_mulcore_ary1_a1_I0_p0_l[50]), .Y(n7048));
AND2X1 mul_U20150(.A(dpath_mulcore_b10[1]), .B(n13233), .Y(dpath_mulcore_ary1_a1_I0_p2_l[49]));
INVX1 mul_U20151(.A(dpath_mulcore_ary1_a1_I0_p2_l[49]), .Y(n7049));
AND2X1 mul_U20152(.A(dpath_mulcore_b9[1]), .B(n13236), .Y(dpath_mulcore_ary1_a1_I0_p1_l[49]));
INVX1 mul_U20153(.A(dpath_mulcore_ary1_a1_I0_p1_l[49]), .Y(n7050));
AND2X1 mul_U20154(.A(dpath_mulcore_b8[1]), .B(n13239), .Y(dpath_mulcore_ary1_a1_I0_p0_l[49]));
INVX1 mul_U20155(.A(dpath_mulcore_ary1_a1_I0_p0_l[49]), .Y(n7051));
AND2X1 mul_U20156(.A(dpath_mulcore_b10[1]), .B(n13242), .Y(dpath_mulcore_ary1_a1_I0_p2_l[48]));
INVX1 mul_U20157(.A(dpath_mulcore_ary1_a1_I0_p2_l[48]), .Y(n7052));
AND2X1 mul_U20158(.A(dpath_mulcore_b9[1]), .B(n13245), .Y(dpath_mulcore_ary1_a1_I0_p1_l[48]));
INVX1 mul_U20159(.A(dpath_mulcore_ary1_a1_I0_p1_l[48]), .Y(n7053));
AND2X1 mul_U20160(.A(dpath_mulcore_b8[1]), .B(n13248), .Y(dpath_mulcore_ary1_a1_I0_p0_l[48]));
INVX1 mul_U20161(.A(dpath_mulcore_ary1_a1_I0_p0_l[48]), .Y(n7054));
AND2X1 mul_U20162(.A(dpath_mulcore_b10[1]), .B(n13251), .Y(dpath_mulcore_ary1_a1_I0_p2_l[47]));
INVX1 mul_U20163(.A(dpath_mulcore_ary1_a1_I0_p2_l[47]), .Y(n7055));
AND2X1 mul_U20164(.A(dpath_mulcore_b9[1]), .B(n13254), .Y(dpath_mulcore_ary1_a1_I0_p1_l[47]));
INVX1 mul_U20165(.A(dpath_mulcore_ary1_a1_I0_p1_l[47]), .Y(n7056));
AND2X1 mul_U20166(.A(dpath_mulcore_b8[1]), .B(n13257), .Y(dpath_mulcore_ary1_a1_I0_p0_l[47]));
INVX1 mul_U20167(.A(dpath_mulcore_ary1_a1_I0_p0_l[47]), .Y(n7057));
AND2X1 mul_U20168(.A(dpath_mulcore_b10[1]), .B(n13260), .Y(dpath_mulcore_ary1_a1_I0_p2_l[46]));
INVX1 mul_U20169(.A(dpath_mulcore_ary1_a1_I0_p2_l[46]), .Y(n7058));
AND2X1 mul_U20170(.A(dpath_mulcore_b9[1]), .B(n13263), .Y(dpath_mulcore_ary1_a1_I0_p1_l[46]));
INVX1 mul_U20171(.A(dpath_mulcore_ary1_a1_I0_p1_l[46]), .Y(n7059));
AND2X1 mul_U20172(.A(dpath_mulcore_b8[1]), .B(n13266), .Y(dpath_mulcore_ary1_a1_I0_p0_l[46]));
INVX1 mul_U20173(.A(dpath_mulcore_ary1_a1_I0_p0_l[46]), .Y(n7060));
AND2X1 mul_U20174(.A(dpath_mulcore_b10[1]), .B(n13269), .Y(dpath_mulcore_ary1_a1_I0_p2_l[45]));
INVX1 mul_U20175(.A(dpath_mulcore_ary1_a1_I0_p2_l[45]), .Y(n7061));
AND2X1 mul_U20176(.A(dpath_mulcore_b9[1]), .B(n13272), .Y(dpath_mulcore_ary1_a1_I0_p1_l[45]));
INVX1 mul_U20177(.A(dpath_mulcore_ary1_a1_I0_p1_l[45]), .Y(n7062));
AND2X1 mul_U20178(.A(dpath_mulcore_b8[1]), .B(n13275), .Y(dpath_mulcore_ary1_a1_I0_p0_l[45]));
INVX1 mul_U20179(.A(dpath_mulcore_ary1_a1_I0_p0_l[45]), .Y(n7063));
AND2X1 mul_U20180(.A(dpath_mulcore_b10[1]), .B(n13278), .Y(dpath_mulcore_ary1_a1_I0_p2_l[44]));
INVX1 mul_U20181(.A(dpath_mulcore_ary1_a1_I0_p2_l[44]), .Y(n7064));
AND2X1 mul_U20182(.A(dpath_mulcore_b9[1]), .B(n13281), .Y(dpath_mulcore_ary1_a1_I0_p1_l[44]));
INVX1 mul_U20183(.A(dpath_mulcore_ary1_a1_I0_p1_l[44]), .Y(n7065));
AND2X1 mul_U20184(.A(dpath_mulcore_b8[1]), .B(n13284), .Y(dpath_mulcore_ary1_a1_I0_p0_l[44]));
INVX1 mul_U20185(.A(dpath_mulcore_ary1_a1_I0_p0_l[44]), .Y(n7066));
AND2X1 mul_U20186(.A(dpath_mulcore_b10[1]), .B(n13287), .Y(dpath_mulcore_ary1_a1_I0_p2_l[43]));
INVX1 mul_U20187(.A(dpath_mulcore_ary1_a1_I0_p2_l[43]), .Y(n7067));
AND2X1 mul_U20188(.A(dpath_mulcore_b9[1]), .B(n13290), .Y(dpath_mulcore_ary1_a1_I0_p1_l[43]));
INVX1 mul_U20189(.A(dpath_mulcore_ary1_a1_I0_p1_l[43]), .Y(n7068));
AND2X1 mul_U20190(.A(dpath_mulcore_b8[1]), .B(n13293), .Y(dpath_mulcore_ary1_a1_I0_p0_l[43]));
INVX1 mul_U20191(.A(dpath_mulcore_ary1_a1_I0_p0_l[43]), .Y(n7069));
AND2X1 mul_U20192(.A(dpath_mulcore_b10[1]), .B(n13296), .Y(dpath_mulcore_ary1_a1_I0_p2_l[42]));
INVX1 mul_U20193(.A(dpath_mulcore_ary1_a1_I0_p2_l[42]), .Y(n7070));
AND2X1 mul_U20194(.A(dpath_mulcore_b9[1]), .B(n13299), .Y(dpath_mulcore_ary1_a1_I0_p1_l[42]));
INVX1 mul_U20195(.A(dpath_mulcore_ary1_a1_I0_p1_l[42]), .Y(n7071));
AND2X1 mul_U20196(.A(dpath_mulcore_b8[1]), .B(n13302), .Y(dpath_mulcore_ary1_a1_I0_p0_l[42]));
INVX1 mul_U20197(.A(dpath_mulcore_ary1_a1_I0_p0_l[42]), .Y(n7072));
AND2X1 mul_U20198(.A(dpath_mulcore_b10[1]), .B(n13305), .Y(dpath_mulcore_ary1_a1_I0_p2_l[41]));
INVX1 mul_U20199(.A(dpath_mulcore_ary1_a1_I0_p2_l[41]), .Y(n7073));
AND2X1 mul_U20200(.A(dpath_mulcore_b9[1]), .B(n13308), .Y(dpath_mulcore_ary1_a1_I0_p1_l[41]));
INVX1 mul_U20201(.A(dpath_mulcore_ary1_a1_I0_p1_l[41]), .Y(n7074));
AND2X1 mul_U20202(.A(dpath_mulcore_b8[1]), .B(n13311), .Y(dpath_mulcore_ary1_a1_I0_p0_l[41]));
INVX1 mul_U20203(.A(dpath_mulcore_ary1_a1_I0_p0_l[41]), .Y(n7075));
AND2X1 mul_U20204(.A(dpath_mulcore_b10[1]), .B(n13314), .Y(dpath_mulcore_ary1_a1_I0_p2_l[40]));
INVX1 mul_U20205(.A(dpath_mulcore_ary1_a1_I0_p2_l[40]), .Y(n7076));
AND2X1 mul_U20206(.A(dpath_mulcore_b9[1]), .B(n13317), .Y(dpath_mulcore_ary1_a1_I0_p1_l[40]));
INVX1 mul_U20207(.A(dpath_mulcore_ary1_a1_I0_p1_l[40]), .Y(n7077));
AND2X1 mul_U20208(.A(dpath_mulcore_b8[1]), .B(n13320), .Y(dpath_mulcore_ary1_a1_I0_p0_l[40]));
INVX1 mul_U20209(.A(dpath_mulcore_ary1_a1_I0_p0_l[40]), .Y(n7078));
AND2X1 mul_U20210(.A(dpath_mulcore_b10[1]), .B(n13323), .Y(dpath_mulcore_ary1_a1_I0_p2_l[39]));
INVX1 mul_U20211(.A(dpath_mulcore_ary1_a1_I0_p2_l[39]), .Y(n7079));
AND2X1 mul_U20212(.A(dpath_mulcore_b9[1]), .B(n13326), .Y(dpath_mulcore_ary1_a1_I0_p1_l[39]));
INVX1 mul_U20213(.A(dpath_mulcore_ary1_a1_I0_p1_l[39]), .Y(n7080));
AND2X1 mul_U20214(.A(dpath_mulcore_b8[1]), .B(n13329), .Y(dpath_mulcore_ary1_a1_I0_p0_l[39]));
INVX1 mul_U20215(.A(dpath_mulcore_ary1_a1_I0_p0_l[39]), .Y(n7081));
AND2X1 mul_U20216(.A(dpath_mulcore_b10[1]), .B(n13332), .Y(dpath_mulcore_ary1_a1_I0_p2_l[38]));
INVX1 mul_U20217(.A(dpath_mulcore_ary1_a1_I0_p2_l[38]), .Y(n7082));
AND2X1 mul_U20218(.A(dpath_mulcore_b9[1]), .B(n13335), .Y(dpath_mulcore_ary1_a1_I0_p1_l[38]));
INVX1 mul_U20219(.A(dpath_mulcore_ary1_a1_I0_p1_l[38]), .Y(n7083));
AND2X1 mul_U20220(.A(dpath_mulcore_b8[1]), .B(n13338), .Y(dpath_mulcore_ary1_a1_I0_p0_l[38]));
INVX1 mul_U20221(.A(dpath_mulcore_ary1_a1_I0_p0_l[38]), .Y(n7084));
AND2X1 mul_U20222(.A(dpath_mulcore_b10[1]), .B(n13341), .Y(dpath_mulcore_ary1_a1_I0_p2_l[37]));
INVX1 mul_U20223(.A(dpath_mulcore_ary1_a1_I0_p2_l[37]), .Y(n7085));
AND2X1 mul_U20224(.A(dpath_mulcore_b9[1]), .B(n13344), .Y(dpath_mulcore_ary1_a1_I0_p1_l[37]));
INVX1 mul_U20225(.A(dpath_mulcore_ary1_a1_I0_p1_l[37]), .Y(n7086));
AND2X1 mul_U20226(.A(dpath_mulcore_b8[1]), .B(n13347), .Y(dpath_mulcore_ary1_a1_I0_p0_l[37]));
INVX1 mul_U20227(.A(dpath_mulcore_ary1_a1_I0_p0_l[37]), .Y(n7087));
AND2X1 mul_U20228(.A(dpath_mulcore_b10[1]), .B(n13350), .Y(dpath_mulcore_ary1_a1_I0_p2_l[36]));
INVX1 mul_U20229(.A(dpath_mulcore_ary1_a1_I0_p2_l[36]), .Y(n7088));
AND2X1 mul_U20230(.A(dpath_mulcore_b9[1]), .B(n13353), .Y(dpath_mulcore_ary1_a1_I0_p1_l[36]));
INVX1 mul_U20231(.A(dpath_mulcore_ary1_a1_I0_p1_l[36]), .Y(n7089));
AND2X1 mul_U20232(.A(dpath_mulcore_b8[1]), .B(n13356), .Y(dpath_mulcore_ary1_a1_I0_p0_l[36]));
INVX1 mul_U20233(.A(dpath_mulcore_ary1_a1_I0_p0_l[36]), .Y(n7090));
AND2X1 mul_U20234(.A(dpath_mulcore_b10[1]), .B(n13359), .Y(dpath_mulcore_ary1_a1_I0_p2_l[35]));
INVX1 mul_U20235(.A(dpath_mulcore_ary1_a1_I0_p2_l[35]), .Y(n7091));
AND2X1 mul_U20236(.A(dpath_mulcore_b9[1]), .B(n13362), .Y(dpath_mulcore_ary1_a1_I0_p1_l[35]));
INVX1 mul_U20237(.A(dpath_mulcore_ary1_a1_I0_p1_l[35]), .Y(n7092));
AND2X1 mul_U20238(.A(dpath_mulcore_b8[1]), .B(n13365), .Y(dpath_mulcore_ary1_a1_I0_p0_l[35]));
INVX1 mul_U20239(.A(dpath_mulcore_ary1_a1_I0_p0_l[35]), .Y(n7093));
AND2X1 mul_U20240(.A(dpath_mulcore_b10[1]), .B(n13368), .Y(dpath_mulcore_ary1_a1_I0_p2_l[34]));
INVX1 mul_U20241(.A(dpath_mulcore_ary1_a1_I0_p2_l[34]), .Y(n7094));
AND2X1 mul_U20242(.A(dpath_mulcore_b9[1]), .B(n13371), .Y(dpath_mulcore_ary1_a1_I0_p1_l[34]));
INVX1 mul_U20243(.A(dpath_mulcore_ary1_a1_I0_p1_l[34]), .Y(n7095));
AND2X1 mul_U20244(.A(dpath_mulcore_b8[1]), .B(n13374), .Y(dpath_mulcore_ary1_a1_I0_p0_l[34]));
INVX1 mul_U20245(.A(dpath_mulcore_ary1_a1_I0_p0_l[34]), .Y(n7096));
AND2X1 mul_U20246(.A(dpath_mulcore_b10[1]), .B(n13377), .Y(dpath_mulcore_ary1_a1_I0_p2_l[33]));
INVX1 mul_U20247(.A(dpath_mulcore_ary1_a1_I0_p2_l[33]), .Y(n7097));
AND2X1 mul_U20248(.A(dpath_mulcore_b9[1]), .B(n13380), .Y(dpath_mulcore_ary1_a1_I0_p1_l[33]));
INVX1 mul_U20249(.A(dpath_mulcore_ary1_a1_I0_p1_l[33]), .Y(n7098));
AND2X1 mul_U20250(.A(dpath_mulcore_b8[1]), .B(n13383), .Y(dpath_mulcore_ary1_a1_I0_p0_l[33]));
INVX1 mul_U20251(.A(dpath_mulcore_ary1_a1_I0_p0_l[33]), .Y(n7099));
AND2X1 mul_U20252(.A(dpath_mulcore_b10[1]), .B(n13386), .Y(dpath_mulcore_ary1_a1_I0_p2_l[32]));
INVX1 mul_U20253(.A(dpath_mulcore_ary1_a1_I0_p2_l[32]), .Y(n7100));
AND2X1 mul_U20254(.A(dpath_mulcore_b9[1]), .B(n13389), .Y(dpath_mulcore_ary1_a1_I0_p1_l[32]));
INVX1 mul_U20255(.A(dpath_mulcore_ary1_a1_I0_p1_l[32]), .Y(n7101));
AND2X1 mul_U20256(.A(dpath_mulcore_b8[1]), .B(n13392), .Y(dpath_mulcore_ary1_a1_I0_p0_l[32]));
INVX1 mul_U20257(.A(dpath_mulcore_ary1_a1_I0_p0_l[32]), .Y(n7102));
AND2X1 mul_U20258(.A(dpath_mulcore_b10[1]), .B(n13395), .Y(dpath_mulcore_ary1_a1_I0_p2_l[31]));
INVX1 mul_U20259(.A(dpath_mulcore_ary1_a1_I0_p2_l[31]), .Y(n7103));
AND2X1 mul_U20260(.A(dpath_mulcore_b9[1]), .B(n13398), .Y(dpath_mulcore_ary1_a1_I0_p1_l[31]));
INVX1 mul_U20261(.A(dpath_mulcore_ary1_a1_I0_p1_l[31]), .Y(n7104));
AND2X1 mul_U20262(.A(dpath_mulcore_b8[1]), .B(n13401), .Y(dpath_mulcore_ary1_a1_I0_p0_l[31]));
INVX1 mul_U20263(.A(dpath_mulcore_ary1_a1_I0_p0_l[31]), .Y(n7105));
AND2X1 mul_U20264(.A(dpath_mulcore_b10[1]), .B(n13404), .Y(dpath_mulcore_ary1_a1_I0_p2_l[30]));
INVX1 mul_U20265(.A(dpath_mulcore_ary1_a1_I0_p2_l[30]), .Y(n7106));
AND2X1 mul_U20266(.A(dpath_mulcore_b9[1]), .B(n13407), .Y(dpath_mulcore_ary1_a1_I0_p1_l[30]));
INVX1 mul_U20267(.A(dpath_mulcore_ary1_a1_I0_p1_l[30]), .Y(n7107));
AND2X1 mul_U20268(.A(dpath_mulcore_b8[1]), .B(n13410), .Y(dpath_mulcore_ary1_a1_I0_p0_l[30]));
INVX1 mul_U20269(.A(dpath_mulcore_ary1_a1_I0_p0_l[30]), .Y(n7108));
AND2X1 mul_U20270(.A(dpath_mulcore_b10[1]), .B(n13413), .Y(dpath_mulcore_ary1_a1_I0_p2_l[29]));
INVX1 mul_U20271(.A(dpath_mulcore_ary1_a1_I0_p2_l[29]), .Y(n7109));
AND2X1 mul_U20272(.A(dpath_mulcore_b9[1]), .B(n13416), .Y(dpath_mulcore_ary1_a1_I0_p1_l[29]));
INVX1 mul_U20273(.A(dpath_mulcore_ary1_a1_I0_p1_l[29]), .Y(n7110));
AND2X1 mul_U20274(.A(dpath_mulcore_b8[1]), .B(n13419), .Y(dpath_mulcore_ary1_a1_I0_p0_l[29]));
INVX1 mul_U20275(.A(dpath_mulcore_ary1_a1_I0_p0_l[29]), .Y(n7111));
AND2X1 mul_U20276(.A(dpath_mulcore_b10[1]), .B(n13422), .Y(dpath_mulcore_ary1_a1_I0_p2_l[28]));
INVX1 mul_U20277(.A(dpath_mulcore_ary1_a1_I0_p2_l[28]), .Y(n7112));
AND2X1 mul_U20278(.A(dpath_mulcore_b9[1]), .B(n13425), .Y(dpath_mulcore_ary1_a1_I0_p1_l[28]));
INVX1 mul_U20279(.A(dpath_mulcore_ary1_a1_I0_p1_l[28]), .Y(n7113));
AND2X1 mul_U20280(.A(dpath_mulcore_b8[1]), .B(n13428), .Y(dpath_mulcore_ary1_a1_I0_p0_l[28]));
INVX1 mul_U20281(.A(dpath_mulcore_ary1_a1_I0_p0_l[28]), .Y(n7114));
AND2X1 mul_U20282(.A(dpath_mulcore_b10[1]), .B(n13431), .Y(dpath_mulcore_ary1_a1_I0_p2_l[27]));
INVX1 mul_U20283(.A(dpath_mulcore_ary1_a1_I0_p2_l[27]), .Y(n7115));
AND2X1 mul_U20284(.A(dpath_mulcore_b9[1]), .B(n13434), .Y(dpath_mulcore_ary1_a1_I0_p1_l[27]));
INVX1 mul_U20285(.A(dpath_mulcore_ary1_a1_I0_p1_l[27]), .Y(n7116));
AND2X1 mul_U20286(.A(dpath_mulcore_b8[1]), .B(n13437), .Y(dpath_mulcore_ary1_a1_I0_p0_l[27]));
INVX1 mul_U20287(.A(dpath_mulcore_ary1_a1_I0_p0_l[27]), .Y(n7117));
AND2X1 mul_U20288(.A(dpath_mulcore_b10[1]), .B(n13440), .Y(dpath_mulcore_ary1_a1_I0_p2_l[26]));
INVX1 mul_U20289(.A(dpath_mulcore_ary1_a1_I0_p2_l[26]), .Y(n7118));
AND2X1 mul_U20290(.A(dpath_mulcore_b9[1]), .B(n13443), .Y(dpath_mulcore_ary1_a1_I0_p1_l[26]));
INVX1 mul_U20291(.A(dpath_mulcore_ary1_a1_I0_p1_l[26]), .Y(n7119));
AND2X1 mul_U20292(.A(dpath_mulcore_b8[1]), .B(n13446), .Y(dpath_mulcore_ary1_a1_I0_p0_l[26]));
INVX1 mul_U20293(.A(dpath_mulcore_ary1_a1_I0_p0_l[26]), .Y(n7120));
AND2X1 mul_U20294(.A(dpath_mulcore_b10[1]), .B(n13449), .Y(dpath_mulcore_ary1_a1_I0_p2_l[25]));
INVX1 mul_U20295(.A(dpath_mulcore_ary1_a1_I0_p2_l[25]), .Y(n7121));
AND2X1 mul_U20296(.A(dpath_mulcore_b9[1]), .B(n13452), .Y(dpath_mulcore_ary1_a1_I0_p1_l[25]));
INVX1 mul_U20297(.A(dpath_mulcore_ary1_a1_I0_p1_l[25]), .Y(n7122));
AND2X1 mul_U20298(.A(dpath_mulcore_b8[1]), .B(n13455), .Y(dpath_mulcore_ary1_a1_I0_p0_l[25]));
INVX1 mul_U20299(.A(dpath_mulcore_ary1_a1_I0_p0_l[25]), .Y(n7123));
AND2X1 mul_U20300(.A(dpath_mulcore_b10[1]), .B(n13458), .Y(dpath_mulcore_ary1_a1_I0_p2_l[24]));
INVX1 mul_U20301(.A(dpath_mulcore_ary1_a1_I0_p2_l[24]), .Y(n7124));
AND2X1 mul_U20302(.A(dpath_mulcore_b9[1]), .B(n13461), .Y(dpath_mulcore_ary1_a1_I0_p1_l[24]));
INVX1 mul_U20303(.A(dpath_mulcore_ary1_a1_I0_p1_l[24]), .Y(n7125));
AND2X1 mul_U20304(.A(dpath_mulcore_b8[1]), .B(n13464), .Y(dpath_mulcore_ary1_a1_I0_p0_l[24]));
INVX1 mul_U20305(.A(dpath_mulcore_ary1_a1_I0_p0_l[24]), .Y(n7126));
AND2X1 mul_U20306(.A(dpath_mulcore_b10[1]), .B(n13467), .Y(dpath_mulcore_ary1_a1_I0_p2_l[23]));
INVX1 mul_U20307(.A(dpath_mulcore_ary1_a1_I0_p2_l[23]), .Y(n7127));
AND2X1 mul_U20308(.A(dpath_mulcore_b9[1]), .B(n13470), .Y(dpath_mulcore_ary1_a1_I0_p1_l[23]));
INVX1 mul_U20309(.A(dpath_mulcore_ary1_a1_I0_p1_l[23]), .Y(n7128));
AND2X1 mul_U20310(.A(dpath_mulcore_b8[1]), .B(n13473), .Y(dpath_mulcore_ary1_a1_I0_p0_l[23]));
INVX1 mul_U20311(.A(dpath_mulcore_ary1_a1_I0_p0_l[23]), .Y(n7129));
AND2X1 mul_U20312(.A(dpath_mulcore_b10[1]), .B(n13476), .Y(dpath_mulcore_ary1_a1_I0_p2_l[22]));
INVX1 mul_U20313(.A(dpath_mulcore_ary1_a1_I0_p2_l[22]), .Y(n7130));
AND2X1 mul_U20314(.A(dpath_mulcore_b9[1]), .B(n13479), .Y(dpath_mulcore_ary1_a1_I0_p1_l[22]));
INVX1 mul_U20315(.A(dpath_mulcore_ary1_a1_I0_p1_l[22]), .Y(n7131));
AND2X1 mul_U20316(.A(dpath_mulcore_b8[1]), .B(n13482), .Y(dpath_mulcore_ary1_a1_I0_p0_l[22]));
INVX1 mul_U20317(.A(dpath_mulcore_ary1_a1_I0_p0_l[22]), .Y(n7132));
AND2X1 mul_U20318(.A(dpath_mulcore_b10[1]), .B(n13485), .Y(dpath_mulcore_ary1_a1_I0_p2_l[21]));
INVX1 mul_U20319(.A(dpath_mulcore_ary1_a1_I0_p2_l[21]), .Y(n7133));
AND2X1 mul_U20320(.A(dpath_mulcore_b9[1]), .B(n13488), .Y(dpath_mulcore_ary1_a1_I0_p1_l[21]));
INVX1 mul_U20321(.A(dpath_mulcore_ary1_a1_I0_p1_l[21]), .Y(n7134));
AND2X1 mul_U20322(.A(dpath_mulcore_b8[1]), .B(n13491), .Y(dpath_mulcore_ary1_a1_I0_p0_l[21]));
INVX1 mul_U20323(.A(dpath_mulcore_ary1_a1_I0_p0_l[21]), .Y(n7135));
AND2X1 mul_U20324(.A(dpath_mulcore_b10[1]), .B(n13494), .Y(dpath_mulcore_ary1_a1_I0_p2_l[20]));
INVX1 mul_U20325(.A(dpath_mulcore_ary1_a1_I0_p2_l[20]), .Y(n7136));
AND2X1 mul_U20326(.A(dpath_mulcore_b9[1]), .B(n13497), .Y(dpath_mulcore_ary1_a1_I0_p1_l[20]));
INVX1 mul_U20327(.A(dpath_mulcore_ary1_a1_I0_p1_l[20]), .Y(n7137));
AND2X1 mul_U20328(.A(dpath_mulcore_b8[1]), .B(n13500), .Y(dpath_mulcore_ary1_a1_I0_p0_l[20]));
INVX1 mul_U20329(.A(dpath_mulcore_ary1_a1_I0_p0_l[20]), .Y(n7138));
AND2X1 mul_U20330(.A(dpath_mulcore_b10[1]), .B(n13503), .Y(dpath_mulcore_ary1_a1_I0_p2_l[19]));
INVX1 mul_U20331(.A(dpath_mulcore_ary1_a1_I0_p2_l[19]), .Y(n7139));
AND2X1 mul_U20332(.A(dpath_mulcore_b9[1]), .B(n13506), .Y(dpath_mulcore_ary1_a1_I0_p1_l[19]));
INVX1 mul_U20333(.A(dpath_mulcore_ary1_a1_I0_p1_l[19]), .Y(n7140));
AND2X1 mul_U20334(.A(dpath_mulcore_b8[1]), .B(n13509), .Y(dpath_mulcore_ary1_a1_I0_p0_l[19]));
INVX1 mul_U20335(.A(dpath_mulcore_ary1_a1_I0_p0_l[19]), .Y(n7141));
AND2X1 mul_U20336(.A(dpath_mulcore_b10[1]), .B(n13512), .Y(dpath_mulcore_ary1_a1_I0_p2_l[18]));
INVX1 mul_U20337(.A(dpath_mulcore_ary1_a1_I0_p2_l[18]), .Y(n7142));
AND2X1 mul_U20338(.A(dpath_mulcore_b9[1]), .B(n13515), .Y(dpath_mulcore_ary1_a1_I0_p1_l[18]));
INVX1 mul_U20339(.A(dpath_mulcore_ary1_a1_I0_p1_l[18]), .Y(n7143));
AND2X1 mul_U20340(.A(dpath_mulcore_b8[1]), .B(n13518), .Y(dpath_mulcore_ary1_a1_I0_p0_l[18]));
INVX1 mul_U20341(.A(dpath_mulcore_ary1_a1_I0_p0_l[18]), .Y(n7144));
AND2X1 mul_U20342(.A(dpath_mulcore_b10[1]), .B(n13521), .Y(dpath_mulcore_ary1_a1_I0_p2_l[17]));
INVX1 mul_U20343(.A(dpath_mulcore_ary1_a1_I0_p2_l[17]), .Y(n7145));
AND2X1 mul_U20344(.A(dpath_mulcore_b9[1]), .B(n13524), .Y(dpath_mulcore_ary1_a1_I0_p1_l[17]));
INVX1 mul_U20345(.A(dpath_mulcore_ary1_a1_I0_p1_l[17]), .Y(n7146));
AND2X1 mul_U20346(.A(dpath_mulcore_b8[1]), .B(n13527), .Y(dpath_mulcore_ary1_a1_I0_p0_l[17]));
INVX1 mul_U20347(.A(dpath_mulcore_ary1_a1_I0_p0_l[17]), .Y(n7147));
AND2X1 mul_U20348(.A(dpath_mulcore_b10[1]), .B(n13530), .Y(dpath_mulcore_ary1_a1_I0_p2_l[16]));
INVX1 mul_U20349(.A(dpath_mulcore_ary1_a1_I0_p2_l[16]), .Y(n7148));
AND2X1 mul_U20350(.A(dpath_mulcore_b9[1]), .B(n13533), .Y(dpath_mulcore_ary1_a1_I0_p1_l[16]));
INVX1 mul_U20351(.A(dpath_mulcore_ary1_a1_I0_p1_l[16]), .Y(n7149));
AND2X1 mul_U20352(.A(dpath_mulcore_b8[1]), .B(n13536), .Y(dpath_mulcore_ary1_a1_I0_p0_l[16]));
INVX1 mul_U20353(.A(dpath_mulcore_ary1_a1_I0_p0_l[16]), .Y(n7150));
AND2X1 mul_U20354(.A(dpath_mulcore_b10[1]), .B(n13539), .Y(dpath_mulcore_ary1_a1_I0_p2_l[15]));
INVX1 mul_U20355(.A(dpath_mulcore_ary1_a1_I0_p2_l[15]), .Y(n7151));
AND2X1 mul_U20356(.A(dpath_mulcore_b9[1]), .B(n13542), .Y(dpath_mulcore_ary1_a1_I0_p1_l[15]));
INVX1 mul_U20357(.A(dpath_mulcore_ary1_a1_I0_p1_l[15]), .Y(n7152));
AND2X1 mul_U20358(.A(dpath_mulcore_b8[1]), .B(n13545), .Y(dpath_mulcore_ary1_a1_I0_p0_l[15]));
INVX1 mul_U20359(.A(dpath_mulcore_ary1_a1_I0_p0_l[15]), .Y(n7153));
AND2X1 mul_U20360(.A(dpath_mulcore_b10[1]), .B(n13548), .Y(dpath_mulcore_ary1_a1_I0_p2_l[14]));
INVX1 mul_U20361(.A(dpath_mulcore_ary1_a1_I0_p2_l[14]), .Y(n7154));
AND2X1 mul_U20362(.A(dpath_mulcore_b9[1]), .B(n13551), .Y(dpath_mulcore_ary1_a1_I0_p1_l[14]));
INVX1 mul_U20363(.A(dpath_mulcore_ary1_a1_I0_p1_l[14]), .Y(n7155));
AND2X1 mul_U20364(.A(dpath_mulcore_b8[1]), .B(n13554), .Y(dpath_mulcore_ary1_a1_I0_p0_l[14]));
INVX1 mul_U20365(.A(dpath_mulcore_ary1_a1_I0_p0_l[14]), .Y(n7156));
AND2X1 mul_U20366(.A(dpath_mulcore_b10[1]), .B(n13557), .Y(dpath_mulcore_ary1_a1_I0_p2_l[13]));
INVX1 mul_U20367(.A(dpath_mulcore_ary1_a1_I0_p2_l[13]), .Y(n7157));
AND2X1 mul_U20368(.A(dpath_mulcore_b9[1]), .B(n13560), .Y(dpath_mulcore_ary1_a1_I0_p1_l[13]));
INVX1 mul_U20369(.A(dpath_mulcore_ary1_a1_I0_p1_l[13]), .Y(n7158));
AND2X1 mul_U20370(.A(dpath_mulcore_b8[1]), .B(n13563), .Y(dpath_mulcore_ary1_a1_I0_p0_l[13]));
INVX1 mul_U20371(.A(dpath_mulcore_ary1_a1_I0_p0_l[13]), .Y(n7159));
AND2X1 mul_U20372(.A(dpath_mulcore_b10[1]), .B(n13566), .Y(dpath_mulcore_ary1_a1_I0_p2_l[12]));
INVX1 mul_U20373(.A(dpath_mulcore_ary1_a1_I0_p2_l[12]), .Y(n7160));
AND2X1 mul_U20374(.A(dpath_mulcore_b9[1]), .B(n13569), .Y(dpath_mulcore_ary1_a1_I0_p1_l[12]));
INVX1 mul_U20375(.A(dpath_mulcore_ary1_a1_I0_p1_l[12]), .Y(n7161));
AND2X1 mul_U20376(.A(dpath_mulcore_b8[1]), .B(n13572), .Y(dpath_mulcore_ary1_a1_I0_p0_l[12]));
INVX1 mul_U20377(.A(dpath_mulcore_ary1_a1_I0_p0_l[12]), .Y(n7162));
AND2X1 mul_U20378(.A(dpath_mulcore_b10[1]), .B(n13575), .Y(dpath_mulcore_ary1_a1_I0_p2_l[11]));
INVX1 mul_U20379(.A(dpath_mulcore_ary1_a1_I0_p2_l[11]), .Y(n7163));
AND2X1 mul_U20380(.A(dpath_mulcore_b9[1]), .B(n13578), .Y(dpath_mulcore_ary1_a1_I0_p1_l[11]));
INVX1 mul_U20381(.A(dpath_mulcore_ary1_a1_I0_p1_l[11]), .Y(n7164));
AND2X1 mul_U20382(.A(dpath_mulcore_b8[1]), .B(n13581), .Y(dpath_mulcore_ary1_a1_I0_p0_l[11]));
INVX1 mul_U20383(.A(dpath_mulcore_ary1_a1_I0_p0_l[11]), .Y(n7165));
AND2X1 mul_U20384(.A(dpath_mulcore_b10[1]), .B(n13584), .Y(dpath_mulcore_ary1_a1_I0_p2_l[10]));
INVX1 mul_U20385(.A(dpath_mulcore_ary1_a1_I0_p2_l[10]), .Y(n7166));
AND2X1 mul_U20386(.A(dpath_mulcore_b9[1]), .B(n13587), .Y(dpath_mulcore_ary1_a1_I0_p1_l[10]));
INVX1 mul_U20387(.A(dpath_mulcore_ary1_a1_I0_p1_l[10]), .Y(n7167));
AND2X1 mul_U20388(.A(dpath_mulcore_b8[1]), .B(n13590), .Y(dpath_mulcore_ary1_a1_I0_p0_l[10]));
INVX1 mul_U20389(.A(dpath_mulcore_ary1_a1_I0_p0_l[10]), .Y(n7168));
AND2X1 mul_U20390(.A(dpath_mulcore_b10[1]), .B(n13593), .Y(dpath_mulcore_ary1_a1_I0_p2_l[9]));
INVX1 mul_U20391(.A(dpath_mulcore_ary1_a1_I0_p2_l[9]), .Y(n7169));
AND2X1 mul_U20392(.A(dpath_mulcore_b9[1]), .B(n13596), .Y(dpath_mulcore_ary1_a1_I0_p1_l[9]));
INVX1 mul_U20393(.A(dpath_mulcore_ary1_a1_I0_p1_l[9]), .Y(n7170));
AND2X1 mul_U20394(.A(dpath_mulcore_b8[1]), .B(n13599), .Y(dpath_mulcore_ary1_a1_I0_p0_l[9]));
INVX1 mul_U20395(.A(dpath_mulcore_ary1_a1_I0_p0_l[9]), .Y(n7171));
AND2X1 mul_U20396(.A(dpath_mulcore_b10[1]), .B(n13602), .Y(dpath_mulcore_ary1_a1_I0_p2_l[8]));
INVX1 mul_U20397(.A(dpath_mulcore_ary1_a1_I0_p2_l[8]), .Y(n7172));
AND2X1 mul_U20398(.A(dpath_mulcore_b9[1]), .B(n13605), .Y(dpath_mulcore_ary1_a1_I0_p1_l[8]));
INVX1 mul_U20399(.A(dpath_mulcore_ary1_a1_I0_p1_l[8]), .Y(n7173));
AND2X1 mul_U20400(.A(dpath_mulcore_b8[1]), .B(n13608), .Y(dpath_mulcore_ary1_a1_I0_p0_l[8]));
INVX1 mul_U20401(.A(dpath_mulcore_ary1_a1_I0_p0_l[8]), .Y(n7174));
AND2X1 mul_U20402(.A(dpath_mulcore_b10[1]), .B(n13611), .Y(dpath_mulcore_ary1_a1_I0_p2_l[7]));
INVX1 mul_U20403(.A(dpath_mulcore_ary1_a1_I0_p2_l[7]), .Y(n7175));
AND2X1 mul_U20404(.A(dpath_mulcore_b9[1]), .B(n13614), .Y(dpath_mulcore_ary1_a1_I0_p1_l[7]));
INVX1 mul_U20405(.A(dpath_mulcore_ary1_a1_I0_p1_l[7]), .Y(n7176));
AND2X1 mul_U20406(.A(dpath_mulcore_b8[1]), .B(n13617), .Y(dpath_mulcore_ary1_a1_I0_p0_l[7]));
INVX1 mul_U20407(.A(dpath_mulcore_ary1_a1_I0_p0_l[7]), .Y(n7177));
AND2X1 mul_U20408(.A(dpath_mulcore_b10[1]), .B(n13620), .Y(dpath_mulcore_ary1_a1_I0_p2_l[6]));
INVX1 mul_U20409(.A(dpath_mulcore_ary1_a1_I0_p2_l[6]), .Y(n7178));
AND2X1 mul_U20410(.A(dpath_mulcore_b9[1]), .B(n13623), .Y(dpath_mulcore_ary1_a1_I0_p1_l[6]));
INVX1 mul_U20411(.A(dpath_mulcore_ary1_a1_I0_p1_l[6]), .Y(n7179));
AND2X1 mul_U20412(.A(dpath_mulcore_b8[1]), .B(n13626), .Y(dpath_mulcore_ary1_a1_I0_p0_l[6]));
INVX1 mul_U20413(.A(dpath_mulcore_ary1_a1_I0_p0_l[6]), .Y(n7180));
AND2X1 mul_U20414(.A(dpath_mulcore_b10[1]), .B(n13629), .Y(dpath_mulcore_ary1_a1_I0_p2_l[5]));
INVX1 mul_U20415(.A(dpath_mulcore_ary1_a1_I0_p2_l[5]), .Y(n7181));
AND2X1 mul_U20416(.A(dpath_mulcore_b9[1]), .B(n13632), .Y(dpath_mulcore_ary1_a1_I0_p1_l[5]));
INVX1 mul_U20417(.A(dpath_mulcore_ary1_a1_I0_p1_l[5]), .Y(n7182));
AND2X1 mul_U20418(.A(dpath_mulcore_b8[1]), .B(n13635), .Y(dpath_mulcore_ary1_a1_I0_p0_l[5]));
INVX1 mul_U20419(.A(dpath_mulcore_ary1_a1_I0_p0_l[5]), .Y(n7183));
AND2X1 mul_U20420(.A(dpath_mulcore_b10[1]), .B(n13637), .Y(dpath_mulcore_ary1_a1_I0_p2_l[4]));
INVX1 mul_U20421(.A(dpath_mulcore_ary1_a1_I0_p2_l[4]), .Y(n7184));
AND2X1 mul_U20422(.A(dpath_mulcore_b9[1]), .B(n13640), .Y(dpath_mulcore_ary1_a1_I0_p1_l[4]));
INVX1 mul_U20423(.A(dpath_mulcore_ary1_a1_I0_p1_l[4]), .Y(n7185));
AND2X1 mul_U20424(.A(dpath_mulcore_b8[1]), .B(n13643), .Y(dpath_mulcore_ary1_a1_I0_p0_l[4]));
INVX1 mul_U20425(.A(dpath_mulcore_ary1_a1_I0_p0_l[4]), .Y(n7186));
AND2X1 mul_U20426(.A(dpath_mulcore_b8[1]), .B(n13646), .Y(dpath_mulcore_ary1_a1_I0_p0_l[3]));
INVX1 mul_U20427(.A(dpath_mulcore_ary1_a1_I0_p0_l[3]), .Y(n7187));
AND2X1 mul_U20428(.A(dpath_mulcore_b9[1]), .B(n13649), .Y(dpath_mulcore_ary1_a1_I0_p1_l[3]));
INVX1 mul_U20429(.A(dpath_mulcore_ary1_a1_I0_p1_l[3]), .Y(n7188));
AND2X1 mul_U20430(.A(dpath_mulcore_b8[1]), .B(n13652), .Y(dpath_mulcore_ary1_a1_I0_I0_p0_l_2));
INVX1 mul_U20431(.A(dpath_mulcore_ary1_a1_I0_I0_p0_l_2), .Y(n7189));
AND2X1 mul_U20432(.A(dpath_mulcore_b8[1]), .B(n13655), .Y(dpath_mulcore_ary1_a1_I0_I0_p0_l_1));
INVX1 mul_U20433(.A(dpath_mulcore_ary1_a1_I0_I0_p0_l_1), .Y(n7190));
AND2X1 mul_U20434(.A(dpath_mulcore_b8[1]), .B(n13657), .Y(dpath_mulcore_ary1_a1_I0_I0_p0_l_0));
INVX1 mul_U20435(.A(dpath_mulcore_ary1_a1_I0_I0_p0_l_0), .Y(n7191));
AND2X1 mul_U20436(.A(dpath_mulcore_b9[1]), .B(n13659), .Y(dpath_mulcore_ary1_a1_I0_I0_p1_l_2));
INVX1 mul_U20437(.A(dpath_mulcore_ary1_a1_I0_I0_p1_l_2), .Y(n7192));
AND2X1 mul_U20438(.A(dpath_n980), .B(acc_imm), .Y(dpath_n979));
INVX1 mul_U20439(.A(dpath_n979), .Y(n7193));
AND2X1 mul_U20440(.A(n9214), .B(dpath_n980), .Y(dpath_n984));
INVX1 mul_U20441(.A(dpath_n984), .Y(n7194));
OR2X1 mul_U20442(.A(se), .B(acc_reg_rst), .Y(dpath_accum_n3));
INVX1 mul_U20443(.A(dpath_accum_n3), .Y(n7195));
OR2X1 mul_U20444(.A(n9215), .B(byp_imm), .Y(dpath_n144));
INVX1 mul_U20445(.A(dpath_n144), .Y(n7196));
INVX1 mul_U20446(.A(dpath_n657), .Y(n7197));
INVX1 mul_U20447(.A(control_n7), .Y(n7198));
INVX1 mul_U20448(.A(n7198), .Y(n9775));
OR2X1 mul_U20449(.A(n9815), .B(n9774), .Y(n18339));
INVX1 mul_U20450(.A(n18339), .Y(mul_spu_ack));
INVX1 mul_U20451(.A(dpath_mulcore_ary1_a0_c0[12]), .Y(n7200));
INVX1 mul_U20452(.A(dpath_mulcore_ary1_a0_c0[11]), .Y(n7201));
INVX1 mul_U20453(.A(dpath_mulcore_ary1_a0_c0[10]), .Y(n7202));
INVX1 mul_U20454(.A(dpath_mulcore_ary1_a0_c0[9]), .Y(n7203));
INVX1 mul_U20455(.A(dpath_mulcore_ary1_a1_c0[12]), .Y(n7204));
INVX1 mul_U20456(.A(dpath_mulcore_ary1_a1_c0[11]), .Y(n7205));
INVX1 mul_U20457(.A(dpath_mulcore_ary1_a1_c0[10]), .Y(n7206));
INVX1 mul_U20458(.A(dpath_mulcore_ary1_a1_c0[9]), .Y(n7207));
INVX1 mul_U20459(.A(dpath_mulcore_ary1_a1_c2[65]), .Y(n7208));
INVX1 mul_U20460(.A(dpath_mulcore_ary1_a1_c2[66]), .Y(n7209));
INVX1 mul_U20461(.A(dpath_mulcore_array2_c1[3]), .Y(n7210));
INVX1 mul_U20462(.A(dpath_mulcore_array2_c1[2]), .Y(n7211));
INVX1 mul_U20463(.A(dpath_mulcore_array2_c1[1]), .Y(n7212));
INVX1 mul_U20464(.A(dpath_mulcore_array2_c2[80]), .Y(n7213));
INVX1 mul_U20465(.A(dpath_mulcore_array2_c2[79]), .Y(n7214));
INVX1 mul_U20466(.A(dpath_mulcore_array2_c2[78]), .Y(n7215));
INVX1 mul_U20467(.A(dpath_mulcore_array2_c2[77]), .Y(n7216));
INVX1 mul_U20468(.A(dpath_mulcore_array2_c2[76]), .Y(n7217));
INVX1 mul_U20469(.A(dpath_mulcore_array2_c2[75]), .Y(n7218));
INVX1 mul_U20470(.A(dpath_mulcore_array2_c2[74]), .Y(n7219));
INVX1 mul_U20471(.A(dpath_mulcore_array2_c2[73]), .Y(n7220));
INVX1 mul_U20472(.A(dpath_mulcore_array2_c2[72]), .Y(n7221));
INVX1 mul_U20473(.A(dpath_mulcore_array2_c2[71]), .Y(n7222));
INVX1 mul_U20474(.A(dpath_mulcore_array2_c2[70]), .Y(n7223));
INVX1 mul_U20475(.A(dpath_mulcore_array2_c2[69]), .Y(n7224));
INVX1 mul_U20476(.A(dpath_mulcore_array2_c2[68]), .Y(n7225));
INVX1 mul_U20477(.A(dpath_mulcore_array2_c1[0]), .Y(n7226));
INVX1 mul_U20478(.A(dpath_mulcore_ary1_a0_co[70]), .Y(n7227));
INVX1 mul_U20479(.A(dpath_mulcore_ary1_a0_co[69]), .Y(n7228));
INVX1 mul_U20480(.A(dpath_mulcore_ary1_a0_co[68]), .Y(n7229));
INVX1 mul_U20481(.A(dpath_mulcore_ary1_a0_co[67]), .Y(n7230));
INVX1 mul_U20482(.A(dpath_mulcore_ary1_a0_co[66]), .Y(n7231));
INVX1 mul_U20483(.A(dpath_mulcore_ary1_a0_co[65]), .Y(n7232));
INVX1 mul_U20484(.A(dpath_mulcore_ary1_a0_co[64]), .Y(n7233));
INVX1 mul_U20485(.A(dpath_mulcore_ary1_a0_co[63]), .Y(n7234));
INVX1 mul_U20486(.A(dpath_mulcore_ary1_a0_co[62]), .Y(n7235));
INVX1 mul_U20487(.A(dpath_mulcore_ary1_a0_co[61]), .Y(n7236));
INVX1 mul_U20488(.A(dpath_mulcore_ary1_a0_co[60]), .Y(n7237));
INVX1 mul_U20489(.A(dpath_mulcore_ary1_a0_co[59]), .Y(n7238));
INVX1 mul_U20490(.A(dpath_mulcore_ary1_a0_co[58]), .Y(n7239));
INVX1 mul_U20491(.A(dpath_mulcore_ary1_a0_co[57]), .Y(n7240));
INVX1 mul_U20492(.A(dpath_mulcore_ary1_a0_co[56]), .Y(n7241));
INVX1 mul_U20493(.A(dpath_mulcore_ary1_a0_co[55]), .Y(n7242));
INVX1 mul_U20494(.A(dpath_mulcore_ary1_a0_co[54]), .Y(n7243));
INVX1 mul_U20495(.A(dpath_mulcore_ary1_a0_co[53]), .Y(n7244));
INVX1 mul_U20496(.A(dpath_mulcore_ary1_a0_co[52]), .Y(n7245));
INVX1 mul_U20497(.A(dpath_mulcore_ary1_a0_co[51]), .Y(n7246));
INVX1 mul_U20498(.A(dpath_mulcore_ary1_a0_co[50]), .Y(n7247));
INVX1 mul_U20499(.A(dpath_mulcore_ary1_a0_co[49]), .Y(n7248));
INVX1 mul_U20500(.A(dpath_mulcore_ary1_a0_co[48]), .Y(n7249));
INVX1 mul_U20501(.A(dpath_mulcore_ary1_a0_co[47]), .Y(n7250));
INVX1 mul_U20502(.A(dpath_mulcore_ary1_a0_co[46]), .Y(n7251));
INVX1 mul_U20503(.A(dpath_mulcore_ary1_a0_co[45]), .Y(n7252));
INVX1 mul_U20504(.A(dpath_mulcore_ary1_a0_co[44]), .Y(n7253));
INVX1 mul_U20505(.A(dpath_mulcore_ary1_a0_co[43]), .Y(n7254));
INVX1 mul_U20506(.A(dpath_mulcore_ary1_a0_co[42]), .Y(n7255));
INVX1 mul_U20507(.A(dpath_mulcore_ary1_a0_co[41]), .Y(n7256));
INVX1 mul_U20508(.A(dpath_mulcore_ary1_a0_co[40]), .Y(n7257));
INVX1 mul_U20509(.A(dpath_mulcore_ary1_a0_co[39]), .Y(n7258));
INVX1 mul_U20510(.A(dpath_mulcore_ary1_a0_co[38]), .Y(n7259));
INVX1 mul_U20511(.A(dpath_mulcore_ary1_a0_co[37]), .Y(n7260));
INVX1 mul_U20512(.A(dpath_mulcore_ary1_a0_co[36]), .Y(n7261));
INVX1 mul_U20513(.A(dpath_mulcore_ary1_a0_co[35]), .Y(n7262));
INVX1 mul_U20514(.A(dpath_mulcore_ary1_a0_co[34]), .Y(n7263));
INVX1 mul_U20515(.A(dpath_mulcore_ary1_a0_co[33]), .Y(n7264));
INVX1 mul_U20516(.A(dpath_mulcore_ary1_a0_co[32]), .Y(n7265));
INVX1 mul_U20517(.A(dpath_mulcore_ary1_a0_co[31]), .Y(n7266));
INVX1 mul_U20518(.A(dpath_mulcore_ary1_a0_co[30]), .Y(n7267));
INVX1 mul_U20519(.A(dpath_mulcore_ary1_a0_co[29]), .Y(n7268));
INVX1 mul_U20520(.A(dpath_mulcore_ary1_a0_co[28]), .Y(n7269));
INVX1 mul_U20521(.A(dpath_mulcore_ary1_a0_co[27]), .Y(n7270));
INVX1 mul_U20522(.A(dpath_mulcore_ary1_a0_co[26]), .Y(n7271));
INVX1 mul_U20523(.A(dpath_mulcore_ary1_a0_co[25]), .Y(n7272));
INVX1 mul_U20524(.A(dpath_mulcore_ary1_a0_co[24]), .Y(n7273));
INVX1 mul_U20525(.A(dpath_mulcore_ary1_a0_co[23]), .Y(n7274));
INVX1 mul_U20526(.A(dpath_mulcore_ary1_a0_co[22]), .Y(n7275));
INVX1 mul_U20527(.A(dpath_mulcore_ary1_a0_co[21]), .Y(n7276));
INVX1 mul_U20528(.A(dpath_mulcore_ary1_a0_co[20]), .Y(n7277));
INVX1 mul_U20529(.A(dpath_mulcore_ary1_a0_co[19]), .Y(n7278));
INVX1 mul_U20530(.A(dpath_mulcore_ary1_a0_co[18]), .Y(n7279));
INVX1 mul_U20531(.A(dpath_mulcore_ary1_a0_co[17]), .Y(n7280));
INVX1 mul_U20532(.A(dpath_mulcore_ary1_a0_co[16]), .Y(n7281));
INVX1 mul_U20533(.A(dpath_mulcore_ary1_a0_co[15]), .Y(n7282));
INVX1 mul_U20534(.A(dpath_mulcore_ary1_a0_co[14]), .Y(n7283));
INVX1 mul_U20535(.A(dpath_mulcore_ary1_a0_co[13]), .Y(n7284));
INVX1 mul_U20536(.A(dpath_mulcore_ary1_a0_co[12]), .Y(n7285));
INVX1 mul_U20537(.A(dpath_mulcore_ary1_a0_co[11]), .Y(n7286));
INVX1 mul_U20538(.A(dpath_mulcore_ary1_a1_co[71]), .Y(n7287));
INVX1 mul_U20539(.A(dpath_mulcore_ary1_a1_co[70]), .Y(n7288));
INVX1 mul_U20540(.A(dpath_mulcore_ary1_a1_co[69]), .Y(n7289));
INVX1 mul_U20541(.A(dpath_mulcore_ary1_a1_co[68]), .Y(n7290));
INVX1 mul_U20542(.A(dpath_mulcore_ary1_a1_co[67]), .Y(n7291));
INVX1 mul_U20543(.A(dpath_mulcore_ary1_a1_co[66]), .Y(n7292));
INVX1 mul_U20544(.A(dpath_mulcore_ary1_a1_co[65]), .Y(n7293));
INVX1 mul_U20545(.A(dpath_mulcore_ary1_a1_co[64]), .Y(n7294));
INVX1 mul_U20546(.A(dpath_mulcore_ary1_a1_co[63]), .Y(n7295));
INVX1 mul_U20547(.A(dpath_mulcore_ary1_a1_co[62]), .Y(n7296));
INVX1 mul_U20548(.A(dpath_mulcore_ary1_a1_co[61]), .Y(n7297));
INVX1 mul_U20549(.A(dpath_mulcore_ary1_a1_co[60]), .Y(n7298));
INVX1 mul_U20550(.A(dpath_mulcore_ary1_a1_co[59]), .Y(n7299));
INVX1 mul_U20551(.A(dpath_mulcore_ary1_a1_co[58]), .Y(n7300));
INVX1 mul_U20552(.A(dpath_mulcore_ary1_a1_co[57]), .Y(n7301));
INVX1 mul_U20553(.A(dpath_mulcore_ary1_a1_co[56]), .Y(n7302));
INVX1 mul_U20554(.A(dpath_mulcore_ary1_a1_co[55]), .Y(n7303));
INVX1 mul_U20555(.A(dpath_mulcore_ary1_a1_co[54]), .Y(n7304));
INVX1 mul_U20556(.A(dpath_mulcore_ary1_a1_co[53]), .Y(n7305));
INVX1 mul_U20557(.A(dpath_mulcore_ary1_a1_co[52]), .Y(n7306));
INVX1 mul_U20558(.A(dpath_mulcore_ary1_a1_co[51]), .Y(n7307));
INVX1 mul_U20559(.A(dpath_mulcore_ary1_a1_co[50]), .Y(n7308));
INVX1 mul_U20560(.A(dpath_mulcore_ary1_a1_co[49]), .Y(n7309));
INVX1 mul_U20561(.A(dpath_mulcore_ary1_a1_co[48]), .Y(n7310));
INVX1 mul_U20562(.A(dpath_mulcore_ary1_a1_co[47]), .Y(n7311));
INVX1 mul_U20563(.A(dpath_mulcore_ary1_a1_co[46]), .Y(n7312));
INVX1 mul_U20564(.A(dpath_mulcore_ary1_a1_co[45]), .Y(n7313));
INVX1 mul_U20565(.A(dpath_mulcore_ary1_a1_co[44]), .Y(n7314));
INVX1 mul_U20566(.A(dpath_mulcore_ary1_a1_co[43]), .Y(n7315));
INVX1 mul_U20567(.A(dpath_mulcore_ary1_a1_co[42]), .Y(n7316));
INVX1 mul_U20568(.A(dpath_mulcore_ary1_a1_co[41]), .Y(n7317));
INVX1 mul_U20569(.A(dpath_mulcore_ary1_a1_co[40]), .Y(n7318));
INVX1 mul_U20570(.A(dpath_mulcore_ary1_a1_co[39]), .Y(n7319));
INVX1 mul_U20571(.A(dpath_mulcore_ary1_a1_co[38]), .Y(n7320));
INVX1 mul_U20572(.A(dpath_mulcore_ary1_a1_co[37]), .Y(n7321));
INVX1 mul_U20573(.A(dpath_mulcore_ary1_a1_co[36]), .Y(n7322));
INVX1 mul_U20574(.A(dpath_mulcore_ary1_a1_co[35]), .Y(n7323));
INVX1 mul_U20575(.A(dpath_mulcore_ary1_a1_co[34]), .Y(n7324));
INVX1 mul_U20576(.A(dpath_mulcore_ary1_a1_co[33]), .Y(n7325));
INVX1 mul_U20577(.A(dpath_mulcore_ary1_a1_co[32]), .Y(n7326));
INVX1 mul_U20578(.A(dpath_mulcore_ary1_a1_co[31]), .Y(n7327));
INVX1 mul_U20579(.A(dpath_mulcore_ary1_a1_co[30]), .Y(n7328));
INVX1 mul_U20580(.A(dpath_mulcore_ary1_a1_co[29]), .Y(n7329));
INVX1 mul_U20581(.A(dpath_mulcore_ary1_a1_co[28]), .Y(n7330));
INVX1 mul_U20582(.A(dpath_mulcore_ary1_a1_co[27]), .Y(n7331));
INVX1 mul_U20583(.A(dpath_mulcore_ary1_a1_co[26]), .Y(n7332));
INVX1 mul_U20584(.A(dpath_mulcore_ary1_a1_co[25]), .Y(n7333));
INVX1 mul_U20585(.A(dpath_mulcore_ary1_a1_co[24]), .Y(n7334));
INVX1 mul_U20586(.A(dpath_mulcore_ary1_a1_co[23]), .Y(n7335));
INVX1 mul_U20587(.A(dpath_mulcore_ary1_a1_co[22]), .Y(n7336));
INVX1 mul_U20588(.A(dpath_mulcore_ary1_a1_co[21]), .Y(n7337));
INVX1 mul_U20589(.A(dpath_mulcore_ary1_a1_co[20]), .Y(n7338));
INVX1 mul_U20590(.A(dpath_mulcore_ary1_a1_co[19]), .Y(n7339));
INVX1 mul_U20591(.A(dpath_mulcore_ary1_a1_co[18]), .Y(n7340));
INVX1 mul_U20592(.A(dpath_mulcore_ary1_a1_co[17]), .Y(n7341));
INVX1 mul_U20593(.A(dpath_mulcore_ary1_a1_co[16]), .Y(n7342));
INVX1 mul_U20594(.A(dpath_mulcore_ary1_a1_co[15]), .Y(n7343));
INVX1 mul_U20595(.A(dpath_mulcore_ary1_a1_co[14]), .Y(n7344));
INVX1 mul_U20596(.A(dpath_mulcore_ary1_a1_co[13]), .Y(n7345));
INVX1 mul_U20597(.A(dpath_mulcore_ary1_a1_co[12]), .Y(n7346));
INVX1 mul_U20598(.A(dpath_mulcore_ary1_a1_co[11]), .Y(n7347));
INVX1 mul_U20599(.A(dpath_mulcore_array2_co[66]), .Y(n7348));
INVX1 mul_U20600(.A(dpath_mulcore_array2_co[65]), .Y(n7349));
INVX1 mul_U20601(.A(dpath_mulcore_array2_co[64]), .Y(n7350));
INVX1 mul_U20602(.A(dpath_mulcore_array2_co[63]), .Y(n7351));
INVX1 mul_U20603(.A(dpath_mulcore_array2_co[62]), .Y(n7352));
INVX1 mul_U20604(.A(dpath_mulcore_array2_co[61]), .Y(n7353));
INVX1 mul_U20605(.A(dpath_mulcore_array2_co[60]), .Y(n7354));
INVX1 mul_U20606(.A(dpath_mulcore_array2_co[59]), .Y(n7355));
INVX1 mul_U20607(.A(dpath_mulcore_array2_co[58]), .Y(n7356));
INVX1 mul_U20608(.A(dpath_mulcore_array2_co[57]), .Y(n7357));
INVX1 mul_U20609(.A(dpath_mulcore_array2_co[56]), .Y(n7358));
INVX1 mul_U20610(.A(dpath_mulcore_array2_co[55]), .Y(n7359));
INVX1 mul_U20611(.A(dpath_mulcore_array2_co[54]), .Y(n7360));
INVX1 mul_U20612(.A(dpath_mulcore_array2_co[53]), .Y(n7361));
INVX1 mul_U20613(.A(dpath_mulcore_array2_co[52]), .Y(n7362));
INVX1 mul_U20614(.A(dpath_mulcore_array2_co[51]), .Y(n7363));
INVX1 mul_U20615(.A(dpath_mulcore_array2_co[50]), .Y(n7364));
INVX1 mul_U20616(.A(dpath_mulcore_array2_co[49]), .Y(n7365));
INVX1 mul_U20617(.A(dpath_mulcore_array2_co[48]), .Y(n7366));
INVX1 mul_U20618(.A(dpath_mulcore_array2_co[47]), .Y(n7367));
INVX1 mul_U20619(.A(dpath_mulcore_array2_co[46]), .Y(n7368));
INVX1 mul_U20620(.A(dpath_mulcore_array2_co[45]), .Y(n7369));
INVX1 mul_U20621(.A(dpath_mulcore_array2_co[44]), .Y(n7370));
INVX1 mul_U20622(.A(dpath_mulcore_array2_co[43]), .Y(n7371));
INVX1 mul_U20623(.A(dpath_mulcore_array2_co[42]), .Y(n7372));
INVX1 mul_U20624(.A(dpath_mulcore_array2_co[41]), .Y(n7373));
INVX1 mul_U20625(.A(dpath_mulcore_array2_co[40]), .Y(n7374));
INVX1 mul_U20626(.A(dpath_mulcore_array2_co[39]), .Y(n7375));
INVX1 mul_U20627(.A(dpath_mulcore_array2_co[38]), .Y(n7376));
INVX1 mul_U20628(.A(dpath_mulcore_array2_co[37]), .Y(n7377));
INVX1 mul_U20629(.A(dpath_mulcore_array2_co[36]), .Y(n7378));
INVX1 mul_U20630(.A(dpath_mulcore_array2_co[35]), .Y(n7379));
INVX1 mul_U20631(.A(dpath_mulcore_array2_co[34]), .Y(n7380));
INVX1 mul_U20632(.A(dpath_mulcore_array2_co[33]), .Y(n7381));
INVX1 mul_U20633(.A(dpath_mulcore_array2_co[32]), .Y(n7382));
INVX1 mul_U20634(.A(dpath_mulcore_array2_co[31]), .Y(n7383));
INVX1 mul_U20635(.A(dpath_mulcore_array2_co[30]), .Y(n7384));
INVX1 mul_U20636(.A(dpath_mulcore_array2_co[29]), .Y(n7385));
INVX1 mul_U20637(.A(dpath_mulcore_array2_co[28]), .Y(n7386));
INVX1 mul_U20638(.A(dpath_mulcore_array2_co[27]), .Y(n7387));
INVX1 mul_U20639(.A(dpath_mulcore_array2_co[26]), .Y(n7388));
INVX1 mul_U20640(.A(dpath_mulcore_array2_co[25]), .Y(n7389));
INVX1 mul_U20641(.A(dpath_mulcore_array2_co[24]), .Y(n7390));
INVX1 mul_U20642(.A(dpath_mulcore_array2_co[23]), .Y(n7391));
INVX1 mul_U20643(.A(dpath_mulcore_array2_co[22]), .Y(n7392));
INVX1 mul_U20644(.A(dpath_mulcore_array2_co[21]), .Y(n7393));
INVX1 mul_U20645(.A(dpath_mulcore_array2_co[20]), .Y(n7394));
INVX1 mul_U20646(.A(dpath_mulcore_ary1_a0_co[71]), .Y(n7395));
INVX1 mul_U20647(.A(dpath_mulcore_ary1_a0_I2_I0_p0_1), .Y(n7396));
INVX1 mul_U20648(.A(dpath_mulcore_ary1_a0_I1_I0_p0_1), .Y(n7397));
INVX1 mul_U20649(.A(dpath_mulcore_ary1_a0_I0_I0_p0_1), .Y(n7398));
INVX1 mul_U20650(.A(dpath_mulcore_ary1_a1_I2_I0_p0_1), .Y(n7399));
INVX1 mul_U20651(.A(dpath_mulcore_ary1_a1_I1_I0_p0_1), .Y(n7400));
INVX1 mul_U20652(.A(dpath_mulcore_ary1_a1_I0_I0_p0_1), .Y(n7401));
INVX1 mul_U20653(.A(dpath_mulcore_ary1_a0_I1_I0_b0n_0), .Y(n7402));
INVX1 mul_U20654(.A(dpath_mulcore_ary1_a0_I0_I0_b0n_0), .Y(n7403));
INVX1 mul_U20655(.A(dpath_mulcore_ary1_a1_I2_I0_b0n_0), .Y(n7404));
INVX1 mul_U20656(.A(dpath_mulcore_ary1_a1_I1_I0_b0n_0), .Y(n7405));
INVX1 mul_U20657(.A(dpath_mulcore_ary1_a1_I0_I0_b0n_0), .Y(n7406));
INVX1 mul_U20658(.A(dpath_mulcore_array2_ain[0]), .Y(n7407));
INVX1 mul_U20659(.A(dpath_mulcore_ary1_a0_c_1[3]), .Y(n7408));
INVX1 mul_U20660(.A(dpath_mulcore_ary1_a0_c_1[6]), .Y(n7409));
INVX1 mul_U20661(.A(dpath_mulcore_ary1_a0_c_1[5]), .Y(n7410));
INVX1 mul_U20662(.A(dpath_mulcore_ary1_a0_c_1[4]), .Y(n7411));
INVX1 mul_U20663(.A(dpath_mulcore_ary1_a1_c_1[3]), .Y(n7412));
INVX1 mul_U20664(.A(dpath_mulcore_ary1_a1_c_1[6]), .Y(n7413));
INVX1 mul_U20665(.A(dpath_mulcore_ary1_a1_c_1[5]), .Y(n7414));
INVX1 mul_U20666(.A(dpath_mulcore_ary1_a1_c_1[4]), .Y(n7415));
INVX1 mul_U20667(.A(dpath_mulcore_ary1_a0_I2_I0_b0n_0), .Y(n7416));
INVX1 mul_U20668(.A(dpath_mulcore_ary1_a0_I2_I2_net43), .Y(n7417));
INVX1 mul_U20669(.A(dpath_mulcore_ary1_a0_I2_I2_net48), .Y(n7418));
INVX1 mul_U20670(.A(dpath_mulcore_ary1_a0_I2_I1_63__net046), .Y(n7419));
INVX1 mul_U20671(.A(dpath_mulcore_ary1_a0_I2_I1_62__net046), .Y(n7420));
INVX1 mul_U20672(.A(dpath_mulcore_ary1_a0_I2_I1_61__net046), .Y(n7421));
INVX1 mul_U20673(.A(dpath_mulcore_ary1_a0_I2_I1_60__net046), .Y(n7422));
INVX1 mul_U20674(.A(dpath_mulcore_ary1_a0_I2_I1_59__net046), .Y(n7423));
INVX1 mul_U20675(.A(dpath_mulcore_ary1_a0_I2_I1_58__net046), .Y(n7424));
INVX1 mul_U20676(.A(dpath_mulcore_ary1_a0_I2_I1_57__net046), .Y(n7425));
INVX1 mul_U20677(.A(dpath_mulcore_ary1_a0_I2_I1_56__net046), .Y(n7426));
INVX1 mul_U20678(.A(dpath_mulcore_ary1_a0_I2_I1_55__net046), .Y(n7427));
INVX1 mul_U20679(.A(dpath_mulcore_ary1_a0_I2_I1_54__net046), .Y(n7428));
INVX1 mul_U20680(.A(dpath_mulcore_ary1_a0_I2_I1_53__net046), .Y(n7429));
INVX1 mul_U20681(.A(dpath_mulcore_ary1_a0_I2_I1_52__net046), .Y(n7430));
INVX1 mul_U20682(.A(dpath_mulcore_ary1_a0_I2_I1_51__net046), .Y(n7431));
INVX1 mul_U20683(.A(dpath_mulcore_ary1_a0_I2_I1_50__net046), .Y(n7432));
INVX1 mul_U20684(.A(dpath_mulcore_ary1_a0_I2_I1_49__net046), .Y(n7433));
INVX1 mul_U20685(.A(dpath_mulcore_ary1_a0_I2_I1_48__net046), .Y(n7434));
INVX1 mul_U20686(.A(dpath_mulcore_ary1_a0_I2_I1_47__net046), .Y(n7435));
INVX1 mul_U20687(.A(dpath_mulcore_ary1_a0_I2_I1_46__net046), .Y(n7436));
INVX1 mul_U20688(.A(dpath_mulcore_ary1_a0_I2_I1_45__net046), .Y(n7437));
INVX1 mul_U20689(.A(dpath_mulcore_ary1_a0_I2_I1_44__net046), .Y(n7438));
INVX1 mul_U20690(.A(dpath_mulcore_ary1_a0_I2_I1_43__net046), .Y(n7439));
INVX1 mul_U20691(.A(dpath_mulcore_ary1_a0_I2_I1_42__net046), .Y(n7440));
INVX1 mul_U20692(.A(dpath_mulcore_ary1_a0_I2_I1_41__net046), .Y(n7441));
INVX1 mul_U20693(.A(dpath_mulcore_ary1_a0_I2_I1_40__net046), .Y(n7442));
INVX1 mul_U20694(.A(dpath_mulcore_ary1_a0_I2_I1_39__net046), .Y(n7443));
INVX1 mul_U20695(.A(dpath_mulcore_ary1_a0_I2_I1_38__net046), .Y(n7444));
INVX1 mul_U20696(.A(dpath_mulcore_ary1_a0_I2_I1_37__net046), .Y(n7445));
INVX1 mul_U20697(.A(dpath_mulcore_ary1_a0_I2_I1_36__net046), .Y(n7446));
INVX1 mul_U20698(.A(dpath_mulcore_ary1_a0_I2_I1_35__net046), .Y(n7447));
INVX1 mul_U20699(.A(dpath_mulcore_ary1_a0_I2_I1_34__net046), .Y(n7448));
INVX1 mul_U20700(.A(dpath_mulcore_ary1_a0_I2_I1_33__net046), .Y(n7449));
INVX1 mul_U20701(.A(dpath_mulcore_ary1_a0_I2_I1_32__net046), .Y(n7450));
INVX1 mul_U20702(.A(dpath_mulcore_ary1_a0_I2_I1_31__net046), .Y(n7451));
INVX1 mul_U20703(.A(dpath_mulcore_ary1_a0_I2_I1_30__net046), .Y(n7452));
INVX1 mul_U20704(.A(dpath_mulcore_ary1_a0_I2_I1_29__net046), .Y(n7453));
INVX1 mul_U20705(.A(dpath_mulcore_ary1_a0_I2_I1_28__net046), .Y(n7454));
INVX1 mul_U20706(.A(dpath_mulcore_ary1_a0_I2_I1_27__net046), .Y(n7455));
INVX1 mul_U20707(.A(dpath_mulcore_ary1_a0_I2_I1_26__net046), .Y(n7456));
INVX1 mul_U20708(.A(dpath_mulcore_ary1_a0_I2_I1_25__net046), .Y(n7457));
INVX1 mul_U20709(.A(dpath_mulcore_ary1_a0_I2_I1_24__net046), .Y(n7458));
INVX1 mul_U20710(.A(dpath_mulcore_ary1_a0_I2_I1_23__net046), .Y(n7459));
INVX1 mul_U20711(.A(dpath_mulcore_ary1_a0_I2_I1_22__net046), .Y(n7460));
INVX1 mul_U20712(.A(dpath_mulcore_ary1_a0_I2_I1_21__net046), .Y(n7461));
INVX1 mul_U20713(.A(dpath_mulcore_ary1_a0_I2_I1_20__net046), .Y(n7462));
INVX1 mul_U20714(.A(dpath_mulcore_ary1_a0_I2_I1_19__net046), .Y(n7463));
INVX1 mul_U20715(.A(dpath_mulcore_ary1_a0_I2_I1_18__net046), .Y(n7464));
INVX1 mul_U20716(.A(dpath_mulcore_ary1_a0_I2_I1_17__net046), .Y(n7465));
INVX1 mul_U20717(.A(dpath_mulcore_ary1_a0_I2_I1_16__net046), .Y(n7466));
INVX1 mul_U20718(.A(dpath_mulcore_ary1_a0_I2_I1_15__net046), .Y(n7467));
INVX1 mul_U20719(.A(dpath_mulcore_ary1_a0_I2_I1_14__net046), .Y(n7468));
INVX1 mul_U20720(.A(dpath_mulcore_ary1_a0_I2_I1_13__net046), .Y(n7469));
INVX1 mul_U20721(.A(dpath_mulcore_ary1_a0_I2_I1_12__net046), .Y(n7470));
INVX1 mul_U20722(.A(dpath_mulcore_ary1_a0_I2_I1_11__net046), .Y(n7471));
INVX1 mul_U20723(.A(dpath_mulcore_ary1_a0_I2_I1_10__net046), .Y(n7472));
INVX1 mul_U20724(.A(dpath_mulcore_ary1_a0_I2_I1_9__net046), .Y(n7473));
INVX1 mul_U20725(.A(dpath_mulcore_ary1_a0_I2_I1_8__net046), .Y(n7474));
INVX1 mul_U20726(.A(dpath_mulcore_ary1_a0_I2_I1_7__net046), .Y(n7475));
INVX1 mul_U20727(.A(dpath_mulcore_ary1_a0_I2_I1_6__net046), .Y(n7476));
INVX1 mul_U20728(.A(dpath_mulcore_ary1_a0_I2_I1_5__net046), .Y(n7477));
INVX1 mul_U20729(.A(dpath_mulcore_ary1_a0_I2_I1_4__net046), .Y(n7478));
INVX1 mul_U20730(.A(dpath_mulcore_ary1_a0_I2_I0_p0_3), .Y(n7479));
INVX1 mul_U20731(.A(dpath_mulcore_ary1_a0_I2_I0_p0_2), .Y(n7480));
INVX1 mul_U20732(.A(dpath_mulcore_ary1_a0_I1_I2_net078), .Y(n7481));
INVX1 mul_U20733(.A(dpath_mulcore_ary1_a0_I1_I2_net8), .Y(n7482));
INVX1 mul_U20734(.A(dpath_mulcore_ary1_a0_I1_I2_net15), .Y(n7483));
INVX1 mul_U20735(.A(dpath_mulcore_ary1_a0_I1_I2_net43), .Y(n7484));
INVX1 mul_U20736(.A(dpath_mulcore_ary1_a0_I1_I2_net48), .Y(n7485));
INVX1 mul_U20737(.A(dpath_mulcore_ary1_a0_I1_I2_net35), .Y(n7486));
INVX1 mul_U20738(.A(dpath_mulcore_ary1_a0_I1_I1_63__net043), .Y(n7487));
INVX1 mul_U20739(.A(dpath_mulcore_ary1_a0_I1_I1_63__net046), .Y(n7488));
INVX1 mul_U20740(.A(dpath_mulcore_ary1_a0_I1_I1_62__net043), .Y(n7489));
INVX1 mul_U20741(.A(dpath_mulcore_ary1_a0_I1_I1_62__net046), .Y(n7490));
INVX1 mul_U20742(.A(dpath_mulcore_ary1_a0_I1_I1_61__net043), .Y(n7491));
INVX1 mul_U20743(.A(dpath_mulcore_ary1_a0_I1_I1_61__net046), .Y(n7492));
INVX1 mul_U20744(.A(dpath_mulcore_ary1_a0_I1_I1_60__net043), .Y(n7493));
INVX1 mul_U20745(.A(dpath_mulcore_ary1_a0_I1_I1_60__net046), .Y(n7494));
INVX1 mul_U20746(.A(dpath_mulcore_ary1_a0_I1_I1_59__net043), .Y(n7495));
INVX1 mul_U20747(.A(dpath_mulcore_ary1_a0_I1_I1_59__net046), .Y(n7496));
INVX1 mul_U20748(.A(dpath_mulcore_ary1_a0_I1_I1_58__net043), .Y(n7497));
INVX1 mul_U20749(.A(dpath_mulcore_ary1_a0_I1_I1_58__net046), .Y(n7498));
INVX1 mul_U20750(.A(dpath_mulcore_ary1_a0_I1_I1_57__net043), .Y(n7499));
INVX1 mul_U20751(.A(dpath_mulcore_ary1_a0_I1_I1_57__net046), .Y(n7500));
INVX1 mul_U20752(.A(dpath_mulcore_ary1_a0_I1_I1_56__net043), .Y(n7501));
INVX1 mul_U20753(.A(dpath_mulcore_ary1_a0_I1_I1_56__net046), .Y(n7502));
INVX1 mul_U20754(.A(dpath_mulcore_ary1_a0_I1_I1_55__net043), .Y(n7503));
INVX1 mul_U20755(.A(dpath_mulcore_ary1_a0_I1_I1_55__net046), .Y(n7504));
INVX1 mul_U20756(.A(dpath_mulcore_ary1_a0_I1_I1_54__net043), .Y(n7505));
INVX1 mul_U20757(.A(dpath_mulcore_ary1_a0_I1_I1_54__net046), .Y(n7506));
INVX1 mul_U20758(.A(dpath_mulcore_ary1_a0_I1_I1_53__net043), .Y(n7507));
INVX1 mul_U20759(.A(dpath_mulcore_ary1_a0_I1_I1_53__net046), .Y(n7508));
INVX1 mul_U20760(.A(dpath_mulcore_ary1_a0_I1_I1_52__net043), .Y(n7509));
INVX1 mul_U20761(.A(dpath_mulcore_ary1_a0_I1_I1_52__net046), .Y(n7510));
INVX1 mul_U20762(.A(dpath_mulcore_ary1_a0_I1_I1_51__net043), .Y(n7511));
INVX1 mul_U20763(.A(dpath_mulcore_ary1_a0_I1_I1_51__net046), .Y(n7512));
INVX1 mul_U20764(.A(dpath_mulcore_ary1_a0_I1_I1_50__net043), .Y(n7513));
INVX1 mul_U20765(.A(dpath_mulcore_ary1_a0_I1_I1_50__net046), .Y(n7514));
INVX1 mul_U20766(.A(dpath_mulcore_ary1_a0_I1_I1_49__net043), .Y(n7515));
INVX1 mul_U20767(.A(dpath_mulcore_ary1_a0_I1_I1_49__net046), .Y(n7516));
INVX1 mul_U20768(.A(dpath_mulcore_ary1_a0_I1_I1_48__net043), .Y(n7517));
INVX1 mul_U20769(.A(dpath_mulcore_ary1_a0_I1_I1_48__net046), .Y(n7518));
INVX1 mul_U20770(.A(dpath_mulcore_ary1_a0_I1_I1_47__net043), .Y(n7519));
INVX1 mul_U20771(.A(dpath_mulcore_ary1_a0_I1_I1_47__net046), .Y(n7520));
INVX1 mul_U20772(.A(dpath_mulcore_ary1_a0_I1_I1_46__net043), .Y(n7521));
INVX1 mul_U20773(.A(dpath_mulcore_ary1_a0_I1_I1_46__net046), .Y(n7522));
INVX1 mul_U20774(.A(dpath_mulcore_ary1_a0_I1_I1_45__net043), .Y(n7523));
INVX1 mul_U20775(.A(dpath_mulcore_ary1_a0_I1_I1_45__net046), .Y(n7524));
INVX1 mul_U20776(.A(dpath_mulcore_ary1_a0_I1_I1_44__net043), .Y(n7525));
INVX1 mul_U20777(.A(dpath_mulcore_ary1_a0_I1_I1_44__net046), .Y(n7526));
INVX1 mul_U20778(.A(dpath_mulcore_ary1_a0_I1_I1_43__net043), .Y(n7527));
INVX1 mul_U20779(.A(dpath_mulcore_ary1_a0_I1_I1_43__net046), .Y(n7528));
INVX1 mul_U20780(.A(dpath_mulcore_ary1_a0_I1_I1_42__net043), .Y(n7529));
INVX1 mul_U20781(.A(dpath_mulcore_ary1_a0_I1_I1_42__net046), .Y(n7530));
INVX1 mul_U20782(.A(dpath_mulcore_ary1_a0_I1_I1_41__net043), .Y(n7531));
INVX1 mul_U20783(.A(dpath_mulcore_ary1_a0_I1_I1_41__net046), .Y(n7532));
INVX1 mul_U20784(.A(dpath_mulcore_ary1_a0_I1_I1_40__net043), .Y(n7533));
INVX1 mul_U20785(.A(dpath_mulcore_ary1_a0_I1_I1_40__net046), .Y(n7534));
INVX1 mul_U20786(.A(dpath_mulcore_ary1_a0_I1_I1_39__net043), .Y(n7535));
INVX1 mul_U20787(.A(dpath_mulcore_ary1_a0_I1_I1_39__net046), .Y(n7536));
INVX1 mul_U20788(.A(dpath_mulcore_ary1_a0_I1_I1_38__net043), .Y(n7537));
INVX1 mul_U20789(.A(dpath_mulcore_ary1_a0_I1_I1_38__net046), .Y(n7538));
INVX1 mul_U20790(.A(dpath_mulcore_ary1_a0_I1_I1_37__net043), .Y(n7539));
INVX1 mul_U20791(.A(dpath_mulcore_ary1_a0_I1_I1_37__net046), .Y(n7540));
INVX1 mul_U20792(.A(dpath_mulcore_ary1_a0_I1_I1_36__net043), .Y(n7541));
INVX1 mul_U20793(.A(dpath_mulcore_ary1_a0_I1_I1_36__net046), .Y(n7542));
INVX1 mul_U20794(.A(dpath_mulcore_ary1_a0_I1_I1_35__net043), .Y(n7543));
INVX1 mul_U20795(.A(dpath_mulcore_ary1_a0_I1_I1_35__net046), .Y(n7544));
INVX1 mul_U20796(.A(dpath_mulcore_ary1_a0_I1_I1_34__net043), .Y(n7545));
INVX1 mul_U20797(.A(dpath_mulcore_ary1_a0_I1_I1_34__net046), .Y(n7546));
INVX1 mul_U20798(.A(dpath_mulcore_ary1_a0_I1_I1_33__net043), .Y(n7547));
INVX1 mul_U20799(.A(dpath_mulcore_ary1_a0_I1_I1_33__net046), .Y(n7548));
INVX1 mul_U20800(.A(dpath_mulcore_ary1_a0_I1_I1_32__net043), .Y(n7549));
INVX1 mul_U20801(.A(dpath_mulcore_ary1_a0_I1_I1_32__net046), .Y(n7550));
INVX1 mul_U20802(.A(dpath_mulcore_ary1_a0_I1_I1_31__net043), .Y(n7551));
INVX1 mul_U20803(.A(dpath_mulcore_ary1_a0_I1_I1_31__net046), .Y(n7552));
INVX1 mul_U20804(.A(dpath_mulcore_ary1_a0_I1_I1_30__net043), .Y(n7553));
INVX1 mul_U20805(.A(dpath_mulcore_ary1_a0_I1_I1_30__net046), .Y(n7554));
INVX1 mul_U20806(.A(dpath_mulcore_ary1_a0_I1_I1_29__net043), .Y(n7555));
INVX1 mul_U20807(.A(dpath_mulcore_ary1_a0_I1_I1_29__net046), .Y(n7556));
INVX1 mul_U20808(.A(dpath_mulcore_ary1_a0_I1_I1_28__net043), .Y(n7557));
INVX1 mul_U20809(.A(dpath_mulcore_ary1_a0_I1_I1_28__net046), .Y(n7558));
INVX1 mul_U20810(.A(dpath_mulcore_ary1_a0_I1_I1_27__net043), .Y(n7559));
INVX1 mul_U20811(.A(dpath_mulcore_ary1_a0_I1_I1_27__net046), .Y(n7560));
INVX1 mul_U20812(.A(dpath_mulcore_ary1_a0_I1_I1_26__net043), .Y(n7561));
INVX1 mul_U20813(.A(dpath_mulcore_ary1_a0_I1_I1_26__net046), .Y(n7562));
INVX1 mul_U20814(.A(dpath_mulcore_ary1_a0_I1_I1_25__net043), .Y(n7563));
INVX1 mul_U20815(.A(dpath_mulcore_ary1_a0_I1_I1_25__net046), .Y(n7564));
INVX1 mul_U20816(.A(dpath_mulcore_ary1_a0_I1_I1_24__net043), .Y(n7565));
INVX1 mul_U20817(.A(dpath_mulcore_ary1_a0_I1_I1_24__net046), .Y(n7566));
INVX1 mul_U20818(.A(dpath_mulcore_ary1_a0_I1_I1_23__net043), .Y(n7567));
INVX1 mul_U20819(.A(dpath_mulcore_ary1_a0_I1_I1_23__net046), .Y(n7568));
INVX1 mul_U20820(.A(dpath_mulcore_ary1_a0_I1_I1_22__net043), .Y(n7569));
INVX1 mul_U20821(.A(dpath_mulcore_ary1_a0_I1_I1_22__net046), .Y(n7570));
INVX1 mul_U20822(.A(dpath_mulcore_ary1_a0_I1_I1_21__net043), .Y(n7571));
INVX1 mul_U20823(.A(dpath_mulcore_ary1_a0_I1_I1_21__net046), .Y(n7572));
INVX1 mul_U20824(.A(dpath_mulcore_ary1_a0_I1_I1_20__net043), .Y(n7573));
INVX1 mul_U20825(.A(dpath_mulcore_ary1_a0_I1_I1_20__net046), .Y(n7574));
INVX1 mul_U20826(.A(dpath_mulcore_ary1_a0_I1_I1_19__net043), .Y(n7575));
INVX1 mul_U20827(.A(dpath_mulcore_ary1_a0_I1_I1_19__net046), .Y(n7576));
INVX1 mul_U20828(.A(dpath_mulcore_ary1_a0_I1_I1_18__net043), .Y(n7577));
INVX1 mul_U20829(.A(dpath_mulcore_ary1_a0_I1_I1_18__net046), .Y(n7578));
INVX1 mul_U20830(.A(dpath_mulcore_ary1_a0_I1_I1_17__net043), .Y(n7579));
INVX1 mul_U20831(.A(dpath_mulcore_ary1_a0_I1_I1_17__net046), .Y(n7580));
INVX1 mul_U20832(.A(dpath_mulcore_ary1_a0_I1_I1_16__net043), .Y(n7581));
INVX1 mul_U20833(.A(dpath_mulcore_ary1_a0_I1_I1_16__net046), .Y(n7582));
INVX1 mul_U20834(.A(dpath_mulcore_ary1_a0_I1_I1_15__net043), .Y(n7583));
INVX1 mul_U20835(.A(dpath_mulcore_ary1_a0_I1_I1_15__net046), .Y(n7584));
INVX1 mul_U20836(.A(dpath_mulcore_ary1_a0_I1_I1_14__net043), .Y(n7585));
INVX1 mul_U20837(.A(dpath_mulcore_ary1_a0_I1_I1_14__net046), .Y(n7586));
INVX1 mul_U20838(.A(dpath_mulcore_ary1_a0_I1_I1_13__net043), .Y(n7587));
INVX1 mul_U20839(.A(dpath_mulcore_ary1_a0_I1_I1_13__net046), .Y(n7588));
INVX1 mul_U20840(.A(dpath_mulcore_ary1_a0_I1_I1_12__net043), .Y(n7589));
INVX1 mul_U20841(.A(dpath_mulcore_ary1_a0_I1_I1_12__net046), .Y(n7590));
INVX1 mul_U20842(.A(dpath_mulcore_ary1_a0_I1_I1_11__net043), .Y(n7591));
INVX1 mul_U20843(.A(dpath_mulcore_ary1_a0_I1_I1_11__net046), .Y(n7592));
INVX1 mul_U20844(.A(dpath_mulcore_ary1_a0_I1_I1_10__net043), .Y(n7593));
INVX1 mul_U20845(.A(dpath_mulcore_ary1_a0_I1_I1_10__net046), .Y(n7594));
INVX1 mul_U20846(.A(dpath_mulcore_ary1_a0_I1_I1_9__net043), .Y(n7595));
INVX1 mul_U20847(.A(dpath_mulcore_ary1_a0_I1_I1_9__net046), .Y(n7596));
INVX1 mul_U20848(.A(dpath_mulcore_ary1_a0_I1_I1_8__net043), .Y(n7597));
INVX1 mul_U20849(.A(dpath_mulcore_ary1_a0_I1_I1_8__net046), .Y(n7598));
INVX1 mul_U20850(.A(dpath_mulcore_ary1_a0_I1_I1_7__net043), .Y(n7599));
INVX1 mul_U20851(.A(dpath_mulcore_ary1_a0_I1_I1_7__net046), .Y(n7600));
INVX1 mul_U20852(.A(dpath_mulcore_ary1_a0_I1_I1_6__net043), .Y(n7601));
INVX1 mul_U20853(.A(dpath_mulcore_ary1_a0_I1_I1_6__net046), .Y(n7602));
INVX1 mul_U20854(.A(dpath_mulcore_ary1_a0_I1_I1_5__net043), .Y(n7603));
INVX1 mul_U20855(.A(dpath_mulcore_ary1_a0_I1_I1_5__net046), .Y(n7604));
INVX1 mul_U20856(.A(dpath_mulcore_ary1_a0_I1_I1_4__net046), .Y(n7605));
INVX1 mul_U20857(.A(dpath_mulcore_ary1_a0_I1_I0_p0_3), .Y(n7606));
INVX1 mul_U20858(.A(dpath_mulcore_ary1_a0_I1_I0_p0_2), .Y(n7607));
INVX1 mul_U20859(.A(dpath_mulcore_ary1_a0_I0_I2_net078), .Y(n7608));
INVX1 mul_U20860(.A(dpath_mulcore_ary1_a0_I0_I2_net8), .Y(n7609));
INVX1 mul_U20861(.A(dpath_mulcore_ary1_a0_I0_I2_net15), .Y(n7610));
INVX1 mul_U20862(.A(dpath_mulcore_ary1_a0_I0_I2_net43), .Y(n7611));
INVX1 mul_U20863(.A(dpath_mulcore_ary1_a0_I0_I2_net48), .Y(n7612));
INVX1 mul_U20864(.A(dpath_mulcore_ary1_a0_I0_I2_net35), .Y(n7613));
INVX1 mul_U20865(.A(dpath_mulcore_ary1_a0_I0_I1_63__net043), .Y(n7614));
INVX1 mul_U20866(.A(dpath_mulcore_ary1_a0_I0_I1_63__net046), .Y(n7615));
INVX1 mul_U20867(.A(dpath_mulcore_ary1_a0_I0_I1_62__net043), .Y(n7616));
INVX1 mul_U20868(.A(dpath_mulcore_ary1_a0_I0_I1_62__net046), .Y(n7617));
INVX1 mul_U20869(.A(dpath_mulcore_ary1_a0_I0_I1_61__net043), .Y(n7618));
INVX1 mul_U20870(.A(dpath_mulcore_ary1_a0_I0_I1_61__net046), .Y(n7619));
INVX1 mul_U20871(.A(dpath_mulcore_ary1_a0_I0_I1_60__net043), .Y(n7620));
INVX1 mul_U20872(.A(dpath_mulcore_ary1_a0_I0_I1_60__net046), .Y(n7621));
INVX1 mul_U20873(.A(dpath_mulcore_ary1_a0_I0_I1_59__net043), .Y(n7622));
INVX1 mul_U20874(.A(dpath_mulcore_ary1_a0_I0_I1_59__net046), .Y(n7623));
INVX1 mul_U20875(.A(dpath_mulcore_ary1_a0_I0_I1_58__net043), .Y(n7624));
INVX1 mul_U20876(.A(dpath_mulcore_ary1_a0_I0_I1_58__net046), .Y(n7625));
INVX1 mul_U20877(.A(dpath_mulcore_ary1_a0_I0_I1_57__net043), .Y(n7626));
INVX1 mul_U20878(.A(dpath_mulcore_ary1_a0_I0_I1_57__net046), .Y(n7627));
INVX1 mul_U20879(.A(dpath_mulcore_ary1_a0_I0_I1_56__net043), .Y(n7628));
INVX1 mul_U20880(.A(dpath_mulcore_ary1_a0_I0_I1_56__net046), .Y(n7629));
INVX1 mul_U20881(.A(dpath_mulcore_ary1_a0_I0_I1_55__net043), .Y(n7630));
INVX1 mul_U20882(.A(dpath_mulcore_ary1_a0_I0_I1_55__net046), .Y(n7631));
INVX1 mul_U20883(.A(dpath_mulcore_ary1_a0_I0_I1_54__net043), .Y(n7632));
INVX1 mul_U20884(.A(dpath_mulcore_ary1_a0_I0_I1_54__net046), .Y(n7633));
INVX1 mul_U20885(.A(dpath_mulcore_ary1_a0_I0_I1_53__net043), .Y(n7634));
INVX1 mul_U20886(.A(dpath_mulcore_ary1_a0_I0_I1_53__net046), .Y(n7635));
INVX1 mul_U20887(.A(dpath_mulcore_ary1_a0_I0_I1_52__net043), .Y(n7636));
INVX1 mul_U20888(.A(dpath_mulcore_ary1_a0_I0_I1_52__net046), .Y(n7637));
INVX1 mul_U20889(.A(dpath_mulcore_ary1_a0_I0_I1_51__net043), .Y(n7638));
INVX1 mul_U20890(.A(dpath_mulcore_ary1_a0_I0_I1_51__net046), .Y(n7639));
INVX1 mul_U20891(.A(dpath_mulcore_ary1_a0_I0_I1_50__net043), .Y(n7640));
INVX1 mul_U20892(.A(dpath_mulcore_ary1_a0_I0_I1_50__net046), .Y(n7641));
INVX1 mul_U20893(.A(dpath_mulcore_ary1_a0_I0_I1_49__net043), .Y(n7642));
INVX1 mul_U20894(.A(dpath_mulcore_ary1_a0_I0_I1_49__net046), .Y(n7643));
INVX1 mul_U20895(.A(dpath_mulcore_ary1_a0_I0_I1_48__net043), .Y(n7644));
INVX1 mul_U20896(.A(dpath_mulcore_ary1_a0_I0_I1_48__net046), .Y(n7645));
INVX1 mul_U20897(.A(dpath_mulcore_ary1_a0_I0_I1_47__net043), .Y(n7646));
INVX1 mul_U20898(.A(dpath_mulcore_ary1_a0_I0_I1_47__net046), .Y(n7647));
INVX1 mul_U20899(.A(dpath_mulcore_ary1_a0_I0_I1_46__net043), .Y(n7648));
INVX1 mul_U20900(.A(dpath_mulcore_ary1_a0_I0_I1_46__net046), .Y(n7649));
INVX1 mul_U20901(.A(dpath_mulcore_ary1_a0_I0_I1_45__net043), .Y(n7650));
INVX1 mul_U20902(.A(dpath_mulcore_ary1_a0_I0_I1_45__net046), .Y(n7651));
INVX1 mul_U20903(.A(dpath_mulcore_ary1_a0_I0_I1_44__net043), .Y(n7652));
INVX1 mul_U20904(.A(dpath_mulcore_ary1_a0_I0_I1_44__net046), .Y(n7653));
INVX1 mul_U20905(.A(dpath_mulcore_ary1_a0_I0_I1_43__net043), .Y(n7654));
INVX1 mul_U20906(.A(dpath_mulcore_ary1_a0_I0_I1_43__net046), .Y(n7655));
INVX1 mul_U20907(.A(dpath_mulcore_ary1_a0_I0_I1_42__net043), .Y(n7656));
INVX1 mul_U20908(.A(dpath_mulcore_ary1_a0_I0_I1_42__net046), .Y(n7657));
INVX1 mul_U20909(.A(dpath_mulcore_ary1_a0_I0_I1_41__net043), .Y(n7658));
INVX1 mul_U20910(.A(dpath_mulcore_ary1_a0_I0_I1_41__net046), .Y(n7659));
INVX1 mul_U20911(.A(dpath_mulcore_ary1_a0_I0_I1_40__net043), .Y(n7660));
INVX1 mul_U20912(.A(dpath_mulcore_ary1_a0_I0_I1_40__net046), .Y(n7661));
INVX1 mul_U20913(.A(dpath_mulcore_ary1_a0_I0_I1_39__net043), .Y(n7662));
INVX1 mul_U20914(.A(dpath_mulcore_ary1_a0_I0_I1_39__net046), .Y(n7663));
INVX1 mul_U20915(.A(dpath_mulcore_ary1_a0_I0_I1_38__net043), .Y(n7664));
INVX1 mul_U20916(.A(dpath_mulcore_ary1_a0_I0_I1_38__net046), .Y(n7665));
INVX1 mul_U20917(.A(dpath_mulcore_ary1_a0_I0_I1_37__net043), .Y(n7666));
INVX1 mul_U20918(.A(dpath_mulcore_ary1_a0_I0_I1_37__net046), .Y(n7667));
INVX1 mul_U20919(.A(dpath_mulcore_ary1_a0_I0_I1_36__net043), .Y(n7668));
INVX1 mul_U20920(.A(dpath_mulcore_ary1_a0_I0_I1_36__net046), .Y(n7669));
INVX1 mul_U20921(.A(dpath_mulcore_ary1_a0_I0_I1_35__net043), .Y(n7670));
INVX1 mul_U20922(.A(dpath_mulcore_ary1_a0_I0_I1_35__net046), .Y(n7671));
INVX1 mul_U20923(.A(dpath_mulcore_ary1_a0_I0_I1_34__net043), .Y(n7672));
INVX1 mul_U20924(.A(dpath_mulcore_ary1_a0_I0_I1_34__net046), .Y(n7673));
INVX1 mul_U20925(.A(dpath_mulcore_ary1_a0_I0_I1_33__net043), .Y(n7674));
INVX1 mul_U20926(.A(dpath_mulcore_ary1_a0_I0_I1_33__net046), .Y(n7675));
INVX1 mul_U20927(.A(dpath_mulcore_ary1_a0_I0_I1_32__net043), .Y(n7676));
INVX1 mul_U20928(.A(dpath_mulcore_ary1_a0_I0_I1_32__net046), .Y(n7677));
INVX1 mul_U20929(.A(dpath_mulcore_ary1_a0_I0_I1_31__net043), .Y(n7678));
INVX1 mul_U20930(.A(dpath_mulcore_ary1_a0_I0_I1_31__net046), .Y(n7679));
INVX1 mul_U20931(.A(dpath_mulcore_ary1_a0_I0_I1_30__net043), .Y(n7680));
INVX1 mul_U20932(.A(dpath_mulcore_ary1_a0_I0_I1_30__net046), .Y(n7681));
INVX1 mul_U20933(.A(dpath_mulcore_ary1_a0_I0_I1_29__net043), .Y(n7682));
INVX1 mul_U20934(.A(dpath_mulcore_ary1_a0_I0_I1_29__net046), .Y(n7683));
INVX1 mul_U20935(.A(dpath_mulcore_ary1_a0_I0_I1_28__net043), .Y(n7684));
INVX1 mul_U20936(.A(dpath_mulcore_ary1_a0_I0_I1_28__net046), .Y(n7685));
INVX1 mul_U20937(.A(dpath_mulcore_ary1_a0_I0_I1_27__net043), .Y(n7686));
INVX1 mul_U20938(.A(dpath_mulcore_ary1_a0_I0_I1_27__net046), .Y(n7687));
INVX1 mul_U20939(.A(dpath_mulcore_ary1_a0_I0_I1_26__net043), .Y(n7688));
INVX1 mul_U20940(.A(dpath_mulcore_ary1_a0_I0_I1_26__net046), .Y(n7689));
INVX1 mul_U20941(.A(dpath_mulcore_ary1_a0_I0_I1_25__net043), .Y(n7690));
INVX1 mul_U20942(.A(dpath_mulcore_ary1_a0_I0_I1_25__net046), .Y(n7691));
INVX1 mul_U20943(.A(dpath_mulcore_ary1_a0_I0_I1_24__net043), .Y(n7692));
INVX1 mul_U20944(.A(dpath_mulcore_ary1_a0_I0_I1_24__net046), .Y(n7693));
INVX1 mul_U20945(.A(dpath_mulcore_ary1_a0_I0_I1_23__net043), .Y(n7694));
INVX1 mul_U20946(.A(dpath_mulcore_ary1_a0_I0_I1_23__net046), .Y(n7695));
INVX1 mul_U20947(.A(dpath_mulcore_ary1_a0_I0_I1_22__net043), .Y(n7696));
INVX1 mul_U20948(.A(dpath_mulcore_ary1_a0_I0_I1_22__net046), .Y(n7697));
INVX1 mul_U20949(.A(dpath_mulcore_ary1_a0_I0_I1_21__net043), .Y(n7698));
INVX1 mul_U20950(.A(dpath_mulcore_ary1_a0_I0_I1_21__net046), .Y(n7699));
INVX1 mul_U20951(.A(dpath_mulcore_ary1_a0_I0_I1_20__net043), .Y(n7700));
INVX1 mul_U20952(.A(dpath_mulcore_ary1_a0_I0_I1_20__net046), .Y(n7701));
INVX1 mul_U20953(.A(dpath_mulcore_ary1_a0_I0_I1_19__net043), .Y(n7702));
INVX1 mul_U20954(.A(dpath_mulcore_ary1_a0_I0_I1_19__net046), .Y(n7703));
INVX1 mul_U20955(.A(dpath_mulcore_ary1_a0_I0_I1_18__net043), .Y(n7704));
INVX1 mul_U20956(.A(dpath_mulcore_ary1_a0_I0_I1_18__net046), .Y(n7705));
INVX1 mul_U20957(.A(dpath_mulcore_ary1_a0_I0_I1_17__net043), .Y(n7706));
INVX1 mul_U20958(.A(dpath_mulcore_ary1_a0_I0_I1_17__net046), .Y(n7707));
INVX1 mul_U20959(.A(dpath_mulcore_ary1_a0_I0_I1_16__net043), .Y(n7708));
INVX1 mul_U20960(.A(dpath_mulcore_ary1_a0_I0_I1_16__net046), .Y(n7709));
INVX1 mul_U20961(.A(dpath_mulcore_ary1_a0_I0_I1_15__net043), .Y(n7710));
INVX1 mul_U20962(.A(dpath_mulcore_ary1_a0_I0_I1_15__net046), .Y(n7711));
INVX1 mul_U20963(.A(dpath_mulcore_ary1_a0_I0_I1_14__net043), .Y(n7712));
INVX1 mul_U20964(.A(dpath_mulcore_ary1_a0_I0_I1_14__net046), .Y(n7713));
INVX1 mul_U20965(.A(dpath_mulcore_ary1_a0_I0_I1_13__net043), .Y(n7714));
INVX1 mul_U20966(.A(dpath_mulcore_ary1_a0_I0_I1_13__net046), .Y(n7715));
INVX1 mul_U20967(.A(dpath_mulcore_ary1_a0_I0_I1_12__net043), .Y(n7716));
INVX1 mul_U20968(.A(dpath_mulcore_ary1_a0_I0_I1_12__net046), .Y(n7717));
INVX1 mul_U20969(.A(dpath_mulcore_ary1_a0_I0_I1_11__net043), .Y(n7718));
INVX1 mul_U20970(.A(dpath_mulcore_ary1_a0_I0_I1_11__net046), .Y(n7719));
INVX1 mul_U20971(.A(dpath_mulcore_ary1_a0_I0_I1_10__net043), .Y(n7720));
INVX1 mul_U20972(.A(dpath_mulcore_ary1_a0_I0_I1_10__net046), .Y(n7721));
INVX1 mul_U20973(.A(dpath_mulcore_ary1_a0_I0_I1_9__net043), .Y(n7722));
INVX1 mul_U20974(.A(dpath_mulcore_ary1_a0_I0_I1_9__net046), .Y(n7723));
INVX1 mul_U20975(.A(dpath_mulcore_ary1_a0_I0_I1_8__net043), .Y(n7724));
INVX1 mul_U20976(.A(dpath_mulcore_ary1_a0_I0_I1_8__net046), .Y(n7725));
INVX1 mul_U20977(.A(dpath_mulcore_ary1_a0_I0_I1_7__net043), .Y(n7726));
INVX1 mul_U20978(.A(dpath_mulcore_ary1_a0_I0_I1_7__net046), .Y(n7727));
INVX1 mul_U20979(.A(dpath_mulcore_ary1_a0_I0_I1_6__net043), .Y(n7728));
INVX1 mul_U20980(.A(dpath_mulcore_ary1_a0_I0_I1_6__net046), .Y(n7729));
INVX1 mul_U20981(.A(dpath_mulcore_ary1_a0_I0_I1_5__net043), .Y(n7730));
INVX1 mul_U20982(.A(dpath_mulcore_ary1_a0_I0_I1_5__net046), .Y(n7731));
INVX1 mul_U20983(.A(dpath_mulcore_ary1_a0_I0_I1_4__net046), .Y(n7732));
INVX1 mul_U20984(.A(dpath_mulcore_ary1_a0_I0_I0_p0_3), .Y(n7733));
INVX1 mul_U20985(.A(dpath_mulcore_ary1_a0_I0_I0_p0_2), .Y(n7734));
INVX1 mul_U20986(.A(dpath_mulcore_ary1_a1_I2_I2_net43), .Y(n7735));
INVX1 mul_U20987(.A(dpath_mulcore_ary1_a1_I2_I2_net48), .Y(n7736));
INVX1 mul_U20988(.A(dpath_mulcore_ary1_a1_I2_I1_63__net046), .Y(n7737));
INVX1 mul_U20989(.A(dpath_mulcore_ary1_a1_I2_I1_62__net046), .Y(n7738));
INVX1 mul_U20990(.A(dpath_mulcore_ary1_a1_I2_I1_61__net046), .Y(n7739));
INVX1 mul_U20991(.A(dpath_mulcore_ary1_a1_I2_I1_60__net046), .Y(n7740));
INVX1 mul_U20992(.A(dpath_mulcore_ary1_a1_I2_I1_59__net046), .Y(n7741));
INVX1 mul_U20993(.A(dpath_mulcore_ary1_a1_I2_I1_58__net046), .Y(n7742));
INVX1 mul_U20994(.A(dpath_mulcore_ary1_a1_I2_I1_57__net046), .Y(n7743));
INVX1 mul_U20995(.A(dpath_mulcore_ary1_a1_I2_I1_56__net046), .Y(n7744));
INVX1 mul_U20996(.A(dpath_mulcore_ary1_a1_I2_I1_55__net046), .Y(n7745));
INVX1 mul_U20997(.A(dpath_mulcore_ary1_a1_I2_I1_54__net046), .Y(n7746));
INVX1 mul_U20998(.A(dpath_mulcore_ary1_a1_I2_I1_53__net046), .Y(n7747));
INVX1 mul_U20999(.A(dpath_mulcore_ary1_a1_I2_I1_52__net046), .Y(n7748));
INVX1 mul_U21000(.A(dpath_mulcore_ary1_a1_I2_I1_51__net046), .Y(n7749));
INVX1 mul_U21001(.A(dpath_mulcore_ary1_a1_I2_I1_50__net046), .Y(n7750));
INVX1 mul_U21002(.A(dpath_mulcore_ary1_a1_I2_I1_49__net046), .Y(n7751));
INVX1 mul_U21003(.A(dpath_mulcore_ary1_a1_I2_I1_48__net046), .Y(n7752));
INVX1 mul_U21004(.A(dpath_mulcore_ary1_a1_I2_I1_47__net046), .Y(n7753));
INVX1 mul_U21005(.A(dpath_mulcore_ary1_a1_I2_I1_46__net046), .Y(n7754));
INVX1 mul_U21006(.A(dpath_mulcore_ary1_a1_I2_I1_45__net046), .Y(n7755));
INVX1 mul_U21007(.A(dpath_mulcore_ary1_a1_I2_I1_44__net046), .Y(n7756));
INVX1 mul_U21008(.A(dpath_mulcore_ary1_a1_I2_I1_43__net046), .Y(n7757));
INVX1 mul_U21009(.A(dpath_mulcore_ary1_a1_I2_I1_42__net046), .Y(n7758));
INVX1 mul_U21010(.A(dpath_mulcore_ary1_a1_I2_I1_41__net046), .Y(n7759));
INVX1 mul_U21011(.A(dpath_mulcore_ary1_a1_I2_I1_40__net046), .Y(n7760));
INVX1 mul_U21012(.A(dpath_mulcore_ary1_a1_I2_I1_39__net046), .Y(n7761));
INVX1 mul_U21013(.A(dpath_mulcore_ary1_a1_I2_I1_38__net046), .Y(n7762));
INVX1 mul_U21014(.A(dpath_mulcore_ary1_a1_I2_I1_37__net046), .Y(n7763));
INVX1 mul_U21015(.A(dpath_mulcore_ary1_a1_I2_I1_36__net046), .Y(n7764));
INVX1 mul_U21016(.A(dpath_mulcore_ary1_a1_I2_I1_35__net046), .Y(n7765));
INVX1 mul_U21017(.A(dpath_mulcore_ary1_a1_I2_I1_34__net046), .Y(n7766));
INVX1 mul_U21018(.A(dpath_mulcore_ary1_a1_I2_I1_33__net046), .Y(n7767));
INVX1 mul_U21019(.A(dpath_mulcore_ary1_a1_I2_I1_32__net046), .Y(n7768));
INVX1 mul_U21020(.A(dpath_mulcore_ary1_a1_I2_I1_31__net046), .Y(n7769));
INVX1 mul_U21021(.A(dpath_mulcore_ary1_a1_I2_I1_30__net046), .Y(n7770));
INVX1 mul_U21022(.A(dpath_mulcore_ary1_a1_I2_I1_29__net046), .Y(n7771));
INVX1 mul_U21023(.A(dpath_mulcore_ary1_a1_I2_I1_28__net046), .Y(n7772));
INVX1 mul_U21024(.A(dpath_mulcore_ary1_a1_I2_I1_27__net046), .Y(n7773));
INVX1 mul_U21025(.A(dpath_mulcore_ary1_a1_I2_I1_26__net046), .Y(n7774));
INVX1 mul_U21026(.A(dpath_mulcore_ary1_a1_I2_I1_25__net046), .Y(n7775));
INVX1 mul_U21027(.A(dpath_mulcore_ary1_a1_I2_I1_24__net046), .Y(n7776));
INVX1 mul_U21028(.A(dpath_mulcore_ary1_a1_I2_I1_23__net046), .Y(n7777));
INVX1 mul_U21029(.A(dpath_mulcore_ary1_a1_I2_I1_22__net046), .Y(n7778));
INVX1 mul_U21030(.A(dpath_mulcore_ary1_a1_I2_I1_21__net046), .Y(n7779));
INVX1 mul_U21031(.A(dpath_mulcore_ary1_a1_I2_I1_20__net046), .Y(n7780));
INVX1 mul_U21032(.A(dpath_mulcore_ary1_a1_I2_I1_19__net046), .Y(n7781));
INVX1 mul_U21033(.A(dpath_mulcore_ary1_a1_I2_I1_18__net046), .Y(n7782));
INVX1 mul_U21034(.A(dpath_mulcore_ary1_a1_I2_I1_17__net046), .Y(n7783));
INVX1 mul_U21035(.A(dpath_mulcore_ary1_a1_I2_I1_16__net046), .Y(n7784));
INVX1 mul_U21036(.A(dpath_mulcore_ary1_a1_I2_I1_15__net046), .Y(n7785));
INVX1 mul_U21037(.A(dpath_mulcore_ary1_a1_I2_I1_14__net046), .Y(n7786));
INVX1 mul_U21038(.A(dpath_mulcore_ary1_a1_I2_I1_13__net046), .Y(n7787));
INVX1 mul_U21039(.A(dpath_mulcore_ary1_a1_I2_I1_12__net046), .Y(n7788));
INVX1 mul_U21040(.A(dpath_mulcore_ary1_a1_I2_I1_11__net046), .Y(n7789));
INVX1 mul_U21041(.A(dpath_mulcore_ary1_a1_I2_I1_10__net046), .Y(n7790));
INVX1 mul_U21042(.A(dpath_mulcore_ary1_a1_I2_I1_9__net046), .Y(n7791));
INVX1 mul_U21043(.A(dpath_mulcore_ary1_a1_I2_I1_8__net046), .Y(n7792));
INVX1 mul_U21044(.A(dpath_mulcore_ary1_a1_I2_I1_7__net046), .Y(n7793));
INVX1 mul_U21045(.A(dpath_mulcore_ary1_a1_I2_I1_6__net046), .Y(n7794));
INVX1 mul_U21046(.A(dpath_mulcore_ary1_a1_I2_I1_5__net046), .Y(n7795));
INVX1 mul_U21047(.A(dpath_mulcore_ary1_a1_I2_I1_4__net046), .Y(n7796));
INVX1 mul_U21048(.A(dpath_mulcore_ary1_a1_I2_I0_p0_3), .Y(n7797));
INVX1 mul_U21049(.A(dpath_mulcore_ary1_a1_I2_I0_p0_2), .Y(n7798));
INVX1 mul_U21050(.A(dpath_mulcore_ary1_a1_I1_I2_net078), .Y(n7799));
INVX1 mul_U21051(.A(dpath_mulcore_ary1_a1_I1_I2_net8), .Y(n7800));
INVX1 mul_U21052(.A(dpath_mulcore_ary1_a1_I1_I2_net15), .Y(n7801));
INVX1 mul_U21053(.A(dpath_mulcore_ary1_a1_I1_I2_net43), .Y(n7802));
INVX1 mul_U21054(.A(dpath_mulcore_ary1_a1_I1_I2_net48), .Y(n7803));
INVX1 mul_U21055(.A(dpath_mulcore_ary1_a1_I1_I2_net35), .Y(n7804));
INVX1 mul_U21056(.A(dpath_mulcore_ary1_a1_I1_I1_63__net043), .Y(n7805));
INVX1 mul_U21057(.A(dpath_mulcore_ary1_a1_I1_I1_63__net046), .Y(n7806));
INVX1 mul_U21058(.A(dpath_mulcore_ary1_a1_I1_I1_62__net043), .Y(n7807));
INVX1 mul_U21059(.A(dpath_mulcore_ary1_a1_I1_I1_62__net046), .Y(n7808));
INVX1 mul_U21060(.A(dpath_mulcore_ary1_a1_I1_I1_61__net043), .Y(n7809));
INVX1 mul_U21061(.A(dpath_mulcore_ary1_a1_I1_I1_61__net046), .Y(n7810));
INVX1 mul_U21062(.A(dpath_mulcore_ary1_a1_I1_I1_60__net043), .Y(n7811));
INVX1 mul_U21063(.A(dpath_mulcore_ary1_a1_I1_I1_60__net046), .Y(n7812));
INVX1 mul_U21064(.A(dpath_mulcore_ary1_a1_I1_I1_59__net043), .Y(n7813));
INVX1 mul_U21065(.A(dpath_mulcore_ary1_a1_I1_I1_59__net046), .Y(n7814));
INVX1 mul_U21066(.A(dpath_mulcore_ary1_a1_I1_I1_58__net043), .Y(n7815));
INVX1 mul_U21067(.A(dpath_mulcore_ary1_a1_I1_I1_58__net046), .Y(n7816));
INVX1 mul_U21068(.A(dpath_mulcore_ary1_a1_I1_I1_57__net043), .Y(n7817));
INVX1 mul_U21069(.A(dpath_mulcore_ary1_a1_I1_I1_57__net046), .Y(n7818));
INVX1 mul_U21070(.A(dpath_mulcore_ary1_a1_I1_I1_56__net043), .Y(n7819));
INVX1 mul_U21071(.A(dpath_mulcore_ary1_a1_I1_I1_56__net046), .Y(n7820));
INVX1 mul_U21072(.A(dpath_mulcore_ary1_a1_I1_I1_55__net043), .Y(n7821));
INVX1 mul_U21073(.A(dpath_mulcore_ary1_a1_I1_I1_55__net046), .Y(n7822));
INVX1 mul_U21074(.A(dpath_mulcore_ary1_a1_I1_I1_54__net043), .Y(n7823));
INVX1 mul_U21075(.A(dpath_mulcore_ary1_a1_I1_I1_54__net046), .Y(n7824));
INVX1 mul_U21076(.A(dpath_mulcore_ary1_a1_I1_I1_53__net043), .Y(n7825));
INVX1 mul_U21077(.A(dpath_mulcore_ary1_a1_I1_I1_53__net046), .Y(n7826));
INVX1 mul_U21078(.A(dpath_mulcore_ary1_a1_I1_I1_52__net043), .Y(n7827));
INVX1 mul_U21079(.A(dpath_mulcore_ary1_a1_I1_I1_52__net046), .Y(n7828));
INVX1 mul_U21080(.A(dpath_mulcore_ary1_a1_I1_I1_51__net043), .Y(n7829));
INVX1 mul_U21081(.A(dpath_mulcore_ary1_a1_I1_I1_51__net046), .Y(n7830));
INVX1 mul_U21082(.A(dpath_mulcore_ary1_a1_I1_I1_50__net043), .Y(n7831));
INVX1 mul_U21083(.A(dpath_mulcore_ary1_a1_I1_I1_50__net046), .Y(n7832));
INVX1 mul_U21084(.A(dpath_mulcore_ary1_a1_I1_I1_49__net043), .Y(n7833));
INVX1 mul_U21085(.A(dpath_mulcore_ary1_a1_I1_I1_49__net046), .Y(n7834));
INVX1 mul_U21086(.A(dpath_mulcore_ary1_a1_I1_I1_48__net043), .Y(n7835));
INVX1 mul_U21087(.A(dpath_mulcore_ary1_a1_I1_I1_48__net046), .Y(n7836));
INVX1 mul_U21088(.A(dpath_mulcore_ary1_a1_I1_I1_47__net043), .Y(n7837));
INVX1 mul_U21089(.A(dpath_mulcore_ary1_a1_I1_I1_47__net046), .Y(n7838));
INVX1 mul_U21090(.A(dpath_mulcore_ary1_a1_I1_I1_46__net043), .Y(n7839));
INVX1 mul_U21091(.A(dpath_mulcore_ary1_a1_I1_I1_46__net046), .Y(n7840));
INVX1 mul_U21092(.A(dpath_mulcore_ary1_a1_I1_I1_45__net043), .Y(n7841));
INVX1 mul_U21093(.A(dpath_mulcore_ary1_a1_I1_I1_45__net046), .Y(n7842));
INVX1 mul_U21094(.A(dpath_mulcore_ary1_a1_I1_I1_44__net043), .Y(n7843));
INVX1 mul_U21095(.A(dpath_mulcore_ary1_a1_I1_I1_44__net046), .Y(n7844));
INVX1 mul_U21096(.A(dpath_mulcore_ary1_a1_I1_I1_43__net043), .Y(n7845));
INVX1 mul_U21097(.A(dpath_mulcore_ary1_a1_I1_I1_43__net046), .Y(n7846));
INVX1 mul_U21098(.A(dpath_mulcore_ary1_a1_I1_I1_42__net043), .Y(n7847));
INVX1 mul_U21099(.A(dpath_mulcore_ary1_a1_I1_I1_42__net046), .Y(n7848));
INVX1 mul_U21100(.A(dpath_mulcore_ary1_a1_I1_I1_41__net043), .Y(n7849));
INVX1 mul_U21101(.A(dpath_mulcore_ary1_a1_I1_I1_41__net046), .Y(n7850));
INVX1 mul_U21102(.A(dpath_mulcore_ary1_a1_I1_I1_40__net043), .Y(n7851));
INVX1 mul_U21103(.A(dpath_mulcore_ary1_a1_I1_I1_40__net046), .Y(n7852));
INVX1 mul_U21104(.A(dpath_mulcore_ary1_a1_I1_I1_39__net043), .Y(n7853));
INVX1 mul_U21105(.A(dpath_mulcore_ary1_a1_I1_I1_39__net046), .Y(n7854));
INVX1 mul_U21106(.A(dpath_mulcore_ary1_a1_I1_I1_38__net043), .Y(n7855));
INVX1 mul_U21107(.A(dpath_mulcore_ary1_a1_I1_I1_38__net046), .Y(n7856));
INVX1 mul_U21108(.A(dpath_mulcore_ary1_a1_I1_I1_37__net043), .Y(n7857));
INVX1 mul_U21109(.A(dpath_mulcore_ary1_a1_I1_I1_37__net046), .Y(n7858));
INVX1 mul_U21110(.A(dpath_mulcore_ary1_a1_I1_I1_36__net043), .Y(n7859));
INVX1 mul_U21111(.A(dpath_mulcore_ary1_a1_I1_I1_36__net046), .Y(n7860));
INVX1 mul_U21112(.A(dpath_mulcore_ary1_a1_I1_I1_35__net043), .Y(n7861));
INVX1 mul_U21113(.A(dpath_mulcore_ary1_a1_I1_I1_35__net046), .Y(n7862));
INVX1 mul_U21114(.A(dpath_mulcore_ary1_a1_I1_I1_34__net043), .Y(n7863));
INVX1 mul_U21115(.A(dpath_mulcore_ary1_a1_I1_I1_34__net046), .Y(n7864));
INVX1 mul_U21116(.A(dpath_mulcore_ary1_a1_I1_I1_33__net043), .Y(n7865));
INVX1 mul_U21117(.A(dpath_mulcore_ary1_a1_I1_I1_33__net046), .Y(n7866));
INVX1 mul_U21118(.A(dpath_mulcore_ary1_a1_I1_I1_32__net043), .Y(n7867));
INVX1 mul_U21119(.A(dpath_mulcore_ary1_a1_I1_I1_32__net046), .Y(n7868));
INVX1 mul_U21120(.A(dpath_mulcore_ary1_a1_I1_I1_31__net043), .Y(n7869));
INVX1 mul_U21121(.A(dpath_mulcore_ary1_a1_I1_I1_31__net046), .Y(n7870));
INVX1 mul_U21122(.A(dpath_mulcore_ary1_a1_I1_I1_30__net043), .Y(n7871));
INVX1 mul_U21123(.A(dpath_mulcore_ary1_a1_I1_I1_30__net046), .Y(n7872));
INVX1 mul_U21124(.A(dpath_mulcore_ary1_a1_I1_I1_29__net043), .Y(n7873));
INVX1 mul_U21125(.A(dpath_mulcore_ary1_a1_I1_I1_29__net046), .Y(n7874));
INVX1 mul_U21126(.A(dpath_mulcore_ary1_a1_I1_I1_28__net043), .Y(n7875));
INVX1 mul_U21127(.A(dpath_mulcore_ary1_a1_I1_I1_28__net046), .Y(n7876));
INVX1 mul_U21128(.A(dpath_mulcore_ary1_a1_I1_I1_27__net043), .Y(n7877));
INVX1 mul_U21129(.A(dpath_mulcore_ary1_a1_I1_I1_27__net046), .Y(n7878));
INVX1 mul_U21130(.A(dpath_mulcore_ary1_a1_I1_I1_26__net043), .Y(n7879));
INVX1 mul_U21131(.A(dpath_mulcore_ary1_a1_I1_I1_26__net046), .Y(n7880));
INVX1 mul_U21132(.A(dpath_mulcore_ary1_a1_I1_I1_25__net043), .Y(n7881));
INVX1 mul_U21133(.A(dpath_mulcore_ary1_a1_I1_I1_25__net046), .Y(n7882));
INVX1 mul_U21134(.A(dpath_mulcore_ary1_a1_I1_I1_24__net043), .Y(n7883));
INVX1 mul_U21135(.A(dpath_mulcore_ary1_a1_I1_I1_24__net046), .Y(n7884));
INVX1 mul_U21136(.A(dpath_mulcore_ary1_a1_I1_I1_23__net043), .Y(n7885));
INVX1 mul_U21137(.A(dpath_mulcore_ary1_a1_I1_I1_23__net046), .Y(n7886));
INVX1 mul_U21138(.A(dpath_mulcore_ary1_a1_I1_I1_22__net043), .Y(n7887));
INVX1 mul_U21139(.A(dpath_mulcore_ary1_a1_I1_I1_22__net046), .Y(n7888));
INVX1 mul_U21140(.A(dpath_mulcore_ary1_a1_I1_I1_21__net043), .Y(n7889));
INVX1 mul_U21141(.A(dpath_mulcore_ary1_a1_I1_I1_21__net046), .Y(n7890));
INVX1 mul_U21142(.A(dpath_mulcore_ary1_a1_I1_I1_20__net043), .Y(n7891));
INVX1 mul_U21143(.A(dpath_mulcore_ary1_a1_I1_I1_20__net046), .Y(n7892));
INVX1 mul_U21144(.A(dpath_mulcore_ary1_a1_I1_I1_19__net043), .Y(n7893));
INVX1 mul_U21145(.A(dpath_mulcore_ary1_a1_I1_I1_19__net046), .Y(n7894));
INVX1 mul_U21146(.A(dpath_mulcore_ary1_a1_I1_I1_18__net043), .Y(n7895));
INVX1 mul_U21147(.A(dpath_mulcore_ary1_a1_I1_I1_18__net046), .Y(n7896));
INVX1 mul_U21148(.A(dpath_mulcore_ary1_a1_I1_I1_17__net043), .Y(n7897));
INVX1 mul_U21149(.A(dpath_mulcore_ary1_a1_I1_I1_17__net046), .Y(n7898));
INVX1 mul_U21150(.A(dpath_mulcore_ary1_a1_I1_I1_16__net043), .Y(n7899));
INVX1 mul_U21151(.A(dpath_mulcore_ary1_a1_I1_I1_16__net046), .Y(n7900));
INVX1 mul_U21152(.A(dpath_mulcore_ary1_a1_I1_I1_15__net043), .Y(n7901));
INVX1 mul_U21153(.A(dpath_mulcore_ary1_a1_I1_I1_15__net046), .Y(n7902));
INVX1 mul_U21154(.A(dpath_mulcore_ary1_a1_I1_I1_14__net043), .Y(n7903));
INVX1 mul_U21155(.A(dpath_mulcore_ary1_a1_I1_I1_14__net046), .Y(n7904));
INVX1 mul_U21156(.A(dpath_mulcore_ary1_a1_I1_I1_13__net043), .Y(n7905));
INVX1 mul_U21157(.A(dpath_mulcore_ary1_a1_I1_I1_13__net046), .Y(n7906));
INVX1 mul_U21158(.A(dpath_mulcore_ary1_a1_I1_I1_12__net043), .Y(n7907));
INVX1 mul_U21159(.A(dpath_mulcore_ary1_a1_I1_I1_12__net046), .Y(n7908));
INVX1 mul_U21160(.A(dpath_mulcore_ary1_a1_I1_I1_11__net043), .Y(n7909));
INVX1 mul_U21161(.A(dpath_mulcore_ary1_a1_I1_I1_11__net046), .Y(n7910));
INVX1 mul_U21162(.A(dpath_mulcore_ary1_a1_I1_I1_10__net043), .Y(n7911));
INVX1 mul_U21163(.A(dpath_mulcore_ary1_a1_I1_I1_10__net046), .Y(n7912));
INVX1 mul_U21164(.A(dpath_mulcore_ary1_a1_I1_I1_9__net043), .Y(n7913));
INVX1 mul_U21165(.A(dpath_mulcore_ary1_a1_I1_I1_9__net046), .Y(n7914));
INVX1 mul_U21166(.A(dpath_mulcore_ary1_a1_I1_I1_8__net043), .Y(n7915));
INVX1 mul_U21167(.A(dpath_mulcore_ary1_a1_I1_I1_8__net046), .Y(n7916));
INVX1 mul_U21168(.A(dpath_mulcore_ary1_a1_I1_I1_7__net043), .Y(n7917));
INVX1 mul_U21169(.A(dpath_mulcore_ary1_a1_I1_I1_7__net046), .Y(n7918));
INVX1 mul_U21170(.A(dpath_mulcore_ary1_a1_I1_I1_6__net043), .Y(n7919));
INVX1 mul_U21171(.A(dpath_mulcore_ary1_a1_I1_I1_6__net046), .Y(n7920));
INVX1 mul_U21172(.A(dpath_mulcore_ary1_a1_I1_I1_5__net043), .Y(n7921));
INVX1 mul_U21173(.A(dpath_mulcore_ary1_a1_I1_I1_5__net046), .Y(n7922));
INVX1 mul_U21174(.A(dpath_mulcore_ary1_a1_I1_I1_4__net046), .Y(n7923));
INVX1 mul_U21175(.A(dpath_mulcore_ary1_a1_I1_I0_p0_3), .Y(n7924));
INVX1 mul_U21176(.A(dpath_mulcore_ary1_a1_I1_I0_p0_2), .Y(n7925));
INVX1 mul_U21177(.A(dpath_mulcore_ary1_a1_I0_I2_net078), .Y(n7926));
INVX1 mul_U21178(.A(dpath_mulcore_ary1_a1_I0_I2_net8), .Y(n7927));
INVX1 mul_U21179(.A(dpath_mulcore_ary1_a1_I0_I2_net15), .Y(n7928));
INVX1 mul_U21180(.A(dpath_mulcore_ary1_a1_I0_I2_net43), .Y(n7929));
INVX1 mul_U21181(.A(dpath_mulcore_ary1_a1_I0_I2_net48), .Y(n7930));
INVX1 mul_U21182(.A(dpath_mulcore_ary1_a1_I0_I2_net35), .Y(n7931));
INVX1 mul_U21183(.A(dpath_mulcore_ary1_a1_I0_I1_63__net043), .Y(n7932));
INVX1 mul_U21184(.A(dpath_mulcore_ary1_a1_I0_I1_63__net046), .Y(n7933));
INVX1 mul_U21185(.A(dpath_mulcore_ary1_a1_I0_I1_62__net043), .Y(n7934));
INVX1 mul_U21186(.A(dpath_mulcore_ary1_a1_I0_I1_62__net046), .Y(n7935));
INVX1 mul_U21187(.A(dpath_mulcore_ary1_a1_I0_I1_61__net043), .Y(n7936));
INVX1 mul_U21188(.A(dpath_mulcore_ary1_a1_I0_I1_61__net046), .Y(n7937));
INVX1 mul_U21189(.A(dpath_mulcore_ary1_a1_I0_I1_60__net043), .Y(n7938));
INVX1 mul_U21190(.A(dpath_mulcore_ary1_a1_I0_I1_60__net046), .Y(n7939));
INVX1 mul_U21191(.A(dpath_mulcore_ary1_a1_I0_I1_59__net043), .Y(n7940));
INVX1 mul_U21192(.A(dpath_mulcore_ary1_a1_I0_I1_59__net046), .Y(n7941));
INVX1 mul_U21193(.A(dpath_mulcore_ary1_a1_I0_I1_58__net043), .Y(n7942));
INVX1 mul_U21194(.A(dpath_mulcore_ary1_a1_I0_I1_58__net046), .Y(n7943));
INVX1 mul_U21195(.A(dpath_mulcore_ary1_a1_I0_I1_57__net043), .Y(n7944));
INVX1 mul_U21196(.A(dpath_mulcore_ary1_a1_I0_I1_57__net046), .Y(n7945));
INVX1 mul_U21197(.A(dpath_mulcore_ary1_a1_I0_I1_56__net043), .Y(n7946));
INVX1 mul_U21198(.A(dpath_mulcore_ary1_a1_I0_I1_56__net046), .Y(n7947));
INVX1 mul_U21199(.A(dpath_mulcore_ary1_a1_I0_I1_55__net043), .Y(n7948));
INVX1 mul_U21200(.A(dpath_mulcore_ary1_a1_I0_I1_55__net046), .Y(n7949));
INVX1 mul_U21201(.A(dpath_mulcore_ary1_a1_I0_I1_54__net043), .Y(n7950));
INVX1 mul_U21202(.A(dpath_mulcore_ary1_a1_I0_I1_54__net046), .Y(n7951));
INVX1 mul_U21203(.A(dpath_mulcore_ary1_a1_I0_I1_53__net043), .Y(n7952));
INVX1 mul_U21204(.A(dpath_mulcore_ary1_a1_I0_I1_53__net046), .Y(n7953));
INVX1 mul_U21205(.A(dpath_mulcore_ary1_a1_I0_I1_52__net043), .Y(n7954));
INVX1 mul_U21206(.A(dpath_mulcore_ary1_a1_I0_I1_52__net046), .Y(n7955));
INVX1 mul_U21207(.A(dpath_mulcore_ary1_a1_I0_I1_51__net043), .Y(n7956));
INVX1 mul_U21208(.A(dpath_mulcore_ary1_a1_I0_I1_51__net046), .Y(n7957));
INVX1 mul_U21209(.A(dpath_mulcore_ary1_a1_I0_I1_50__net043), .Y(n7958));
INVX1 mul_U21210(.A(dpath_mulcore_ary1_a1_I0_I1_50__net046), .Y(n7959));
INVX1 mul_U21211(.A(dpath_mulcore_ary1_a1_I0_I1_49__net043), .Y(n7960));
INVX1 mul_U21212(.A(dpath_mulcore_ary1_a1_I0_I1_49__net046), .Y(n7961));
INVX1 mul_U21213(.A(dpath_mulcore_ary1_a1_I0_I1_48__net043), .Y(n7962));
INVX1 mul_U21214(.A(dpath_mulcore_ary1_a1_I0_I1_48__net046), .Y(n7963));
INVX1 mul_U21215(.A(dpath_mulcore_ary1_a1_I0_I1_47__net043), .Y(n7964));
INVX1 mul_U21216(.A(dpath_mulcore_ary1_a1_I0_I1_47__net046), .Y(n7965));
INVX1 mul_U21217(.A(dpath_mulcore_ary1_a1_I0_I1_46__net043), .Y(n7966));
INVX1 mul_U21218(.A(dpath_mulcore_ary1_a1_I0_I1_46__net046), .Y(n7967));
INVX1 mul_U21219(.A(dpath_mulcore_ary1_a1_I0_I1_45__net043), .Y(n7968));
INVX1 mul_U21220(.A(dpath_mulcore_ary1_a1_I0_I1_45__net046), .Y(n7969));
INVX1 mul_U21221(.A(dpath_mulcore_ary1_a1_I0_I1_44__net043), .Y(n7970));
INVX1 mul_U21222(.A(dpath_mulcore_ary1_a1_I0_I1_44__net046), .Y(n7971));
INVX1 mul_U21223(.A(dpath_mulcore_ary1_a1_I0_I1_43__net043), .Y(n7972));
INVX1 mul_U21224(.A(dpath_mulcore_ary1_a1_I0_I1_43__net046), .Y(n7973));
INVX1 mul_U21225(.A(dpath_mulcore_ary1_a1_I0_I1_42__net043), .Y(n7974));
INVX1 mul_U21226(.A(dpath_mulcore_ary1_a1_I0_I1_42__net046), .Y(n7975));
INVX1 mul_U21227(.A(dpath_mulcore_ary1_a1_I0_I1_41__net043), .Y(n7976));
INVX1 mul_U21228(.A(dpath_mulcore_ary1_a1_I0_I1_41__net046), .Y(n7977));
INVX1 mul_U21229(.A(dpath_mulcore_ary1_a1_I0_I1_40__net043), .Y(n7978));
INVX1 mul_U21230(.A(dpath_mulcore_ary1_a1_I0_I1_40__net046), .Y(n7979));
INVX1 mul_U21231(.A(dpath_mulcore_ary1_a1_I0_I1_39__net043), .Y(n7980));
INVX1 mul_U21232(.A(dpath_mulcore_ary1_a1_I0_I1_39__net046), .Y(n7981));
INVX1 mul_U21233(.A(dpath_mulcore_ary1_a1_I0_I1_38__net043), .Y(n7982));
INVX1 mul_U21234(.A(dpath_mulcore_ary1_a1_I0_I1_38__net046), .Y(n7983));
INVX1 mul_U21235(.A(dpath_mulcore_ary1_a1_I0_I1_37__net043), .Y(n7984));
INVX1 mul_U21236(.A(dpath_mulcore_ary1_a1_I0_I1_37__net046), .Y(n7985));
INVX1 mul_U21237(.A(dpath_mulcore_ary1_a1_I0_I1_36__net043), .Y(n7986));
INVX1 mul_U21238(.A(dpath_mulcore_ary1_a1_I0_I1_36__net046), .Y(n7987));
INVX1 mul_U21239(.A(dpath_mulcore_ary1_a1_I0_I1_35__net043), .Y(n7988));
INVX1 mul_U21240(.A(dpath_mulcore_ary1_a1_I0_I1_35__net046), .Y(n7989));
INVX1 mul_U21241(.A(dpath_mulcore_ary1_a1_I0_I1_34__net043), .Y(n7990));
INVX1 mul_U21242(.A(dpath_mulcore_ary1_a1_I0_I1_34__net046), .Y(n7991));
INVX1 mul_U21243(.A(dpath_mulcore_ary1_a1_I0_I1_33__net043), .Y(n7992));
INVX1 mul_U21244(.A(dpath_mulcore_ary1_a1_I0_I1_33__net046), .Y(n7993));
INVX1 mul_U21245(.A(dpath_mulcore_ary1_a1_I0_I1_32__net043), .Y(n7994));
INVX1 mul_U21246(.A(dpath_mulcore_ary1_a1_I0_I1_32__net046), .Y(n7995));
INVX1 mul_U21247(.A(dpath_mulcore_ary1_a1_I0_I1_31__net043), .Y(n7996));
INVX1 mul_U21248(.A(dpath_mulcore_ary1_a1_I0_I1_31__net046), .Y(n7997));
INVX1 mul_U21249(.A(dpath_mulcore_ary1_a1_I0_I1_30__net043), .Y(n7998));
INVX1 mul_U21250(.A(dpath_mulcore_ary1_a1_I0_I1_30__net046), .Y(n7999));
INVX1 mul_U21251(.A(dpath_mulcore_ary1_a1_I0_I1_29__net043), .Y(n8000));
INVX1 mul_U21252(.A(dpath_mulcore_ary1_a1_I0_I1_29__net046), .Y(n8001));
INVX1 mul_U21253(.A(dpath_mulcore_ary1_a1_I0_I1_28__net043), .Y(n8002));
INVX1 mul_U21254(.A(dpath_mulcore_ary1_a1_I0_I1_28__net046), .Y(n8003));
INVX1 mul_U21255(.A(dpath_mulcore_ary1_a1_I0_I1_27__net043), .Y(n8004));
INVX1 mul_U21256(.A(dpath_mulcore_ary1_a1_I0_I1_27__net046), .Y(n8005));
INVX1 mul_U21257(.A(dpath_mulcore_ary1_a1_I0_I1_26__net043), .Y(n8006));
INVX1 mul_U21258(.A(dpath_mulcore_ary1_a1_I0_I1_26__net046), .Y(n8007));
INVX1 mul_U21259(.A(dpath_mulcore_ary1_a1_I0_I1_25__net043), .Y(n8008));
INVX1 mul_U21260(.A(dpath_mulcore_ary1_a1_I0_I1_25__net046), .Y(n8009));
INVX1 mul_U21261(.A(dpath_mulcore_ary1_a1_I0_I1_24__net043), .Y(n8010));
INVX1 mul_U21262(.A(dpath_mulcore_ary1_a1_I0_I1_24__net046), .Y(n8011));
INVX1 mul_U21263(.A(dpath_mulcore_ary1_a1_I0_I1_23__net043), .Y(n8012));
INVX1 mul_U21264(.A(dpath_mulcore_ary1_a1_I0_I1_23__net046), .Y(n8013));
INVX1 mul_U21265(.A(dpath_mulcore_ary1_a1_I0_I1_22__net043), .Y(n8014));
INVX1 mul_U21266(.A(dpath_mulcore_ary1_a1_I0_I1_22__net046), .Y(n8015));
INVX1 mul_U21267(.A(dpath_mulcore_ary1_a1_I0_I1_21__net043), .Y(n8016));
INVX1 mul_U21268(.A(dpath_mulcore_ary1_a1_I0_I1_21__net046), .Y(n8017));
INVX1 mul_U21269(.A(dpath_mulcore_ary1_a1_I0_I1_20__net043), .Y(n8018));
INVX1 mul_U21270(.A(dpath_mulcore_ary1_a1_I0_I1_20__net046), .Y(n8019));
INVX1 mul_U21271(.A(dpath_mulcore_ary1_a1_I0_I1_19__net043), .Y(n8020));
INVX1 mul_U21272(.A(dpath_mulcore_ary1_a1_I0_I1_19__net046), .Y(n8021));
INVX1 mul_U21273(.A(dpath_mulcore_ary1_a1_I0_I1_18__net043), .Y(n8022));
INVX1 mul_U21274(.A(dpath_mulcore_ary1_a1_I0_I1_18__net046), .Y(n8023));
INVX1 mul_U21275(.A(dpath_mulcore_ary1_a1_I0_I1_17__net043), .Y(n8024));
INVX1 mul_U21276(.A(dpath_mulcore_ary1_a1_I0_I1_17__net046), .Y(n8025));
INVX1 mul_U21277(.A(dpath_mulcore_ary1_a1_I0_I1_16__net043), .Y(n8026));
INVX1 mul_U21278(.A(dpath_mulcore_ary1_a1_I0_I1_16__net046), .Y(n8027));
INVX1 mul_U21279(.A(dpath_mulcore_ary1_a1_I0_I1_15__net043), .Y(n8028));
INVX1 mul_U21280(.A(dpath_mulcore_ary1_a1_I0_I1_15__net046), .Y(n8029));
INVX1 mul_U21281(.A(dpath_mulcore_ary1_a1_I0_I1_14__net043), .Y(n8030));
INVX1 mul_U21282(.A(dpath_mulcore_ary1_a1_I0_I1_14__net046), .Y(n8031));
INVX1 mul_U21283(.A(dpath_mulcore_ary1_a1_I0_I1_13__net043), .Y(n8032));
INVX1 mul_U21284(.A(dpath_mulcore_ary1_a1_I0_I1_13__net046), .Y(n8033));
INVX1 mul_U21285(.A(dpath_mulcore_ary1_a1_I0_I1_12__net043), .Y(n8034));
INVX1 mul_U21286(.A(dpath_mulcore_ary1_a1_I0_I1_12__net046), .Y(n8035));
INVX1 mul_U21287(.A(dpath_mulcore_ary1_a1_I0_I1_11__net043), .Y(n8036));
INVX1 mul_U21288(.A(dpath_mulcore_ary1_a1_I0_I1_11__net046), .Y(n8037));
INVX1 mul_U21289(.A(dpath_mulcore_ary1_a1_I0_I1_10__net043), .Y(n8038));
INVX1 mul_U21290(.A(dpath_mulcore_ary1_a1_I0_I1_10__net046), .Y(n8039));
INVX1 mul_U21291(.A(dpath_mulcore_ary1_a1_I0_I1_9__net043), .Y(n8040));
INVX1 mul_U21292(.A(dpath_mulcore_ary1_a1_I0_I1_9__net046), .Y(n8041));
INVX1 mul_U21293(.A(dpath_mulcore_ary1_a1_I0_I1_8__net043), .Y(n8042));
INVX1 mul_U21294(.A(dpath_mulcore_ary1_a1_I0_I1_8__net046), .Y(n8043));
INVX1 mul_U21295(.A(dpath_mulcore_ary1_a1_I0_I1_7__net043), .Y(n8044));
INVX1 mul_U21296(.A(dpath_mulcore_ary1_a1_I0_I1_7__net046), .Y(n8045));
INVX1 mul_U21297(.A(dpath_mulcore_ary1_a1_I0_I1_6__net043), .Y(n8046));
INVX1 mul_U21298(.A(dpath_mulcore_ary1_a1_I0_I1_6__net046), .Y(n8047));
INVX1 mul_U21299(.A(dpath_mulcore_ary1_a1_I0_I1_5__net043), .Y(n8048));
INVX1 mul_U21300(.A(dpath_mulcore_ary1_a1_I0_I1_5__net046), .Y(n8049));
INVX1 mul_U21301(.A(dpath_mulcore_ary1_a1_I0_I1_4__net046), .Y(n8050));
INVX1 mul_U21302(.A(dpath_mulcore_ary1_a1_I0_I0_p0_3), .Y(n8051));
INVX1 mul_U21303(.A(dpath_mulcore_ary1_a1_I0_I0_p0_2), .Y(n8052));
INVX1 mul_U21304(.A(dpath_mulcore_ary1_a0_I0_I2_net38), .Y(n8053));
INVX1 mul_U21305(.A(dpath_mulcore_ary1_a0_I1_I0_b1n_0), .Y(n8054));
INVX1 mul_U21306(.A(dpath_mulcore_ary1_a0_I1_I0_b1n_1), .Y(n8055));
INVX1 mul_U21307(.A(dpath_mulcore_ary1_a0_c1[3]), .Y(n8056));
INVX1 mul_U21308(.A(dpath_mulcore_ary1_a0_c1[2]), .Y(n8057));
INVX1 mul_U21309(.A(dpath_mulcore_ary1_a0_I0_I0_b1n_0), .Y(n8058));
INVX1 mul_U21310(.A(dpath_mulcore_ary1_a0_I0_I0_b1n_1), .Y(n8059));
INVX1 mul_U21311(.A(dpath_mulcore_ary1_a1_I2_I0_b1n_0), .Y(n8060));
INVX1 mul_U21312(.A(dpath_mulcore_ary1_a1_I2_I0_b1n_1), .Y(n8061));
INVX1 mul_U21313(.A(dpath_mulcore_ary1_a1_I1_I0_b1n_0), .Y(n8062));
INVX1 mul_U21314(.A(dpath_mulcore_ary1_a1_I1_I0_b1n_1), .Y(n8063));
INVX1 mul_U21315(.A(dpath_mulcore_ary1_a1_c1[3]), .Y(n8064));
INVX1 mul_U21316(.A(dpath_mulcore_ary1_a1_c1[2]), .Y(n8065));
INVX1 mul_U21317(.A(dpath_mulcore_ary1_a1_I0_I0_b1n_0), .Y(n8066));
INVX1 mul_U21318(.A(dpath_mulcore_ary1_a1_I0_I0_b1n_1), .Y(n8067));
INVX1 mul_U21319(.A(dpath_mulcore_ary1_a0_c1[63]), .Y(n8068));
INVX1 mul_U21320(.A(dpath_mulcore_ary1_a0_c1[62]), .Y(n8069));
INVX1 mul_U21321(.A(dpath_mulcore_ary1_a0_c1[61]), .Y(n8070));
INVX1 mul_U21322(.A(dpath_mulcore_ary1_a0_c1[60]), .Y(n8071));
INVX1 mul_U21323(.A(dpath_mulcore_ary1_a0_c1[59]), .Y(n8072));
INVX1 mul_U21324(.A(dpath_mulcore_ary1_a0_c1[58]), .Y(n8073));
INVX1 mul_U21325(.A(dpath_mulcore_ary1_a0_c1[57]), .Y(n8074));
INVX1 mul_U21326(.A(dpath_mulcore_ary1_a0_c1[56]), .Y(n8075));
INVX1 mul_U21327(.A(dpath_mulcore_ary1_a0_c1[55]), .Y(n8076));
INVX1 mul_U21328(.A(dpath_mulcore_ary1_a0_c1[54]), .Y(n8077));
INVX1 mul_U21329(.A(dpath_mulcore_ary1_a0_c1[53]), .Y(n8078));
INVX1 mul_U21330(.A(dpath_mulcore_ary1_a0_c1[52]), .Y(n8079));
INVX1 mul_U21331(.A(dpath_mulcore_ary1_a0_c1[51]), .Y(n8080));
INVX1 mul_U21332(.A(dpath_mulcore_ary1_a0_c1[50]), .Y(n8081));
INVX1 mul_U21333(.A(dpath_mulcore_ary1_a0_c1[49]), .Y(n8082));
INVX1 mul_U21334(.A(dpath_mulcore_ary1_a0_c1[48]), .Y(n8083));
INVX1 mul_U21335(.A(dpath_mulcore_ary1_a0_c1[47]), .Y(n8084));
INVX1 mul_U21336(.A(dpath_mulcore_ary1_a0_c1[46]), .Y(n8085));
INVX1 mul_U21337(.A(dpath_mulcore_ary1_a0_c1[45]), .Y(n8086));
INVX1 mul_U21338(.A(dpath_mulcore_ary1_a0_c1[44]), .Y(n8087));
INVX1 mul_U21339(.A(dpath_mulcore_ary1_a0_c1[43]), .Y(n8088));
INVX1 mul_U21340(.A(dpath_mulcore_ary1_a0_c1[42]), .Y(n8089));
INVX1 mul_U21341(.A(dpath_mulcore_ary1_a0_c1[41]), .Y(n8090));
INVX1 mul_U21342(.A(dpath_mulcore_ary1_a0_c1[40]), .Y(n8091));
INVX1 mul_U21343(.A(dpath_mulcore_ary1_a0_c1[39]), .Y(n8092));
INVX1 mul_U21344(.A(dpath_mulcore_ary1_a0_c1[38]), .Y(n8093));
INVX1 mul_U21345(.A(dpath_mulcore_ary1_a0_c1[37]), .Y(n8094));
INVX1 mul_U21346(.A(dpath_mulcore_ary1_a0_c1[36]), .Y(n8095));
INVX1 mul_U21347(.A(dpath_mulcore_ary1_a0_c1[35]), .Y(n8096));
INVX1 mul_U21348(.A(dpath_mulcore_ary1_a0_c1[34]), .Y(n8097));
INVX1 mul_U21349(.A(dpath_mulcore_ary1_a0_c1[33]), .Y(n8098));
INVX1 mul_U21350(.A(dpath_mulcore_ary1_a0_c1[32]), .Y(n8099));
INVX1 mul_U21351(.A(dpath_mulcore_ary1_a0_c1[31]), .Y(n8100));
INVX1 mul_U21352(.A(dpath_mulcore_ary1_a0_c1[30]), .Y(n8101));
INVX1 mul_U21353(.A(dpath_mulcore_ary1_a0_c1[29]), .Y(n8102));
INVX1 mul_U21354(.A(dpath_mulcore_ary1_a0_c1[28]), .Y(n8103));
INVX1 mul_U21355(.A(dpath_mulcore_ary1_a0_c1[27]), .Y(n8104));
INVX1 mul_U21356(.A(dpath_mulcore_ary1_a0_c1[26]), .Y(n8105));
INVX1 mul_U21357(.A(dpath_mulcore_ary1_a0_c1[25]), .Y(n8106));
INVX1 mul_U21358(.A(dpath_mulcore_ary1_a0_c1[24]), .Y(n8107));
INVX1 mul_U21359(.A(dpath_mulcore_ary1_a0_c1[23]), .Y(n8108));
INVX1 mul_U21360(.A(dpath_mulcore_ary1_a0_c1[22]), .Y(n8109));
INVX1 mul_U21361(.A(dpath_mulcore_ary1_a0_c1[21]), .Y(n8110));
INVX1 mul_U21362(.A(dpath_mulcore_ary1_a0_c1[20]), .Y(n8111));
INVX1 mul_U21363(.A(dpath_mulcore_ary1_a0_c1[19]), .Y(n8112));
INVX1 mul_U21364(.A(dpath_mulcore_ary1_a0_c1[18]), .Y(n8113));
INVX1 mul_U21365(.A(dpath_mulcore_ary1_a0_c1[17]), .Y(n8114));
INVX1 mul_U21366(.A(dpath_mulcore_ary1_a0_c1[16]), .Y(n8115));
INVX1 mul_U21367(.A(dpath_mulcore_ary1_a0_c1[15]), .Y(n8116));
INVX1 mul_U21368(.A(dpath_mulcore_ary1_a0_c1[14]), .Y(n8117));
INVX1 mul_U21369(.A(dpath_mulcore_ary1_a0_c1[13]), .Y(n8118));
INVX1 mul_U21370(.A(dpath_mulcore_ary1_a0_c1[12]), .Y(n8119));
INVX1 mul_U21371(.A(dpath_mulcore_ary1_a0_c1[11]), .Y(n8120));
INVX1 mul_U21372(.A(dpath_mulcore_ary1_a0_c1[10]), .Y(n8121));
INVX1 mul_U21373(.A(dpath_mulcore_ary1_a0_c1[9]), .Y(n8122));
INVX1 mul_U21374(.A(dpath_mulcore_ary1_a0_c1[8]), .Y(n8123));
INVX1 mul_U21375(.A(dpath_mulcore_ary1_a0_c1[7]), .Y(n8124));
INVX1 mul_U21376(.A(dpath_mulcore_ary1_a0_c1[6]), .Y(n8125));
INVX1 mul_U21377(.A(dpath_mulcore_ary1_a0_c1[5]), .Y(n8126));
INVX1 mul_U21378(.A(dpath_mulcore_ary1_a0_c1[4]), .Y(n8127));
INVX1 mul_U21379(.A(dpath_mulcore_ary1_a1_c1[63]), .Y(n8128));
INVX1 mul_U21380(.A(dpath_mulcore_ary1_a1_c1[62]), .Y(n8129));
INVX1 mul_U21381(.A(dpath_mulcore_ary1_a1_c1[61]), .Y(n8130));
INVX1 mul_U21382(.A(dpath_mulcore_ary1_a1_c1[60]), .Y(n8131));
INVX1 mul_U21383(.A(dpath_mulcore_ary1_a1_c1[59]), .Y(n8132));
INVX1 mul_U21384(.A(dpath_mulcore_ary1_a1_c1[58]), .Y(n8133));
INVX1 mul_U21385(.A(dpath_mulcore_ary1_a1_c1[57]), .Y(n8134));
INVX1 mul_U21386(.A(dpath_mulcore_ary1_a1_c1[56]), .Y(n8135));
INVX1 mul_U21387(.A(dpath_mulcore_ary1_a1_c1[55]), .Y(n8136));
INVX1 mul_U21388(.A(dpath_mulcore_ary1_a1_c1[54]), .Y(n8137));
INVX1 mul_U21389(.A(dpath_mulcore_ary1_a1_c1[53]), .Y(n8138));
INVX1 mul_U21390(.A(dpath_mulcore_ary1_a1_c1[52]), .Y(n8139));
INVX1 mul_U21391(.A(dpath_mulcore_ary1_a1_c1[51]), .Y(n8140));
INVX1 mul_U21392(.A(dpath_mulcore_ary1_a1_c1[50]), .Y(n8141));
INVX1 mul_U21393(.A(dpath_mulcore_ary1_a1_c1[49]), .Y(n8142));
INVX1 mul_U21394(.A(dpath_mulcore_ary1_a1_c1[48]), .Y(n8143));
INVX1 mul_U21395(.A(dpath_mulcore_ary1_a1_c1[47]), .Y(n8144));
INVX1 mul_U21396(.A(dpath_mulcore_ary1_a1_c1[46]), .Y(n8145));
INVX1 mul_U21397(.A(dpath_mulcore_ary1_a1_c1[45]), .Y(n8146));
INVX1 mul_U21398(.A(dpath_mulcore_ary1_a1_c1[44]), .Y(n8147));
INVX1 mul_U21399(.A(dpath_mulcore_ary1_a1_c1[43]), .Y(n8148));
INVX1 mul_U21400(.A(dpath_mulcore_ary1_a1_c1[42]), .Y(n8149));
INVX1 mul_U21401(.A(dpath_mulcore_ary1_a1_c1[41]), .Y(n8150));
INVX1 mul_U21402(.A(dpath_mulcore_ary1_a1_c1[40]), .Y(n8151));
INVX1 mul_U21403(.A(dpath_mulcore_ary1_a1_c1[39]), .Y(n8152));
INVX1 mul_U21404(.A(dpath_mulcore_ary1_a1_c1[38]), .Y(n8153));
INVX1 mul_U21405(.A(dpath_mulcore_ary1_a1_c1[37]), .Y(n8154));
INVX1 mul_U21406(.A(dpath_mulcore_ary1_a1_c1[36]), .Y(n8155));
INVX1 mul_U21407(.A(dpath_mulcore_ary1_a1_c1[35]), .Y(n8156));
INVX1 mul_U21408(.A(dpath_mulcore_ary1_a1_c1[34]), .Y(n8157));
INVX1 mul_U21409(.A(dpath_mulcore_ary1_a1_c1[33]), .Y(n8158));
INVX1 mul_U21410(.A(dpath_mulcore_ary1_a1_c1[32]), .Y(n8159));
INVX1 mul_U21411(.A(dpath_mulcore_ary1_a1_c1[31]), .Y(n8160));
INVX1 mul_U21412(.A(dpath_mulcore_ary1_a1_c1[30]), .Y(n8161));
INVX1 mul_U21413(.A(dpath_mulcore_ary1_a1_c1[29]), .Y(n8162));
INVX1 mul_U21414(.A(dpath_mulcore_ary1_a1_c1[28]), .Y(n8163));
INVX1 mul_U21415(.A(dpath_mulcore_ary1_a1_c1[27]), .Y(n8164));
INVX1 mul_U21416(.A(dpath_mulcore_ary1_a1_c1[26]), .Y(n8165));
INVX1 mul_U21417(.A(dpath_mulcore_ary1_a1_c1[25]), .Y(n8166));
INVX1 mul_U21418(.A(dpath_mulcore_ary1_a1_c1[24]), .Y(n8167));
INVX1 mul_U21419(.A(dpath_mulcore_ary1_a1_c1[23]), .Y(n8168));
INVX1 mul_U21420(.A(dpath_mulcore_ary1_a1_c1[22]), .Y(n8169));
INVX1 mul_U21421(.A(dpath_mulcore_ary1_a1_c1[21]), .Y(n8170));
INVX1 mul_U21422(.A(dpath_mulcore_ary1_a1_c1[20]), .Y(n8171));
INVX1 mul_U21423(.A(dpath_mulcore_ary1_a1_c1[19]), .Y(n8172));
INVX1 mul_U21424(.A(dpath_mulcore_ary1_a1_c1[18]), .Y(n8173));
INVX1 mul_U21425(.A(dpath_mulcore_ary1_a1_c1[17]), .Y(n8174));
INVX1 mul_U21426(.A(dpath_mulcore_ary1_a1_c1[16]), .Y(n8175));
INVX1 mul_U21427(.A(dpath_mulcore_ary1_a1_c1[15]), .Y(n8176));
INVX1 mul_U21428(.A(dpath_mulcore_ary1_a1_c1[14]), .Y(n8177));
INVX1 mul_U21429(.A(dpath_mulcore_ary1_a1_c1[13]), .Y(n8178));
INVX1 mul_U21430(.A(dpath_mulcore_ary1_a1_c1[12]), .Y(n8179));
INVX1 mul_U21431(.A(dpath_mulcore_ary1_a1_c1[11]), .Y(n8180));
INVX1 mul_U21432(.A(dpath_mulcore_ary1_a1_c1[10]), .Y(n8181));
INVX1 mul_U21433(.A(dpath_mulcore_ary1_a1_c1[9]), .Y(n8182));
INVX1 mul_U21434(.A(dpath_mulcore_ary1_a1_c1[8]), .Y(n8183));
INVX1 mul_U21435(.A(dpath_mulcore_ary1_a1_c1[7]), .Y(n8184));
INVX1 mul_U21436(.A(dpath_mulcore_ary1_a1_c1[6]), .Y(n8185));
INVX1 mul_U21437(.A(dpath_mulcore_ary1_a1_c1[5]), .Y(n8186));
INVX1 mul_U21438(.A(dpath_mulcore_ary1_a1_c1[4]), .Y(n8187));
INVX1 mul_U21439(.A(dpath_mulcore_ary1_a1_c1[64]), .Y(n8188));
INVX1 mul_U21440(.A(dpath_mulcore_ary1_a1_c1[65]), .Y(n8189));
INVX1 mul_U21441(.A(dpath_mulcore_ary1_a1_c1[66]), .Y(n8190));
INVX1 mul_U21442(.A(dpath_mulcore_array2_ain[68]), .Y(n8191));
INVX1 mul_U21443(.A(dpath_mulcore_array2_ain[67]), .Y(n8192));
INVX1 mul_U21444(.A(dpath_mulcore_array2_ain[66]), .Y(n8193));
INVX1 mul_U21445(.A(dpath_mulcore_array2_ain[65]), .Y(n8194));
INVX1 mul_U21446(.A(dpath_mulcore_array2_ain[64]), .Y(n8195));
INVX1 mul_U21447(.A(dpath_mulcore_array2_ain[63]), .Y(n8196));
INVX1 mul_U21448(.A(dpath_mulcore_array2_ain[62]), .Y(n8197));
INVX1 mul_U21449(.A(dpath_mulcore_array2_ain[61]), .Y(n8198));
INVX1 mul_U21450(.A(dpath_mulcore_array2_ain[60]), .Y(n8199));
INVX1 mul_U21451(.A(dpath_mulcore_array2_ain[59]), .Y(n8200));
INVX1 mul_U21452(.A(dpath_mulcore_array2_ain[58]), .Y(n8201));
INVX1 mul_U21453(.A(dpath_mulcore_array2_ain[57]), .Y(n8202));
INVX1 mul_U21454(.A(dpath_mulcore_array2_ain[56]), .Y(n8203));
INVX1 mul_U21455(.A(dpath_mulcore_array2_ain[55]), .Y(n8204));
INVX1 mul_U21456(.A(dpath_mulcore_array2_ain[54]), .Y(n8205));
INVX1 mul_U21457(.A(dpath_mulcore_array2_ain[53]), .Y(n8206));
INVX1 mul_U21458(.A(dpath_mulcore_array2_ain[52]), .Y(n8207));
INVX1 mul_U21459(.A(dpath_mulcore_array2_ain[51]), .Y(n8208));
INVX1 mul_U21460(.A(dpath_mulcore_array2_ain[50]), .Y(n8209));
INVX1 mul_U21461(.A(dpath_mulcore_array2_ain[49]), .Y(n8210));
INVX1 mul_U21462(.A(dpath_mulcore_array2_ain[48]), .Y(n8211));
INVX1 mul_U21463(.A(dpath_mulcore_array2_ain[47]), .Y(n8212));
INVX1 mul_U21464(.A(dpath_mulcore_array2_ain[46]), .Y(n8213));
INVX1 mul_U21465(.A(dpath_mulcore_array2_ain[45]), .Y(n8214));
INVX1 mul_U21466(.A(dpath_mulcore_array2_ain[44]), .Y(n8215));
INVX1 mul_U21467(.A(dpath_mulcore_array2_ain[43]), .Y(n8216));
INVX1 mul_U21468(.A(dpath_mulcore_array2_ain[42]), .Y(n8217));
INVX1 mul_U21469(.A(dpath_mulcore_array2_ain[41]), .Y(n8218));
INVX1 mul_U21470(.A(dpath_mulcore_array2_ain[40]), .Y(n8219));
INVX1 mul_U21471(.A(dpath_mulcore_array2_ain[39]), .Y(n8220));
INVX1 mul_U21472(.A(dpath_mulcore_array2_ain[38]), .Y(n8221));
INVX1 mul_U21473(.A(dpath_mulcore_array2_ain[37]), .Y(n8222));
INVX1 mul_U21474(.A(dpath_mulcore_array2_ain[36]), .Y(n8223));
INVX1 mul_U21475(.A(dpath_mulcore_array2_ain[35]), .Y(n8224));
INVX1 mul_U21476(.A(dpath_mulcore_array2_ain[34]), .Y(n8225));
INVX1 mul_U21477(.A(dpath_mulcore_array2_ain[33]), .Y(n8226));
INVX1 mul_U21478(.A(dpath_mulcore_array2_ain[32]), .Y(n8227));
INVX1 mul_U21479(.A(dpath_mulcore_array2_ain[31]), .Y(n8228));
INVX1 mul_U21480(.A(dpath_mulcore_array2_ain[30]), .Y(n8229));
INVX1 mul_U21481(.A(dpath_mulcore_array2_ain[29]), .Y(n8230));
INVX1 mul_U21482(.A(dpath_mulcore_array2_ain[28]), .Y(n8231));
INVX1 mul_U21483(.A(dpath_mulcore_array2_ain[27]), .Y(n8232));
INVX1 mul_U21484(.A(dpath_mulcore_array2_ain[26]), .Y(n8233));
INVX1 mul_U21485(.A(dpath_mulcore_array2_ain[25]), .Y(n8234));
INVX1 mul_U21486(.A(dpath_mulcore_array2_ain[24]), .Y(n8235));
INVX1 mul_U21487(.A(dpath_mulcore_array2_ain[23]), .Y(n8236));
INVX1 mul_U21488(.A(dpath_mulcore_array2_ain[22]), .Y(n8237));
INVX1 mul_U21489(.A(dpath_mulcore_array2_ain[21]), .Y(n8238));
INVX1 mul_U21490(.A(dpath_mulcore_array2_ain[20]), .Y(n8239));
INVX1 mul_U21491(.A(dpath_mulcore_array2_ain[95]), .Y(n8240));
INVX1 mul_U21492(.A(dpath_mulcore_array2_ain[94]), .Y(n8241));
INVX1 mul_U21493(.A(dpath_mulcore_array2_ain[93]), .Y(n8242));
INVX1 mul_U21494(.A(dpath_mulcore_array2_ain[92]), .Y(n8243));
INVX1 mul_U21495(.A(dpath_mulcore_array2_ain[91]), .Y(n8244));
INVX1 mul_U21496(.A(dpath_mulcore_array2_ain[90]), .Y(n8245));
INVX1 mul_U21497(.A(dpath_mulcore_array2_ain[89]), .Y(n8246));
INVX1 mul_U21498(.A(dpath_mulcore_array2_ain[88]), .Y(n8247));
INVX1 mul_U21499(.A(dpath_mulcore_array2_ain[87]), .Y(n8248));
INVX1 mul_U21500(.A(dpath_mulcore_array2_ain[86]), .Y(n8249));
INVX1 mul_U21501(.A(dpath_mulcore_array2_ain[85]), .Y(n8250));
INVX1 mul_U21502(.A(dpath_mulcore_array2_ain[84]), .Y(n8251));
INVX1 mul_U21503(.A(dpath_mulcore_array2_ain[81]), .Y(n8252));
INVX1 mul_U21504(.A(dpath_mulcore_array2_ain[80]), .Y(n8253));
INVX1 mul_U21505(.A(dpath_mulcore_array2_ain[79]), .Y(n8254));
INVX1 mul_U21506(.A(dpath_mulcore_array2_ain[78]), .Y(n8255));
INVX1 mul_U21507(.A(dpath_mulcore_array2_ain[77]), .Y(n8256));
INVX1 mul_U21508(.A(dpath_mulcore_array2_ain[76]), .Y(n8257));
INVX1 mul_U21509(.A(dpath_mulcore_array2_ain[75]), .Y(n8258));
INVX1 mul_U21510(.A(dpath_mulcore_array2_ain[74]), .Y(n8259));
INVX1 mul_U21511(.A(dpath_mulcore_array2_ain[73]), .Y(n8260));
INVX1 mul_U21512(.A(dpath_mulcore_array2_ain[72]), .Y(n8261));
INVX1 mul_U21513(.A(dpath_mulcore_array2_ain[71]), .Y(n8262));
INVX1 mul_U21514(.A(dpath_mulcore_array2_ain[70]), .Y(n8263));
INVX1 mul_U21515(.A(dpath_mulcore_array2_ain[69]), .Y(n8264));
INVX1 mul_U21516(.A(dpath_mulcore_array2_ain[19]), .Y(n8265));
INVX1 mul_U21517(.A(dpath_mulcore_array2_ain[18]), .Y(n8266));
INVX1 mul_U21518(.A(dpath_mulcore_array2_ain[17]), .Y(n8267));
INVX1 mul_U21519(.A(dpath_mulcore_array2_ain[16]), .Y(n8268));
INVX1 mul_U21520(.A(dpath_mulcore_array2_ain[15]), .Y(n8269));
INVX1 mul_U21521(.A(dpath_mulcore_array2_ain[4]), .Y(n8270));
INVX1 mul_U21522(.A(dpath_mulcore_array2_ain[3]), .Y(n8271));
INVX1 mul_U21523(.A(dpath_mulcore_array2_ain[2]), .Y(n8272));
INVX1 mul_U21524(.A(dpath_mulcore_array2_ain[1]), .Y(n8273));
INVX1 mul_U21525(.A(dpath_mulcore_array2_ain[83]), .Y(n8274));
INVX1 mul_U21526(.A(dpath_mulcore_array2_ain[14]), .Y(n8275));
INVX1 mul_U21527(.A(dpath_mulcore_array2_ain[13]), .Y(n8276));
INVX1 mul_U21528(.A(dpath_mulcore_array2_ain[12]), .Y(n8277));
INVX1 mul_U21529(.A(dpath_mulcore_array2_ain[11]), .Y(n8278));
INVX1 mul_U21530(.A(dpath_mulcore_array2_ain[10]), .Y(n8279));
INVX1 mul_U21531(.A(dpath_mulcore_array2_ain[9]), .Y(n8280));
INVX1 mul_U21532(.A(dpath_mulcore_array2_ain[8]), .Y(n8281));
INVX1 mul_U21533(.A(dpath_mulcore_array2_ain[7]), .Y(n8282));
INVX1 mul_U21534(.A(dpath_mulcore_array2_ain[6]), .Y(n8283));
INVX1 mul_U21535(.A(dpath_mulcore_array2_ain[5]), .Y(n8284));
INVX1 mul_U21536(.A(dpath_mulcore_ary1_a0_c_2[76]), .Y(n8285));
INVX1 mul_U21537(.A(dpath_mulcore_ary1_a0_c_1[9]), .Y(n8286));
INVX1 mul_U21538(.A(dpath_mulcore_ary1_a0_c_1[8]), .Y(n8287));
INVX1 mul_U21539(.A(dpath_mulcore_ary1_a0_c_2[71]), .Y(n8288));
INVX1 mul_U21540(.A(dpath_mulcore_ary1_a0_c_2[75]), .Y(n8289));
INVX1 mul_U21541(.A(dpath_mulcore_ary1_a0_c_2[74]), .Y(n8290));
INVX1 mul_U21542(.A(dpath_mulcore_ary1_a0_c_2[73]), .Y(n8291));
INVX1 mul_U21543(.A(dpath_mulcore_ary1_a0_c_2[72]), .Y(n8292));
INVX1 mul_U21544(.A(dpath_mulcore_ary1_a0_c_1[7]), .Y(n8293));
INVX1 mul_U21545(.A(dpath_mulcore_ary1_a1_c_2[76]), .Y(n8294));
INVX1 mul_U21546(.A(dpath_mulcore_ary1_a1_c_1[9]), .Y(n8295));
INVX1 mul_U21547(.A(dpath_mulcore_ary1_a1_c_1[8]), .Y(n8296));
INVX1 mul_U21548(.A(dpath_mulcore_ary1_a1_c_2[71]), .Y(n8297));
INVX1 mul_U21549(.A(dpath_mulcore_ary1_a1_c_2[75]), .Y(n8298));
INVX1 mul_U21550(.A(dpath_mulcore_ary1_a1_c_2[74]), .Y(n8299));
INVX1 mul_U21551(.A(dpath_mulcore_ary1_a1_c_2[73]), .Y(n8300));
INVX1 mul_U21552(.A(dpath_mulcore_ary1_a1_c_2[72]), .Y(n8301));
INVX1 mul_U21553(.A(dpath_mulcore_ary1_a1_c_1[7]), .Y(n8302));
INVX1 mul_U21554(.A(dpath_mulcore_array2_c2[83]), .Y(n8303));
INVX1 mul_U21555(.A(dpath_mulcore_array2_c2[18]), .Y(n8304));
INVX1 mul_U21556(.A(dpath_mulcore_array2_c2[17]), .Y(n8305));
INVX1 mul_U21557(.A(dpath_mulcore_array2_c2[16]), .Y(n8306));
INVX1 mul_U21558(.A(dpath_mulcore_array2_c2[15]), .Y(n8307));
INVX1 mul_U21559(.A(dpath_mulcore_array2_c3[19]), .Y(n8308));
INVX1 mul_U21560(.A(dpath_mulcore_array2_c3[18]), .Y(n8309));
INVX1 mul_U21561(.A(dpath_mulcore_array2_c3[17]), .Y(n8310));
INVX1 mul_U21562(.A(dpath_mulcore_array2_c3[16]), .Y(n8311));
INVX1 mul_U21563(.A(dpath_mulcore_array2_c3[15]), .Y(n8312));
INVX1 mul_U21564(.A(dpath_mulcore_array2_c1[82]), .Y(n8313));
INVX1 mul_U21565(.A(dpath_mulcore_array2_c2[14]), .Y(n8314));
INVX1 mul_U21566(.A(dpath_mulcore_array2_c2[13]), .Y(n8315));
INVX1 mul_U21567(.A(dpath_mulcore_array2_c2[12]), .Y(n8316));
INVX1 mul_U21568(.A(dpath_mulcore_array2_c2[11]), .Y(n8317));
INVX1 mul_U21569(.A(dpath_mulcore_array2_c2[10]), .Y(n8318));
INVX1 mul_U21570(.A(dpath_mulcore_array2_c2[9]), .Y(n8319));
INVX1 mul_U21571(.A(dpath_mulcore_array2_c2[8]), .Y(n8320));
INVX1 mul_U21572(.A(dpath_mulcore_array2_c2[7]), .Y(n8321));
INVX1 mul_U21573(.A(dpath_mulcore_array2_c2[6]), .Y(n8322));
INVX1 mul_U21574(.A(dpath_mulcore_array2_c2[5]), .Y(n8323));
INVX1 mul_U21575(.A(dpath_mulcore_array2_c2[82]), .Y(n8324));
INVX1 mul_U21576(.A(dpath_mulcore_array2_c2[81]), .Y(n8325));
INVX1 mul_U21577(.A(dpath_mulcore_ary1_a0_c1[66]), .Y(n8326));
INVX1 mul_U21578(.A(dpath_mulcore_ary1_a0_c1[65]), .Y(n8327));
INVX1 mul_U21579(.A(dpath_mulcore_ary1_a0_c1[64]), .Y(n8328));
INVX1 mul_U21580(.A(dpath_mulcore_array2_c3[68]), .Y(n8329));
INVX1 mul_U21581(.A(dpath_mulcore_array2_c3[67]), .Y(n8330));
INVX1 mul_U21582(.A(dpath_mulcore_array2_c3[66]), .Y(n8331));
INVX1 mul_U21583(.A(dpath_mulcore_array2_c3[65]), .Y(n8332));
INVX1 mul_U21584(.A(dpath_mulcore_array2_c3[64]), .Y(n8333));
INVX1 mul_U21585(.A(dpath_mulcore_array2_c3[63]), .Y(n8334));
INVX1 mul_U21586(.A(dpath_mulcore_array2_c3[62]), .Y(n8335));
INVX1 mul_U21587(.A(dpath_mulcore_array2_c3[61]), .Y(n8336));
INVX1 mul_U21588(.A(dpath_mulcore_array2_c3[60]), .Y(n8337));
INVX1 mul_U21589(.A(dpath_mulcore_array2_c3[59]), .Y(n8338));
INVX1 mul_U21590(.A(dpath_mulcore_array2_c3[58]), .Y(n8339));
INVX1 mul_U21591(.A(dpath_mulcore_array2_c3[57]), .Y(n8340));
INVX1 mul_U21592(.A(dpath_mulcore_array2_c3[56]), .Y(n8341));
INVX1 mul_U21593(.A(dpath_mulcore_array2_c3[55]), .Y(n8342));
INVX1 mul_U21594(.A(dpath_mulcore_array2_c3[54]), .Y(n8343));
INVX1 mul_U21595(.A(dpath_mulcore_array2_c3[53]), .Y(n8344));
INVX1 mul_U21596(.A(dpath_mulcore_array2_c3[52]), .Y(n8345));
INVX1 mul_U21597(.A(dpath_mulcore_array2_c3[51]), .Y(n8346));
INVX1 mul_U21598(.A(dpath_mulcore_array2_c3[50]), .Y(n8347));
INVX1 mul_U21599(.A(dpath_mulcore_array2_c3[49]), .Y(n8348));
INVX1 mul_U21600(.A(dpath_mulcore_array2_c3[48]), .Y(n8349));
INVX1 mul_U21601(.A(dpath_mulcore_array2_c3[47]), .Y(n8350));
INVX1 mul_U21602(.A(dpath_mulcore_array2_c3[46]), .Y(n8351));
INVX1 mul_U21603(.A(dpath_mulcore_array2_c3[45]), .Y(n8352));
INVX1 mul_U21604(.A(dpath_mulcore_array2_c3[44]), .Y(n8353));
INVX1 mul_U21605(.A(dpath_mulcore_array2_c3[43]), .Y(n8354));
INVX1 mul_U21606(.A(dpath_mulcore_array2_c3[42]), .Y(n8355));
INVX1 mul_U21607(.A(dpath_mulcore_array2_c3[41]), .Y(n8356));
INVX1 mul_U21608(.A(dpath_mulcore_array2_c3[40]), .Y(n8357));
INVX1 mul_U21609(.A(dpath_mulcore_array2_c3[39]), .Y(n8358));
INVX1 mul_U21610(.A(dpath_mulcore_array2_c3[38]), .Y(n8359));
INVX1 mul_U21611(.A(dpath_mulcore_array2_c3[37]), .Y(n8360));
INVX1 mul_U21612(.A(dpath_mulcore_array2_c3[36]), .Y(n8361));
INVX1 mul_U21613(.A(dpath_mulcore_array2_c3[35]), .Y(n8362));
INVX1 mul_U21614(.A(dpath_mulcore_array2_c3[34]), .Y(n8363));
INVX1 mul_U21615(.A(dpath_mulcore_array2_c3[33]), .Y(n8364));
INVX1 mul_U21616(.A(dpath_mulcore_array2_c3[32]), .Y(n8365));
INVX1 mul_U21617(.A(dpath_mulcore_array2_c3[31]), .Y(n8366));
INVX1 mul_U21618(.A(dpath_mulcore_array2_c3[30]), .Y(n8367));
INVX1 mul_U21619(.A(dpath_mulcore_array2_c3[29]), .Y(n8368));
INVX1 mul_U21620(.A(dpath_mulcore_array2_c3[28]), .Y(n8369));
INVX1 mul_U21621(.A(dpath_mulcore_array2_c3[27]), .Y(n8370));
INVX1 mul_U21622(.A(dpath_mulcore_array2_c3[26]), .Y(n8371));
INVX1 mul_U21623(.A(dpath_mulcore_array2_c3[25]), .Y(n8372));
INVX1 mul_U21624(.A(dpath_mulcore_array2_c3[24]), .Y(n8373));
INVX1 mul_U21625(.A(dpath_mulcore_array2_c3[23]), .Y(n8374));
INVX1 mul_U21626(.A(dpath_mulcore_array2_c3[22]), .Y(n8375));
INVX1 mul_U21627(.A(dpath_mulcore_array2_c3[21]), .Y(n8376));
INVX1 mul_U21628(.A(dpath_mulcore_ary1_a0_b2n[1]), .Y(n8377));
INVX1 mul_U21629(.A(dpath_mulcore_ary1_a0_b2n[0]), .Y(n8378));
INVX1 mul_U21630(.A(dpath_mulcore_ary1_a1_b5n[1]), .Y(n8379));
INVX1 mul_U21631(.A(dpath_mulcore_ary1_a1_b5n[0]), .Y(n8380));
INVX1 mul_U21632(.A(dpath_mulcore_ary1_a1_b2n[1]), .Y(n8381));
INVX1 mul_U21633(.A(dpath_mulcore_ary1_a1_b2n[0]), .Y(n8382));
INVX1 mul_U21634(.A(dpath_mulcore_ary1_a0_I2_I0_b1n_1), .Y(n8383));
INVX1 mul_U21635(.A(dpath_mulcore_ary1_a0_I2_I0_b1n_0), .Y(n8384));
INVX1 mul_U21636(.A(dpath_mulcore_array2_ain[82]), .Y(n8385));
INVX1 mul_U21637(.A(dpath_mulcore_ary1_a0_b5n[1]), .Y(n8386));
INVX1 mul_U21638(.A(dpath_mulcore_ary1_a0_b5n[0]), .Y(n8387));
INVX1 mul_U21639(.A(dpath_mulcore_ary1_a0_I2_I1_63__net32), .Y(n8388));
INVX1 mul_U21640(.A(dpath_mulcore_ary1_a0_I2_I1_62__net32), .Y(n8389));
INVX1 mul_U21641(.A(dpath_mulcore_ary1_a0_I2_I1_61__net32), .Y(n8390));
INVX1 mul_U21642(.A(dpath_mulcore_ary1_a0_I2_I1_60__net32), .Y(n8391));
INVX1 mul_U21643(.A(dpath_mulcore_ary1_a0_I2_I1_59__net32), .Y(n8392));
INVX1 mul_U21644(.A(dpath_mulcore_ary1_a0_I2_I1_58__net32), .Y(n8393));
INVX1 mul_U21645(.A(dpath_mulcore_ary1_a0_I2_I1_57__net32), .Y(n8394));
INVX1 mul_U21646(.A(dpath_mulcore_ary1_a0_I2_I1_56__net32), .Y(n8395));
INVX1 mul_U21647(.A(dpath_mulcore_ary1_a0_I2_I1_55__net32), .Y(n8396));
INVX1 mul_U21648(.A(dpath_mulcore_ary1_a0_I2_I1_54__net32), .Y(n8397));
INVX1 mul_U21649(.A(dpath_mulcore_ary1_a0_I2_I1_53__net32), .Y(n8398));
INVX1 mul_U21650(.A(dpath_mulcore_ary1_a0_I2_I1_52__net32), .Y(n8399));
INVX1 mul_U21651(.A(dpath_mulcore_ary1_a0_I2_I1_51__net32), .Y(n8400));
INVX1 mul_U21652(.A(dpath_mulcore_ary1_a0_I2_I1_50__net32), .Y(n8401));
INVX1 mul_U21653(.A(dpath_mulcore_ary1_a0_I2_I1_49__net32), .Y(n8402));
INVX1 mul_U21654(.A(dpath_mulcore_ary1_a0_I2_I1_48__net32), .Y(n8403));
INVX1 mul_U21655(.A(dpath_mulcore_ary1_a0_I2_I1_47__net32), .Y(n8404));
INVX1 mul_U21656(.A(dpath_mulcore_ary1_a0_I2_I1_46__net32), .Y(n8405));
INVX1 mul_U21657(.A(dpath_mulcore_ary1_a0_I2_I1_45__net32), .Y(n8406));
INVX1 mul_U21658(.A(dpath_mulcore_ary1_a0_I2_I1_44__net32), .Y(n8407));
INVX1 mul_U21659(.A(dpath_mulcore_ary1_a0_I2_I1_43__net32), .Y(n8408));
INVX1 mul_U21660(.A(dpath_mulcore_ary1_a0_I2_I1_42__net32), .Y(n8409));
INVX1 mul_U21661(.A(dpath_mulcore_ary1_a0_I2_I1_41__net32), .Y(n8410));
INVX1 mul_U21662(.A(dpath_mulcore_ary1_a0_I2_I1_40__net32), .Y(n8411));
INVX1 mul_U21663(.A(dpath_mulcore_ary1_a0_I2_I1_39__net32), .Y(n8412));
INVX1 mul_U21664(.A(dpath_mulcore_ary1_a0_I2_I1_38__net32), .Y(n8413));
INVX1 mul_U21665(.A(dpath_mulcore_ary1_a0_I2_I1_37__net32), .Y(n8414));
INVX1 mul_U21666(.A(dpath_mulcore_ary1_a0_I2_I1_36__net32), .Y(n8415));
INVX1 mul_U21667(.A(dpath_mulcore_ary1_a0_I2_I1_35__net32), .Y(n8416));
INVX1 mul_U21668(.A(dpath_mulcore_ary1_a0_I2_I1_34__net32), .Y(n8417));
INVX1 mul_U21669(.A(dpath_mulcore_ary1_a0_I2_I1_33__net32), .Y(n8418));
INVX1 mul_U21670(.A(dpath_mulcore_ary1_a0_I2_I1_32__net32), .Y(n8419));
INVX1 mul_U21671(.A(dpath_mulcore_ary1_a0_I2_I1_31__net32), .Y(n8420));
INVX1 mul_U21672(.A(dpath_mulcore_ary1_a0_I2_I1_30__net32), .Y(n8421));
INVX1 mul_U21673(.A(dpath_mulcore_ary1_a0_I2_I1_29__net32), .Y(n8422));
INVX1 mul_U21674(.A(dpath_mulcore_ary1_a0_I2_I1_28__net32), .Y(n8423));
INVX1 mul_U21675(.A(dpath_mulcore_ary1_a0_I2_I1_27__net32), .Y(n8424));
INVX1 mul_U21676(.A(dpath_mulcore_ary1_a0_I2_I1_26__net32), .Y(n8425));
INVX1 mul_U21677(.A(dpath_mulcore_ary1_a0_I2_I1_25__net32), .Y(n8426));
INVX1 mul_U21678(.A(dpath_mulcore_ary1_a0_I2_I1_24__net32), .Y(n8427));
INVX1 mul_U21679(.A(dpath_mulcore_ary1_a0_I2_I1_23__net32), .Y(n8428));
INVX1 mul_U21680(.A(dpath_mulcore_ary1_a0_I2_I1_22__net32), .Y(n8429));
INVX1 mul_U21681(.A(dpath_mulcore_ary1_a0_I2_I1_21__net32), .Y(n8430));
INVX1 mul_U21682(.A(dpath_mulcore_ary1_a0_I2_I1_20__net32), .Y(n8431));
INVX1 mul_U21683(.A(dpath_mulcore_ary1_a0_I2_I1_19__net32), .Y(n8432));
INVX1 mul_U21684(.A(dpath_mulcore_ary1_a0_I2_I1_18__net32), .Y(n8433));
INVX1 mul_U21685(.A(dpath_mulcore_ary1_a0_I2_I1_17__net32), .Y(n8434));
INVX1 mul_U21686(.A(dpath_mulcore_ary1_a0_I2_I1_16__net32), .Y(n8435));
INVX1 mul_U21687(.A(dpath_mulcore_ary1_a0_I2_I1_15__net32), .Y(n8436));
INVX1 mul_U21688(.A(dpath_mulcore_ary1_a0_I2_I1_14__net32), .Y(n8437));
INVX1 mul_U21689(.A(dpath_mulcore_ary1_a0_I2_I1_13__net32), .Y(n8438));
INVX1 mul_U21690(.A(dpath_mulcore_ary1_a0_I2_I1_12__net32), .Y(n8439));
INVX1 mul_U21691(.A(dpath_mulcore_ary1_a0_I2_I1_11__net32), .Y(n8440));
INVX1 mul_U21692(.A(dpath_mulcore_ary1_a0_I2_I1_10__net32), .Y(n8441));
INVX1 mul_U21693(.A(dpath_mulcore_ary1_a0_I2_I1_9__net32), .Y(n8442));
INVX1 mul_U21694(.A(dpath_mulcore_ary1_a0_I2_I1_8__net32), .Y(n8443));
INVX1 mul_U21695(.A(dpath_mulcore_ary1_a0_I2_I1_7__net32), .Y(n8444));
INVX1 mul_U21696(.A(dpath_mulcore_ary1_a0_I2_I1_6__net32), .Y(n8445));
INVX1 mul_U21697(.A(dpath_mulcore_ary1_a0_I2_I1_5__net32), .Y(n8446));
INVX1 mul_U21698(.A(dpath_mulcore_ary1_a0_I2_I1_4__net32), .Y(n8447));
INVX1 mul_U21699(.A(dpath_mulcore_ary1_a0_I2_I0_p1_3), .Y(n8448));
INVX1 mul_U21700(.A(dpath_mulcore_ary1_a0_I1_I1_63__net32), .Y(n8449));
INVX1 mul_U21701(.A(dpath_mulcore_ary1_a0_I1_I1_62__net32), .Y(n8450));
INVX1 mul_U21702(.A(dpath_mulcore_ary1_a0_I1_I1_61__net32), .Y(n8451));
INVX1 mul_U21703(.A(dpath_mulcore_ary1_a0_I1_I1_60__net32), .Y(n8452));
INVX1 mul_U21704(.A(dpath_mulcore_ary1_a0_I1_I1_59__net32), .Y(n8453));
INVX1 mul_U21705(.A(dpath_mulcore_ary1_a0_I1_I1_58__net32), .Y(n8454));
INVX1 mul_U21706(.A(dpath_mulcore_ary1_a0_I1_I1_57__net32), .Y(n8455));
INVX1 mul_U21707(.A(dpath_mulcore_ary1_a0_I1_I1_56__net32), .Y(n8456));
INVX1 mul_U21708(.A(dpath_mulcore_ary1_a0_I1_I1_55__net32), .Y(n8457));
INVX1 mul_U21709(.A(dpath_mulcore_ary1_a0_I1_I1_54__net32), .Y(n8458));
INVX1 mul_U21710(.A(dpath_mulcore_ary1_a0_I1_I1_53__net32), .Y(n8459));
INVX1 mul_U21711(.A(dpath_mulcore_ary1_a0_I1_I1_52__net32), .Y(n8460));
INVX1 mul_U21712(.A(dpath_mulcore_ary1_a0_I1_I1_51__net32), .Y(n8461));
INVX1 mul_U21713(.A(dpath_mulcore_ary1_a0_I1_I1_50__net32), .Y(n8462));
INVX1 mul_U21714(.A(dpath_mulcore_ary1_a0_I1_I1_49__net32), .Y(n8463));
INVX1 mul_U21715(.A(dpath_mulcore_ary1_a0_I1_I1_48__net32), .Y(n8464));
INVX1 mul_U21716(.A(dpath_mulcore_ary1_a0_I1_I1_47__net32), .Y(n8465));
INVX1 mul_U21717(.A(dpath_mulcore_ary1_a0_I1_I1_46__net32), .Y(n8466));
INVX1 mul_U21718(.A(dpath_mulcore_ary1_a0_I1_I1_45__net32), .Y(n8467));
INVX1 mul_U21719(.A(dpath_mulcore_ary1_a0_I1_I1_44__net32), .Y(n8468));
INVX1 mul_U21720(.A(dpath_mulcore_ary1_a0_I1_I1_43__net32), .Y(n8469));
INVX1 mul_U21721(.A(dpath_mulcore_ary1_a0_I1_I1_42__net32), .Y(n8470));
INVX1 mul_U21722(.A(dpath_mulcore_ary1_a0_I1_I1_41__net32), .Y(n8471));
INVX1 mul_U21723(.A(dpath_mulcore_ary1_a0_I1_I1_40__net32), .Y(n8472));
INVX1 mul_U21724(.A(dpath_mulcore_ary1_a0_I1_I1_39__net32), .Y(n8473));
INVX1 mul_U21725(.A(dpath_mulcore_ary1_a0_I1_I1_38__net32), .Y(n8474));
INVX1 mul_U21726(.A(dpath_mulcore_ary1_a0_I1_I1_37__net32), .Y(n8475));
INVX1 mul_U21727(.A(dpath_mulcore_ary1_a0_I1_I1_36__net32), .Y(n8476));
INVX1 mul_U21728(.A(dpath_mulcore_ary1_a0_I1_I1_35__net32), .Y(n8477));
INVX1 mul_U21729(.A(dpath_mulcore_ary1_a0_I1_I1_34__net32), .Y(n8478));
INVX1 mul_U21730(.A(dpath_mulcore_ary1_a0_I1_I1_33__net32), .Y(n8479));
INVX1 mul_U21731(.A(dpath_mulcore_ary1_a0_I1_I1_32__net32), .Y(n8480));
INVX1 mul_U21732(.A(dpath_mulcore_ary1_a0_I1_I1_31__net32), .Y(n8481));
INVX1 mul_U21733(.A(dpath_mulcore_ary1_a0_I1_I1_30__net32), .Y(n8482));
INVX1 mul_U21734(.A(dpath_mulcore_ary1_a0_I1_I1_29__net32), .Y(n8483));
INVX1 mul_U21735(.A(dpath_mulcore_ary1_a0_I1_I1_28__net32), .Y(n8484));
INVX1 mul_U21736(.A(dpath_mulcore_ary1_a0_I1_I1_27__net32), .Y(n8485));
INVX1 mul_U21737(.A(dpath_mulcore_ary1_a0_I1_I1_26__net32), .Y(n8486));
INVX1 mul_U21738(.A(dpath_mulcore_ary1_a0_I1_I1_25__net32), .Y(n8487));
INVX1 mul_U21739(.A(dpath_mulcore_ary1_a0_I1_I1_24__net32), .Y(n8488));
INVX1 mul_U21740(.A(dpath_mulcore_ary1_a0_I1_I1_23__net32), .Y(n8489));
INVX1 mul_U21741(.A(dpath_mulcore_ary1_a0_I1_I1_22__net32), .Y(n8490));
INVX1 mul_U21742(.A(dpath_mulcore_ary1_a0_I1_I1_21__net32), .Y(n8491));
INVX1 mul_U21743(.A(dpath_mulcore_ary1_a0_I1_I1_20__net32), .Y(n8492));
INVX1 mul_U21744(.A(dpath_mulcore_ary1_a0_I1_I1_19__net32), .Y(n8493));
INVX1 mul_U21745(.A(dpath_mulcore_ary1_a0_I1_I1_18__net32), .Y(n8494));
INVX1 mul_U21746(.A(dpath_mulcore_ary1_a0_I1_I1_17__net32), .Y(n8495));
INVX1 mul_U21747(.A(dpath_mulcore_ary1_a0_I1_I1_16__net32), .Y(n8496));
INVX1 mul_U21748(.A(dpath_mulcore_ary1_a0_I1_I1_15__net32), .Y(n8497));
INVX1 mul_U21749(.A(dpath_mulcore_ary1_a0_I1_I1_14__net32), .Y(n8498));
INVX1 mul_U21750(.A(dpath_mulcore_ary1_a0_I1_I1_13__net32), .Y(n8499));
INVX1 mul_U21751(.A(dpath_mulcore_ary1_a0_I1_I1_12__net32), .Y(n8500));
INVX1 mul_U21752(.A(dpath_mulcore_ary1_a0_I1_I1_11__net32), .Y(n8501));
INVX1 mul_U21753(.A(dpath_mulcore_ary1_a0_I1_I1_10__net32), .Y(n8502));
INVX1 mul_U21754(.A(dpath_mulcore_ary1_a0_I1_I1_9__net32), .Y(n8503));
INVX1 mul_U21755(.A(dpath_mulcore_ary1_a0_I1_I1_8__net32), .Y(n8504));
INVX1 mul_U21756(.A(dpath_mulcore_ary1_a0_I1_I1_7__net32), .Y(n8505));
INVX1 mul_U21757(.A(dpath_mulcore_ary1_a0_I1_I1_6__net32), .Y(n8506));
INVX1 mul_U21758(.A(dpath_mulcore_ary1_a0_I1_I1_5__net32), .Y(n8507));
INVX1 mul_U21759(.A(dpath_mulcore_ary1_a0_I1_I1_4__net32), .Y(n8508));
INVX1 mul_U21760(.A(dpath_mulcore_ary1_a0_I1_I0_p1_3), .Y(n8509));
INVX1 mul_U21761(.A(dpath_mulcore_ary1_a0_I0_I1_63__net32), .Y(n8510));
INVX1 mul_U21762(.A(dpath_mulcore_ary1_a0_I0_I1_62__net32), .Y(n8511));
INVX1 mul_U21763(.A(dpath_mulcore_ary1_a0_I0_I1_61__net32), .Y(n8512));
INVX1 mul_U21764(.A(dpath_mulcore_ary1_a0_I0_I1_60__net32), .Y(n8513));
INVX1 mul_U21765(.A(dpath_mulcore_ary1_a0_I0_I1_59__net32), .Y(n8514));
INVX1 mul_U21766(.A(dpath_mulcore_ary1_a0_I0_I1_58__net32), .Y(n8515));
INVX1 mul_U21767(.A(dpath_mulcore_ary1_a0_I0_I1_57__net32), .Y(n8516));
INVX1 mul_U21768(.A(dpath_mulcore_ary1_a0_I0_I1_56__net32), .Y(n8517));
INVX1 mul_U21769(.A(dpath_mulcore_ary1_a0_I0_I1_55__net32), .Y(n8518));
INVX1 mul_U21770(.A(dpath_mulcore_ary1_a0_I0_I1_54__net32), .Y(n8519));
INVX1 mul_U21771(.A(dpath_mulcore_ary1_a0_I0_I1_53__net32), .Y(n8520));
INVX1 mul_U21772(.A(dpath_mulcore_ary1_a0_I0_I1_52__net32), .Y(n8521));
INVX1 mul_U21773(.A(dpath_mulcore_ary1_a0_I0_I1_51__net32), .Y(n8522));
INVX1 mul_U21774(.A(dpath_mulcore_ary1_a0_I0_I1_50__net32), .Y(n8523));
INVX1 mul_U21775(.A(dpath_mulcore_ary1_a0_I0_I1_49__net32), .Y(n8524));
INVX1 mul_U21776(.A(dpath_mulcore_ary1_a0_I0_I1_48__net32), .Y(n8525));
INVX1 mul_U21777(.A(dpath_mulcore_ary1_a0_I0_I1_47__net32), .Y(n8526));
INVX1 mul_U21778(.A(dpath_mulcore_ary1_a0_I0_I1_46__net32), .Y(n8527));
INVX1 mul_U21779(.A(dpath_mulcore_ary1_a0_I0_I1_45__net32), .Y(n8528));
INVX1 mul_U21780(.A(dpath_mulcore_ary1_a0_I0_I1_44__net32), .Y(n8529));
INVX1 mul_U21781(.A(dpath_mulcore_ary1_a0_I0_I1_43__net32), .Y(n8530));
INVX1 mul_U21782(.A(dpath_mulcore_ary1_a0_I0_I1_42__net32), .Y(n8531));
INVX1 mul_U21783(.A(dpath_mulcore_ary1_a0_I0_I1_41__net32), .Y(n8532));
INVX1 mul_U21784(.A(dpath_mulcore_ary1_a0_I0_I1_40__net32), .Y(n8533));
INVX1 mul_U21785(.A(dpath_mulcore_ary1_a0_I0_I1_39__net32), .Y(n8534));
INVX1 mul_U21786(.A(dpath_mulcore_ary1_a0_I0_I1_38__net32), .Y(n8535));
INVX1 mul_U21787(.A(dpath_mulcore_ary1_a0_I0_I1_37__net32), .Y(n8536));
INVX1 mul_U21788(.A(dpath_mulcore_ary1_a0_I0_I1_36__net32), .Y(n8537));
INVX1 mul_U21789(.A(dpath_mulcore_ary1_a0_I0_I1_35__net32), .Y(n8538));
INVX1 mul_U21790(.A(dpath_mulcore_ary1_a0_I0_I1_34__net32), .Y(n8539));
INVX1 mul_U21791(.A(dpath_mulcore_ary1_a0_I0_I1_33__net32), .Y(n8540));
INVX1 mul_U21792(.A(dpath_mulcore_ary1_a0_I0_I1_32__net32), .Y(n8541));
INVX1 mul_U21793(.A(dpath_mulcore_ary1_a0_I0_I1_31__net32), .Y(n8542));
INVX1 mul_U21794(.A(dpath_mulcore_ary1_a0_I0_I1_30__net32), .Y(n8543));
INVX1 mul_U21795(.A(dpath_mulcore_ary1_a0_I0_I1_29__net32), .Y(n8544));
INVX1 mul_U21796(.A(dpath_mulcore_ary1_a0_I0_I1_28__net32), .Y(n8545));
INVX1 mul_U21797(.A(dpath_mulcore_ary1_a0_I0_I1_27__net32), .Y(n8546));
INVX1 mul_U21798(.A(dpath_mulcore_ary1_a0_I0_I1_26__net32), .Y(n8547));
INVX1 mul_U21799(.A(dpath_mulcore_ary1_a0_I0_I1_25__net32), .Y(n8548));
INVX1 mul_U21800(.A(dpath_mulcore_ary1_a0_I0_I1_24__net32), .Y(n8549));
INVX1 mul_U21801(.A(dpath_mulcore_ary1_a0_I0_I1_23__net32), .Y(n8550));
INVX1 mul_U21802(.A(dpath_mulcore_ary1_a0_I0_I1_22__net32), .Y(n8551));
INVX1 mul_U21803(.A(dpath_mulcore_ary1_a0_I0_I1_21__net32), .Y(n8552));
INVX1 mul_U21804(.A(dpath_mulcore_ary1_a0_I0_I1_20__net32), .Y(n8553));
INVX1 mul_U21805(.A(dpath_mulcore_ary1_a0_I0_I1_19__net32), .Y(n8554));
INVX1 mul_U21806(.A(dpath_mulcore_ary1_a0_I0_I1_18__net32), .Y(n8555));
INVX1 mul_U21807(.A(dpath_mulcore_ary1_a0_I0_I1_17__net32), .Y(n8556));
INVX1 mul_U21808(.A(dpath_mulcore_ary1_a0_I0_I1_16__net32), .Y(n8557));
INVX1 mul_U21809(.A(dpath_mulcore_ary1_a0_I0_I1_15__net32), .Y(n8558));
INVX1 mul_U21810(.A(dpath_mulcore_ary1_a0_I0_I1_14__net32), .Y(n8559));
INVX1 mul_U21811(.A(dpath_mulcore_ary1_a0_I0_I1_13__net32), .Y(n8560));
INVX1 mul_U21812(.A(dpath_mulcore_ary1_a0_I0_I1_12__net32), .Y(n8561));
INVX1 mul_U21813(.A(dpath_mulcore_ary1_a0_I0_I1_11__net32), .Y(n8562));
INVX1 mul_U21814(.A(dpath_mulcore_ary1_a0_I0_I1_10__net32), .Y(n8563));
INVX1 mul_U21815(.A(dpath_mulcore_ary1_a0_I0_I1_9__net32), .Y(n8564));
INVX1 mul_U21816(.A(dpath_mulcore_ary1_a0_I0_I1_8__net32), .Y(n8565));
INVX1 mul_U21817(.A(dpath_mulcore_ary1_a0_I0_I1_7__net32), .Y(n8566));
INVX1 mul_U21818(.A(dpath_mulcore_ary1_a0_I0_I1_6__net32), .Y(n8567));
INVX1 mul_U21819(.A(dpath_mulcore_ary1_a0_I0_I1_5__net32), .Y(n8568));
INVX1 mul_U21820(.A(dpath_mulcore_ary1_a0_I0_I1_4__net32), .Y(n8569));
INVX1 mul_U21821(.A(dpath_mulcore_ary1_a0_I0_I0_p1_3), .Y(n8570));
INVX1 mul_U21822(.A(dpath_mulcore_ary1_a1_I2_I1_63__net32), .Y(n8571));
INVX1 mul_U21823(.A(dpath_mulcore_ary1_a1_I2_I1_62__net32), .Y(n8572));
INVX1 mul_U21824(.A(dpath_mulcore_ary1_a1_I2_I1_61__net32), .Y(n8573));
INVX1 mul_U21825(.A(dpath_mulcore_ary1_a1_I2_I1_60__net32), .Y(n8574));
INVX1 mul_U21826(.A(dpath_mulcore_ary1_a1_I2_I1_59__net32), .Y(n8575));
INVX1 mul_U21827(.A(dpath_mulcore_ary1_a1_I2_I1_58__net32), .Y(n8576));
INVX1 mul_U21828(.A(dpath_mulcore_ary1_a1_I2_I1_57__net32), .Y(n8577));
INVX1 mul_U21829(.A(dpath_mulcore_ary1_a1_I2_I1_56__net32), .Y(n8578));
INVX1 mul_U21830(.A(dpath_mulcore_ary1_a1_I2_I1_55__net32), .Y(n8579));
INVX1 mul_U21831(.A(dpath_mulcore_ary1_a1_I2_I1_54__net32), .Y(n8580));
INVX1 mul_U21832(.A(dpath_mulcore_ary1_a1_I2_I1_53__net32), .Y(n8581));
INVX1 mul_U21833(.A(dpath_mulcore_ary1_a1_I2_I1_52__net32), .Y(n8582));
INVX1 mul_U21834(.A(dpath_mulcore_ary1_a1_I2_I1_51__net32), .Y(n8583));
INVX1 mul_U21835(.A(dpath_mulcore_ary1_a1_I2_I1_50__net32), .Y(n8584));
INVX1 mul_U21836(.A(dpath_mulcore_ary1_a1_I2_I1_49__net32), .Y(n8585));
INVX1 mul_U21837(.A(dpath_mulcore_ary1_a1_I2_I1_48__net32), .Y(n8586));
INVX1 mul_U21838(.A(dpath_mulcore_ary1_a1_I2_I1_47__net32), .Y(n8587));
INVX1 mul_U21839(.A(dpath_mulcore_ary1_a1_I2_I1_46__net32), .Y(n8588));
INVX1 mul_U21840(.A(dpath_mulcore_ary1_a1_I2_I1_45__net32), .Y(n8589));
INVX1 mul_U21841(.A(dpath_mulcore_ary1_a1_I2_I1_44__net32), .Y(n8590));
INVX1 mul_U21842(.A(dpath_mulcore_ary1_a1_I2_I1_43__net32), .Y(n8591));
INVX1 mul_U21843(.A(dpath_mulcore_ary1_a1_I2_I1_42__net32), .Y(n8592));
INVX1 mul_U21844(.A(dpath_mulcore_ary1_a1_I2_I1_41__net32), .Y(n8593));
INVX1 mul_U21845(.A(dpath_mulcore_ary1_a1_I2_I1_40__net32), .Y(n8594));
INVX1 mul_U21846(.A(dpath_mulcore_ary1_a1_I2_I1_39__net32), .Y(n8595));
INVX1 mul_U21847(.A(dpath_mulcore_ary1_a1_I2_I1_38__net32), .Y(n8596));
INVX1 mul_U21848(.A(dpath_mulcore_ary1_a1_I2_I1_37__net32), .Y(n8597));
INVX1 mul_U21849(.A(dpath_mulcore_ary1_a1_I2_I1_36__net32), .Y(n8598));
INVX1 mul_U21850(.A(dpath_mulcore_ary1_a1_I2_I1_35__net32), .Y(n8599));
INVX1 mul_U21851(.A(dpath_mulcore_ary1_a1_I2_I1_34__net32), .Y(n8600));
INVX1 mul_U21852(.A(dpath_mulcore_ary1_a1_I2_I1_33__net32), .Y(n8601));
INVX1 mul_U21853(.A(dpath_mulcore_ary1_a1_I2_I1_32__net32), .Y(n8602));
INVX1 mul_U21854(.A(dpath_mulcore_ary1_a1_I2_I1_31__net32), .Y(n8603));
INVX1 mul_U21855(.A(dpath_mulcore_ary1_a1_I2_I1_30__net32), .Y(n8604));
INVX1 mul_U21856(.A(dpath_mulcore_ary1_a1_I2_I1_29__net32), .Y(n8605));
INVX1 mul_U21857(.A(dpath_mulcore_ary1_a1_I2_I1_28__net32), .Y(n8606));
INVX1 mul_U21858(.A(dpath_mulcore_ary1_a1_I2_I1_27__net32), .Y(n8607));
INVX1 mul_U21859(.A(dpath_mulcore_ary1_a1_I2_I1_26__net32), .Y(n8608));
INVX1 mul_U21860(.A(dpath_mulcore_ary1_a1_I2_I1_25__net32), .Y(n8609));
INVX1 mul_U21861(.A(dpath_mulcore_ary1_a1_I2_I1_24__net32), .Y(n8610));
INVX1 mul_U21862(.A(dpath_mulcore_ary1_a1_I2_I1_23__net32), .Y(n8611));
INVX1 mul_U21863(.A(dpath_mulcore_ary1_a1_I2_I1_22__net32), .Y(n8612));
INVX1 mul_U21864(.A(dpath_mulcore_ary1_a1_I2_I1_21__net32), .Y(n8613));
INVX1 mul_U21865(.A(dpath_mulcore_ary1_a1_I2_I1_20__net32), .Y(n8614));
INVX1 mul_U21866(.A(dpath_mulcore_ary1_a1_I2_I1_19__net32), .Y(n8615));
INVX1 mul_U21867(.A(dpath_mulcore_ary1_a1_I2_I1_18__net32), .Y(n8616));
INVX1 mul_U21868(.A(dpath_mulcore_ary1_a1_I2_I1_17__net32), .Y(n8617));
INVX1 mul_U21869(.A(dpath_mulcore_ary1_a1_I2_I1_16__net32), .Y(n8618));
INVX1 mul_U21870(.A(dpath_mulcore_ary1_a1_I2_I1_15__net32), .Y(n8619));
INVX1 mul_U21871(.A(dpath_mulcore_ary1_a1_I2_I1_14__net32), .Y(n8620));
INVX1 mul_U21872(.A(dpath_mulcore_ary1_a1_I2_I1_13__net32), .Y(n8621));
INVX1 mul_U21873(.A(dpath_mulcore_ary1_a1_I2_I1_12__net32), .Y(n8622));
INVX1 mul_U21874(.A(dpath_mulcore_ary1_a1_I2_I1_11__net32), .Y(n8623));
INVX1 mul_U21875(.A(dpath_mulcore_ary1_a1_I2_I1_10__net32), .Y(n8624));
INVX1 mul_U21876(.A(dpath_mulcore_ary1_a1_I2_I1_9__net32), .Y(n8625));
INVX1 mul_U21877(.A(dpath_mulcore_ary1_a1_I2_I1_8__net32), .Y(n8626));
INVX1 mul_U21878(.A(dpath_mulcore_ary1_a1_I2_I1_7__net32), .Y(n8627));
INVX1 mul_U21879(.A(dpath_mulcore_ary1_a1_I2_I1_6__net32), .Y(n8628));
INVX1 mul_U21880(.A(dpath_mulcore_ary1_a1_I2_I1_5__net32), .Y(n8629));
INVX1 mul_U21881(.A(dpath_mulcore_ary1_a1_I2_I1_4__net32), .Y(n8630));
INVX1 mul_U21882(.A(dpath_mulcore_ary1_a1_I2_I0_p1_3), .Y(n8631));
INVX1 mul_U21883(.A(dpath_mulcore_ary1_a1_I1_I1_63__net32), .Y(n8632));
INVX1 mul_U21884(.A(dpath_mulcore_ary1_a1_I1_I1_62__net32), .Y(n8633));
INVX1 mul_U21885(.A(dpath_mulcore_ary1_a1_I1_I1_61__net32), .Y(n8634));
INVX1 mul_U21886(.A(dpath_mulcore_ary1_a1_I1_I1_60__net32), .Y(n8635));
INVX1 mul_U21887(.A(dpath_mulcore_ary1_a1_I1_I1_59__net32), .Y(n8636));
INVX1 mul_U21888(.A(dpath_mulcore_ary1_a1_I1_I1_58__net32), .Y(n8637));
INVX1 mul_U21889(.A(dpath_mulcore_ary1_a1_I1_I1_57__net32), .Y(n8638));
INVX1 mul_U21890(.A(dpath_mulcore_ary1_a1_I1_I1_56__net32), .Y(n8639));
INVX1 mul_U21891(.A(dpath_mulcore_ary1_a1_I1_I1_55__net32), .Y(n8640));
INVX1 mul_U21892(.A(dpath_mulcore_ary1_a1_I1_I1_54__net32), .Y(n8641));
INVX1 mul_U21893(.A(dpath_mulcore_ary1_a1_I1_I1_53__net32), .Y(n8642));
INVX1 mul_U21894(.A(dpath_mulcore_ary1_a1_I1_I1_52__net32), .Y(n8643));
INVX1 mul_U21895(.A(dpath_mulcore_ary1_a1_I1_I1_51__net32), .Y(n8644));
INVX1 mul_U21896(.A(dpath_mulcore_ary1_a1_I1_I1_50__net32), .Y(n8645));
INVX1 mul_U21897(.A(dpath_mulcore_ary1_a1_I1_I1_49__net32), .Y(n8646));
INVX1 mul_U21898(.A(dpath_mulcore_ary1_a1_I1_I1_48__net32), .Y(n8647));
INVX1 mul_U21899(.A(dpath_mulcore_ary1_a1_I1_I1_47__net32), .Y(n8648));
INVX1 mul_U21900(.A(dpath_mulcore_ary1_a1_I1_I1_46__net32), .Y(n8649));
INVX1 mul_U21901(.A(dpath_mulcore_ary1_a1_I1_I1_45__net32), .Y(n8650));
INVX1 mul_U21902(.A(dpath_mulcore_ary1_a1_I1_I1_44__net32), .Y(n8651));
INVX1 mul_U21903(.A(dpath_mulcore_ary1_a1_I1_I1_43__net32), .Y(n8652));
INVX1 mul_U21904(.A(dpath_mulcore_ary1_a1_I1_I1_42__net32), .Y(n8653));
INVX1 mul_U21905(.A(dpath_mulcore_ary1_a1_I1_I1_41__net32), .Y(n8654));
INVX1 mul_U21906(.A(dpath_mulcore_ary1_a1_I1_I1_40__net32), .Y(n8655));
INVX1 mul_U21907(.A(dpath_mulcore_ary1_a1_I1_I1_39__net32), .Y(n8656));
INVX1 mul_U21908(.A(dpath_mulcore_ary1_a1_I1_I1_38__net32), .Y(n8657));
INVX1 mul_U21909(.A(dpath_mulcore_ary1_a1_I1_I1_37__net32), .Y(n8658));
INVX1 mul_U21910(.A(dpath_mulcore_ary1_a1_I1_I1_36__net32), .Y(n8659));
INVX1 mul_U21911(.A(dpath_mulcore_ary1_a1_I1_I1_35__net32), .Y(n8660));
INVX1 mul_U21912(.A(dpath_mulcore_ary1_a1_I1_I1_34__net32), .Y(n8661));
INVX1 mul_U21913(.A(dpath_mulcore_ary1_a1_I1_I1_33__net32), .Y(n8662));
INVX1 mul_U21914(.A(dpath_mulcore_ary1_a1_I1_I1_32__net32), .Y(n8663));
INVX1 mul_U21915(.A(dpath_mulcore_ary1_a1_I1_I1_31__net32), .Y(n8664));
INVX1 mul_U21916(.A(dpath_mulcore_ary1_a1_I1_I1_30__net32), .Y(n8665));
INVX1 mul_U21917(.A(dpath_mulcore_ary1_a1_I1_I1_29__net32), .Y(n8666));
INVX1 mul_U21918(.A(dpath_mulcore_ary1_a1_I1_I1_28__net32), .Y(n8667));
INVX1 mul_U21919(.A(dpath_mulcore_ary1_a1_I1_I1_27__net32), .Y(n8668));
INVX1 mul_U21920(.A(dpath_mulcore_ary1_a1_I1_I1_26__net32), .Y(n8669));
INVX1 mul_U21921(.A(dpath_mulcore_ary1_a1_I1_I1_25__net32), .Y(n8670));
INVX1 mul_U21922(.A(dpath_mulcore_ary1_a1_I1_I1_24__net32), .Y(n8671));
INVX1 mul_U21923(.A(dpath_mulcore_ary1_a1_I1_I1_23__net32), .Y(n8672));
INVX1 mul_U21924(.A(dpath_mulcore_ary1_a1_I1_I1_22__net32), .Y(n8673));
INVX1 mul_U21925(.A(dpath_mulcore_ary1_a1_I1_I1_21__net32), .Y(n8674));
INVX1 mul_U21926(.A(dpath_mulcore_ary1_a1_I1_I1_20__net32), .Y(n8675));
INVX1 mul_U21927(.A(dpath_mulcore_ary1_a1_I1_I1_19__net32), .Y(n8676));
INVX1 mul_U21928(.A(dpath_mulcore_ary1_a1_I1_I1_18__net32), .Y(n8677));
INVX1 mul_U21929(.A(dpath_mulcore_ary1_a1_I1_I1_17__net32), .Y(n8678));
INVX1 mul_U21930(.A(dpath_mulcore_ary1_a1_I1_I1_16__net32), .Y(n8679));
INVX1 mul_U21931(.A(dpath_mulcore_ary1_a1_I1_I1_15__net32), .Y(n8680));
INVX1 mul_U21932(.A(dpath_mulcore_ary1_a1_I1_I1_14__net32), .Y(n8681));
INVX1 mul_U21933(.A(dpath_mulcore_ary1_a1_I1_I1_13__net32), .Y(n8682));
INVX1 mul_U21934(.A(dpath_mulcore_ary1_a1_I1_I1_12__net32), .Y(n8683));
INVX1 mul_U21935(.A(dpath_mulcore_ary1_a1_I1_I1_11__net32), .Y(n8684));
INVX1 mul_U21936(.A(dpath_mulcore_ary1_a1_I1_I1_10__net32), .Y(n8685));
INVX1 mul_U21937(.A(dpath_mulcore_ary1_a1_I1_I1_9__net32), .Y(n8686));
INVX1 mul_U21938(.A(dpath_mulcore_ary1_a1_I1_I1_8__net32), .Y(n8687));
INVX1 mul_U21939(.A(dpath_mulcore_ary1_a1_I1_I1_7__net32), .Y(n8688));
INVX1 mul_U21940(.A(dpath_mulcore_ary1_a1_I1_I1_6__net32), .Y(n8689));
INVX1 mul_U21941(.A(dpath_mulcore_ary1_a1_I1_I1_5__net32), .Y(n8690));
INVX1 mul_U21942(.A(dpath_mulcore_ary1_a1_I1_I1_4__net32), .Y(n8691));
INVX1 mul_U21943(.A(dpath_mulcore_ary1_a1_I1_I0_p1_3), .Y(n8692));
INVX1 mul_U21944(.A(dpath_mulcore_ary1_a1_I0_I1_63__net32), .Y(n8693));
INVX1 mul_U21945(.A(dpath_mulcore_ary1_a1_I0_I1_62__net32), .Y(n8694));
INVX1 mul_U21946(.A(dpath_mulcore_ary1_a1_I0_I1_61__net32), .Y(n8695));
INVX1 mul_U21947(.A(dpath_mulcore_ary1_a1_I0_I1_60__net32), .Y(n8696));
INVX1 mul_U21948(.A(dpath_mulcore_ary1_a1_I0_I1_59__net32), .Y(n8697));
INVX1 mul_U21949(.A(dpath_mulcore_ary1_a1_I0_I1_58__net32), .Y(n8698));
INVX1 mul_U21950(.A(dpath_mulcore_ary1_a1_I0_I1_57__net32), .Y(n8699));
INVX1 mul_U21951(.A(dpath_mulcore_ary1_a1_I0_I1_56__net32), .Y(n8700));
INVX1 mul_U21952(.A(dpath_mulcore_ary1_a1_I0_I1_55__net32), .Y(n8701));
INVX1 mul_U21953(.A(dpath_mulcore_ary1_a1_I0_I1_54__net32), .Y(n8702));
INVX1 mul_U21954(.A(dpath_mulcore_ary1_a1_I0_I1_53__net32), .Y(n8703));
INVX1 mul_U21955(.A(dpath_mulcore_ary1_a1_I0_I1_52__net32), .Y(n8704));
INVX1 mul_U21956(.A(dpath_mulcore_ary1_a1_I0_I1_51__net32), .Y(n8705));
INVX1 mul_U21957(.A(dpath_mulcore_ary1_a1_I0_I1_50__net32), .Y(n8706));
INVX1 mul_U21958(.A(dpath_mulcore_ary1_a1_I0_I1_49__net32), .Y(n8707));
INVX1 mul_U21959(.A(dpath_mulcore_ary1_a1_I0_I1_48__net32), .Y(n8708));
INVX1 mul_U21960(.A(dpath_mulcore_ary1_a1_I0_I1_47__net32), .Y(n8709));
INVX1 mul_U21961(.A(dpath_mulcore_ary1_a1_I0_I1_46__net32), .Y(n8710));
INVX1 mul_U21962(.A(dpath_mulcore_ary1_a1_I0_I1_45__net32), .Y(n8711));
INVX1 mul_U21963(.A(dpath_mulcore_ary1_a1_I0_I1_44__net32), .Y(n8712));
INVX1 mul_U21964(.A(dpath_mulcore_ary1_a1_I0_I1_43__net32), .Y(n8713));
INVX1 mul_U21965(.A(dpath_mulcore_ary1_a1_I0_I1_42__net32), .Y(n8714));
INVX1 mul_U21966(.A(dpath_mulcore_ary1_a1_I0_I1_41__net32), .Y(n8715));
INVX1 mul_U21967(.A(dpath_mulcore_ary1_a1_I0_I1_40__net32), .Y(n8716));
INVX1 mul_U21968(.A(dpath_mulcore_ary1_a1_I0_I1_39__net32), .Y(n8717));
INVX1 mul_U21969(.A(dpath_mulcore_ary1_a1_I0_I1_38__net32), .Y(n8718));
INVX1 mul_U21970(.A(dpath_mulcore_ary1_a1_I0_I1_37__net32), .Y(n8719));
INVX1 mul_U21971(.A(dpath_mulcore_ary1_a1_I0_I1_36__net32), .Y(n8720));
INVX1 mul_U21972(.A(dpath_mulcore_ary1_a1_I0_I1_35__net32), .Y(n8721));
INVX1 mul_U21973(.A(dpath_mulcore_ary1_a1_I0_I1_34__net32), .Y(n8722));
INVX1 mul_U21974(.A(dpath_mulcore_ary1_a1_I0_I1_33__net32), .Y(n8723));
INVX1 mul_U21975(.A(dpath_mulcore_ary1_a1_I0_I1_32__net32), .Y(n8724));
INVX1 mul_U21976(.A(dpath_mulcore_ary1_a1_I0_I1_31__net32), .Y(n8725));
INVX1 mul_U21977(.A(dpath_mulcore_ary1_a1_I0_I1_30__net32), .Y(n8726));
INVX1 mul_U21978(.A(dpath_mulcore_ary1_a1_I0_I1_29__net32), .Y(n8727));
INVX1 mul_U21979(.A(dpath_mulcore_ary1_a1_I0_I1_28__net32), .Y(n8728));
INVX1 mul_U21980(.A(dpath_mulcore_ary1_a1_I0_I1_27__net32), .Y(n8729));
INVX1 mul_U21981(.A(dpath_mulcore_ary1_a1_I0_I1_26__net32), .Y(n8730));
INVX1 mul_U21982(.A(dpath_mulcore_ary1_a1_I0_I1_25__net32), .Y(n8731));
INVX1 mul_U21983(.A(dpath_mulcore_ary1_a1_I0_I1_24__net32), .Y(n8732));
INVX1 mul_U21984(.A(dpath_mulcore_ary1_a1_I0_I1_23__net32), .Y(n8733));
INVX1 mul_U21985(.A(dpath_mulcore_ary1_a1_I0_I1_22__net32), .Y(n8734));
INVX1 mul_U21986(.A(dpath_mulcore_ary1_a1_I0_I1_21__net32), .Y(n8735));
INVX1 mul_U21987(.A(dpath_mulcore_ary1_a1_I0_I1_20__net32), .Y(n8736));
INVX1 mul_U21988(.A(dpath_mulcore_ary1_a1_I0_I1_19__net32), .Y(n8737));
INVX1 mul_U21989(.A(dpath_mulcore_ary1_a1_I0_I1_18__net32), .Y(n8738));
INVX1 mul_U21990(.A(dpath_mulcore_ary1_a1_I0_I1_17__net32), .Y(n8739));
INVX1 mul_U21991(.A(dpath_mulcore_ary1_a1_I0_I1_16__net32), .Y(n8740));
INVX1 mul_U21992(.A(dpath_mulcore_ary1_a1_I0_I1_15__net32), .Y(n8741));
INVX1 mul_U21993(.A(dpath_mulcore_ary1_a1_I0_I1_14__net32), .Y(n8742));
INVX1 mul_U21994(.A(dpath_mulcore_ary1_a1_I0_I1_13__net32), .Y(n8743));
INVX1 mul_U21995(.A(dpath_mulcore_ary1_a1_I0_I1_12__net32), .Y(n8744));
INVX1 mul_U21996(.A(dpath_mulcore_ary1_a1_I0_I1_11__net32), .Y(n8745));
INVX1 mul_U21997(.A(dpath_mulcore_ary1_a1_I0_I1_10__net32), .Y(n8746));
INVX1 mul_U21998(.A(dpath_mulcore_ary1_a1_I0_I1_9__net32), .Y(n8747));
INVX1 mul_U21999(.A(dpath_mulcore_ary1_a1_I0_I1_8__net32), .Y(n8748));
INVX1 mul_U22000(.A(dpath_mulcore_ary1_a1_I0_I1_7__net32), .Y(n8749));
INVX1 mul_U22001(.A(dpath_mulcore_ary1_a1_I0_I1_6__net32), .Y(n8750));
INVX1 mul_U22002(.A(dpath_mulcore_ary1_a1_I0_I1_5__net32), .Y(n8751));
INVX1 mul_U22003(.A(dpath_mulcore_ary1_a1_I0_I1_4__net32), .Y(n8752));
INVX1 mul_U22004(.A(dpath_mulcore_ary1_a1_I0_I0_p1_3), .Y(n8753));
INVX1 mul_U22005(.A(dpath_mulcore_ary1_a0_I1_I2_net47), .Y(n8754));
INVX1 mul_U22006(.A(dpath_mulcore_ary1_a0_I0_I2_net47), .Y(n8755));
INVX1 mul_U22007(.A(dpath_mulcore_ary1_a1_I2_I2_net47), .Y(n8756));
INVX1 mul_U22008(.A(dpath_mulcore_ary1_a1_I1_I2_net47), .Y(n8757));
INVX1 mul_U22009(.A(dpath_mulcore_ary1_a1_I0_I2_net47), .Y(n8758));
INVX1 mul_U22010(.A(dpath_mulcore_ary1_a0_c0[3]), .Y(n8759));
INVX1 mul_U22011(.A(dpath_mulcore_ary1_a0_c0[2]), .Y(n8760));
INVX1 mul_U22012(.A(dpath_mulcore_ary1_a1_c2[3]), .Y(n8761));
INVX1 mul_U22013(.A(dpath_mulcore_ary1_a1_c2[2]), .Y(n8762));
INVX1 mul_U22014(.A(dpath_mulcore_ary1_a1_c0[3]), .Y(n8763));
INVX1 mul_U22015(.A(dpath_mulcore_ary1_a1_c0[2]), .Y(n8764));
INVX1 mul_U22016(.A(dpath_mulcore_ary1_a0_c0[63]), .Y(n8765));
INVX1 mul_U22017(.A(dpath_mulcore_ary1_a0_c0[62]), .Y(n8766));
INVX1 mul_U22018(.A(dpath_mulcore_ary1_a0_c0[61]), .Y(n8767));
INVX1 mul_U22019(.A(dpath_mulcore_ary1_a0_c0[60]), .Y(n8768));
INVX1 mul_U22020(.A(dpath_mulcore_ary1_a0_c0[59]), .Y(n8769));
INVX1 mul_U22021(.A(dpath_mulcore_ary1_a0_c0[58]), .Y(n8770));
INVX1 mul_U22022(.A(dpath_mulcore_ary1_a0_c0[57]), .Y(n8771));
INVX1 mul_U22023(.A(dpath_mulcore_ary1_a0_c0[56]), .Y(n8772));
INVX1 mul_U22024(.A(dpath_mulcore_ary1_a0_c0[55]), .Y(n8773));
INVX1 mul_U22025(.A(dpath_mulcore_ary1_a0_c0[54]), .Y(n8774));
INVX1 mul_U22026(.A(dpath_mulcore_ary1_a0_c0[53]), .Y(n8775));
INVX1 mul_U22027(.A(dpath_mulcore_ary1_a0_c0[52]), .Y(n8776));
INVX1 mul_U22028(.A(dpath_mulcore_ary1_a0_c0[51]), .Y(n8777));
INVX1 mul_U22029(.A(dpath_mulcore_ary1_a0_c0[50]), .Y(n8778));
INVX1 mul_U22030(.A(dpath_mulcore_ary1_a0_c0[49]), .Y(n8779));
INVX1 mul_U22031(.A(dpath_mulcore_ary1_a0_c0[48]), .Y(n8780));
INVX1 mul_U22032(.A(dpath_mulcore_ary1_a0_c0[47]), .Y(n8781));
INVX1 mul_U22033(.A(dpath_mulcore_ary1_a0_c0[46]), .Y(n8782));
INVX1 mul_U22034(.A(dpath_mulcore_ary1_a0_c0[45]), .Y(n8783));
INVX1 mul_U22035(.A(dpath_mulcore_ary1_a0_c0[44]), .Y(n8784));
INVX1 mul_U22036(.A(dpath_mulcore_ary1_a0_c0[43]), .Y(n8785));
INVX1 mul_U22037(.A(dpath_mulcore_ary1_a0_c0[42]), .Y(n8786));
INVX1 mul_U22038(.A(dpath_mulcore_ary1_a0_c0[41]), .Y(n8787));
INVX1 mul_U22039(.A(dpath_mulcore_ary1_a0_c0[40]), .Y(n8788));
INVX1 mul_U22040(.A(dpath_mulcore_ary1_a0_c0[39]), .Y(n8789));
INVX1 mul_U22041(.A(dpath_mulcore_ary1_a0_c0[38]), .Y(n8790));
INVX1 mul_U22042(.A(dpath_mulcore_ary1_a0_c0[37]), .Y(n8791));
INVX1 mul_U22043(.A(dpath_mulcore_ary1_a0_c0[36]), .Y(n8792));
INVX1 mul_U22044(.A(dpath_mulcore_ary1_a0_c0[35]), .Y(n8793));
INVX1 mul_U22045(.A(dpath_mulcore_ary1_a0_c0[34]), .Y(n8794));
INVX1 mul_U22046(.A(dpath_mulcore_ary1_a0_c0[33]), .Y(n8795));
INVX1 mul_U22047(.A(dpath_mulcore_ary1_a0_c0[32]), .Y(n8796));
INVX1 mul_U22048(.A(dpath_mulcore_ary1_a0_c0[31]), .Y(n8797));
INVX1 mul_U22049(.A(dpath_mulcore_ary1_a0_c0[30]), .Y(n8798));
INVX1 mul_U22050(.A(dpath_mulcore_ary1_a0_c0[29]), .Y(n8799));
INVX1 mul_U22051(.A(dpath_mulcore_ary1_a0_c0[28]), .Y(n8800));
INVX1 mul_U22052(.A(dpath_mulcore_ary1_a0_c0[27]), .Y(n8801));
INVX1 mul_U22053(.A(dpath_mulcore_ary1_a0_c0[26]), .Y(n8802));
INVX1 mul_U22054(.A(dpath_mulcore_ary1_a0_c0[25]), .Y(n8803));
INVX1 mul_U22055(.A(dpath_mulcore_ary1_a0_c0[24]), .Y(n8804));
INVX1 mul_U22056(.A(dpath_mulcore_ary1_a0_c0[23]), .Y(n8805));
INVX1 mul_U22057(.A(dpath_mulcore_ary1_a0_c0[22]), .Y(n8806));
INVX1 mul_U22058(.A(dpath_mulcore_ary1_a0_c0[21]), .Y(n8807));
INVX1 mul_U22059(.A(dpath_mulcore_ary1_a0_c0[20]), .Y(n8808));
INVX1 mul_U22060(.A(dpath_mulcore_ary1_a0_c0[19]), .Y(n8809));
INVX1 mul_U22061(.A(dpath_mulcore_ary1_a0_c0[18]), .Y(n8810));
INVX1 mul_U22062(.A(dpath_mulcore_ary1_a0_c0[17]), .Y(n8811));
INVX1 mul_U22063(.A(dpath_mulcore_ary1_a0_c0[16]), .Y(n8812));
INVX1 mul_U22064(.A(dpath_mulcore_ary1_a0_c0[15]), .Y(n8813));
INVX1 mul_U22065(.A(dpath_mulcore_ary1_a0_c0[14]), .Y(n8814));
INVX1 mul_U22066(.A(dpath_mulcore_ary1_a0_c0[13]), .Y(n8815));
INVX1 mul_U22067(.A(dpath_mulcore_ary1_a0_c0[8]), .Y(n8816));
INVX1 mul_U22068(.A(dpath_mulcore_ary1_a0_c0[7]), .Y(n8817));
INVX1 mul_U22069(.A(dpath_mulcore_ary1_a0_c0[6]), .Y(n8818));
INVX1 mul_U22070(.A(dpath_mulcore_ary1_a0_c0[5]), .Y(n8819));
INVX1 mul_U22071(.A(dpath_mulcore_ary1_a0_c0[4]), .Y(n8820));
INVX1 mul_U22072(.A(dpath_mulcore_ary1_a1_c2[63]), .Y(n8821));
INVX1 mul_U22073(.A(dpath_mulcore_ary1_a1_c2[62]), .Y(n8822));
INVX1 mul_U22074(.A(dpath_mulcore_ary1_a1_c2[61]), .Y(n8823));
INVX1 mul_U22075(.A(dpath_mulcore_ary1_a1_c2[60]), .Y(n8824));
INVX1 mul_U22076(.A(dpath_mulcore_ary1_a1_c2[59]), .Y(n8825));
INVX1 mul_U22077(.A(dpath_mulcore_ary1_a1_c2[58]), .Y(n8826));
INVX1 mul_U22078(.A(dpath_mulcore_ary1_a1_c2[57]), .Y(n8827));
INVX1 mul_U22079(.A(dpath_mulcore_ary1_a1_c2[56]), .Y(n8828));
INVX1 mul_U22080(.A(dpath_mulcore_ary1_a1_c2[55]), .Y(n8829));
INVX1 mul_U22081(.A(dpath_mulcore_ary1_a1_c2[54]), .Y(n8830));
INVX1 mul_U22082(.A(dpath_mulcore_ary1_a1_c2[53]), .Y(n8831));
INVX1 mul_U22083(.A(dpath_mulcore_ary1_a1_c2[52]), .Y(n8832));
INVX1 mul_U22084(.A(dpath_mulcore_ary1_a1_c2[51]), .Y(n8833));
INVX1 mul_U22085(.A(dpath_mulcore_ary1_a1_c2[50]), .Y(n8834));
INVX1 mul_U22086(.A(dpath_mulcore_ary1_a1_c2[49]), .Y(n8835));
INVX1 mul_U22087(.A(dpath_mulcore_ary1_a1_c2[48]), .Y(n8836));
INVX1 mul_U22088(.A(dpath_mulcore_ary1_a1_c2[47]), .Y(n8837));
INVX1 mul_U22089(.A(dpath_mulcore_ary1_a1_c2[46]), .Y(n8838));
INVX1 mul_U22090(.A(dpath_mulcore_ary1_a1_c2[45]), .Y(n8839));
INVX1 mul_U22091(.A(dpath_mulcore_ary1_a1_c2[44]), .Y(n8840));
INVX1 mul_U22092(.A(dpath_mulcore_ary1_a1_c2[43]), .Y(n8841));
INVX1 mul_U22093(.A(dpath_mulcore_ary1_a1_c2[42]), .Y(n8842));
INVX1 mul_U22094(.A(dpath_mulcore_ary1_a1_c2[41]), .Y(n8843));
INVX1 mul_U22095(.A(dpath_mulcore_ary1_a1_c2[40]), .Y(n8844));
INVX1 mul_U22096(.A(dpath_mulcore_ary1_a1_c2[39]), .Y(n8845));
INVX1 mul_U22097(.A(dpath_mulcore_ary1_a1_c2[38]), .Y(n8846));
INVX1 mul_U22098(.A(dpath_mulcore_ary1_a1_c2[37]), .Y(n8847));
INVX1 mul_U22099(.A(dpath_mulcore_ary1_a1_c2[36]), .Y(n8848));
INVX1 mul_U22100(.A(dpath_mulcore_ary1_a1_c2[35]), .Y(n8849));
INVX1 mul_U22101(.A(dpath_mulcore_ary1_a1_c2[34]), .Y(n8850));
INVX1 mul_U22102(.A(dpath_mulcore_ary1_a1_c2[33]), .Y(n8851));
INVX1 mul_U22103(.A(dpath_mulcore_ary1_a1_c2[32]), .Y(n8852));
INVX1 mul_U22104(.A(dpath_mulcore_ary1_a1_c2[31]), .Y(n8853));
INVX1 mul_U22105(.A(dpath_mulcore_ary1_a1_c2[30]), .Y(n8854));
INVX1 mul_U22106(.A(dpath_mulcore_ary1_a1_c2[29]), .Y(n8855));
INVX1 mul_U22107(.A(dpath_mulcore_ary1_a1_c2[28]), .Y(n8856));
INVX1 mul_U22108(.A(dpath_mulcore_ary1_a1_c2[27]), .Y(n8857));
INVX1 mul_U22109(.A(dpath_mulcore_ary1_a1_c2[26]), .Y(n8858));
INVX1 mul_U22110(.A(dpath_mulcore_ary1_a1_c2[25]), .Y(n8859));
INVX1 mul_U22111(.A(dpath_mulcore_ary1_a1_c2[24]), .Y(n8860));
INVX1 mul_U22112(.A(dpath_mulcore_ary1_a1_c2[23]), .Y(n8861));
INVX1 mul_U22113(.A(dpath_mulcore_ary1_a1_c2[22]), .Y(n8862));
INVX1 mul_U22114(.A(dpath_mulcore_ary1_a1_c2[21]), .Y(n8863));
INVX1 mul_U22115(.A(dpath_mulcore_ary1_a1_c2[20]), .Y(n8864));
INVX1 mul_U22116(.A(dpath_mulcore_ary1_a1_c2[19]), .Y(n8865));
INVX1 mul_U22117(.A(dpath_mulcore_ary1_a1_c2[18]), .Y(n8866));
INVX1 mul_U22118(.A(dpath_mulcore_ary1_a1_c2[17]), .Y(n8867));
INVX1 mul_U22119(.A(dpath_mulcore_ary1_a1_c2[16]), .Y(n8868));
INVX1 mul_U22120(.A(dpath_mulcore_ary1_a1_c2[15]), .Y(n8869));
INVX1 mul_U22121(.A(dpath_mulcore_ary1_a1_c2[14]), .Y(n8870));
INVX1 mul_U22122(.A(dpath_mulcore_ary1_a1_c2[13]), .Y(n8871));
INVX1 mul_U22123(.A(dpath_mulcore_ary1_a1_c2[12]), .Y(n8872));
INVX1 mul_U22124(.A(dpath_mulcore_ary1_a1_c2[11]), .Y(n8873));
INVX1 mul_U22125(.A(dpath_mulcore_ary1_a1_c2[10]), .Y(n8874));
INVX1 mul_U22126(.A(dpath_mulcore_ary1_a1_c2[9]), .Y(n8875));
INVX1 mul_U22127(.A(dpath_mulcore_ary1_a1_c2[8]), .Y(n8876));
INVX1 mul_U22128(.A(dpath_mulcore_ary1_a1_c2[7]), .Y(n8877));
INVX1 mul_U22129(.A(dpath_mulcore_ary1_a1_c2[6]), .Y(n8878));
INVX1 mul_U22130(.A(dpath_mulcore_ary1_a1_c2[5]), .Y(n8879));
INVX1 mul_U22131(.A(dpath_mulcore_ary1_a1_c2[4]), .Y(n8880));
INVX1 mul_U22132(.A(dpath_mulcore_ary1_a1_c0[63]), .Y(n8881));
INVX1 mul_U22133(.A(dpath_mulcore_ary1_a1_c0[62]), .Y(n8882));
INVX1 mul_U22134(.A(dpath_mulcore_ary1_a1_c0[61]), .Y(n8883));
INVX1 mul_U22135(.A(dpath_mulcore_ary1_a1_c0[60]), .Y(n8884));
INVX1 mul_U22136(.A(dpath_mulcore_ary1_a1_c0[59]), .Y(n8885));
INVX1 mul_U22137(.A(dpath_mulcore_ary1_a1_c0[58]), .Y(n8886));
INVX1 mul_U22138(.A(dpath_mulcore_ary1_a1_c0[57]), .Y(n8887));
INVX1 mul_U22139(.A(dpath_mulcore_ary1_a1_c0[56]), .Y(n8888));
INVX1 mul_U22140(.A(dpath_mulcore_ary1_a1_c0[55]), .Y(n8889));
INVX1 mul_U22141(.A(dpath_mulcore_ary1_a1_c0[54]), .Y(n8890));
INVX1 mul_U22142(.A(dpath_mulcore_ary1_a1_c0[53]), .Y(n8891));
INVX1 mul_U22143(.A(dpath_mulcore_ary1_a1_c0[52]), .Y(n8892));
INVX1 mul_U22144(.A(dpath_mulcore_ary1_a1_c0[51]), .Y(n8893));
INVX1 mul_U22145(.A(dpath_mulcore_ary1_a1_c0[50]), .Y(n8894));
INVX1 mul_U22146(.A(dpath_mulcore_ary1_a1_c0[49]), .Y(n8895));
INVX1 mul_U22147(.A(dpath_mulcore_ary1_a1_c0[48]), .Y(n8896));
INVX1 mul_U22148(.A(dpath_mulcore_ary1_a1_c0[47]), .Y(n8897));
INVX1 mul_U22149(.A(dpath_mulcore_ary1_a1_c0[46]), .Y(n8898));
INVX1 mul_U22150(.A(dpath_mulcore_ary1_a1_c0[45]), .Y(n8899));
INVX1 mul_U22151(.A(dpath_mulcore_ary1_a1_c0[44]), .Y(n8900));
INVX1 mul_U22152(.A(dpath_mulcore_ary1_a1_c0[43]), .Y(n8901));
INVX1 mul_U22153(.A(dpath_mulcore_ary1_a1_c0[42]), .Y(n8902));
INVX1 mul_U22154(.A(dpath_mulcore_ary1_a1_c0[41]), .Y(n8903));
INVX1 mul_U22155(.A(dpath_mulcore_ary1_a1_c0[40]), .Y(n8904));
INVX1 mul_U22156(.A(dpath_mulcore_ary1_a1_c0[39]), .Y(n8905));
INVX1 mul_U22157(.A(dpath_mulcore_ary1_a1_c0[38]), .Y(n8906));
INVX1 mul_U22158(.A(dpath_mulcore_ary1_a1_c0[37]), .Y(n8907));
INVX1 mul_U22159(.A(dpath_mulcore_ary1_a1_c0[36]), .Y(n8908));
INVX1 mul_U22160(.A(dpath_mulcore_ary1_a1_c0[35]), .Y(n8909));
INVX1 mul_U22161(.A(dpath_mulcore_ary1_a1_c0[34]), .Y(n8910));
INVX1 mul_U22162(.A(dpath_mulcore_ary1_a1_c0[33]), .Y(n8911));
INVX1 mul_U22163(.A(dpath_mulcore_ary1_a1_c0[32]), .Y(n8912));
INVX1 mul_U22164(.A(dpath_mulcore_ary1_a1_c0[31]), .Y(n8913));
INVX1 mul_U22165(.A(dpath_mulcore_ary1_a1_c0[30]), .Y(n8914));
INVX1 mul_U22166(.A(dpath_mulcore_ary1_a1_c0[29]), .Y(n8915));
INVX1 mul_U22167(.A(dpath_mulcore_ary1_a1_c0[28]), .Y(n8916));
INVX1 mul_U22168(.A(dpath_mulcore_ary1_a1_c0[27]), .Y(n8917));
INVX1 mul_U22169(.A(dpath_mulcore_ary1_a1_c0[26]), .Y(n8918));
INVX1 mul_U22170(.A(dpath_mulcore_ary1_a1_c0[25]), .Y(n8919));
INVX1 mul_U22171(.A(dpath_mulcore_ary1_a1_c0[24]), .Y(n8920));
INVX1 mul_U22172(.A(dpath_mulcore_ary1_a1_c0[23]), .Y(n8921));
INVX1 mul_U22173(.A(dpath_mulcore_ary1_a1_c0[22]), .Y(n8922));
INVX1 mul_U22174(.A(dpath_mulcore_ary1_a1_c0[21]), .Y(n8923));
INVX1 mul_U22175(.A(dpath_mulcore_ary1_a1_c0[20]), .Y(n8924));
INVX1 mul_U22176(.A(dpath_mulcore_ary1_a1_c0[19]), .Y(n8925));
INVX1 mul_U22177(.A(dpath_mulcore_ary1_a1_c0[18]), .Y(n8926));
INVX1 mul_U22178(.A(dpath_mulcore_ary1_a1_c0[17]), .Y(n8927));
INVX1 mul_U22179(.A(dpath_mulcore_ary1_a1_c0[16]), .Y(n8928));
INVX1 mul_U22180(.A(dpath_mulcore_ary1_a1_c0[15]), .Y(n8929));
INVX1 mul_U22181(.A(dpath_mulcore_ary1_a1_c0[14]), .Y(n8930));
INVX1 mul_U22182(.A(dpath_mulcore_ary1_a1_c0[13]), .Y(n8931));
INVX1 mul_U22183(.A(dpath_mulcore_ary1_a1_c0[8]), .Y(n8932));
INVX1 mul_U22184(.A(dpath_mulcore_ary1_a1_c0[7]), .Y(n8933));
INVX1 mul_U22185(.A(dpath_mulcore_ary1_a1_c0[6]), .Y(n8934));
INVX1 mul_U22186(.A(dpath_mulcore_ary1_a1_c0[5]), .Y(n8935));
INVX1 mul_U22187(.A(dpath_mulcore_ary1_a1_c0[4]), .Y(n8936));
INVX1 mul_U22188(.A(dpath_mulcore_ary1_a0_c0[64]), .Y(n8937));
INVX1 mul_U22189(.A(dpath_mulcore_ary1_a0_c0[65]), .Y(n8938));
INVX1 mul_U22190(.A(dpath_mulcore_ary1_a0_c0[66]), .Y(n8939));
INVX1 mul_U22191(.A(dpath_mulcore_ary1_a0_c0[67]), .Y(n8940));
INVX1 mul_U22192(.A(dpath_mulcore_ary1_a1_c2[64]), .Y(n8941));
INVX1 mul_U22193(.A(dpath_mulcore_ary1_a1_c0[64]), .Y(n8942));
INVX1 mul_U22194(.A(dpath_mulcore_ary1_a1_c0[65]), .Y(n8943));
INVX1 mul_U22195(.A(dpath_mulcore_ary1_a1_c0[66]), .Y(n8944));
INVX1 mul_U22196(.A(dpath_mulcore_array2_c1[18]), .Y(n8945));
INVX1 mul_U22197(.A(dpath_mulcore_array2_c1[17]), .Y(n8946));
INVX1 mul_U22198(.A(dpath_mulcore_array2_c1[16]), .Y(n8947));
INVX1 mul_U22199(.A(dpath_mulcore_array2_c1[81]), .Y(n8948));
INVX1 mul_U22200(.A(dpath_mulcore_array2_c1[80]), .Y(n8949));
INVX1 mul_U22201(.A(dpath_mulcore_array2_c1[79]), .Y(n8950));
INVX1 mul_U22202(.A(dpath_mulcore_array2_c1[78]), .Y(n8951));
INVX1 mul_U22203(.A(dpath_mulcore_array2_c1[77]), .Y(n8952));
INVX1 mul_U22204(.A(dpath_mulcore_array2_c1[76]), .Y(n8953));
INVX1 mul_U22205(.A(dpath_mulcore_array2_c1[75]), .Y(n8954));
INVX1 mul_U22206(.A(dpath_mulcore_array2_c1[74]), .Y(n8955));
INVX1 mul_U22207(.A(dpath_mulcore_array2_c1[73]), .Y(n8956));
INVX1 mul_U22208(.A(dpath_mulcore_array2_c1[72]), .Y(n8957));
INVX1 mul_U22209(.A(dpath_mulcore_array2_c1[71]), .Y(n8958));
INVX1 mul_U22210(.A(dpath_mulcore_array2_c1[70]), .Y(n8959));
INVX1 mul_U22211(.A(dpath_mulcore_array2_c1[69]), .Y(n8960));
INVX1 mul_U22212(.A(dpath_mulcore_array2_c1[68]), .Y(n8961));
INVX1 mul_U22213(.A(dpath_mulcore_array2_c1[14]), .Y(n8962));
INVX1 mul_U22214(.A(dpath_mulcore_array2_c1[13]), .Y(n8963));
INVX1 mul_U22215(.A(dpath_mulcore_array2_c1[12]), .Y(n8964));
INVX1 mul_U22216(.A(dpath_mulcore_array2_c1[11]), .Y(n8965));
INVX1 mul_U22217(.A(dpath_mulcore_array2_c1[10]), .Y(n8966));
INVX1 mul_U22218(.A(dpath_mulcore_array2_c1[9]), .Y(n8967));
INVX1 mul_U22219(.A(dpath_mulcore_array2_c1[8]), .Y(n8968));
INVX1 mul_U22220(.A(dpath_mulcore_array2_c1[7]), .Y(n8969));
INVX1 mul_U22221(.A(dpath_mulcore_array2_c1[6]), .Y(n8970));
INVX1 mul_U22222(.A(dpath_mulcore_array2_c1[5]), .Y(n8971));
INVX1 mul_U22223(.A(dpath_mulcore_array2_c1[4]), .Y(n8972));
INVX1 mul_U22224(.A(dpath_mulcore_array2_c1[66]), .Y(n8973));
INVX1 mul_U22225(.A(dpath_mulcore_array2_c1[67]), .Y(n8974));
INVX1 mul_U22226(.A(dpath_mulcore_ary1_a0_c2[2]), .Y(n8975));
INVX1 mul_U22227(.A(dpath_mulcore_ary1_a0_c2[3]), .Y(n8976));
INVX1 mul_U22228(.A(dpath_mulcore_ary1_a0_I2_I2_net47), .Y(n8977));
INVX1 mul_U22229(.A(dpath_mulcore_ary1_a0_c_2[69]), .Y(n8978));
INVX1 mul_U22230(.A(dpath_mulcore_ary1_a0_c_2[68]), .Y(n8979));
INVX1 mul_U22231(.A(dpath_mulcore_ary1_a0_c_2[67]), .Y(n8980));
INVX1 mul_U22232(.A(dpath_mulcore_ary1_a0_c_2[66]), .Y(n8981));
INVX1 mul_U22233(.A(dpath_mulcore_ary1_a0_c_2[65]), .Y(n8982));
INVX1 mul_U22234(.A(dpath_mulcore_ary1_a0_c_2[64]), .Y(n8983));
INVX1 mul_U22235(.A(dpath_mulcore_ary1_a0_c_2[63]), .Y(n8984));
INVX1 mul_U22236(.A(dpath_mulcore_ary1_a0_c_2[62]), .Y(n8985));
INVX1 mul_U22237(.A(dpath_mulcore_ary1_a0_c_2[61]), .Y(n8986));
INVX1 mul_U22238(.A(dpath_mulcore_ary1_a0_c_2[60]), .Y(n8987));
INVX1 mul_U22239(.A(dpath_mulcore_ary1_a0_c_2[59]), .Y(n8988));
INVX1 mul_U22240(.A(dpath_mulcore_ary1_a0_c_2[58]), .Y(n8989));
INVX1 mul_U22241(.A(dpath_mulcore_ary1_a0_c_2[57]), .Y(n8990));
INVX1 mul_U22242(.A(dpath_mulcore_ary1_a0_c_2[56]), .Y(n8991));
INVX1 mul_U22243(.A(dpath_mulcore_ary1_a0_c_2[55]), .Y(n8992));
INVX1 mul_U22244(.A(dpath_mulcore_ary1_a0_c_2[54]), .Y(n8993));
INVX1 mul_U22245(.A(dpath_mulcore_ary1_a0_c_2[53]), .Y(n8994));
INVX1 mul_U22246(.A(dpath_mulcore_ary1_a0_c_2[52]), .Y(n8995));
INVX1 mul_U22247(.A(dpath_mulcore_ary1_a0_c_2[51]), .Y(n8996));
INVX1 mul_U22248(.A(dpath_mulcore_ary1_a0_c_2[50]), .Y(n8997));
INVX1 mul_U22249(.A(dpath_mulcore_ary1_a0_c_2[49]), .Y(n8998));
INVX1 mul_U22250(.A(dpath_mulcore_ary1_a0_c_2[48]), .Y(n8999));
INVX1 mul_U22251(.A(dpath_mulcore_ary1_a0_c_2[47]), .Y(n9000));
INVX1 mul_U22252(.A(dpath_mulcore_ary1_a0_c_2[46]), .Y(n9001));
INVX1 mul_U22253(.A(dpath_mulcore_ary1_a0_c_2[45]), .Y(n9002));
INVX1 mul_U22254(.A(dpath_mulcore_ary1_a0_c_2[44]), .Y(n9003));
INVX1 mul_U22255(.A(dpath_mulcore_ary1_a0_c_2[43]), .Y(n9004));
INVX1 mul_U22256(.A(dpath_mulcore_ary1_a0_c_2[42]), .Y(n9005));
INVX1 mul_U22257(.A(dpath_mulcore_ary1_a0_c_2[41]), .Y(n9006));
INVX1 mul_U22258(.A(dpath_mulcore_ary1_a0_c_2[40]), .Y(n9007));
INVX1 mul_U22259(.A(dpath_mulcore_ary1_a0_c_2[39]), .Y(n9008));
INVX1 mul_U22260(.A(dpath_mulcore_ary1_a0_c_2[38]), .Y(n9009));
INVX1 mul_U22261(.A(dpath_mulcore_ary1_a0_c_2[37]), .Y(n9010));
INVX1 mul_U22262(.A(dpath_mulcore_ary1_a0_c_2[36]), .Y(n9011));
INVX1 mul_U22263(.A(dpath_mulcore_ary1_a0_c_2[35]), .Y(n9012));
INVX1 mul_U22264(.A(dpath_mulcore_ary1_a0_c_2[34]), .Y(n9013));
INVX1 mul_U22265(.A(dpath_mulcore_ary1_a0_c_2[33]), .Y(n9014));
INVX1 mul_U22266(.A(dpath_mulcore_ary1_a0_c_2[32]), .Y(n9015));
INVX1 mul_U22267(.A(dpath_mulcore_ary1_a0_c_2[31]), .Y(n9016));
INVX1 mul_U22268(.A(dpath_mulcore_ary1_a0_c_2[30]), .Y(n9017));
INVX1 mul_U22269(.A(dpath_mulcore_ary1_a0_c_2[29]), .Y(n9018));
INVX1 mul_U22270(.A(dpath_mulcore_ary1_a0_c_2[28]), .Y(n9019));
INVX1 mul_U22271(.A(dpath_mulcore_ary1_a0_c_2[27]), .Y(n9020));
INVX1 mul_U22272(.A(dpath_mulcore_ary1_a0_c_2[26]), .Y(n9021));
INVX1 mul_U22273(.A(dpath_mulcore_ary1_a0_c_2[25]), .Y(n9022));
INVX1 mul_U22274(.A(dpath_mulcore_ary1_a0_c_2[24]), .Y(n9023));
INVX1 mul_U22275(.A(dpath_mulcore_ary1_a0_c_2[23]), .Y(n9024));
INVX1 mul_U22276(.A(dpath_mulcore_ary1_a0_c_2[22]), .Y(n9025));
INVX1 mul_U22277(.A(dpath_mulcore_ary1_a0_c_2[21]), .Y(n9026));
INVX1 mul_U22278(.A(dpath_mulcore_ary1_a0_c_2[20]), .Y(n9027));
INVX1 mul_U22279(.A(dpath_mulcore_ary1_a0_c_2[19]), .Y(n9028));
INVX1 mul_U22280(.A(dpath_mulcore_ary1_a0_c_2[18]), .Y(n9029));
INVX1 mul_U22281(.A(dpath_mulcore_ary1_a0_c_2[17]), .Y(n9030));
INVX1 mul_U22282(.A(dpath_mulcore_ary1_a0_c_2[16]), .Y(n9031));
INVX1 mul_U22283(.A(dpath_mulcore_ary1_a0_c_2[15]), .Y(n9032));
INVX1 mul_U22284(.A(dpath_mulcore_ary1_a0_c_2[14]), .Y(n9033));
INVX1 mul_U22285(.A(dpath_mulcore_ary1_a0_c_2[13]), .Y(n9034));
INVX1 mul_U22286(.A(dpath_mulcore_ary1_a0_c_2[12]), .Y(n9035));
INVX1 mul_U22287(.A(dpath_mulcore_ary1_a0_c_2[11]), .Y(n9036));
INVX1 mul_U22288(.A(dpath_mulcore_ary1_a0_c_2[10]), .Y(n9037));
INVX1 mul_U22289(.A(dpath_mulcore_ary1_a1_c_2[70]), .Y(n9038));
INVX1 mul_U22290(.A(dpath_mulcore_ary1_a1_c_2[69]), .Y(n9039));
INVX1 mul_U22291(.A(dpath_mulcore_ary1_a1_c_2[68]), .Y(n9040));
INVX1 mul_U22292(.A(dpath_mulcore_ary1_a1_c_2[67]), .Y(n9041));
INVX1 mul_U22293(.A(dpath_mulcore_ary1_a1_c_2[66]), .Y(n9042));
INVX1 mul_U22294(.A(dpath_mulcore_ary1_a1_c_2[65]), .Y(n9043));
INVX1 mul_U22295(.A(dpath_mulcore_ary1_a1_c_2[64]), .Y(n9044));
INVX1 mul_U22296(.A(dpath_mulcore_ary1_a1_c_2[63]), .Y(n9045));
INVX1 mul_U22297(.A(dpath_mulcore_ary1_a1_c_2[62]), .Y(n9046));
INVX1 mul_U22298(.A(dpath_mulcore_ary1_a1_c_2[61]), .Y(n9047));
INVX1 mul_U22299(.A(dpath_mulcore_ary1_a1_c_2[60]), .Y(n9048));
INVX1 mul_U22300(.A(dpath_mulcore_ary1_a1_c_2[59]), .Y(n9049));
INVX1 mul_U22301(.A(dpath_mulcore_ary1_a1_c_2[58]), .Y(n9050));
INVX1 mul_U22302(.A(dpath_mulcore_ary1_a1_c_2[57]), .Y(n9051));
INVX1 mul_U22303(.A(dpath_mulcore_ary1_a1_c_2[56]), .Y(n9052));
INVX1 mul_U22304(.A(dpath_mulcore_ary1_a1_c_2[55]), .Y(n9053));
INVX1 mul_U22305(.A(dpath_mulcore_ary1_a1_c_2[54]), .Y(n9054));
INVX1 mul_U22306(.A(dpath_mulcore_ary1_a1_c_2[53]), .Y(n9055));
INVX1 mul_U22307(.A(dpath_mulcore_ary1_a1_c_2[52]), .Y(n9056));
INVX1 mul_U22308(.A(dpath_mulcore_ary1_a1_c_2[51]), .Y(n9057));
INVX1 mul_U22309(.A(dpath_mulcore_ary1_a1_c_2[50]), .Y(n9058));
INVX1 mul_U22310(.A(dpath_mulcore_ary1_a1_c_2[49]), .Y(n9059));
INVX1 mul_U22311(.A(dpath_mulcore_ary1_a1_c_2[48]), .Y(n9060));
INVX1 mul_U22312(.A(dpath_mulcore_ary1_a1_c_2[47]), .Y(n9061));
INVX1 mul_U22313(.A(dpath_mulcore_ary1_a1_c_2[46]), .Y(n9062));
INVX1 mul_U22314(.A(dpath_mulcore_ary1_a1_c_2[45]), .Y(n9063));
INVX1 mul_U22315(.A(dpath_mulcore_ary1_a1_c_2[44]), .Y(n9064));
INVX1 mul_U22316(.A(dpath_mulcore_ary1_a1_c_2[43]), .Y(n9065));
INVX1 mul_U22317(.A(dpath_mulcore_ary1_a1_c_2[42]), .Y(n9066));
INVX1 mul_U22318(.A(dpath_mulcore_ary1_a1_c_2[41]), .Y(n9067));
INVX1 mul_U22319(.A(dpath_mulcore_ary1_a1_c_2[40]), .Y(n9068));
INVX1 mul_U22320(.A(dpath_mulcore_ary1_a1_c_2[39]), .Y(n9069));
INVX1 mul_U22321(.A(dpath_mulcore_ary1_a1_c_2[38]), .Y(n9070));
INVX1 mul_U22322(.A(dpath_mulcore_ary1_a1_c_2[37]), .Y(n9071));
INVX1 mul_U22323(.A(dpath_mulcore_ary1_a1_c_2[36]), .Y(n9072));
INVX1 mul_U22324(.A(dpath_mulcore_ary1_a1_c_2[35]), .Y(n9073));
INVX1 mul_U22325(.A(dpath_mulcore_ary1_a1_c_2[34]), .Y(n9074));
INVX1 mul_U22326(.A(dpath_mulcore_ary1_a1_c_2[33]), .Y(n9075));
INVX1 mul_U22327(.A(dpath_mulcore_ary1_a1_c_2[32]), .Y(n9076));
INVX1 mul_U22328(.A(dpath_mulcore_ary1_a1_c_2[31]), .Y(n9077));
INVX1 mul_U22329(.A(dpath_mulcore_ary1_a1_c_2[30]), .Y(n9078));
INVX1 mul_U22330(.A(dpath_mulcore_ary1_a1_c_2[29]), .Y(n9079));
INVX1 mul_U22331(.A(dpath_mulcore_ary1_a1_c_2[28]), .Y(n9080));
INVX1 mul_U22332(.A(dpath_mulcore_ary1_a1_c_2[27]), .Y(n9081));
INVX1 mul_U22333(.A(dpath_mulcore_ary1_a1_c_2[26]), .Y(n9082));
INVX1 mul_U22334(.A(dpath_mulcore_ary1_a1_c_2[25]), .Y(n9083));
INVX1 mul_U22335(.A(dpath_mulcore_ary1_a1_c_2[24]), .Y(n9084));
INVX1 mul_U22336(.A(dpath_mulcore_ary1_a1_c_2[23]), .Y(n9085));
INVX1 mul_U22337(.A(dpath_mulcore_ary1_a1_c_2[22]), .Y(n9086));
INVX1 mul_U22338(.A(dpath_mulcore_ary1_a1_c_2[21]), .Y(n9087));
INVX1 mul_U22339(.A(dpath_mulcore_ary1_a1_c_2[20]), .Y(n9088));
INVX1 mul_U22340(.A(dpath_mulcore_ary1_a1_c_2[19]), .Y(n9089));
INVX1 mul_U22341(.A(dpath_mulcore_ary1_a1_c_2[18]), .Y(n9090));
INVX1 mul_U22342(.A(dpath_mulcore_ary1_a1_c_2[17]), .Y(n9091));
INVX1 mul_U22343(.A(dpath_mulcore_ary1_a1_c_2[16]), .Y(n9092));
INVX1 mul_U22344(.A(dpath_mulcore_ary1_a1_c_2[15]), .Y(n9093));
INVX1 mul_U22345(.A(dpath_mulcore_ary1_a1_c_2[14]), .Y(n9094));
INVX1 mul_U22346(.A(dpath_mulcore_ary1_a1_c_2[13]), .Y(n9095));
INVX1 mul_U22347(.A(dpath_mulcore_ary1_a1_c_2[12]), .Y(n9096));
INVX1 mul_U22348(.A(dpath_mulcore_ary1_a1_c_2[11]), .Y(n9097));
INVX1 mul_U22349(.A(dpath_mulcore_ary1_a1_c_2[10]), .Y(n9098));
INVX1 mul_U22350(.A(dpath_mulcore_array2_c1[19]), .Y(n9099));
INVX1 mul_U22351(.A(dpath_mulcore_array2_c2[66]), .Y(n9100));
INVX1 mul_U22352(.A(dpath_mulcore_array2_c1[65]), .Y(n9101));
INVX1 mul_U22353(.A(dpath_mulcore_array2_c1[64]), .Y(n9102));
INVX1 mul_U22354(.A(dpath_mulcore_array2_c1[63]), .Y(n9103));
INVX1 mul_U22355(.A(dpath_mulcore_array2_c1[62]), .Y(n9104));
INVX1 mul_U22356(.A(dpath_mulcore_array2_c1[61]), .Y(n9105));
INVX1 mul_U22357(.A(dpath_mulcore_array2_c1[60]), .Y(n9106));
INVX1 mul_U22358(.A(dpath_mulcore_array2_c1[59]), .Y(n9107));
INVX1 mul_U22359(.A(dpath_mulcore_array2_c1[58]), .Y(n9108));
INVX1 mul_U22360(.A(dpath_mulcore_array2_c1[57]), .Y(n9109));
INVX1 mul_U22361(.A(dpath_mulcore_array2_c1[56]), .Y(n9110));
INVX1 mul_U22362(.A(dpath_mulcore_array2_c1[55]), .Y(n9111));
INVX1 mul_U22363(.A(dpath_mulcore_array2_c1[54]), .Y(n9112));
INVX1 mul_U22364(.A(dpath_mulcore_array2_c1[53]), .Y(n9113));
INVX1 mul_U22365(.A(dpath_mulcore_array2_c1[52]), .Y(n9114));
INVX1 mul_U22366(.A(dpath_mulcore_array2_c1[51]), .Y(n9115));
INVX1 mul_U22367(.A(dpath_mulcore_array2_c1[50]), .Y(n9116));
INVX1 mul_U22368(.A(dpath_mulcore_array2_c1[49]), .Y(n9117));
INVX1 mul_U22369(.A(dpath_mulcore_array2_c1[48]), .Y(n9118));
INVX1 mul_U22370(.A(dpath_mulcore_array2_c1[47]), .Y(n9119));
INVX1 mul_U22371(.A(dpath_mulcore_array2_c1[46]), .Y(n9120));
INVX1 mul_U22372(.A(dpath_mulcore_array2_c1[45]), .Y(n9121));
INVX1 mul_U22373(.A(dpath_mulcore_array2_c1[44]), .Y(n9122));
INVX1 mul_U22374(.A(dpath_mulcore_array2_c1[43]), .Y(n9123));
INVX1 mul_U22375(.A(dpath_mulcore_array2_c1[42]), .Y(n9124));
INVX1 mul_U22376(.A(dpath_mulcore_array2_c1[41]), .Y(n9125));
INVX1 mul_U22377(.A(dpath_mulcore_array2_c1[40]), .Y(n9126));
INVX1 mul_U22378(.A(dpath_mulcore_array2_c1[39]), .Y(n9127));
INVX1 mul_U22379(.A(dpath_mulcore_array2_c1[38]), .Y(n9128));
INVX1 mul_U22380(.A(dpath_mulcore_array2_c1[37]), .Y(n9129));
INVX1 mul_U22381(.A(dpath_mulcore_array2_c1[36]), .Y(n9130));
INVX1 mul_U22382(.A(dpath_mulcore_array2_c1[35]), .Y(n9131));
INVX1 mul_U22383(.A(dpath_mulcore_array2_c1[34]), .Y(n9132));
INVX1 mul_U22384(.A(dpath_mulcore_array2_c1[33]), .Y(n9133));
INVX1 mul_U22385(.A(dpath_mulcore_array2_c1[32]), .Y(n9134));
INVX1 mul_U22386(.A(dpath_mulcore_array2_c1[31]), .Y(n9135));
INVX1 mul_U22387(.A(dpath_mulcore_array2_c1[30]), .Y(n9136));
INVX1 mul_U22388(.A(dpath_mulcore_array2_c1[29]), .Y(n9137));
INVX1 mul_U22389(.A(dpath_mulcore_array2_c1[28]), .Y(n9138));
INVX1 mul_U22390(.A(dpath_mulcore_array2_c1[27]), .Y(n9139));
INVX1 mul_U22391(.A(dpath_mulcore_array2_c1[26]), .Y(n9140));
INVX1 mul_U22392(.A(dpath_mulcore_array2_c1[25]), .Y(n9141));
INVX1 mul_U22393(.A(dpath_mulcore_array2_c1[24]), .Y(n9142));
INVX1 mul_U22394(.A(dpath_mulcore_array2_c1[23]), .Y(n9143));
INVX1 mul_U22395(.A(dpath_mulcore_array2_c1[22]), .Y(n9144));
INVX1 mul_U22396(.A(dpath_mulcore_array2_c1[21]), .Y(n9145));
INVX1 mul_U22397(.A(dpath_mulcore_array2_c1[20]), .Y(n9146));
INVX1 mul_U22398(.A(dpath_mulcore_ary1_a0_c_2[70]), .Y(n9147));
INVX1 mul_U22399(.A(dpath_mulcore_pcout[82]), .Y(n9148));
INVX1 mul_U22400(.A(dpath_mulcore_pcout[68]), .Y(n9149));
INVX1 mul_U22401(.A(dpath_mulcore_pcout[67]), .Y(n9150));
INVX1 mul_U22402(.A(dpath_mulcore_pcout[66]), .Y(n9151));
INVX1 mul_U22403(.A(dpath_mulcore_pcout[65]), .Y(n9152));
INVX1 mul_U22404(.A(dpath_mulcore_pcout[64]), .Y(n9153));
INVX1 mul_U22405(.A(dpath_mulcore_pcout[63]), .Y(n9154));
INVX1 mul_U22406(.A(dpath_mulcore_pcout[62]), .Y(n9155));
INVX1 mul_U22407(.A(dpath_mulcore_pcout[61]), .Y(n9156));
INVX1 mul_U22408(.A(dpath_mulcore_pcout[60]), .Y(n9157));
INVX1 mul_U22409(.A(dpath_mulcore_pcout[59]), .Y(n9158));
INVX1 mul_U22410(.A(dpath_mulcore_pcout[58]), .Y(n9159));
INVX1 mul_U22411(.A(dpath_mulcore_pcout[57]), .Y(n9160));
INVX1 mul_U22412(.A(dpath_mulcore_pcout[56]), .Y(n9161));
INVX1 mul_U22413(.A(dpath_mulcore_pcout[55]), .Y(n9162));
INVX1 mul_U22414(.A(dpath_mulcore_pcout[54]), .Y(n9163));
INVX1 mul_U22415(.A(dpath_mulcore_pcout[53]), .Y(n9164));
INVX1 mul_U22416(.A(dpath_mulcore_pcout[52]), .Y(n9165));
INVX1 mul_U22417(.A(dpath_mulcore_pcout[51]), .Y(n9166));
INVX1 mul_U22418(.A(dpath_mulcore_pcout[50]), .Y(n9167));
INVX1 mul_U22419(.A(dpath_mulcore_pcout[49]), .Y(n9168));
INVX1 mul_U22420(.A(dpath_mulcore_pcout[48]), .Y(n9169));
INVX1 mul_U22421(.A(dpath_mulcore_pcout[47]), .Y(n9170));
INVX1 mul_U22422(.A(dpath_mulcore_pcout[46]), .Y(n9171));
INVX1 mul_U22423(.A(dpath_mulcore_pcout[45]), .Y(n9172));
INVX1 mul_U22424(.A(dpath_mulcore_pcout[44]), .Y(n9173));
INVX1 mul_U22425(.A(dpath_mulcore_pcout[43]), .Y(n9174));
INVX1 mul_U22426(.A(dpath_mulcore_pcout[42]), .Y(n9175));
INVX1 mul_U22427(.A(dpath_mulcore_pcout[41]), .Y(n9176));
INVX1 mul_U22428(.A(dpath_mulcore_pcout[40]), .Y(n9177));
INVX1 mul_U22429(.A(dpath_mulcore_pcout[39]), .Y(n9178));
INVX1 mul_U22430(.A(dpath_mulcore_pcout[38]), .Y(n9179));
INVX1 mul_U22431(.A(dpath_mulcore_pcout[37]), .Y(n9180));
INVX1 mul_U22432(.A(dpath_mulcore_pcout[36]), .Y(n9181));
INVX1 mul_U22433(.A(dpath_mulcore_pcout[35]), .Y(n9182));
INVX1 mul_U22434(.A(dpath_mulcore_pcout[34]), .Y(n9183));
INVX1 mul_U22435(.A(dpath_mulcore_pcout[33]), .Y(n9184));
INVX1 mul_U22436(.A(dpath_mulcore_pcout[32]), .Y(n9185));
INVX1 mul_U22437(.A(dpath_mulcore_pcout[31]), .Y(n9186));
INVX1 mul_U22438(.A(dpath_mulcore_pcout[30]), .Y(n9187));
INVX1 mul_U22439(.A(dpath_mulcore_pcout[95]), .Y(n9188));
INVX1 mul_U22440(.A(dpath_mulcore_pcout[94]), .Y(n9189));
INVX1 mul_U22441(.A(dpath_mulcore_pcout[93]), .Y(n9190));
INVX1 mul_U22442(.A(dpath_mulcore_pcout[92]), .Y(n9191));
INVX1 mul_U22443(.A(dpath_mulcore_pcout[91]), .Y(n9192));
INVX1 mul_U22444(.A(dpath_mulcore_pcout[90]), .Y(n9193));
INVX1 mul_U22445(.A(dpath_mulcore_pcout[89]), .Y(n9194));
INVX1 mul_U22446(.A(dpath_mulcore_pcout[88]), .Y(n9195));
INVX1 mul_U22447(.A(dpath_mulcore_pcout[87]), .Y(n9196));
INVX1 mul_U22448(.A(dpath_mulcore_pcout[86]), .Y(n9197));
INVX1 mul_U22449(.A(dpath_mulcore_pcout[85]), .Y(n9198));
INVX1 mul_U22450(.A(dpath_mulcore_pcout[84]), .Y(n9199));
INVX1 mul_U22451(.A(dpath_mulcore_pcout[81]), .Y(n9200));
INVX1 mul_U22452(.A(dpath_mulcore_pcout[80]), .Y(n9201));
INVX1 mul_U22453(.A(dpath_mulcore_pcout[79]), .Y(n9202));
INVX1 mul_U22454(.A(dpath_mulcore_pcout[78]), .Y(n9203));
INVX1 mul_U22455(.A(dpath_mulcore_pcout[77]), .Y(n9204));
INVX1 mul_U22456(.A(dpath_mulcore_pcout[76]), .Y(n9205));
INVX1 mul_U22457(.A(dpath_mulcore_pcout[75]), .Y(n9206));
INVX1 mul_U22458(.A(dpath_mulcore_pcout[74]), .Y(n9207));
INVX1 mul_U22459(.A(dpath_mulcore_pcout[73]), .Y(n9208));
INVX1 mul_U22460(.A(dpath_mulcore_pcout[72]), .Y(n9209));
INVX1 mul_U22461(.A(dpath_mulcore_pcout[71]), .Y(n9210));
INVX1 mul_U22462(.A(dpath_mulcore_pcout[70]), .Y(n9211));
INVX1 mul_U22463(.A(dpath_mulcore_pcout[69]), .Y(n9212));
INVX1 mul_U22464(.A(dpath_mulcore_pcout[83]), .Y(n9213));
INVX1 mul_U22465(.A(acc_imm), .Y(n9214));
INVX1 mul_U22466(.A(dpath_n522), .Y(n9215));
INVX1 mul_U22467(.A(dpath_mulcore_add_co31), .Y(n9216));
AND2X1 mul_U22468(.A(dpath_mulcore_b0[2]), .B(dpath_mulcore_b0[1]), .Y(dpath_mulcore_ary1_a0_I0_I2_net088));
INVX1 mul_U22469(.A(dpath_mulcore_ary1_a0_I0_I2_net088), .Y(n9217));
INVX1 mul_U22470(.A(n10236), .Y(n9218));
INVX1 mul_U22471(.A(n10252), .Y(n9219));
INVX1 mul_U22472(.A(n10254), .Y(n9220));
INVX1 mul_U22473(.A(n10256), .Y(n9221));
INVX1 mul_U22474(.A(n10258), .Y(n9222));
INVX1 mul_U22475(.A(n10260), .Y(n9223));
INVX1 mul_U22476(.A(n10262), .Y(n9224));
INVX1 mul_U22477(.A(n10264), .Y(n9225));
INVX1 mul_U22478(.A(n10343), .Y(n9226));
INVX1 mul_U22479(.A(n10395), .Y(n9227));
INVX1 mul_U22480(.A(n10447), .Y(n9228));
INVX1 mul_U22481(.A(n10499), .Y(n9229));
INVX1 mul_U22482(.A(n10551), .Y(n9230));
INVX1 mul_U22483(.A(n10584), .Y(n9231));
INVX1 mul_U22484(.A(n10586), .Y(n9232));
INVX1 mul_U22485(.A(n10588), .Y(n9233));
INVX1 mul_U22486(.A(n10590), .Y(n9234));
INVX1 mul_U22487(.A(n10138), .Y(n9235));
INVX1 mul_U22488(.A(n10143), .Y(n9236));
INVX1 mul_U22489(.A(n10148), .Y(n9237));
INVX1 mul_U22490(.A(n10153), .Y(n9238));
INVX1 mul_U22491(.A(n10158), .Y(n9239));
INVX1 mul_U22492(.A(n10163), .Y(n9240));
INVX1 mul_U22493(.A(n10168), .Y(n9241));
INVX1 mul_U22494(.A(n10173), .Y(n9242));
INVX1 mul_U22495(.A(n10178), .Y(n9243));
INVX1 mul_U22496(.A(n10185), .Y(n9244));
INVX1 mul_U22497(.A(n10190), .Y(n9245));
INVX1 mul_U22498(.A(n10195), .Y(n9246));
INVX1 mul_U22499(.A(n10200), .Y(n9247));
INVX1 mul_U22500(.A(n10205), .Y(n9248));
INVX1 mul_U22501(.A(n10210), .Y(n9249));
INVX1 mul_U22502(.A(n10215), .Y(n9250));
INVX1 mul_U22503(.A(n10220), .Y(n9251));
INVX1 mul_U22504(.A(n10225), .Y(n9252));
INVX1 mul_U22505(.A(n10230), .Y(n9253));
INVX1 mul_U22506(.A(n10237), .Y(n9254));
INVX1 mul_U22507(.A(n10242), .Y(n9255));
INVX1 mul_U22508(.A(n10247), .Y(n9256));
INVX1 mul_U22509(.A(n10297), .Y(n9257));
INVX1 mul_U22510(.A(n10302), .Y(n9258));
INVX1 mul_U22511(.A(n10307), .Y(n9259));
INVX1 mul_U22512(.A(n10312), .Y(n9260));
INVX1 mul_U22513(.A(n10317), .Y(n9261));
INVX1 mul_U22514(.A(n10322), .Y(n9262));
INVX1 mul_U22515(.A(n10327), .Y(n9263));
INVX1 mul_U22516(.A(n10332), .Y(n9264));
INVX1 mul_U22517(.A(n10337), .Y(n9265));
INVX1 mul_U22518(.A(n10344), .Y(n9266));
INVX1 mul_U22519(.A(n10349), .Y(n9267));
INVX1 mul_U22520(.A(n10354), .Y(n9268));
INVX1 mul_U22521(.A(n10359), .Y(n9269));
INVX1 mul_U22522(.A(n10364), .Y(n9270));
INVX1 mul_U22523(.A(n10369), .Y(n9271));
INVX1 mul_U22524(.A(n10374), .Y(n9272));
INVX1 mul_U22525(.A(n10379), .Y(n9273));
INVX1 mul_U22526(.A(n10384), .Y(n9274));
INVX1 mul_U22527(.A(n10389), .Y(n9275));
INVX1 mul_U22528(.A(n10396), .Y(n9276));
INVX1 mul_U22529(.A(n10401), .Y(n9277));
INVX1 mul_U22530(.A(n10406), .Y(n9278));
INVX1 mul_U22531(.A(n10411), .Y(n9279));
INVX1 mul_U22532(.A(n10416), .Y(n9280));
INVX1 mul_U22533(.A(n10421), .Y(n9281));
INVX1 mul_U22534(.A(n10426), .Y(n9282));
INVX1 mul_U22535(.A(n10431), .Y(n9283));
INVX1 mul_U22536(.A(n10436), .Y(n9284));
INVX1 mul_U22537(.A(n10441), .Y(n9285));
INVX1 mul_U22538(.A(n10448), .Y(n9286));
INVX1 mul_U22539(.A(n10453), .Y(n9287));
INVX1 mul_U22540(.A(n10458), .Y(n9288));
INVX1 mul_U22541(.A(n10463), .Y(n9289));
INVX1 mul_U22542(.A(n10468), .Y(n9290));
INVX1 mul_U22543(.A(n10473), .Y(n9291));
INVX1 mul_U22544(.A(n10478), .Y(n9292));
INVX1 mul_U22545(.A(n10483), .Y(n9293));
INVX1 mul_U22546(.A(n10488), .Y(n9294));
INVX1 mul_U22547(.A(n10493), .Y(n9295));
INVX1 mul_U22548(.A(n10500), .Y(n9296));
INVX1 mul_U22549(.A(n10505), .Y(n9297));
INVX1 mul_U22550(.A(n10510), .Y(n9298));
INVX1 mul_U22551(.A(n10515), .Y(n9299));
INVX1 mul_U22552(.A(n10520), .Y(n9300));
INVX1 mul_U22553(.A(n10525), .Y(n9301));
INVX1 mul_U22554(.A(n10530), .Y(n9302));
INVX1 mul_U22555(.A(n10535), .Y(n9303));
INVX1 mul_U22556(.A(n10540), .Y(n9304));
INVX1 mul_U22557(.A(n10545), .Y(n9305));
INVX1 mul_U22558(.A(n10552), .Y(n9306));
INVX1 mul_U22559(.A(n10557), .Y(n9307));
INVX1 mul_U22560(.A(n10562), .Y(n9308));
INVX1 mul_U22561(.A(n10567), .Y(n9309));
INVX1 mul_U22562(.A(n10572), .Y(n9310));
INVX1 mul_U22563(.A(n10577), .Y(n9311));
AND2X1 mul_U22564(.A(dpath_mulcore_b7[2]), .B(dpath_mulcore_b7[1]), .Y(dpath_mulcore_ary1_a0_I2_I2_net0118));
INVX1 mul_U22565(.A(dpath_mulcore_ary1_a0_I2_I2_net0118), .Y(n9312));
INVX1 mul_U22566(.A(dpath_mulcore_ary1_a0_c_1[69]), .Y(n9313));
INVX1 mul_U22567(.A(dpath_mulcore_ary1_a0_c_1[68]), .Y(n9314));
INVX1 mul_U22568(.A(dpath_mulcore_ary1_a0_c_1[67]), .Y(n9315));
INVX1 mul_U22569(.A(dpath_mulcore_ary1_a0_c_1[66]), .Y(n9316));
INVX1 mul_U22570(.A(dpath_mulcore_ary1_a0_c_1[65]), .Y(n9317));
INVX1 mul_U22571(.A(dpath_mulcore_ary1_a0_c_1[64]), .Y(n9318));
INVX1 mul_U22572(.A(dpath_mulcore_ary1_a0_c_1[63]), .Y(n9319));
INVX1 mul_U22573(.A(dpath_mulcore_ary1_a0_c_1[62]), .Y(n9320));
INVX1 mul_U22574(.A(dpath_mulcore_ary1_a0_c_1[61]), .Y(n9321));
INVX1 mul_U22575(.A(dpath_mulcore_ary1_a0_c_1[60]), .Y(n9322));
INVX1 mul_U22576(.A(dpath_mulcore_ary1_a0_c_1[59]), .Y(n9323));
INVX1 mul_U22577(.A(dpath_mulcore_ary1_a0_c_1[58]), .Y(n9324));
INVX1 mul_U22578(.A(dpath_mulcore_ary1_a0_c_1[57]), .Y(n9325));
INVX1 mul_U22579(.A(dpath_mulcore_ary1_a0_c_1[56]), .Y(n9326));
INVX1 mul_U22580(.A(dpath_mulcore_ary1_a0_c_1[55]), .Y(n9327));
INVX1 mul_U22581(.A(dpath_mulcore_ary1_a0_c_1[54]), .Y(n9328));
INVX1 mul_U22582(.A(dpath_mulcore_ary1_a0_c_1[53]), .Y(n9329));
INVX1 mul_U22583(.A(dpath_mulcore_ary1_a0_c_1[52]), .Y(n9330));
INVX1 mul_U22584(.A(dpath_mulcore_ary1_a0_c_1[51]), .Y(n9331));
INVX1 mul_U22585(.A(dpath_mulcore_ary1_a0_c_1[50]), .Y(n9332));
INVX1 mul_U22586(.A(dpath_mulcore_ary1_a0_c_1[49]), .Y(n9333));
INVX1 mul_U22587(.A(dpath_mulcore_ary1_a0_c_1[48]), .Y(n9334));
INVX1 mul_U22588(.A(dpath_mulcore_ary1_a0_c_1[47]), .Y(n9335));
INVX1 mul_U22589(.A(dpath_mulcore_ary1_a0_c_1[46]), .Y(n9336));
INVX1 mul_U22590(.A(dpath_mulcore_ary1_a0_c_1[45]), .Y(n9337));
INVX1 mul_U22591(.A(dpath_mulcore_ary1_a0_c_1[44]), .Y(n9338));
INVX1 mul_U22592(.A(dpath_mulcore_ary1_a0_c_1[43]), .Y(n9339));
INVX1 mul_U22593(.A(dpath_mulcore_ary1_a0_c_1[42]), .Y(n9340));
INVX1 mul_U22594(.A(dpath_mulcore_ary1_a0_c_1[41]), .Y(n9341));
INVX1 mul_U22595(.A(dpath_mulcore_ary1_a0_c_1[40]), .Y(n9342));
INVX1 mul_U22596(.A(dpath_mulcore_ary1_a0_c_1[39]), .Y(n9343));
INVX1 mul_U22597(.A(dpath_mulcore_ary1_a0_c_1[38]), .Y(n9344));
INVX1 mul_U22598(.A(dpath_mulcore_ary1_a0_c_1[37]), .Y(n9345));
INVX1 mul_U22599(.A(dpath_mulcore_ary1_a0_c_1[36]), .Y(n9346));
INVX1 mul_U22600(.A(dpath_mulcore_ary1_a0_c_1[35]), .Y(n9347));
INVX1 mul_U22601(.A(dpath_mulcore_ary1_a0_c_1[34]), .Y(n9348));
INVX1 mul_U22602(.A(dpath_mulcore_ary1_a0_c_1[33]), .Y(n9349));
INVX1 mul_U22603(.A(dpath_mulcore_ary1_a0_c_1[32]), .Y(n9350));
INVX1 mul_U22604(.A(dpath_mulcore_ary1_a0_c_1[31]), .Y(n9351));
INVX1 mul_U22605(.A(dpath_mulcore_ary1_a0_c_1[30]), .Y(n9352));
INVX1 mul_U22606(.A(dpath_mulcore_ary1_a0_c_1[29]), .Y(n9353));
INVX1 mul_U22607(.A(dpath_mulcore_ary1_a0_c_1[28]), .Y(n9354));
INVX1 mul_U22608(.A(dpath_mulcore_ary1_a0_c_1[27]), .Y(n9355));
INVX1 mul_U22609(.A(dpath_mulcore_ary1_a0_c_1[26]), .Y(n9356));
INVX1 mul_U22610(.A(dpath_mulcore_ary1_a0_c_1[25]), .Y(n9357));
INVX1 mul_U22611(.A(dpath_mulcore_ary1_a0_c_1[24]), .Y(n9358));
INVX1 mul_U22612(.A(dpath_mulcore_ary1_a0_c_1[23]), .Y(n9359));
INVX1 mul_U22613(.A(dpath_mulcore_ary1_a0_c_1[22]), .Y(n9360));
INVX1 mul_U22614(.A(dpath_mulcore_ary1_a0_c_1[21]), .Y(n9361));
INVX1 mul_U22615(.A(dpath_mulcore_ary1_a0_c_1[20]), .Y(n9362));
INVX1 mul_U22616(.A(dpath_mulcore_ary1_a0_c_1[19]), .Y(n9363));
INVX1 mul_U22617(.A(dpath_mulcore_ary1_a0_c_1[18]), .Y(n9364));
INVX1 mul_U22618(.A(dpath_mulcore_ary1_a0_c_1[17]), .Y(n9365));
INVX1 mul_U22619(.A(dpath_mulcore_ary1_a0_c_1[16]), .Y(n9366));
INVX1 mul_U22620(.A(dpath_mulcore_ary1_a0_c_1[15]), .Y(n9367));
INVX1 mul_U22621(.A(dpath_mulcore_ary1_a0_c_1[14]), .Y(n9368));
INVX1 mul_U22622(.A(dpath_mulcore_ary1_a1_c_1[69]), .Y(n9369));
INVX1 mul_U22623(.A(dpath_mulcore_ary1_a1_c_1[68]), .Y(n9370));
INVX1 mul_U22624(.A(dpath_mulcore_ary1_a1_c_1[67]), .Y(n9371));
INVX1 mul_U22625(.A(dpath_mulcore_ary1_a1_c_1[66]), .Y(n9372));
INVX1 mul_U22626(.A(dpath_mulcore_ary1_a1_c_1[65]), .Y(n9373));
INVX1 mul_U22627(.A(dpath_mulcore_ary1_a1_c_1[64]), .Y(n9374));
INVX1 mul_U22628(.A(dpath_mulcore_ary1_a1_c_1[63]), .Y(n9375));
INVX1 mul_U22629(.A(dpath_mulcore_ary1_a1_c_1[62]), .Y(n9376));
INVX1 mul_U22630(.A(dpath_mulcore_ary1_a1_c_1[61]), .Y(n9377));
INVX1 mul_U22631(.A(dpath_mulcore_ary1_a1_c_1[60]), .Y(n9378));
INVX1 mul_U22632(.A(dpath_mulcore_ary1_a1_c_1[59]), .Y(n9379));
INVX1 mul_U22633(.A(dpath_mulcore_ary1_a1_c_1[58]), .Y(n9380));
INVX1 mul_U22634(.A(dpath_mulcore_ary1_a1_c_1[57]), .Y(n9381));
INVX1 mul_U22635(.A(dpath_mulcore_ary1_a1_c_1[56]), .Y(n9382));
INVX1 mul_U22636(.A(dpath_mulcore_ary1_a1_c_1[55]), .Y(n9383));
INVX1 mul_U22637(.A(dpath_mulcore_ary1_a1_c_1[54]), .Y(n9384));
INVX1 mul_U22638(.A(dpath_mulcore_ary1_a1_c_1[53]), .Y(n9385));
INVX1 mul_U22639(.A(dpath_mulcore_ary1_a1_c_1[52]), .Y(n9386));
INVX1 mul_U22640(.A(dpath_mulcore_ary1_a1_c_1[51]), .Y(n9387));
INVX1 mul_U22641(.A(dpath_mulcore_ary1_a1_c_1[50]), .Y(n9388));
INVX1 mul_U22642(.A(dpath_mulcore_ary1_a1_c_1[49]), .Y(n9389));
INVX1 mul_U22643(.A(dpath_mulcore_ary1_a1_c_1[48]), .Y(n9390));
INVX1 mul_U22644(.A(dpath_mulcore_ary1_a1_c_1[47]), .Y(n9391));
INVX1 mul_U22645(.A(dpath_mulcore_ary1_a1_c_1[46]), .Y(n9392));
INVX1 mul_U22646(.A(dpath_mulcore_ary1_a1_c_1[45]), .Y(n9393));
INVX1 mul_U22647(.A(dpath_mulcore_ary1_a1_c_1[44]), .Y(n9394));
INVX1 mul_U22648(.A(dpath_mulcore_ary1_a1_c_1[43]), .Y(n9395));
INVX1 mul_U22649(.A(dpath_mulcore_ary1_a1_c_1[42]), .Y(n9396));
INVX1 mul_U22650(.A(dpath_mulcore_ary1_a1_c_1[41]), .Y(n9397));
INVX1 mul_U22651(.A(dpath_mulcore_ary1_a1_c_1[40]), .Y(n9398));
INVX1 mul_U22652(.A(dpath_mulcore_ary1_a1_c_1[39]), .Y(n9399));
INVX1 mul_U22653(.A(dpath_mulcore_ary1_a1_c_1[38]), .Y(n9400));
INVX1 mul_U22654(.A(dpath_mulcore_ary1_a1_c_1[37]), .Y(n9401));
INVX1 mul_U22655(.A(dpath_mulcore_ary1_a1_c_1[36]), .Y(n9402));
INVX1 mul_U22656(.A(dpath_mulcore_ary1_a1_c_1[35]), .Y(n9403));
INVX1 mul_U22657(.A(dpath_mulcore_ary1_a1_c_1[34]), .Y(n9404));
INVX1 mul_U22658(.A(dpath_mulcore_ary1_a1_c_1[33]), .Y(n9405));
INVX1 mul_U22659(.A(dpath_mulcore_ary1_a1_c_1[32]), .Y(n9406));
INVX1 mul_U22660(.A(dpath_mulcore_ary1_a1_c_1[31]), .Y(n9407));
INVX1 mul_U22661(.A(dpath_mulcore_ary1_a1_c_1[30]), .Y(n9408));
INVX1 mul_U22662(.A(dpath_mulcore_ary1_a1_c_1[29]), .Y(n9409));
INVX1 mul_U22663(.A(dpath_mulcore_ary1_a1_c_1[28]), .Y(n9410));
INVX1 mul_U22664(.A(dpath_mulcore_ary1_a1_c_1[27]), .Y(n9411));
INVX1 mul_U22665(.A(dpath_mulcore_ary1_a1_c_1[26]), .Y(n9412));
INVX1 mul_U22666(.A(dpath_mulcore_ary1_a1_c_1[25]), .Y(n9413));
INVX1 mul_U22667(.A(dpath_mulcore_ary1_a1_c_1[24]), .Y(n9414));
INVX1 mul_U22668(.A(dpath_mulcore_ary1_a1_c_1[23]), .Y(n9415));
INVX1 mul_U22669(.A(dpath_mulcore_ary1_a1_c_1[22]), .Y(n9416));
INVX1 mul_U22670(.A(dpath_mulcore_ary1_a1_c_1[21]), .Y(n9417));
INVX1 mul_U22671(.A(dpath_mulcore_ary1_a1_c_1[20]), .Y(n9418));
INVX1 mul_U22672(.A(dpath_mulcore_ary1_a1_c_1[19]), .Y(n9419));
INVX1 mul_U22673(.A(dpath_mulcore_ary1_a1_c_1[18]), .Y(n9420));
INVX1 mul_U22674(.A(dpath_mulcore_ary1_a1_c_1[17]), .Y(n9421));
INVX1 mul_U22675(.A(dpath_mulcore_ary1_a1_c_1[16]), .Y(n9422));
INVX1 mul_U22676(.A(dpath_mulcore_ary1_a1_c_1[15]), .Y(n9423));
INVX1 mul_U22677(.A(dpath_mulcore_ary1_a1_c_1[14]), .Y(n9424));
AND2X1 mul_U22678(.A(dpath_mulcore_b2[2]), .B(dpath_mulcore_b2[1]), .Y(dpath_mulcore_ary1_a0_I0_I2_net075));
INVX1 mul_U22679(.A(dpath_mulcore_ary1_a0_I0_I2_net075), .Y(n9425));
AND2X1 mul_U22680(.A(dpath_mulcore_b1[2]), .B(dpath_mulcore_b1[1]), .Y(dpath_mulcore_ary1_a0_I0_I2_net0118));
INVX1 mul_U22681(.A(dpath_mulcore_ary1_a0_I0_I2_net0118), .Y(n9426));
AND2X1 mul_U22682(.A(dpath_mulcore_b10[2]), .B(dpath_mulcore_b10[1]), .Y(dpath_mulcore_ary1_a1_I0_I2_net075));
INVX1 mul_U22683(.A(dpath_mulcore_ary1_a1_I0_I2_net075), .Y(n9427));
INVX1 mul_U22684(.A(dpath_mulcore_array2_c2[19]), .Y(n9428));
INVX1 mul_U22685(.A(dpath_mulcore_array2_c2[65]), .Y(n9429));
INVX1 mul_U22686(.A(dpath_mulcore_array2_c2[64]), .Y(n9430));
INVX1 mul_U22687(.A(dpath_mulcore_array2_c2[63]), .Y(n9431));
INVX1 mul_U22688(.A(dpath_mulcore_array2_c2[62]), .Y(n9432));
INVX1 mul_U22689(.A(dpath_mulcore_array2_c2[61]), .Y(n9433));
INVX1 mul_U22690(.A(dpath_mulcore_array2_c2[60]), .Y(n9434));
INVX1 mul_U22691(.A(dpath_mulcore_array2_c2[59]), .Y(n9435));
INVX1 mul_U22692(.A(dpath_mulcore_array2_c2[58]), .Y(n9436));
INVX1 mul_U22693(.A(dpath_mulcore_array2_c2[57]), .Y(n9437));
INVX1 mul_U22694(.A(dpath_mulcore_array2_c2[56]), .Y(n9438));
INVX1 mul_U22695(.A(dpath_mulcore_array2_c2[55]), .Y(n9439));
INVX1 mul_U22696(.A(dpath_mulcore_array2_c2[54]), .Y(n9440));
INVX1 mul_U22697(.A(dpath_mulcore_array2_c2[53]), .Y(n9441));
INVX1 mul_U22698(.A(dpath_mulcore_array2_c2[52]), .Y(n9442));
INVX1 mul_U22699(.A(dpath_mulcore_array2_c2[51]), .Y(n9443));
INVX1 mul_U22700(.A(dpath_mulcore_array2_c2[50]), .Y(n9444));
INVX1 mul_U22701(.A(dpath_mulcore_array2_c2[49]), .Y(n9445));
INVX1 mul_U22702(.A(dpath_mulcore_array2_c2[48]), .Y(n9446));
INVX1 mul_U22703(.A(dpath_mulcore_array2_c2[47]), .Y(n9447));
INVX1 mul_U22704(.A(dpath_mulcore_array2_c2[46]), .Y(n9448));
INVX1 mul_U22705(.A(dpath_mulcore_array2_c2[45]), .Y(n9449));
INVX1 mul_U22706(.A(dpath_mulcore_array2_c2[44]), .Y(n9450));
INVX1 mul_U22707(.A(dpath_mulcore_array2_c2[43]), .Y(n9451));
INVX1 mul_U22708(.A(dpath_mulcore_array2_c2[42]), .Y(n9452));
INVX1 mul_U22709(.A(dpath_mulcore_array2_c2[41]), .Y(n9453));
INVX1 mul_U22710(.A(dpath_mulcore_array2_c2[40]), .Y(n9454));
INVX1 mul_U22711(.A(dpath_mulcore_array2_c2[39]), .Y(n9455));
INVX1 mul_U22712(.A(dpath_mulcore_array2_c2[38]), .Y(n9456));
INVX1 mul_U22713(.A(dpath_mulcore_array2_c2[37]), .Y(n9457));
INVX1 mul_U22714(.A(dpath_mulcore_array2_c2[36]), .Y(n9458));
INVX1 mul_U22715(.A(dpath_mulcore_array2_c2[35]), .Y(n9459));
INVX1 mul_U22716(.A(dpath_mulcore_array2_c2[34]), .Y(n9460));
INVX1 mul_U22717(.A(dpath_mulcore_array2_c2[33]), .Y(n9461));
INVX1 mul_U22718(.A(dpath_mulcore_array2_c2[32]), .Y(n9462));
INVX1 mul_U22719(.A(dpath_mulcore_array2_c2[31]), .Y(n9463));
INVX1 mul_U22720(.A(dpath_mulcore_array2_c2[30]), .Y(n9464));
INVX1 mul_U22721(.A(dpath_mulcore_array2_c2[29]), .Y(n9465));
INVX1 mul_U22722(.A(dpath_mulcore_array2_c2[28]), .Y(n9466));
INVX1 mul_U22723(.A(dpath_mulcore_array2_c2[27]), .Y(n9467));
INVX1 mul_U22724(.A(dpath_mulcore_array2_c2[26]), .Y(n9468));
INVX1 mul_U22725(.A(dpath_mulcore_array2_c2[25]), .Y(n9469));
INVX1 mul_U22726(.A(dpath_mulcore_array2_c2[24]), .Y(n9470));
INVX1 mul_U22727(.A(dpath_mulcore_array2_c2[23]), .Y(n9471));
INVX1 mul_U22728(.A(dpath_mulcore_array2_c2[22]), .Y(n9472));
INVX1 mul_U22729(.A(dpath_mulcore_array2_c2[21]), .Y(n9473));
INVX1 mul_U22730(.A(dpath_mulcore_ary1_a0_I2_I2_net38), .Y(n9474));
AND2X1 mul_U22731(.A(dpath_mulcore_b3[2]), .B(dpath_mulcore_b3[1]), .Y(dpath_mulcore_ary1_a0_I1_I2_net088));
INVX1 mul_U22732(.A(dpath_mulcore_ary1_a0_I1_I2_net088), .Y(n9475));
AND2X1 mul_U22733(.A(dpath_mulcore_b4[2]), .B(dpath_mulcore_b4[1]), .Y(dpath_mulcore_ary1_a0_I1_I2_net0118));
INVX1 mul_U22734(.A(dpath_mulcore_ary1_a0_I1_I2_net0118), .Y(n9476));
AND2X1 mul_U22735(.A(dpath_mulcore_b14[2]), .B(dpath_mulcore_b14[1]), .Y(dpath_mulcore_ary1_a1_I2_I2_net088));
INVX1 mul_U22736(.A(dpath_mulcore_ary1_a1_I2_I2_net088), .Y(n9477));
AND2X1 mul_U22737(.A(dpath_mulcore_b15[2]), .B(dpath_mulcore_b15[1]), .Y(dpath_mulcore_ary1_a1_I2_I2_net0118));
INVX1 mul_U22738(.A(dpath_mulcore_ary1_a1_I2_I2_net0118), .Y(n9478));
AND2X1 mul_U22739(.A(dpath_mulcore_b11[2]), .B(dpath_mulcore_b11[1]), .Y(dpath_mulcore_ary1_a1_I1_I2_net088));
INVX1 mul_U22740(.A(dpath_mulcore_ary1_a1_I1_I2_net088), .Y(n9479));
AND2X1 mul_U22741(.A(dpath_mulcore_b12[2]), .B(dpath_mulcore_b12[1]), .Y(dpath_mulcore_ary1_a1_I1_I2_net0118));
INVX1 mul_U22742(.A(dpath_mulcore_ary1_a1_I1_I2_net0118), .Y(n9480));
AND2X1 mul_U22743(.A(dpath_mulcore_b8[2]), .B(dpath_mulcore_b8[1]), .Y(dpath_mulcore_ary1_a1_I0_I2_net088));
INVX1 mul_U22744(.A(dpath_mulcore_ary1_a1_I0_I2_net088), .Y(n9481));
AND2X1 mul_U22745(.A(dpath_mulcore_b9[2]), .B(dpath_mulcore_b9[1]), .Y(dpath_mulcore_ary1_a1_I0_I2_net0118));
INVX1 mul_U22746(.A(dpath_mulcore_ary1_a1_I0_I2_net0118), .Y(n9482));
AND2X1 mul_U22747(.A(dpath_mulcore_b6[2]), .B(dpath_mulcore_b6[1]), .Y(dpath_mulcore_ary1_a0_I2_I2_net088));
INVX1 mul_U22748(.A(dpath_mulcore_ary1_a0_I2_I2_net088), .Y(n9483));
AND2X1 mul_U22749(.A(dpath_mulcore_b5[2]), .B(dpath_mulcore_b5[1]), .Y(dpath_mulcore_ary1_a0_I1_I2_net075));
INVX1 mul_U22750(.A(dpath_mulcore_ary1_a0_I1_I2_net075), .Y(n9484));
AND2X1 mul_U22751(.A(dpath_mulcore_b13[2]), .B(dpath_mulcore_b13[1]), .Y(dpath_mulcore_ary1_a1_I1_I2_net075));
INVX1 mul_U22752(.A(dpath_mulcore_ary1_a1_I1_I2_net075), .Y(n9485));
INVX1 mul_U22753(.A(dpath_mulcore_ary1_a0_I1_I2_net073), .Y(n9486));
INVX1 mul_U22754(.A(dpath_mulcore_ary1_a1_I1_I2_net073), .Y(n9487));
INVX1 mul_U22755(.A(dpath_mulcore_ary1_a0_I0_I2_net073), .Y(n9488));
INVX1 mul_U22756(.A(dpath_mulcore_ary1_a1_I0_I2_net073), .Y(n9489));
INVX1 mul_U22757(.A(dpath_mulcore_ary1_a0_I0_I2_sc1_66__b), .Y(n9490));
BUFX2 mul_U22758(.A(rst_l), .Y(n9491));
XOR2X1 mul_U22759(.A(dpath_mulcore_addin_cin), .B(dpath_mulcore_addin_sum[0]), .Y(dpath_mulcore_addout[0]));
XOR2X1 mul_U22760(.A(dpath_mulcore_addin_cout[9]), .B(dpath_mulcore_addin_sum[10]), .Y(n10137));
XOR2X1 mul_U22761(.A(n9235), .B(n10137), .Y(dpath_mulcore_addout[10]));
XOR2X1 mul_U22762(.A(dpath_mulcore_addin_cout[10]), .B(dpath_mulcore_addin_sum[11]), .Y(n10142));
XOR2X1 mul_U22763(.A(n9236), .B(n10142), .Y(dpath_mulcore_addout[11]));
XOR2X1 mul_U22764(.A(dpath_mulcore_addin_cout[11]), .B(dpath_mulcore_addin_sum[12]), .Y(n10147));
XOR2X1 mul_U22765(.A(n9237), .B(n10147), .Y(dpath_mulcore_addout[12]));
XOR2X1 mul_U22766(.A(dpath_mulcore_addin_cout[12]), .B(dpath_mulcore_addin_sum[13]), .Y(n10152));
XOR2X1 mul_U22767(.A(n9238), .B(n10152), .Y(dpath_mulcore_addout[13]));
XOR2X1 mul_U22768(.A(dpath_mulcore_addin_cout[13]), .B(dpath_mulcore_addin_sum[14]), .Y(n10157));
XOR2X1 mul_U22769(.A(n9239), .B(n10157), .Y(dpath_mulcore_addout[14]));
XOR2X1 mul_U22770(.A(dpath_mulcore_addin_cout[14]), .B(dpath_mulcore_addin_sum[15]), .Y(n10162));
XOR2X1 mul_U22771(.A(n9240), .B(n10162), .Y(dpath_mulcore_addout[15]));
XOR2X1 mul_U22772(.A(dpath_mulcore_addin_cout[15]), .B(dpath_mulcore_addin_sum[16]), .Y(n10167));
XOR2X1 mul_U22773(.A(n9241), .B(n10167), .Y(dpath_mulcore_addout[16]));
XOR2X1 mul_U22774(.A(dpath_mulcore_addin_cout[16]), .B(dpath_mulcore_addin_sum[17]), .Y(n10172));
XOR2X1 mul_U22775(.A(n9242), .B(n10172), .Y(dpath_mulcore_addout[17]));
XOR2X1 mul_U22776(.A(dpath_mulcore_addin_cout[17]), .B(dpath_mulcore_addin_sum[18]), .Y(n10177));
XOR2X1 mul_U22777(.A(n9243), .B(n10177), .Y(dpath_mulcore_addout[18]));
XOR2X1 mul_U22778(.A(dpath_mulcore_addin_cout[18]), .B(dpath_mulcore_addin_sum[19]), .Y(n10182));
XOR2X1 mul_U22779(.A(n9244), .B(n10182), .Y(dpath_mulcore_addout[19]));
XOR2X1 mul_U22780(.A(dpath_mulcore_addin_cout[0]), .B(dpath_mulcore_addin_sum[1]), .Y(n10183));
XOR2X1 mul_U22781(.A(n10184), .B(n10183), .Y(dpath_mulcore_addout[1]));
XOR2X1 mul_U22782(.A(dpath_mulcore_addin_cout[19]), .B(dpath_mulcore_addin_sum[20]), .Y(n10189));
XOR2X1 mul_U22783(.A(n9245), .B(n10189), .Y(dpath_mulcore_addout[20]));
XOR2X1 mul_U22784(.A(dpath_mulcore_addin_cout[20]), .B(dpath_mulcore_addin_sum[21]), .Y(n10194));
XOR2X1 mul_U22785(.A(n9246), .B(n10194), .Y(dpath_mulcore_addout[21]));
XOR2X1 mul_U22786(.A(dpath_mulcore_addin_cout[21]), .B(dpath_mulcore_addin_sum[22]), .Y(n10199));
XOR2X1 mul_U22787(.A(n9247), .B(n10199), .Y(dpath_mulcore_addout[22]));
XOR2X1 mul_U22788(.A(dpath_mulcore_addin_cout[22]), .B(dpath_mulcore_addin_sum[23]), .Y(n10204));
XOR2X1 mul_U22789(.A(n9248), .B(n10204), .Y(dpath_mulcore_addout[23]));
XOR2X1 mul_U22790(.A(dpath_mulcore_addin_cout[23]), .B(dpath_mulcore_addin_sum[24]), .Y(n10209));
XOR2X1 mul_U22791(.A(n9249), .B(n10209), .Y(dpath_mulcore_addout[24]));
XOR2X1 mul_U22792(.A(dpath_mulcore_addin_cout[24]), .B(dpath_mulcore_addin_sum[25]), .Y(n10214));
XOR2X1 mul_U22793(.A(n9250), .B(n10214), .Y(dpath_mulcore_addout[25]));
XOR2X1 mul_U22794(.A(dpath_mulcore_addin_cout[25]), .B(dpath_mulcore_addin_sum[26]), .Y(n10219));
XOR2X1 mul_U22795(.A(n9251), .B(n10219), .Y(dpath_mulcore_addout[26]));
XOR2X1 mul_U22796(.A(dpath_mulcore_addin_cout[26]), .B(dpath_mulcore_addin_sum[27]), .Y(n10224));
XOR2X1 mul_U22797(.A(n9252), .B(n10224), .Y(dpath_mulcore_addout[27]));
XOR2X1 mul_U22798(.A(dpath_mulcore_addin_cout[27]), .B(dpath_mulcore_addin_sum[28]), .Y(n10229));
XOR2X1 mul_U22799(.A(n9253), .B(n10229), .Y(dpath_mulcore_addout[28]));
XOR2X1 mul_U22800(.A(dpath_mulcore_addin_cout[28]), .B(dpath_mulcore_addin_sum[29]), .Y(n10234));
XOR2X1 mul_U22801(.A(n9254), .B(n10234), .Y(dpath_mulcore_addout[29]));
XOR2X1 mul_U22802(.A(dpath_mulcore_addin_cout[1]), .B(dpath_mulcore_addin_sum[2]), .Y(n10235));
XOR2X1 mul_U22803(.A(n9218), .B(n10235), .Y(dpath_mulcore_addout[2]));
XOR2X1 mul_U22804(.A(dpath_mulcore_addin_cout[29]), .B(dpath_mulcore_addin_sum[30]), .Y(n10241));
XOR2X1 mul_U22805(.A(n9255), .B(n10241), .Y(dpath_mulcore_addout[30]));
XOR2X1 mul_U22806(.A(dpath_mulcore_addin_cout[30]), .B(dpath_mulcore_addin_sum[31]), .Y(n10246));
XOR2X1 mul_U22807(.A(n9256), .B(n10246), .Y(dpath_mulcore_addout[31]));
XOR2X1 mul_U22808(.A(dpath_mulcore_addin_cout[2]), .B(dpath_mulcore_addin_sum[3]), .Y(n10251));
XOR2X1 mul_U22809(.A(n9219), .B(n10251), .Y(dpath_mulcore_addout[3]));
XOR2X1 mul_U22810(.A(dpath_mulcore_addin_cout[3]), .B(dpath_mulcore_addin_sum[4]), .Y(n10253));
XOR2X1 mul_U22811(.A(n9220), .B(n10253), .Y(dpath_mulcore_addout[4]));
XOR2X1 mul_U22812(.A(dpath_mulcore_addin_cout[4]), .B(dpath_mulcore_addin_sum[5]), .Y(n10255));
XOR2X1 mul_U22813(.A(n9221), .B(n10255), .Y(dpath_mulcore_addout[5]));
XOR2X1 mul_U22814(.A(dpath_mulcore_addin_cout[5]), .B(dpath_mulcore_addin_sum[6]), .Y(n10257));
XOR2X1 mul_U22815(.A(n9222), .B(n10257), .Y(dpath_mulcore_addout[6]));
XOR2X1 mul_U22816(.A(dpath_mulcore_addin_cout[6]), .B(dpath_mulcore_addin_sum[7]), .Y(n10259));
XOR2X1 mul_U22817(.A(n9223), .B(n10259), .Y(dpath_mulcore_addout[7]));
XOR2X1 mul_U22818(.A(dpath_mulcore_addin_cout[7]), .B(dpath_mulcore_addin_sum[8]), .Y(n10261));
XOR2X1 mul_U22819(.A(n9224), .B(n10261), .Y(dpath_mulcore_addout[8]));
XOR2X1 mul_U22820(.A(dpath_mulcore_addin_cout[8]), .B(dpath_mulcore_addin_sum[9]), .Y(n10263));
XOR2X1 mul_U22821(.A(n9225), .B(n10263), .Y(dpath_mulcore_addout[9]));
XOR2X1 mul_U22822(.A(n9216), .B(dpath_mulcore_addin_cout[31]), .Y(n10265));
XOR2X1 mul_U22823(.A(dpath_mulcore_addin_sum[32]), .B(n10265), .Y(dpath_mulcore_addout[32]));
XOR2X1 mul_U22824(.A(dpath_mulcore_addin_cout[41]), .B(dpath_mulcore_addin_sum[42]), .Y(n10296));
XOR2X1 mul_U22825(.A(n9257), .B(n10296), .Y(dpath_mulcore_addout[42]));
XOR2X1 mul_U22826(.A(dpath_mulcore_addin_cout[42]), .B(dpath_mulcore_addin_sum[43]), .Y(n10301));
XOR2X1 mul_U22827(.A(n9258), .B(n10301), .Y(dpath_mulcore_addout[43]));
XOR2X1 mul_U22828(.A(dpath_mulcore_addin_cout[43]), .B(dpath_mulcore_addin_sum[44]), .Y(n10306));
XOR2X1 mul_U22829(.A(n9259), .B(n10306), .Y(dpath_mulcore_addout[44]));
XOR2X1 mul_U22830(.A(dpath_mulcore_addin_cout[44]), .B(dpath_mulcore_addin_sum[45]), .Y(n10311));
XOR2X1 mul_U22831(.A(n9260), .B(n10311), .Y(dpath_mulcore_addout[45]));
XOR2X1 mul_U22832(.A(dpath_mulcore_addin_cout[45]), .B(dpath_mulcore_addin_sum[46]), .Y(n10316));
XOR2X1 mul_U22833(.A(n9261), .B(n10316), .Y(dpath_mulcore_addout[46]));
XOR2X1 mul_U22834(.A(dpath_mulcore_addin_cout[46]), .B(dpath_mulcore_addin_sum[47]), .Y(n10321));
XOR2X1 mul_U22835(.A(n9262), .B(n10321), .Y(dpath_mulcore_addout[47]));
XOR2X1 mul_U22836(.A(dpath_mulcore_addin_cout[47]), .B(dpath_mulcore_addin_sum[48]), .Y(n10326));
XOR2X1 mul_U22837(.A(n9263), .B(n10326), .Y(dpath_mulcore_addout[48]));
XOR2X1 mul_U22838(.A(dpath_mulcore_addin_cout[48]), .B(dpath_mulcore_addin_sum[49]), .Y(n10331));
XOR2X1 mul_U22839(.A(n9264), .B(n10331), .Y(dpath_mulcore_addout[49]));
XOR2X1 mul_U22840(.A(dpath_mulcore_addin_cout[49]), .B(dpath_mulcore_addin_sum[50]), .Y(n10336));
XOR2X1 mul_U22841(.A(n9265), .B(n10336), .Y(dpath_mulcore_addout[50]));
XOR2X1 mul_U22842(.A(dpath_mulcore_addin_cout[50]), .B(dpath_mulcore_addin_sum[51]), .Y(n10341));
XOR2X1 mul_U22843(.A(n9266), .B(n10341), .Y(dpath_mulcore_addout[51]));
XOR2X1 mul_U22844(.A(dpath_mulcore_addin_cout[32]), .B(dpath_mulcore_addin_sum[33]), .Y(n10342));
XOR2X1 mul_U22845(.A(n9226), .B(n10342), .Y(dpath_mulcore_addout[33]));
XOR2X1 mul_U22846(.A(dpath_mulcore_addin_cout[51]), .B(dpath_mulcore_addin_sum[52]), .Y(n10348));
XOR2X1 mul_U22847(.A(n9267), .B(n10348), .Y(dpath_mulcore_addout[52]));
XOR2X1 mul_U22848(.A(dpath_mulcore_addin_cout[52]), .B(dpath_mulcore_addin_sum[53]), .Y(n10353));
XOR2X1 mul_U22849(.A(n9268), .B(n10353), .Y(dpath_mulcore_addout[53]));
XOR2X1 mul_U22850(.A(dpath_mulcore_addin_cout[53]), .B(dpath_mulcore_addin_sum[54]), .Y(n10358));
XOR2X1 mul_U22851(.A(n9269), .B(n10358), .Y(dpath_mulcore_addout[54]));
XOR2X1 mul_U22852(.A(dpath_mulcore_addin_cout[54]), .B(dpath_mulcore_addin_sum[55]), .Y(n10363));
XOR2X1 mul_U22853(.A(n9270), .B(n10363), .Y(dpath_mulcore_addout[55]));
XOR2X1 mul_U22854(.A(dpath_mulcore_addin_cout[55]), .B(dpath_mulcore_addin_sum[56]), .Y(n10368));
XOR2X1 mul_U22855(.A(n9271), .B(n10368), .Y(dpath_mulcore_addout[56]));
XOR2X1 mul_U22856(.A(dpath_mulcore_addin_cout[56]), .B(dpath_mulcore_addin_sum[57]), .Y(n10373));
XOR2X1 mul_U22857(.A(n9272), .B(n10373), .Y(dpath_mulcore_addout[57]));
XOR2X1 mul_U22858(.A(dpath_mulcore_addin_cout[57]), .B(dpath_mulcore_addin_sum[58]), .Y(n10378));
XOR2X1 mul_U22859(.A(n9273), .B(n10378), .Y(dpath_mulcore_addout[58]));
XOR2X1 mul_U22860(.A(dpath_mulcore_addin_cout[58]), .B(dpath_mulcore_addin_sum[59]), .Y(n10383));
XOR2X1 mul_U22861(.A(n9274), .B(n10383), .Y(dpath_mulcore_addout[59]));
XOR2X1 mul_U22862(.A(dpath_mulcore_addin_cout[59]), .B(dpath_mulcore_addin_sum[60]), .Y(n10388));
XOR2X1 mul_U22863(.A(n9275), .B(n10388), .Y(dpath_mulcore_addout[60]));
XOR2X1 mul_U22864(.A(dpath_mulcore_addin_cout[60]), .B(dpath_mulcore_addin_sum[61]), .Y(n10393));
XOR2X1 mul_U22865(.A(n9276), .B(n10393), .Y(dpath_mulcore_addout[61]));
XOR2X1 mul_U22866(.A(dpath_mulcore_addin_cout[33]), .B(dpath_mulcore_addin_sum[34]), .Y(n10394));
XOR2X1 mul_U22867(.A(n9227), .B(n10394), .Y(dpath_mulcore_addout[34]));
XOR2X1 mul_U22868(.A(dpath_mulcore_addin_cout[61]), .B(dpath_mulcore_addin_sum[62]), .Y(n10400));
XOR2X1 mul_U22869(.A(n9277), .B(n10400), .Y(dpath_mulcore_addout[62]));
XOR2X1 mul_U22870(.A(dpath_mulcore_addin_cout[62]), .B(dpath_mulcore_addin_sum[63]), .Y(n10405));
XOR2X1 mul_U22871(.A(n9278), .B(n10405), .Y(dpath_mulcore_addout[63]));
XOR2X1 mul_U22872(.A(dpath_mulcore_addin_cout[63]), .B(dpath_mulcore_addin_sum[64]), .Y(n10410));
XOR2X1 mul_U22873(.A(n9279), .B(n10410), .Y(dpath_mulcore_addout[64]));
XOR2X1 mul_U22874(.A(dpath_mulcore_addin_cout[64]), .B(dpath_mulcore_addin_sum[65]), .Y(n10415));
XOR2X1 mul_U22875(.A(n9280), .B(n10415), .Y(dpath_mulcore_addout[65]));
XOR2X1 mul_U22876(.A(dpath_mulcore_addin_cout[65]), .B(dpath_mulcore_addin_sum[66]), .Y(n10420));
XOR2X1 mul_U22877(.A(n9281), .B(n10420), .Y(dpath_mulcore_addout[66]));
XOR2X1 mul_U22878(.A(dpath_mulcore_addin_cout[66]), .B(dpath_mulcore_addin_sum[67]), .Y(n10425));
XOR2X1 mul_U22879(.A(n9282), .B(n10425), .Y(dpath_mulcore_addout[67]));
XOR2X1 mul_U22880(.A(dpath_mulcore_addin_cout[67]), .B(dpath_mulcore_addin_sum[68]), .Y(n10430));
XOR2X1 mul_U22881(.A(n9283), .B(n10430), .Y(dpath_mulcore_addout[68]));
XOR2X1 mul_U22882(.A(dpath_mulcore_addin_cout[68]), .B(dpath_mulcore_addin_sum[69]), .Y(n10435));
XOR2X1 mul_U22883(.A(n9284), .B(n10435), .Y(dpath_mulcore_addout[69]));
XOR2X1 mul_U22884(.A(dpath_mulcore_addin_cout[69]), .B(dpath_mulcore_addin_sum[70]), .Y(n10440));
XOR2X1 mul_U22885(.A(n9285), .B(n10440), .Y(dpath_mulcore_addout[70]));
XOR2X1 mul_U22886(.A(dpath_mulcore_addin_cout[70]), .B(dpath_mulcore_addin_sum[71]), .Y(n10445));
XOR2X1 mul_U22887(.A(n9286), .B(n10445), .Y(dpath_mulcore_addout[71]));
XOR2X1 mul_U22888(.A(dpath_mulcore_addin_cout[34]), .B(dpath_mulcore_addin_sum[35]), .Y(n10446));
XOR2X1 mul_U22889(.A(n9228), .B(n10446), .Y(dpath_mulcore_addout[35]));
XOR2X1 mul_U22890(.A(dpath_mulcore_addin_cout[71]), .B(dpath_mulcore_addin_sum[72]), .Y(n10452));
XOR2X1 mul_U22891(.A(n9287), .B(n10452), .Y(dpath_mulcore_addout[72]));
XOR2X1 mul_U22892(.A(dpath_mulcore_addin_cout[72]), .B(dpath_mulcore_addin_sum[73]), .Y(n10457));
XOR2X1 mul_U22893(.A(n9288), .B(n10457), .Y(dpath_mulcore_addout[73]));
XOR2X1 mul_U22894(.A(dpath_mulcore_addin_cout[73]), .B(dpath_mulcore_addin_sum[74]), .Y(n10462));
XOR2X1 mul_U22895(.A(n9289), .B(n10462), .Y(dpath_mulcore_addout[74]));
XOR2X1 mul_U22896(.A(dpath_mulcore_addin_cout[74]), .B(dpath_mulcore_addin_sum[75]), .Y(n10467));
XOR2X1 mul_U22897(.A(n9290), .B(n10467), .Y(dpath_mulcore_addout[75]));
XOR2X1 mul_U22898(.A(dpath_mulcore_addin_cout[75]), .B(dpath_mulcore_addin_sum[76]), .Y(n10472));
XOR2X1 mul_U22899(.A(n9291), .B(n10472), .Y(dpath_mulcore_addout[76]));
XOR2X1 mul_U22900(.A(dpath_mulcore_addin_cout[76]), .B(dpath_mulcore_addin_sum[77]), .Y(n10477));
XOR2X1 mul_U22901(.A(n9292), .B(n10477), .Y(dpath_mulcore_addout[77]));
XOR2X1 mul_U22902(.A(dpath_mulcore_addin_cout[77]), .B(dpath_mulcore_addin_sum[78]), .Y(n10482));
XOR2X1 mul_U22903(.A(n9293), .B(n10482), .Y(dpath_mulcore_addout[78]));
XOR2X1 mul_U22904(.A(dpath_mulcore_addin_cout[78]), .B(dpath_mulcore_addin_sum[79]), .Y(n10487));
XOR2X1 mul_U22905(.A(n9294), .B(n10487), .Y(dpath_mulcore_addout[79]));
XOR2X1 mul_U22906(.A(dpath_mulcore_addin_cout[79]), .B(dpath_mulcore_addin_sum[80]), .Y(n10492));
XOR2X1 mul_U22907(.A(n9295), .B(n10492), .Y(dpath_mulcore_addout[80]));
XOR2X1 mul_U22908(.A(dpath_mulcore_addin_cout[80]), .B(dpath_mulcore_addin_sum[81]), .Y(n10497));
XOR2X1 mul_U22909(.A(n9296), .B(n10497), .Y(dpath_mulcore_addout[81]));
XOR2X1 mul_U22910(.A(dpath_mulcore_addin_cout[35]), .B(dpath_mulcore_addin_sum[36]), .Y(n10498));
XOR2X1 mul_U22911(.A(n9229), .B(n10498), .Y(dpath_mulcore_addout[36]));
XOR2X1 mul_U22912(.A(dpath_mulcore_addin_cout[81]), .B(dpath_mulcore_addin_sum[82]), .Y(n10504));
XOR2X1 mul_U22913(.A(n9297), .B(n10504), .Y(dpath_mulcore_addout[82]));
XOR2X1 mul_U22914(.A(dpath_mulcore_addin_cout[82]), .B(dpath_mulcore_addin_sum[83]), .Y(n10509));
XOR2X1 mul_U22915(.A(n9298), .B(n10509), .Y(dpath_mulcore_addout[83]));
XOR2X1 mul_U22916(.A(dpath_mulcore_addin_cout[83]), .B(dpath_mulcore_addin_sum[84]), .Y(n10514));
XOR2X1 mul_U22917(.A(n9299), .B(n10514), .Y(dpath_mulcore_addout[84]));
XOR2X1 mul_U22918(.A(dpath_mulcore_addin_cout[84]), .B(dpath_mulcore_addin_sum[85]), .Y(n10519));
XOR2X1 mul_U22919(.A(n9300), .B(n10519), .Y(dpath_mulcore_addout[85]));
XOR2X1 mul_U22920(.A(dpath_mulcore_addin_cout[85]), .B(dpath_mulcore_addin_sum[86]), .Y(n10524));
XOR2X1 mul_U22921(.A(n9301), .B(n10524), .Y(dpath_mulcore_addout[86]));
XOR2X1 mul_U22922(.A(dpath_mulcore_addin_cout[86]), .B(dpath_mulcore_addin_sum[87]), .Y(n10529));
XOR2X1 mul_U22923(.A(n9302), .B(n10529), .Y(dpath_mulcore_addout[87]));
XOR2X1 mul_U22924(.A(dpath_mulcore_addin_cout[87]), .B(dpath_mulcore_addin_sum[88]), .Y(n10534));
XOR2X1 mul_U22925(.A(n9303), .B(n10534), .Y(dpath_mulcore_addout[88]));
XOR2X1 mul_U22926(.A(dpath_mulcore_addin_cout[88]), .B(dpath_mulcore_addin_sum[89]), .Y(n10539));
XOR2X1 mul_U22927(.A(n9304), .B(n10539), .Y(dpath_mulcore_addout[89]));
XOR2X1 mul_U22928(.A(dpath_mulcore_addin_cout[89]), .B(dpath_mulcore_addin_sum[90]), .Y(n10544));
XOR2X1 mul_U22929(.A(n9305), .B(n10544), .Y(dpath_mulcore_addout[90]));
XOR2X1 mul_U22930(.A(dpath_mulcore_addin_cout[90]), .B(dpath_mulcore_addin_sum[91]), .Y(n10549));
XOR2X1 mul_U22931(.A(n9306), .B(n10549), .Y(dpath_mulcore_addout[91]));
XOR2X1 mul_U22932(.A(dpath_mulcore_addin_cout[36]), .B(dpath_mulcore_addin_sum[37]), .Y(n10550));
XOR2X1 mul_U22933(.A(n9230), .B(n10550), .Y(dpath_mulcore_addout[37]));
XOR2X1 mul_U22934(.A(dpath_mulcore_addin_cout[91]), .B(dpath_mulcore_addin_sum[92]), .Y(n10556));
XOR2X1 mul_U22935(.A(n9307), .B(n10556), .Y(dpath_mulcore_addout[92]));
XOR2X1 mul_U22936(.A(dpath_mulcore_addin_cout[92]), .B(dpath_mulcore_addin_sum[93]), .Y(n10561));
XOR2X1 mul_U22937(.A(n9308), .B(n10561), .Y(dpath_mulcore_addout[93]));
XOR2X1 mul_U22938(.A(dpath_mulcore_addin_cout[93]), .B(dpath_mulcore_addin_sum[94]), .Y(n10566));
XOR2X1 mul_U22939(.A(n9309), .B(n10566), .Y(dpath_mulcore_addout[94]));
XOR2X1 mul_U22940(.A(dpath_mulcore_addin_cout[94]), .B(dpath_mulcore_addin_sum[95]), .Y(n10571));
XOR2X1 mul_U22941(.A(n9310), .B(n10571), .Y(dpath_mulcore_addout[95]));
XOR2X1 mul_U22942(.A(dpath_mulcore_addin_cout[95]), .B(dpath_mulcore_addin_sum[96]), .Y(n10576));
XOR2X1 mul_U22943(.A(n9311), .B(n10576), .Y(dpath_mulcore_addout[96]));
XOR2X1 mul_U22944(.A(dpath_mulcore_addin_cout[96]), .B(dpath_mulcore_addin_sum[97]), .Y(n10581));
XOR2X1 mul_U22945(.A(n6066), .B(n10581), .Y(dpath_mulcore_add_co96));
XOR2X1 mul_U22946(.A(dpath_mulcore_addin_cout[37]), .B(dpath_mulcore_addin_sum[38]), .Y(n10583));
XOR2X1 mul_U22947(.A(n9231), .B(n10583), .Y(dpath_mulcore_addout[38]));
XOR2X1 mul_U22948(.A(dpath_mulcore_addin_cout[38]), .B(dpath_mulcore_addin_sum[39]), .Y(n10585));
XOR2X1 mul_U22949(.A(n9232), .B(n10585), .Y(dpath_mulcore_addout[39]));
XOR2X1 mul_U22950(.A(dpath_mulcore_addin_cout[39]), .B(dpath_mulcore_addin_sum[40]), .Y(n10587));
XOR2X1 mul_U22951(.A(n9233), .B(n10587), .Y(dpath_mulcore_addout[40]));
XOR2X1 mul_U22952(.A(dpath_mulcore_addin_cout[40]), .B(dpath_mulcore_addin_sum[41]), .Y(n10589));
XOR2X1 mul_U22953(.A(n9234), .B(n10589), .Y(dpath_mulcore_addout[41]));
XOR2X1 mul_U22954(.A(dpath_mulcore_add_co96), .B(dpath_acc_reg[129]), .Y(dpath_mulcore_addout[97]));
XNOR2X1 mul_U22955(.A(dpath_acc_reg[130]), .B(n6067), .Y(dpath_mulcore_addout[98]));
XOR2X1 mul_U22956(.A(dpath_acc_reg[131]), .B(n10594), .Y(dpath_mulcore_addout[99]));
XNOR2X1 mul_U22957(.A(dpath_acc_reg[132]), .B(n6068), .Y(dpath_mulcore_addout[100]));
XOR2X1 mul_U22958(.A(dpath_acc_reg[133]), .B(n10596), .Y(dpath_mulcore_addout[101]));
XNOR2X1 mul_U22959(.A(dpath_acc_reg[134]), .B(n6069), .Y(dpath_mulcore_addout[102]));
XNOR2X1 mul_U22960(.A(dpath_acc_reg[135]), .B(n6070), .Y(dpath_mulcore_addout[103]));
endmodule
