module sparc_exu ( exu_tlu_wsr_data_m, exu_tlu_va_oor_m, 
        exu_tlu_va_oor_jl_ret_m, exu_tlu_ue_trap_m, exu_tlu_ttype_vld_m, 
        exu_tlu_ttype_m, exu_tlu_spill_wtype, exu_tlu_spill_tid, 
        exu_tlu_spill_other, exu_tlu_spill, exu_tlu_misalign_addr_jmpl_rtn_m, 
        exu_tlu_cwp_retry, exu_tlu_cwp_cmplt_tid, exu_tlu_cwp_cmplt, 
        exu_tlu_cwp3_w, exu_tlu_cwp2_w, exu_tlu_cwp1_w, exu_tlu_cwp0_w, 
        exu_tlu_ccr3_w, exu_tlu_ccr2_w, exu_tlu_ccr1_w, exu_tlu_ccr0_w, 
        exu_spu_rs3_data_e, exu_mul_rs2_data, exu_mul_rs1_data, 
        exu_mul_input_vld, exu_mmu_early_va_e, exu_lsu_rs3_data_e, 
        exu_lsu_rs2_data_e, exu_lsu_priority_trap_m, exu_lsu_ldst_va_e, 
        exu_lsu_early_va_e, exu_ifu_va_oor_m, exu_ifu_spill_e, exu_ifu_regz_e, 
        exu_ifu_regn_e, exu_ifu_oddwin_s, exu_ifu_longop_done_g, 
        exu_ifu_inj_ack, exu_ifu_err_reg_m, exu_ifu_ecc_ue_m, exu_ifu_ecc_ce_m, 
        exu_ifu_cc_d, exu_ifu_brpc_e, exu_ffu_wsr_inst_e, short_so0, short_so1, 
        so0, exu_ifu_err_synd_m, tlu_exu_rsr_data_m, tlu_exu_priv_trap_m, 
        tlu_exu_pic_twobelow_m, tlu_exu_pic_onebelow_m, 
        tlu_exu_cwpccr_update_m, tlu_exu_cwp_retry_m, tlu_exu_cwp_m, 
        tlu_exu_ccr_m, tlu_exu_agp_tid, tlu_exu_agp_swap, tlu_exu_agp, sehold, 
        se, rclk, mul_data_out, mul_exu_ack, lsu_exu_thr_m, 
        lsu_exu_st_dtlb_perr_g, lsu_exu_rd_m, lsu_exu_ldxa_m, 
        lsu_exu_ldxa_data_g, lsu_exu_ldst_miss_g2, lsu_exu_flush_pipe_w, 
        lsu_exu_dfill_vld_g, lsu_exu_dfill_data_g, ifu_tlu_wsr_inst_d, 
        ifu_tlu_sraddr_d, ifu_tlu_flush_m, ifu_exu_wen_d, ifu_exu_useimm_d, 
        ifu_exu_usecin_d, ifu_exu_use_rsr_e_l, ifu_exu_tv_d, 
        ifu_exu_ttype_vld_m, ifu_exu_tid_s2, ifu_exu_tcc_e, ifu_exu_tagop_d, 
        ifu_exu_shiftop_d, ifu_exu_sethi_inst_d, ifu_exu_setcc_d, 
        ifu_exu_saved_e, ifu_exu_save_d, ifu_exu_rs3o_vld_d, 
        ifu_exu_rs3e_vld_d, ifu_exu_rs3_s, ifu_exu_rs2_vld_d, ifu_exu_rs2_s, 
        ifu_exu_rs1_vld_d, ifu_exu_rs1_s, ifu_exu_return_d, ifu_exu_restored_e, 
        ifu_exu_restore_d, ifu_exu_ren3_s, ifu_exu_ren2_s, ifu_exu_ren1_s, 
        ifu_exu_rd_ifusr_e, ifu_exu_rd_ffusr_e, ifu_exu_rd_exusr_e, 
        ifu_exu_rd_d, ifu_exu_range_check_other_d, ifu_exu_range_check_jlret_d, 
        ifu_exu_pcver_e, ifu_exu_pc_d, ifu_exu_nceen_e, ifu_exu_muls_d, 
        ifu_exu_muldivop_d, ifu_exu_kill_e, ifu_exu_invert_d, 
        ifu_exu_inst_vld_w, ifu_exu_inst_vld_e, ifu_exu_inj_irferr, 
        ifu_exu_imm_data_d, ifu_exu_ialign_d, ifu_exu_flushw_e, 
        ifu_exu_enshift_d, ifu_exu_ecc_mask, ifu_exu_dontmv_regz1_e, 
        ifu_exu_dontmv_regz0_e, ifu_exu_disable_ce_e, ifu_exu_dbrinst_d, 
        ifu_exu_casa_d, ifu_exu_aluop_d, ifu_exu_addr_mask_d, grst_l, 
        ffu_exu_rsr_data_m, arst_l, mux_drive_disable, mem_write_disable, 
        short_si0, short_si1, si0 );
  output [63:0] exu_tlu_wsr_data_m;
  output [8:0] exu_tlu_ttype_m;
  output [2:0] exu_tlu_spill_wtype;
  output [1:0] exu_tlu_spill_tid;
  output [1:0] exu_tlu_cwp_cmplt_tid;
  output [2:0] exu_tlu_cwp3_w;
  output [2:0] exu_tlu_cwp2_w;
  output [2:0] exu_tlu_cwp1_w;
  output [2:0] exu_tlu_cwp0_w;
  output [7:0] exu_tlu_ccr3_w;
  output [7:0] exu_tlu_ccr2_w;
  output [7:0] exu_tlu_ccr1_w;
  output [7:0] exu_tlu_ccr0_w;
  output [63:0] exu_spu_rs3_data_e;
  output [63:0] exu_mul_rs2_data;
  output [63:0] exu_mul_rs1_data;
  output [7:0] exu_mmu_early_va_e;
  output [63:0] exu_lsu_rs3_data_e;
  output [63:0] exu_lsu_rs2_data_e;
  output [47:0] exu_lsu_ldst_va_e;
  output [10:3] exu_lsu_early_va_e;
  output [3:0] exu_ifu_oddwin_s;
  output [3:0] exu_ifu_longop_done_g;
  output [7:0] exu_ifu_err_reg_m;
  output [7:0] exu_ifu_cc_d;
  output [47:0] exu_ifu_brpc_e;
  output [7:0] exu_ifu_err_synd_m;
  input [63:0] tlu_exu_rsr_data_m;
  input [2:0] tlu_exu_cwp_m;
  input [7:0] tlu_exu_ccr_m;
  input [1:0] tlu_exu_agp_tid;
  input [1:0] tlu_exu_agp;
  input [63:0] mul_data_out;
  input [1:0] lsu_exu_thr_m;
  input [4:0] lsu_exu_rd_m;
  input [63:0] lsu_exu_ldxa_data_g;
  input [63:0] lsu_exu_dfill_data_g;
  input [6:0] ifu_tlu_sraddr_d;
  input [1:0] ifu_exu_tid_s2;
  input [2:0] ifu_exu_shiftop_d;
  input [4:0] ifu_exu_rs3_s;
  input [4:0] ifu_exu_rs2_s;
  input [4:0] ifu_exu_rs1_s;
  input [4:0] ifu_exu_rd_d;
  input [63:0] ifu_exu_pcver_e;
  input [47:0] ifu_exu_pc_d;
  input [4:0] ifu_exu_muldivop_d;
  input [31:0] ifu_exu_imm_data_d;
  input [7:0] ifu_exu_ecc_mask;
  input [2:0] ifu_exu_aluop_d;
  input [63:0] ffu_exu_rsr_data_m;
  input tlu_exu_priv_trap_m, tlu_exu_pic_twobelow_m, tlu_exu_pic_onebelow_m,
         tlu_exu_cwpccr_update_m, tlu_exu_cwp_retry_m, tlu_exu_agp_swap,
         sehold, se, rclk, mul_exu_ack, lsu_exu_st_dtlb_perr_g, lsu_exu_ldxa_m,
         lsu_exu_ldst_miss_g2, lsu_exu_flush_pipe_w, lsu_exu_dfill_vld_g,
         ifu_tlu_wsr_inst_d, ifu_tlu_flush_m, ifu_exu_wen_d, ifu_exu_useimm_d,
         ifu_exu_usecin_d, ifu_exu_use_rsr_e_l, ifu_exu_tv_d,
         ifu_exu_ttype_vld_m, ifu_exu_tcc_e, ifu_exu_tagop_d,
         ifu_exu_sethi_inst_d, ifu_exu_setcc_d, ifu_exu_saved_e,
         ifu_exu_save_d, ifu_exu_rs3o_vld_d, ifu_exu_rs3e_vld_d,
         ifu_exu_rs2_vld_d, ifu_exu_rs1_vld_d, ifu_exu_return_d,
         ifu_exu_restored_e, ifu_exu_restore_d, ifu_exu_ren3_s, ifu_exu_ren2_s,
         ifu_exu_ren1_s, ifu_exu_rd_ifusr_e, ifu_exu_rd_ffusr_e,
         ifu_exu_rd_exusr_e, ifu_exu_range_check_other_d,
         ifu_exu_range_check_jlret_d, ifu_exu_nceen_e, ifu_exu_muls_d,
         ifu_exu_kill_e, ifu_exu_invert_d, ifu_exu_inst_vld_w,
         ifu_exu_inst_vld_e, ifu_exu_inj_irferr, ifu_exu_ialign_d,
         ifu_exu_flushw_e, ifu_exu_enshift_d, ifu_exu_dontmv_regz1_e,
         ifu_exu_dontmv_regz0_e, ifu_exu_disable_ce_e, ifu_exu_dbrinst_d,
         ifu_exu_casa_d, ifu_exu_addr_mask_d, grst_l, arst_l,
         mux_drive_disable, mem_write_disable, short_si0, short_si1, si0;
  output exu_tlu_va_oor_m, exu_tlu_va_oor_jl_ret_m, exu_tlu_ue_trap_m,
         exu_tlu_ttype_vld_m, exu_tlu_spill_other, exu_tlu_spill,
         exu_tlu_misalign_addr_jmpl_rtn_m, exu_tlu_cwp_retry,
         exu_tlu_cwp_cmplt, exu_mul_input_vld, exu_lsu_priority_trap_m,
         exu_ifu_va_oor_m, exu_ifu_spill_e, exu_ifu_regz_e, exu_ifu_regn_e,
         exu_ifu_inj_ack, exu_ifu_ecc_ue_m, exu_ifu_ecc_ce_m,
         exu_ffu_wsr_inst_e, short_so0, short_so1, so0;
  wire   n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712,
         n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720,
         n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728,
         n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736,
         n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744,
         n31745, n31746, n31747, n31748, ecl_byp_rs1_mux2_sel_e,
         ecl_byp_rs1_mux2_sel_rf, ecl_byp_rs1_mux2_sel_ld,
         ecl_byp_rs1_mux2_sel_usemux1, ecl_byp_rs1_mux1_sel_m,
         ecl_byp_rs1_mux1_sel_w, ecl_byp_rs1_mux1_sel_w2,
         ecl_byp_rs1_mux1_sel_other, ecl_byp_rcc_mux2_sel_e,
         ecl_byp_rcc_mux2_sel_rf, ecl_byp_rcc_mux2_sel_ld,
         ecl_byp_rcc_mux2_sel_usemux1, ecl_byp_rcc_mux1_sel_m,
         ecl_byp_rcc_mux1_sel_w, ecl_byp_rcc_mux1_sel_w2,
         ecl_byp_rs2_mux2_sel_e, ecl_byp_rs2_mux2_sel_rf,
         ecl_byp_rs2_mux2_sel_ld, ecl_byp_rs2_mux2_sel_usemux1,
         ecl_byp_rs2_mux1_sel_m, ecl_byp_rs2_mux1_sel_w,
         ecl_byp_rs3_mux2_sel_e, ecl_byp_rs3_mux2_sel_ld,
         ecl_byp_rs3_mux1_sel_m, ecl_byp_rs3_mux1_sel_w,
         ecl_byp_rs3h_mux2_sel_e, ecl_byp_rs3h_mux2_sel_ld,
         ecl_byp_rs3h_mux1_sel_m, ecl_byp_rs3h_mux1_sel_w,
         ecl_byp_rs1_longmux_sel_g2, ecl_byp_rs1_longmux_sel_w2,
         ecl_byp_rs2_longmux_sel_g2, ecl_byp_rs2_longmux_sel_w2,
         ecl_byp_rs3_longmux_sel_g2, ecl_byp_rs3_longmux_sel_w2,
         ecl_byp_rs3h_longmux_sel_g2, ecl_byp_rs3h_longmux_sel_w2,
         ecl_byp_sel_pipe_m, ecl_byp_sel_ecc_m, ecl_byp_sel_muldiv_g,
         ecl_byp_sel_load_g, ecl_byp_ldxa_g, ecl_byp_restore_m,
         ecl_byp_sel_yreg_e, ecl_byp_sel_eclpr_e, ecl_byp_sel_ifusr_e,
         ecl_byp_sel_alu_e, ecl_byp_sel_ifex_m, ecl_byp_sel_ffusr_m,
         ecl_byp_sel_tlusr_m, ecc_ecl_rs1_ce, ecc_ecl_rs1_ue, ecc_ecl_rs2_ce,
         ecc_ecl_rs2_ue, ecc_ecl_rs3_ce, ecc_ecl_rs3_ue, ecl_ecc_rs1_use_rf_e,
         ecl_ecc_rs2_use_rf_e, ecl_ecc_rs3_use_rf_e, ecl_ecc_sel_rs1_m_l,
         ecl_ecc_sel_rs2_m_l, ecl_ecc_sel_rs3_m_l, ecl_ecc_log_rs1_m,
         ecl_ecc_log_rs2_m, ecl_ecc_log_rs3_m, ecl_alu_casa_e, ecl_div_cin,
         ecl_div_dividend_sign, ecl_div_keep_d, ecl_div_last_cycle,
         ecl_div_mul_get_32bit_data, ecl_div_mul_get_new_data,
         ecl_div_mul_sext_rs1_e, ecl_div_mul_sext_rs2_e, ecl_div_newq,
         ecl_div_sel_64b, ecl_div_sel_adder, ecl_div_sel_neg32,
         ecl_div_sel_u32, ecl_div_upper33_zero, ecl_div_xinmask,
         ecl_div_yreg_wen_g[0] , ecl_rml_canrestore_wen_w,
         ecl_rml_cansave_wen_w, ecl_rml_cleanwin_wen_w, ecl_rml_cwp_wen_e,
         ecl_rml_otherwin_wen_w, ecl_rml_wstate_wen_w, ecl_alu_out_sel_rs3_e_l,
         ecl_alu_out_sel_shift_e_l, ecl_alu_out_sel_logic_e_l,
         ecl_alu_log_sel_and_e, ecl_alu_log_sel_or_e, ecl_alu_log_sel_xor_e,
         ecl_alu_log_sel_move_e, ecl_alu_sethi_inst_e, ecl_alu_cin_e,
         ecl_shft_lshift_e_l, ecl_div_ld_inputs, ecl_div_sel_div,
         ecl_div_div64, ecl_shft_extendbit_e, ecl_shft_extend32bit_e_l,
         ecl_div_zero_rs2_e, ecl_div_muls_rs1_31_e_l, ecl_div_yreg_data_31_g,
         ecl_rml_kill_e, ecl_rml_kill_w, ecl_div_mul_wen, ecl_div_muls,
         ecl_rml_early_flush_w, ecl_rml_inst_vld_w, div_ecl_adder_out_31,
         div_ecl_cout32, div_ecl_cout64, div_ecl_d_62, div_ecl_d_msb,
         div_ecl_detect_zero_high, div_ecl_detect_zero_low,
         div_ecl_dividend_msb, div_ecl_gencc_in_31, div_ecl_low32_nonzero,
         div_ecl_x_msb, rml_ecl_kill_m, rml_ecl_rmlop_done_e,
         alu_ecl_add_n64_e, alu_ecl_log_n64_e, alu_ecl_log_n32_e,
         alu_ecl_zhigh_e, alu_ecl_zlow_e, alu_ecl_cout32_e,
         alu_ecl_adderin2_63_e, alu_ecl_adderin2_31_e,
         alu_ecl_mem_addr_invalid_e_l, rml_ecl_clean_window_e, rml_ecl_fill_e,
         rml_ecl_other_e, bypass_rd_synd_w2_l[7] , bypass_rd_synd_w2_l[6] ,
         bypass_rd_synd_w2_l[5] , bypass_rd_synd_w2_l[4] ,
         bypass_rd_synd_w2_l[3] , bypass_rd_synd_w2_l[2] ,
         bypass_rd_synd_w2_l[1] , bypass_rd_synd_w2_l[0] ,
         bypass_rd_synd_w_l[7] , bypass_rd_synd_w_l[6] ,
         bypass_rd_synd_w_l[5] , bypass_rd_synd_w_l[4] ,
         bypass_rd_synd_w_l[3] , bypass_rd_synd_w_l[2] ,
         bypass_rd_synd_w_l[1] , bypass_rd_synd_w_l[0] ,
         bypass_rs3h_data_btwn_mux[31] , bypass_rs3h_data_btwn_mux[30] ,
         bypass_rs3h_data_btwn_mux[29] , bypass_rs3h_data_btwn_mux[28] ,
         bypass_rs3h_data_btwn_mux[27] , bypass_rs3h_data_btwn_mux[26] ,
         bypass_rs3h_data_btwn_mux[25] , bypass_rs3h_data_btwn_mux[24] ,
         bypass_rs3h_data_btwn_mux[23] , bypass_rs3h_data_btwn_mux[22] ,
         bypass_rs3h_data_btwn_mux[21] , bypass_rs3h_data_btwn_mux[20] ,
         bypass_rs3h_data_btwn_mux[19] , bypass_rs3h_data_btwn_mux[18] ,
         bypass_rs3h_data_btwn_mux[17] , bypass_rs3h_data_btwn_mux[16] ,
         bypass_rs3h_data_btwn_mux[15] , bypass_rs3h_data_btwn_mux[14] ,
         bypass_rs3h_data_btwn_mux[13] , bypass_rs3h_data_btwn_mux[12] ,
         bypass_rs3h_data_btwn_mux[11] , bypass_rs3h_data_btwn_mux[10] ,
         bypass_rs3h_data_btwn_mux[9] , bypass_rs3h_data_btwn_mux[8] ,
         bypass_rs3h_data_btwn_mux[7] , bypass_rs3h_data_btwn_mux[6] ,
         bypass_rs3h_data_btwn_mux[5] , bypass_rs3h_data_btwn_mux[4] ,
         bypass_rs3h_data_btwn_mux[3] , bypass_rs3h_data_btwn_mux[2] ,
         bypass_rs3h_data_btwn_mux[1] , bypass_rs3h_data_btwn_mux[0] ,
         bypass_rs3_data_btwn_mux[63] , bypass_rs3_data_btwn_mux[62] ,
         bypass_rs3_data_btwn_mux[61] , bypass_rs3_data_btwn_mux[60] ,
         bypass_rs3_data_btwn_mux[59] , bypass_rs3_data_btwn_mux[58] ,
         bypass_rs3_data_btwn_mux[57] , bypass_rs3_data_btwn_mux[56] ,
         bypass_rs3_data_btwn_mux[55] , bypass_rs3_data_btwn_mux[54] ,
         bypass_rs3_data_btwn_mux[53] , bypass_rs3_data_btwn_mux[52] ,
         bypass_rs3_data_btwn_mux[51] , bypass_rs3_data_btwn_mux[50] ,
         bypass_rs3_data_btwn_mux[49] , bypass_rs3_data_btwn_mux[48] ,
         bypass_rs3_data_btwn_mux[47] , bypass_rs3_data_btwn_mux[46] ,
         bypass_rs3_data_btwn_mux[45] , bypass_rs3_data_btwn_mux[44] ,
         bypass_rs3_data_btwn_mux[43] , bypass_rs3_data_btwn_mux[42] ,
         bypass_rs3_data_btwn_mux[41] , bypass_rs3_data_btwn_mux[40] ,
         bypass_rs3_data_btwn_mux[39] , bypass_rs3_data_btwn_mux[38] ,
         bypass_rs3_data_btwn_mux[37] , bypass_rs3_data_btwn_mux[36] ,
         bypass_rs3_data_btwn_mux[35] , bypass_rs3_data_btwn_mux[34] ,
         bypass_rs3_data_btwn_mux[33] , bypass_rs3_data_btwn_mux[32] ,
         bypass_rs3_data_btwn_mux[31] , bypass_rs3_data_btwn_mux[30] ,
         bypass_rs3_data_btwn_mux[29] , bypass_rs3_data_btwn_mux[28] ,
         bypass_rs3_data_btwn_mux[27] , bypass_rs3_data_btwn_mux[26] ,
         bypass_rs3_data_btwn_mux[25] , bypass_rs3_data_btwn_mux[24] ,
         bypass_rs3_data_btwn_mux[23] , bypass_rs3_data_btwn_mux[22] ,
         bypass_rs3_data_btwn_mux[21] , bypass_rs3_data_btwn_mux[20] ,
         bypass_rs3_data_btwn_mux[19] , bypass_rs3_data_btwn_mux[18] ,
         bypass_rs3_data_btwn_mux[17] , bypass_rs3_data_btwn_mux[16] ,
         bypass_rs3_data_btwn_mux[15] , bypass_rs3_data_btwn_mux[14] ,
         bypass_rs3_data_btwn_mux[13] , bypass_rs3_data_btwn_mux[12] ,
         bypass_rs3_data_btwn_mux[11] , bypass_rs3_data_btwn_mux[10] ,
         bypass_rs3_data_btwn_mux[9] , bypass_rs3_data_btwn_mux[8] ,
         bypass_rs3_data_btwn_mux[7] , bypass_rs3_data_btwn_mux[6] ,
         bypass_rs3_data_btwn_mux[5] , bypass_rs3_data_btwn_mux[4] ,
         bypass_rs3_data_btwn_mux[3] , bypass_rs3_data_btwn_mux[2] ,
         bypass_rs3_data_btwn_mux[1] , bypass_rs3_data_btwn_mux[0] ,
         bypass_rs2_data_btwn_mux[63] , bypass_rs2_data_btwn_mux[62] ,
         bypass_rs2_data_btwn_mux[61] , bypass_rs2_data_btwn_mux[60] ,
         bypass_rs2_data_btwn_mux[59] , bypass_rs2_data_btwn_mux[58] ,
         bypass_rs2_data_btwn_mux[57] , bypass_rs2_data_btwn_mux[56] ,
         bypass_rs2_data_btwn_mux[55] , bypass_rs2_data_btwn_mux[54] ,
         bypass_rs2_data_btwn_mux[53] , bypass_rs2_data_btwn_mux[52] ,
         bypass_rs2_data_btwn_mux[51] , bypass_rs2_data_btwn_mux[50] ,
         bypass_rs2_data_btwn_mux[49] , bypass_rs2_data_btwn_mux[48] ,
         bypass_rs2_data_btwn_mux[47] , bypass_rs2_data_btwn_mux[46] ,
         bypass_rs2_data_btwn_mux[45] , bypass_rs2_data_btwn_mux[44] ,
         bypass_rs2_data_btwn_mux[43] , bypass_rs2_data_btwn_mux[42] ,
         bypass_rs2_data_btwn_mux[41] , bypass_rs2_data_btwn_mux[40] ,
         bypass_rs2_data_btwn_mux[39] , bypass_rs2_data_btwn_mux[38] ,
         bypass_rs2_data_btwn_mux[37] , bypass_rs2_data_btwn_mux[36] ,
         bypass_rs2_data_btwn_mux[35] , bypass_rs2_data_btwn_mux[34] ,
         bypass_rs2_data_btwn_mux[33] , bypass_rs2_data_btwn_mux[32] ,
         bypass_rs2_data_btwn_mux[31] , bypass_rs2_data_btwn_mux[30] ,
         bypass_rs2_data_btwn_mux[29] , bypass_rs2_data_btwn_mux[28] ,
         bypass_rs2_data_btwn_mux[27] , bypass_rs2_data_btwn_mux[26] ,
         bypass_rs2_data_btwn_mux[25] , bypass_rs2_data_btwn_mux[24] ,
         bypass_rs2_data_btwn_mux[23] , bypass_rs2_data_btwn_mux[22] ,
         bypass_rs2_data_btwn_mux[21] , bypass_rs2_data_btwn_mux[20] ,
         bypass_rs2_data_btwn_mux[19] , bypass_rs2_data_btwn_mux[18] ,
         bypass_rs2_data_btwn_mux[17] , bypass_rs2_data_btwn_mux[16] ,
         bypass_rs2_data_btwn_mux[15] , bypass_rs2_data_btwn_mux[14] ,
         bypass_rs2_data_btwn_mux[13] , bypass_rs2_data_btwn_mux[12] ,
         bypass_rs2_data_btwn_mux[11] , bypass_rs2_data_btwn_mux[10] ,
         bypass_rs2_data_btwn_mux[9] , bypass_rs2_data_btwn_mux[8] ,
         bypass_rs2_data_btwn_mux[7] , bypass_rs2_data_btwn_mux[6] ,
         bypass_rs2_data_btwn_mux[5] , bypass_rs2_data_btwn_mux[4] ,
         bypass_rs2_data_btwn_mux[3] , bypass_rs2_data_btwn_mux[2] ,
         bypass_rs2_data_btwn_mux[1] , bypass_rs2_data_btwn_mux[0] ,
         bypass_rcc_data_btwn_mux[63] , bypass_rcc_data_btwn_mux[62] ,
         bypass_rcc_data_btwn_mux[61] , bypass_rcc_data_btwn_mux[60] ,
         bypass_rcc_data_btwn_mux[59] , bypass_rcc_data_btwn_mux[58] ,
         bypass_rcc_data_btwn_mux[57] , bypass_rcc_data_btwn_mux[56] ,
         bypass_rcc_data_btwn_mux[55] , bypass_rcc_data_btwn_mux[54] ,
         bypass_rcc_data_btwn_mux[53] , bypass_rcc_data_btwn_mux[52] ,
         bypass_rcc_data_btwn_mux[51] , bypass_rcc_data_btwn_mux[50] ,
         bypass_rcc_data_btwn_mux[49] , bypass_rcc_data_btwn_mux[48] ,
         bypass_rcc_data_btwn_mux[47] , bypass_rcc_data_btwn_mux[46] ,
         bypass_rcc_data_btwn_mux[45] , bypass_rcc_data_btwn_mux[44] ,
         bypass_rcc_data_btwn_mux[43] , bypass_rcc_data_btwn_mux[42] ,
         bypass_rcc_data_btwn_mux[41] , bypass_rcc_data_btwn_mux[40] ,
         bypass_rcc_data_btwn_mux[39] , bypass_rcc_data_btwn_mux[38] ,
         bypass_rcc_data_btwn_mux[37] , bypass_rcc_data_btwn_mux[36] ,
         bypass_rcc_data_btwn_mux[35] , bypass_rcc_data_btwn_mux[34] ,
         bypass_rcc_data_btwn_mux[33] , bypass_rcc_data_btwn_mux[32] ,
         bypass_rcc_data_btwn_mux[31] , bypass_rcc_data_btwn_mux[30] ,
         bypass_rcc_data_btwn_mux[29] , bypass_rcc_data_btwn_mux[28] ,
         bypass_rcc_data_btwn_mux[27] , bypass_rcc_data_btwn_mux[26] ,
         bypass_rcc_data_btwn_mux[25] , bypass_rcc_data_btwn_mux[24] ,
         bypass_rcc_data_btwn_mux[23] , bypass_rcc_data_btwn_mux[22] ,
         bypass_rcc_data_btwn_mux[21] , bypass_rcc_data_btwn_mux[20] ,
         bypass_rcc_data_btwn_mux[19] , bypass_rcc_data_btwn_mux[18] ,
         bypass_rcc_data_btwn_mux[17] , bypass_rcc_data_btwn_mux[16] ,
         bypass_rcc_data_btwn_mux[15] , bypass_rcc_data_btwn_mux[14] ,
         bypass_rcc_data_btwn_mux[13] , bypass_rcc_data_btwn_mux[12] ,
         bypass_rcc_data_btwn_mux[11] , bypass_rcc_data_btwn_mux[10] ,
         bypass_rcc_data_btwn_mux[9] , bypass_rcc_data_btwn_mux[8] ,
         bypass_rcc_data_btwn_mux[7] , bypass_rcc_data_btwn_mux[6] ,
         bypass_rcc_data_btwn_mux[5] , bypass_rcc_data_btwn_mux[4] ,
         bypass_rcc_data_btwn_mux[3] , bypass_rcc_data_btwn_mux[2] ,
         bypass_rcc_data_btwn_mux[1] , bypass_rcc_data_btwn_mux[0] ,
         bypass_rs1_data_btwn_mux[63] , bypass_rs1_data_btwn_mux[62] ,
         bypass_rs1_data_btwn_mux[61] , bypass_rs1_data_btwn_mux[60] ,
         bypass_rs1_data_btwn_mux[59] , bypass_rs1_data_btwn_mux[58] ,
         bypass_rs1_data_btwn_mux[57] , bypass_rs1_data_btwn_mux[56] ,
         bypass_rs1_data_btwn_mux[55] , bypass_rs1_data_btwn_mux[54] ,
         bypass_rs1_data_btwn_mux[53] , bypass_rs1_data_btwn_mux[52] ,
         bypass_rs1_data_btwn_mux[51] , bypass_rs1_data_btwn_mux[50] ,
         bypass_rs1_data_btwn_mux[49] , bypass_rs1_data_btwn_mux[48] ,
         bypass_rs1_data_btwn_mux[47] , bypass_rs1_data_btwn_mux[46] ,
         bypass_rs1_data_btwn_mux[45] , bypass_rs1_data_btwn_mux[44] ,
         bypass_rs1_data_btwn_mux[43] , bypass_rs1_data_btwn_mux[42] ,
         bypass_rs1_data_btwn_mux[41] , bypass_rs1_data_btwn_mux[40] ,
         bypass_rs1_data_btwn_mux[39] , bypass_rs1_data_btwn_mux[38] ,
         bypass_rs1_data_btwn_mux[37] , bypass_rs1_data_btwn_mux[36] ,
         bypass_rs1_data_btwn_mux[35] , bypass_rs1_data_btwn_mux[34] ,
         bypass_rs1_data_btwn_mux[33] , bypass_rs1_data_btwn_mux[32] ,
         bypass_rs1_data_btwn_mux[31] , bypass_rs1_data_btwn_mux[30] ,
         bypass_rs1_data_btwn_mux[29] , bypass_rs1_data_btwn_mux[28] ,
         bypass_rs1_data_btwn_mux[27] , bypass_rs1_data_btwn_mux[26] ,
         bypass_rs1_data_btwn_mux[25] , bypass_rs1_data_btwn_mux[24] ,
         bypass_rs1_data_btwn_mux[23] , bypass_rs1_data_btwn_mux[22] ,
         bypass_rs1_data_btwn_mux[21] , bypass_rs1_data_btwn_mux[20] ,
         bypass_rs1_data_btwn_mux[19] , bypass_rs1_data_btwn_mux[18] ,
         bypass_rs1_data_btwn_mux[17] , bypass_rs1_data_btwn_mux[16] ,
         bypass_rs1_data_btwn_mux[15] , bypass_rs1_data_btwn_mux[14] ,
         bypass_rs1_data_btwn_mux[13] , bypass_rs1_data_btwn_mux[12] ,
         bypass_rs1_data_btwn_mux[11] , bypass_rs1_data_btwn_mux[10] ,
         bypass_rs1_data_btwn_mux[9] , bypass_rs1_data_btwn_mux[8] ,
         bypass_rs1_data_btwn_mux[7] , bypass_rs1_data_btwn_mux[6] ,
         bypass_rs1_data_btwn_mux[5] , bypass_rs1_data_btwn_mux[4] ,
         bypass_rs1_data_btwn_mux[3] , bypass_rs1_data_btwn_mux[2] ,
         bypass_rs1_data_btwn_mux[1] , bypass_rs1_data_btwn_mux[0] ,
         bypass_rs3h_data_w2[31] , bypass_rs3h_data_w2[30] ,
         bypass_rs3h_data_w2[29] , bypass_rs3h_data_w2[28] ,
         bypass_rs3h_data_w2[27] , bypass_rs3h_data_w2[26] ,
         bypass_rs3h_data_w2[25] , bypass_rs3h_data_w2[24] ,
         bypass_rs3h_data_w2[23] , bypass_rs3h_data_w2[22] ,
         bypass_rs3h_data_w2[21] , bypass_rs3h_data_w2[20] ,
         bypass_rs3h_data_w2[19] , bypass_rs3h_data_w2[18] ,
         bypass_rs3h_data_w2[17] , bypass_rs3h_data_w2[16] ,
         bypass_rs3h_data_w2[15] , bypass_rs3h_data_w2[14] ,
         bypass_rs3h_data_w2[13] , bypass_rs3h_data_w2[12] ,
         bypass_rs3h_data_w2[11] , bypass_rs3h_data_w2[10] ,
         bypass_rs3h_data_w2[9] , bypass_rs3h_data_w2[8] ,
         bypass_rs3h_data_w2[7] , bypass_rs3h_data_w2[6] ,
         bypass_rs3h_data_w2[5] , bypass_rs3h_data_w2[4] ,
         bypass_rs3h_data_w2[3] , bypass_rs3h_data_w2[2] ,
         bypass_rs3h_data_w2[1] , bypass_rs3h_data_w2[0] ,
         bypass_rs3_data_w2[63] , bypass_rs3_data_w2[62] ,
         bypass_rs3_data_w2[61] , bypass_rs3_data_w2[60] ,
         bypass_rs3_data_w2[59] , bypass_rs3_data_w2[58] ,
         bypass_rs3_data_w2[57] , bypass_rs3_data_w2[56] ,
         bypass_rs3_data_w2[55] , bypass_rs3_data_w2[54] ,
         bypass_rs3_data_w2[53] , bypass_rs3_data_w2[52] ,
         bypass_rs3_data_w2[51] , bypass_rs3_data_w2[50] ,
         bypass_rs3_data_w2[49] , bypass_rs3_data_w2[48] ,
         bypass_rs3_data_w2[47] , bypass_rs3_data_w2[46] ,
         bypass_rs3_data_w2[45] , bypass_rs3_data_w2[44] ,
         bypass_rs3_data_w2[43] , bypass_rs3_data_w2[42] ,
         bypass_rs3_data_w2[41] , bypass_rs3_data_w2[40] ,
         bypass_rs3_data_w2[39] , bypass_rs3_data_w2[38] ,
         bypass_rs3_data_w2[37] , bypass_rs3_data_w2[36] ,
         bypass_rs3_data_w2[35] , bypass_rs3_data_w2[34] ,
         bypass_rs3_data_w2[33] , bypass_rs3_data_w2[32] ,
         bypass_rs3_data_w2[31] , bypass_rs3_data_w2[30] ,
         bypass_rs3_data_w2[29] , bypass_rs3_data_w2[28] ,
         bypass_rs3_data_w2[27] , bypass_rs3_data_w2[26] ,
         bypass_rs3_data_w2[25] , bypass_rs3_data_w2[24] ,
         bypass_rs3_data_w2[23] , bypass_rs3_data_w2[22] ,
         bypass_rs3_data_w2[21] , bypass_rs3_data_w2[20] ,
         bypass_rs3_data_w2[19] , bypass_rs3_data_w2[18] ,
         bypass_rs3_data_w2[17] , bypass_rs3_data_w2[16] ,
         bypass_rs3_data_w2[15] , bypass_rs3_data_w2[14] ,
         bypass_rs3_data_w2[13] , bypass_rs3_data_w2[12] ,
         bypass_rs3_data_w2[11] , bypass_rs3_data_w2[10] ,
         bypass_rs3_data_w2[9] , bypass_rs3_data_w2[8] ,
         bypass_rs3_data_w2[7] , bypass_rs3_data_w2[6] ,
         bypass_rs3_data_w2[5] , bypass_rs3_data_w2[4] ,
         bypass_rs3_data_w2[3] , bypass_rs3_data_w2[2] ,
         bypass_rs3_data_w2[1] , bypass_rs3_data_w2[0] ,
         bypass_rs2_data_w2[63] , bypass_rs2_data_w2[62] ,
         bypass_rs2_data_w2[61] , bypass_rs2_data_w2[60] ,
         bypass_rs2_data_w2[59] , bypass_rs2_data_w2[58] ,
         bypass_rs2_data_w2[57] , bypass_rs2_data_w2[56] ,
         bypass_rs2_data_w2[55] , bypass_rs2_data_w2[54] ,
         bypass_rs2_data_w2[53] , bypass_rs2_data_w2[52] ,
         bypass_rs2_data_w2[51] , bypass_rs2_data_w2[50] ,
         bypass_rs2_data_w2[49] , bypass_rs2_data_w2[48] ,
         bypass_rs2_data_w2[47] , bypass_rs2_data_w2[46] ,
         bypass_rs2_data_w2[45] , bypass_rs2_data_w2[44] ,
         bypass_rs2_data_w2[43] , bypass_rs2_data_w2[42] ,
         bypass_rs2_data_w2[41] , bypass_rs2_data_w2[40] ,
         bypass_rs2_data_w2[39] , bypass_rs2_data_w2[38] ,
         bypass_rs2_data_w2[37] , bypass_rs2_data_w2[36] ,
         bypass_rs2_data_w2[35] , bypass_rs2_data_w2[34] ,
         bypass_rs2_data_w2[33] , bypass_rs2_data_w2[32] ,
         bypass_rs2_data_w2[31] , bypass_rs2_data_w2[30] ,
         bypass_rs2_data_w2[29] , bypass_rs2_data_w2[28] ,
         bypass_rs2_data_w2[27] , bypass_rs2_data_w2[26] ,
         bypass_rs2_data_w2[25] , bypass_rs2_data_w2[24] ,
         bypass_rs2_data_w2[23] , bypass_rs2_data_w2[22] ,
         bypass_rs2_data_w2[21] , bypass_rs2_data_w2[20] ,
         bypass_rs2_data_w2[19] , bypass_rs2_data_w2[18] ,
         bypass_rs2_data_w2[17] , bypass_rs2_data_w2[16] ,
         bypass_rs2_data_w2[15] , bypass_rs2_data_w2[14] ,
         bypass_rs2_data_w2[13] , bypass_rs2_data_w2[12] ,
         bypass_rs2_data_w2[11] , bypass_rs2_data_w2[10] ,
         bypass_rs2_data_w2[9] , bypass_rs2_data_w2[8] ,
         bypass_rs2_data_w2[7] , bypass_rs2_data_w2[6] ,
         bypass_rs2_data_w2[5] , bypass_rs2_data_w2[4] ,
         bypass_rs2_data_w2[3] , bypass_rs2_data_w2[2] ,
         bypass_rs2_data_w2[1] , bypass_rs2_data_w2[0] ,
         bypass_rs1_data_w2[0] , bypass_rs1_data_w2[1] ,
         bypass_rs1_data_w2[2] , bypass_rs1_data_w2[3] ,
         bypass_rs1_data_w2[4] , bypass_rs1_data_w2[5] ,
         bypass_rs1_data_w2[6] , bypass_rs1_data_w2[7] ,
         bypass_rs1_data_w2[8] , bypass_rs1_data_w2[9] ,
         bypass_rs1_data_w2[10] , bypass_rs1_data_w2[11] ,
         bypass_rs1_data_w2[12] , bypass_rs1_data_w2[13] ,
         bypass_rs1_data_w2[14] , bypass_rs1_data_w2[15] ,
         bypass_rs1_data_w2[16] , bypass_rs1_data_w2[17] ,
         bypass_rs1_data_w2[18] , bypass_rs1_data_w2[19] ,
         bypass_rs1_data_w2[20] , bypass_rs1_data_w2[21] ,
         bypass_rs1_data_w2[22] , bypass_rs1_data_w2[23] ,
         bypass_rs1_data_w2[24] , bypass_rs1_data_w2[25] ,
         bypass_rs1_data_w2[26] , bypass_rs1_data_w2[27] ,
         bypass_rs1_data_w2[28] , bypass_rs1_data_w2[29] ,
         bypass_rs1_data_w2[30] , bypass_rs1_data_w2[31] ,
         bypass_rs1_data_w2[32] , bypass_rs1_data_w2[33] ,
         bypass_rs1_data_w2[34] , bypass_rs1_data_w2[35] ,
         bypass_rs1_data_w2[36] , bypass_rs1_data_w2[37] ,
         bypass_rs1_data_w2[38] , bypass_rs1_data_w2[39] ,
         bypass_rs1_data_w2[40] , bypass_rs1_data_w2[41] ,
         bypass_rs1_data_w2[42] , bypass_rs1_data_w2[43] ,
         bypass_rs1_data_w2[44] , bypass_rs1_data_w2[45] ,
         bypass_rs1_data_w2[46] , bypass_rs1_data_w2[47] ,
         bypass_rs1_data_w2[48] , bypass_rs1_data_w2[49] ,
         bypass_rs1_data_w2[50] , bypass_rs1_data_w2[51] ,
         bypass_rs1_data_w2[52] , bypass_rs1_data_w2[53] ,
         bypass_rs1_data_w2[54] , bypass_rs1_data_w2[55] ,
         bypass_rs1_data_w2[56] , bypass_rs1_data_w2[57] ,
         bypass_rs1_data_w2[58] , bypass_rs1_data_w2[59] ,
         bypass_rs1_data_w2[60] , bypass_rs1_data_w2[61] ,
         bypass_rs1_data_w2[62] , bypass_rs1_data_w2[63] ,
         bypass_byp_alu_rcc_data_d[63] , bypass_byp_alu_rcc_data_d[62] ,
         bypass_byp_alu_rcc_data_d[61] , bypass_byp_alu_rcc_data_d[60] ,
         bypass_byp_alu_rcc_data_d[59] , bypass_byp_alu_rcc_data_d[58] ,
         bypass_byp_alu_rcc_data_d[57] , bypass_byp_alu_rcc_data_d[56] ,
         bypass_byp_alu_rcc_data_d[55] , bypass_byp_alu_rcc_data_d[54] ,
         bypass_byp_alu_rcc_data_d[53] , bypass_byp_alu_rcc_data_d[52] ,
         bypass_byp_alu_rcc_data_d[51] , bypass_byp_alu_rcc_data_d[50] ,
         bypass_byp_alu_rcc_data_d[49] , bypass_byp_alu_rcc_data_d[48] ,
         bypass_byp_alu_rcc_data_d[47] , bypass_byp_alu_rcc_data_d[46] ,
         bypass_byp_alu_rcc_data_d[45] , bypass_byp_alu_rcc_data_d[44] ,
         bypass_byp_alu_rcc_data_d[43] , bypass_byp_alu_rcc_data_d[42] ,
         bypass_byp_alu_rcc_data_d[41] , bypass_byp_alu_rcc_data_d[40] ,
         bypass_byp_alu_rcc_data_d[39] , bypass_byp_alu_rcc_data_d[38] ,
         bypass_byp_alu_rcc_data_d[37] , bypass_byp_alu_rcc_data_d[36] ,
         bypass_byp_alu_rcc_data_d[35] , bypass_byp_alu_rcc_data_d[34] ,
         bypass_byp_alu_rcc_data_d[33] , bypass_byp_alu_rcc_data_d[32] ,
         bypass_byp_alu_rcc_data_d[31] , bypass_byp_alu_rcc_data_d[30] ,
         bypass_byp_alu_rcc_data_d[29] , bypass_byp_alu_rcc_data_d[28] ,
         bypass_byp_alu_rcc_data_d[27] , bypass_byp_alu_rcc_data_d[26] ,
         bypass_byp_alu_rcc_data_d[25] , bypass_byp_alu_rcc_data_d[24] ,
         bypass_byp_alu_rcc_data_d[23] , bypass_byp_alu_rcc_data_d[22] ,
         bypass_byp_alu_rcc_data_d[21] , bypass_byp_alu_rcc_data_d[20] ,
         bypass_byp_alu_rcc_data_d[19] , bypass_byp_alu_rcc_data_d[18] ,
         bypass_byp_alu_rcc_data_d[17] , bypass_byp_alu_rcc_data_d[16] ,
         bypass_byp_alu_rcc_data_d[15] , bypass_byp_alu_rcc_data_d[14] ,
         bypass_byp_alu_rcc_data_d[13] , bypass_byp_alu_rcc_data_d[12] ,
         bypass_byp_alu_rcc_data_d[11] , bypass_byp_alu_rcc_data_d[10] ,
         bypass_byp_alu_rcc_data_d[9] , bypass_byp_alu_rcc_data_d[8] ,
         bypass_byp_alu_rcc_data_d[7] , bypass_byp_alu_rcc_data_d[6] ,
         bypass_byp_alu_rcc_data_d[5] , bypass_byp_alu_rcc_data_d[4] ,
         bypass_byp_alu_rcc_data_d[3] , bypass_byp_alu_rcc_data_d[2] ,
         bypass_byp_alu_rcc_data_d[1] , bypass_byp_alu_rcc_data_d[0] ,
         bypass_rs3h_data_e[31] , bypass_rs3h_data_e[30] ,
         bypass_rs3h_data_e[29] , bypass_rs3h_data_e[28] ,
         bypass_rs3h_data_e[27] , bypass_rs3h_data_e[26] ,
         bypass_rs3h_data_e[25] , bypass_rs3h_data_e[24] ,
         bypass_rs3h_data_e[23] , bypass_rs3h_data_e[22] ,
         bypass_rs3h_data_e[21] , bypass_rs3h_data_e[20] ,
         bypass_rs3h_data_e[19] , bypass_rs3h_data_e[18] ,
         bypass_rs3h_data_e[17] , bypass_rs3h_data_e[16] ,
         bypass_rs3h_data_e[15] , bypass_rs3h_data_e[14] ,
         bypass_rs3h_data_e[13] , bypass_rs3h_data_e[12] ,
         bypass_rs3h_data_e[11] , bypass_rs3h_data_e[10] ,
         bypass_rs3h_data_e[9] , bypass_rs3h_data_e[8] ,
         bypass_rs3h_data_e[7] , bypass_rs3h_data_e[6] ,
         bypass_rs3h_data_e[5] , bypass_rs3h_data_e[4] ,
         bypass_rs3h_data_e[3] , bypass_rs3h_data_e[2] ,
         bypass_rs3h_data_e[1] , bypass_rs3h_data_e[0] ,
         bypass_rs3h_data_d[31] , bypass_rs3h_data_d[30] ,
         bypass_rs3h_data_d[29] , bypass_rs3h_data_d[28] ,
         bypass_rs3h_data_d[27] , bypass_rs3h_data_d[26] ,
         bypass_rs3h_data_d[25] , bypass_rs3h_data_d[24] ,
         bypass_rs3h_data_d[23] , bypass_rs3h_data_d[22] ,
         bypass_rs3h_data_d[21] , bypass_rs3h_data_d[20] ,
         bypass_rs3h_data_d[19] , bypass_rs3h_data_d[18] ,
         bypass_rs3h_data_d[17] , bypass_rs3h_data_d[16] ,
         bypass_rs3h_data_d[15] , bypass_rs3h_data_d[14] ,
         bypass_rs3h_data_d[13] , bypass_rs3h_data_d[12] ,
         bypass_rs3h_data_d[11] , bypass_rs3h_data_d[10] ,
         bypass_rs3h_data_d[9] , bypass_rs3h_data_d[8] ,
         bypass_rs3h_data_d[7] , bypass_rs3h_data_d[6] ,
         bypass_rs3h_data_d[5] , bypass_rs3h_data_d[4] ,
         bypass_rs3h_data_d[3] , bypass_rs3h_data_d[2] ,
         bypass_rs3h_data_d[1] , bypass_rs3h_data_d[0] ,
         bypass_rs3_data_d[63] , bypass_rs3_data_d[62] ,
         bypass_rs3_data_d[61] , bypass_rs3_data_d[60] ,
         bypass_rs3_data_d[59] , bypass_rs3_data_d[58] ,
         bypass_rs3_data_d[57] , bypass_rs3_data_d[56] ,
         bypass_rs3_data_d[55] , bypass_rs3_data_d[54] ,
         bypass_rs3_data_d[53] , bypass_rs3_data_d[52] ,
         bypass_rs3_data_d[51] , bypass_rs3_data_d[50] ,
         bypass_rs3_data_d[49] , bypass_rs3_data_d[48] ,
         bypass_rs3_data_d[47] , bypass_rs3_data_d[46] ,
         bypass_rs3_data_d[45] , bypass_rs3_data_d[44] ,
         bypass_rs3_data_d[43] , bypass_rs3_data_d[42] ,
         bypass_rs3_data_d[41] , bypass_rs3_data_d[40] ,
         bypass_rs3_data_d[39] , bypass_rs3_data_d[38] ,
         bypass_rs3_data_d[37] , bypass_rs3_data_d[36] ,
         bypass_rs3_data_d[35] , bypass_rs3_data_d[34] ,
         bypass_rs3_data_d[33] , bypass_rs3_data_d[32] ,
         bypass_rs3_data_d[31] , bypass_rs3_data_d[30] ,
         bypass_rs3_data_d[29] , bypass_rs3_data_d[28] ,
         bypass_rs3_data_d[27] , bypass_rs3_data_d[26] ,
         bypass_rs3_data_d[25] , bypass_rs3_data_d[24] ,
         bypass_rs3_data_d[23] , bypass_rs3_data_d[22] ,
         bypass_rs3_data_d[21] , bypass_rs3_data_d[20] ,
         bypass_rs3_data_d[19] , bypass_rs3_data_d[18] ,
         bypass_rs3_data_d[17] , bypass_rs3_data_d[16] ,
         bypass_rs3_data_d[15] , bypass_rs3_data_d[14] ,
         bypass_rs3_data_d[13] , bypass_rs3_data_d[12] ,
         bypass_rs3_data_d[11] , bypass_rs3_data_d[10] ,
         bypass_rs3_data_d[9] , bypass_rs3_data_d[8] ,
         bypass_rs3_data_d[7] , bypass_rs3_data_d[6] ,
         bypass_rs3_data_d[5] , bypass_rs3_data_d[4] ,
         bypass_rs3_data_d[3] , bypass_rs3_data_d[2] ,
         bypass_rs3_data_d[1] , bypass_rs3_data_d[0] ,
         bypass_byp_alu_rs2_data_d[63] , bypass_byp_alu_rs2_data_d[62] ,
         bypass_byp_alu_rs2_data_d[61] , bypass_byp_alu_rs2_data_d[60] ,
         bypass_byp_alu_rs2_data_d[59] , bypass_byp_alu_rs2_data_d[58] ,
         bypass_byp_alu_rs2_data_d[57] , bypass_byp_alu_rs2_data_d[56] ,
         bypass_byp_alu_rs2_data_d[55] , bypass_byp_alu_rs2_data_d[54] ,
         bypass_byp_alu_rs2_data_d[53] , bypass_byp_alu_rs2_data_d[52] ,
         bypass_byp_alu_rs2_data_d[51] , bypass_byp_alu_rs2_data_d[50] ,
         bypass_byp_alu_rs2_data_d[49] , bypass_byp_alu_rs2_data_d[48] ,
         bypass_byp_alu_rs2_data_d[47] , bypass_byp_alu_rs2_data_d[46] ,
         bypass_byp_alu_rs2_data_d[45] , bypass_byp_alu_rs2_data_d[44] ,
         bypass_byp_alu_rs2_data_d[43] , bypass_byp_alu_rs2_data_d[42] ,
         bypass_byp_alu_rs2_data_d[41] , bypass_byp_alu_rs2_data_d[40] ,
         bypass_byp_alu_rs2_data_d[39] , bypass_byp_alu_rs2_data_d[38] ,
         bypass_byp_alu_rs2_data_d[37] , bypass_byp_alu_rs2_data_d[36] ,
         bypass_byp_alu_rs2_data_d[35] , bypass_byp_alu_rs2_data_d[34] ,
         bypass_byp_alu_rs2_data_d[33] , bypass_byp_alu_rs2_data_d[32] ,
         bypass_byp_alu_rs2_data_d[31] , bypass_byp_alu_rs2_data_d[30] ,
         bypass_byp_alu_rs2_data_d[29] , bypass_byp_alu_rs2_data_d[28] ,
         bypass_byp_alu_rs2_data_d[27] , bypass_byp_alu_rs2_data_d[26] ,
         bypass_byp_alu_rs2_data_d[25] , bypass_byp_alu_rs2_data_d[24] ,
         bypass_byp_alu_rs2_data_d[23] , bypass_byp_alu_rs2_data_d[22] ,
         bypass_byp_alu_rs2_data_d[21] , bypass_byp_alu_rs2_data_d[20] ,
         bypass_byp_alu_rs2_data_d[19] , bypass_byp_alu_rs2_data_d[18] ,
         bypass_byp_alu_rs2_data_d[17] , bypass_byp_alu_rs2_data_d[16] ,
         bypass_byp_alu_rs2_data_d[15] , bypass_byp_alu_rs2_data_d[14] ,
         bypass_byp_alu_rs2_data_d[13] , bypass_byp_alu_rs2_data_d[12] ,
         bypass_byp_alu_rs2_data_d[11] , bypass_byp_alu_rs2_data_d[10] ,
         bypass_byp_alu_rs2_data_d[9] , bypass_byp_alu_rs2_data_d[8] ,
         bypass_byp_alu_rs2_data_d[7] , bypass_byp_alu_rs2_data_d[6] ,
         bypass_byp_alu_rs2_data_d[5] , bypass_byp_alu_rs2_data_d[4] ,
         bypass_byp_alu_rs2_data_d[3] , bypass_byp_alu_rs2_data_d[2] ,
         bypass_byp_alu_rs2_data_d[1] , bypass_byp_alu_rs2_data_d[0] ,
         bypass_byp_alu_rs1_data_d[63] , bypass_byp_alu_rs1_data_d[62] ,
         bypass_byp_alu_rs1_data_d[61] , bypass_byp_alu_rs1_data_d[60] ,
         bypass_byp_alu_rs1_data_d[59] , bypass_byp_alu_rs1_data_d[58] ,
         bypass_byp_alu_rs1_data_d[57] , bypass_byp_alu_rs1_data_d[56] ,
         bypass_byp_alu_rs1_data_d[55] , bypass_byp_alu_rs1_data_d[54] ,
         bypass_byp_alu_rs1_data_d[53] , bypass_byp_alu_rs1_data_d[52] ,
         bypass_byp_alu_rs1_data_d[51] , bypass_byp_alu_rs1_data_d[50] ,
         bypass_byp_alu_rs1_data_d[49] , bypass_byp_alu_rs1_data_d[48] ,
         bypass_byp_alu_rs1_data_d[47] , bypass_byp_alu_rs1_data_d[46] ,
         bypass_byp_alu_rs1_data_d[45] , bypass_byp_alu_rs1_data_d[44] ,
         bypass_byp_alu_rs1_data_d[43] , bypass_byp_alu_rs1_data_d[42] ,
         bypass_byp_alu_rs1_data_d[41] , bypass_byp_alu_rs1_data_d[40] ,
         bypass_byp_alu_rs1_data_d[39] , bypass_byp_alu_rs1_data_d[38] ,
         bypass_byp_alu_rs1_data_d[37] , bypass_byp_alu_rs1_data_d[36] ,
         bypass_byp_alu_rs1_data_d[35] , bypass_byp_alu_rs1_data_d[34] ,
         bypass_byp_alu_rs1_data_d[33] , bypass_byp_alu_rs1_data_d[32] ,
         bypass_byp_alu_rs1_data_d[31] , bypass_byp_alu_rs1_data_d[30] ,
         bypass_byp_alu_rs1_data_d[29] , bypass_byp_alu_rs1_data_d[28] ,
         bypass_byp_alu_rs1_data_d[27] , bypass_byp_alu_rs1_data_d[26] ,
         bypass_byp_alu_rs1_data_d[25] , bypass_byp_alu_rs1_data_d[24] ,
         bypass_byp_alu_rs1_data_d[23] , bypass_byp_alu_rs1_data_d[22] ,
         bypass_byp_alu_rs1_data_d[21] , bypass_byp_alu_rs1_data_d[20] ,
         bypass_byp_alu_rs1_data_d[19] , bypass_byp_alu_rs1_data_d[18] ,
         bypass_byp_alu_rs1_data_d[17] , bypass_byp_alu_rs1_data_d[16] ,
         bypass_byp_alu_rs1_data_d[15] , bypass_byp_alu_rs1_data_d[14] ,
         bypass_byp_alu_rs1_data_d[13] , bypass_byp_alu_rs1_data_d[12] ,
         bypass_byp_alu_rs1_data_d[11] , bypass_byp_alu_rs1_data_d[10] ,
         bypass_byp_alu_rs1_data_d[9] , bypass_byp_alu_rs1_data_d[8] ,
         bypass_byp_alu_rs1_data_d[7] , bypass_byp_alu_rs1_data_d[6] ,
         bypass_byp_alu_rs1_data_d[5] , bypass_byp_alu_rs1_data_d[4] ,
         bypass_byp_alu_rs1_data_d[3] , bypass_byp_alu_rs1_data_d[2] ,
         bypass_byp_alu_rs1_data_d[1] , bypass_byp_alu_rs1_data_d[0] ,
         bypass_rd_data_g[0] , bypass_rd_data_g[1] , bypass_rd_data_g[2] ,
         bypass_rd_data_g[3] , bypass_rd_data_g[4] , bypass_rd_data_g[5] ,
         bypass_rd_data_g[6] , bypass_rd_data_g[7] , bypass_rd_data_g[8] ,
         bypass_rd_data_g[9] , bypass_rd_data_g[10] , bypass_rd_data_g[11] ,
         bypass_rd_data_g[12] , bypass_rd_data_g[13] ,
         bypass_rd_data_g[14] , bypass_rd_data_g[15] ,
         bypass_rd_data_g[16] , bypass_rd_data_g[17] ,
         bypass_rd_data_g[18] , bypass_rd_data_g[19] ,
         bypass_rd_data_g[20] , bypass_rd_data_g[21] ,
         bypass_rd_data_g[22] , bypass_rd_data_g[23] ,
         bypass_rd_data_g[24] , bypass_rd_data_g[25] ,
         bypass_rd_data_g[26] , bypass_rd_data_g[27] ,
         bypass_rd_data_g[28] , bypass_rd_data_g[29] ,
         bypass_rd_data_g[30] , bypass_rd_data_g[31] ,
         bypass_rd_data_g[32] , bypass_rd_data_g[33] ,
         bypass_rd_data_g[34] , bypass_rd_data_g[35] ,
         bypass_rd_data_g[36] , bypass_rd_data_g[37] ,
         bypass_rd_data_g[38] , bypass_rd_data_g[39] ,
         bypass_rd_data_g[40] , bypass_rd_data_g[41] ,
         bypass_rd_data_g[42] , bypass_rd_data_g[43] ,
         bypass_rd_data_g[44] , bypass_rd_data_g[45] ,
         bypass_rd_data_g[46] , bypass_rd_data_g[47] ,
         bypass_rd_data_g[48] , bypass_rd_data_g[49] ,
         bypass_rd_data_g[50] , bypass_rd_data_g[51] ,
         bypass_rd_data_g[52] , bypass_rd_data_g[53] ,
         bypass_rd_data_g[54] , bypass_rd_data_g[55] ,
         bypass_rd_data_g[56] , bypass_rd_data_g[57] ,
         bypass_rd_data_g[58] , bypass_rd_data_g[59] ,
         bypass_rd_data_g[60] , bypass_rd_data_g[61] ,
         bypass_rd_data_g[62] , bypass_rd_data_g[63] ,
         bypass_byp_irf_rd_data_m[0] , bypass_byp_irf_rd_data_m[1] ,
         bypass_byp_irf_rd_data_m[2] , bypass_byp_irf_rd_data_m[3] ,
         bypass_byp_irf_rd_data_m[4] , bypass_byp_irf_rd_data_m[5] ,
         bypass_byp_irf_rd_data_m[6] , bypass_byp_irf_rd_data_m[7] ,
         bypass_byp_irf_rd_data_m[8] , bypass_byp_irf_rd_data_m[9] ,
         bypass_byp_irf_rd_data_m[10] , bypass_byp_irf_rd_data_m[11] ,
         bypass_byp_irf_rd_data_m[12] , bypass_byp_irf_rd_data_m[13] ,
         bypass_byp_irf_rd_data_m[14] , bypass_byp_irf_rd_data_m[15] ,
         bypass_byp_irf_rd_data_m[16] , bypass_byp_irf_rd_data_m[17] ,
         bypass_byp_irf_rd_data_m[18] , bypass_byp_irf_rd_data_m[19] ,
         bypass_byp_irf_rd_data_m[20] , bypass_byp_irf_rd_data_m[21] ,
         bypass_byp_irf_rd_data_m[22] , bypass_byp_irf_rd_data_m[23] ,
         bypass_byp_irf_rd_data_m[24] , bypass_byp_irf_rd_data_m[25] ,
         bypass_byp_irf_rd_data_m[26] , bypass_byp_irf_rd_data_m[27] ,
         bypass_byp_irf_rd_data_m[28] , bypass_byp_irf_rd_data_m[29] ,
         bypass_byp_irf_rd_data_m[30] , bypass_byp_irf_rd_data_m[31] ,
         bypass_byp_irf_rd_data_m[32] , bypass_byp_irf_rd_data_m[33] ,
         bypass_byp_irf_rd_data_m[34] , bypass_byp_irf_rd_data_m[35] ,
         bypass_byp_irf_rd_data_m[36] , bypass_byp_irf_rd_data_m[37] ,
         bypass_byp_irf_rd_data_m[38] , bypass_byp_irf_rd_data_m[39] ,
         bypass_byp_irf_rd_data_m[40] , bypass_byp_irf_rd_data_m[41] ,
         bypass_byp_irf_rd_data_m[42] , bypass_byp_irf_rd_data_m[43] ,
         bypass_byp_irf_rd_data_m[44] , bypass_byp_irf_rd_data_m[45] ,
         bypass_byp_irf_rd_data_m[46] , bypass_byp_irf_rd_data_m[47] ,
         bypass_byp_irf_rd_data_m[48] , bypass_byp_irf_rd_data_m[49] ,
         bypass_byp_irf_rd_data_m[50] , bypass_byp_irf_rd_data_m[51] ,
         bypass_byp_irf_rd_data_m[52] , bypass_byp_irf_rd_data_m[53] ,
         bypass_byp_irf_rd_data_m[54] , bypass_byp_irf_rd_data_m[55] ,
         bypass_byp_irf_rd_data_m[56] , bypass_byp_irf_rd_data_m[57] ,
         bypass_byp_irf_rd_data_m[58] , bypass_byp_irf_rd_data_m[59] ,
         bypass_byp_irf_rd_data_m[60] , bypass_byp_irf_rd_data_m[61] ,
         bypass_byp_irf_rd_data_m[62] , bypass_byp_irf_rd_data_m[63] ,
         bypass_restore_rd_data[0] , bypass_restore_rd_data[1] ,
         bypass_restore_rd_data[2] , bypass_restore_rd_data[3] ,
         bypass_restore_rd_data[4] , bypass_restore_rd_data[5] ,
         bypass_restore_rd_data[6] , bypass_restore_rd_data[7] ,
         bypass_restore_rd_data[8] , bypass_restore_rd_data[9] ,
         bypass_restore_rd_data[10] , bypass_restore_rd_data[11] ,
         bypass_restore_rd_data[12] , bypass_restore_rd_data[13] ,
         bypass_restore_rd_data[14] , bypass_restore_rd_data[15] ,
         bypass_restore_rd_data[16] , bypass_restore_rd_data[17] ,
         bypass_restore_rd_data[18] , bypass_restore_rd_data[19] ,
         bypass_restore_rd_data[20] , bypass_restore_rd_data[21] ,
         bypass_restore_rd_data[22] , bypass_restore_rd_data[23] ,
         bypass_restore_rd_data[24] , bypass_restore_rd_data[25] ,
         bypass_restore_rd_data[26] , bypass_restore_rd_data[27] ,
         bypass_restore_rd_data[28] , bypass_restore_rd_data[29] ,
         bypass_restore_rd_data[30] , bypass_restore_rd_data[31] ,
         bypass_restore_rd_data[32] , bypass_restore_rd_data[33] ,
         bypass_restore_rd_data[34] , bypass_restore_rd_data[35] ,
         bypass_restore_rd_data[36] , bypass_restore_rd_data[37] ,
         bypass_restore_rd_data[38] , bypass_restore_rd_data[39] ,
         bypass_restore_rd_data[40] , bypass_restore_rd_data[41] ,
         bypass_restore_rd_data[42] , bypass_restore_rd_data[43] ,
         bypass_restore_rd_data[44] , bypass_restore_rd_data[45] ,
         bypass_restore_rd_data[46] , bypass_restore_rd_data[47] ,
         bypass_restore_rd_data[48] , bypass_restore_rd_data[49] ,
         bypass_restore_rd_data[50] , bypass_restore_rd_data[51] ,
         bypass_restore_rd_data[52] , bypass_restore_rd_data[53] ,
         bypass_restore_rd_data[54] , bypass_restore_rd_data[55] ,
         bypass_restore_rd_data[56] , bypass_restore_rd_data[57] ,
         bypass_restore_rd_data[58] , bypass_restore_rd_data[59] ,
         bypass_restore_rd_data[60] , bypass_restore_rd_data[61] ,
         bypass_restore_rd_data[62] , bypass_restore_rd_data[63] ,
         bypass_restore_rd_data_next[63] , bypass_restore_rd_data_next[62] ,
         bypass_restore_rd_data_next[61] , bypass_restore_rd_data_next[60] ,
         bypass_restore_rd_data_next[59] , bypass_restore_rd_data_next[58] ,
         bypass_restore_rd_data_next[57] , bypass_restore_rd_data_next[56] ,
         bypass_restore_rd_data_next[55] , bypass_restore_rd_data_next[54] ,
         bypass_restore_rd_data_next[53] , bypass_restore_rd_data_next[52] ,
         bypass_restore_rd_data_next[51] , bypass_restore_rd_data_next[50] ,
         bypass_restore_rd_data_next[49] , bypass_restore_rd_data_next[48] ,
         bypass_restore_rd_data_next[47] , bypass_restore_rd_data_next[46] ,
         bypass_restore_rd_data_next[45] , bypass_restore_rd_data_next[44] ,
         bypass_restore_rd_data_next[43] , bypass_restore_rd_data_next[42] ,
         bypass_restore_rd_data_next[41] , bypass_restore_rd_data_next[40] ,
         bypass_restore_rd_data_next[39] , bypass_restore_rd_data_next[38] ,
         bypass_restore_rd_data_next[37] , bypass_restore_rd_data_next[36] ,
         bypass_restore_rd_data_next[35] , bypass_restore_rd_data_next[34] ,
         bypass_restore_rd_data_next[33] , bypass_restore_rd_data_next[32] ,
         bypass_restore_rd_data_next[31] , bypass_restore_rd_data_next[30] ,
         bypass_restore_rd_data_next[29] , bypass_restore_rd_data_next[28] ,
         bypass_restore_rd_data_next[27] , bypass_restore_rd_data_next[26] ,
         bypass_restore_rd_data_next[25] , bypass_restore_rd_data_next[24] ,
         bypass_restore_rd_data_next[23] , bypass_restore_rd_data_next[22] ,
         bypass_restore_rd_data_next[21] , bypass_restore_rd_data_next[20] ,
         bypass_restore_rd_data_next[19] , bypass_restore_rd_data_next[18] ,
         bypass_restore_rd_data_next[17] , bypass_restore_rd_data_next[16] ,
         bypass_restore_rd_data_next[15] , bypass_restore_rd_data_next[14] ,
         bypass_restore_rd_data_next[13] , bypass_restore_rd_data_next[12] ,
         bypass_restore_rd_data_next[11] , bypass_restore_rd_data_next[10] ,
         bypass_restore_rd_data_next[9] , bypass_restore_rd_data_next[8] ,
         bypass_restore_rd_data_next[7] , bypass_restore_rd_data_next[6] ,
         bypass_restore_rd_data_next[5] , bypass_restore_rd_data_next[4] ,
         bypass_restore_rd_data_next[3] , bypass_restore_rd_data_next[2] ,
         bypass_restore_rd_data_next[1] , bypass_restore_rd_data_next[0] ,
         bypass_full_rd_data_m[63] , bypass_full_rd_data_m[62] ,
         bypass_full_rd_data_m[61] , bypass_full_rd_data_m[60] ,
         bypass_full_rd_data_m[59] , bypass_full_rd_data_m[58] ,
         bypass_full_rd_data_m[57] , bypass_full_rd_data_m[56] ,
         bypass_full_rd_data_m[55] , bypass_full_rd_data_m[54] ,
         bypass_full_rd_data_m[53] , bypass_full_rd_data_m[52] ,
         bypass_full_rd_data_m[51] , bypass_full_rd_data_m[50] ,
         bypass_full_rd_data_m[49] , bypass_full_rd_data_m[48] ,
         bypass_full_rd_data_m[47] , bypass_full_rd_data_m[46] ,
         bypass_full_rd_data_m[45] , bypass_full_rd_data_m[44] ,
         bypass_full_rd_data_m[43] , bypass_full_rd_data_m[42] ,
         bypass_full_rd_data_m[41] , bypass_full_rd_data_m[40] ,
         bypass_full_rd_data_m[39] , bypass_full_rd_data_m[38] ,
         bypass_full_rd_data_m[37] , bypass_full_rd_data_m[36] ,
         bypass_full_rd_data_m[35] , bypass_full_rd_data_m[34] ,
         bypass_full_rd_data_m[33] , bypass_full_rd_data_m[32] ,
         bypass_full_rd_data_m[31] , bypass_full_rd_data_m[30] ,
         bypass_full_rd_data_m[29] , bypass_full_rd_data_m[28] ,
         bypass_full_rd_data_m[27] , bypass_full_rd_data_m[26] ,
         bypass_full_rd_data_m[25] , bypass_full_rd_data_m[24] ,
         bypass_full_rd_data_m[23] , bypass_full_rd_data_m[22] ,
         bypass_full_rd_data_m[21] , bypass_full_rd_data_m[20] ,
         bypass_full_rd_data_m[19] , bypass_full_rd_data_m[18] ,
         bypass_full_rd_data_m[17] , bypass_full_rd_data_m[16] ,
         bypass_full_rd_data_m[15] , bypass_full_rd_data_m[14] ,
         bypass_full_rd_data_m[13] , bypass_full_rd_data_m[12] ,
         bypass_full_rd_data_m[11] , bypass_full_rd_data_m[10] ,
         bypass_full_rd_data_m[9] , bypass_full_rd_data_m[8] ,
         bypass_full_rd_data_m[7] , bypass_full_rd_data_m[6] ,
         bypass_full_rd_data_m[5] , bypass_full_rd_data_m[4] ,
         bypass_full_rd_data_m[3] , bypass_full_rd_data_m[2] ,
         bypass_full_rd_data_m[1] , bypass_full_rd_data_m[0] ,
         bypass_rd_data_e[31] , bypass_rd_data_e[30] ,
         bypass_rd_data_e[29] , bypass_rd_data_e[28] ,
         bypass_rd_data_e[27] , bypass_rd_data_e[26] ,
         bypass_rd_data_e[25] , bypass_rd_data_e[24] ,
         bypass_rd_data_e[23] , bypass_rd_data_e[22] ,
         bypass_rd_data_e[21] , bypass_rd_data_e[20] ,
         bypass_rd_data_e[19] , bypass_rd_data_e[18] ,
         bypass_rd_data_e[17] , bypass_rd_data_e[16] ,
         bypass_rd_data_e[15] , bypass_rd_data_e[14] ,
         bypass_rd_data_e[13] , bypass_rd_data_e[12] ,
         bypass_rd_data_e[11] , bypass_rd_data_e[10] , bypass_rd_data_e[9] ,
         bypass_rd_data_e[8] , bypass_rd_data_e[7] , bypass_rd_data_e[6] ,
         bypass_rd_data_e[5] , bypass_rd_data_e[4] , bypass_rd_data_e[3] ,
         bypass_rd_data_e[2] , bypass_rd_data_e[1] , bypass_rd_data_e[0] ,
         bypass_dfill_data_g2[0] , bypass_dfill_data_g2[1] ,
         bypass_dfill_data_g2[2] , bypass_dfill_data_g2[3] ,
         bypass_dfill_data_g2[4] , bypass_dfill_data_g2[5] ,
         bypass_dfill_data_g2[6] , bypass_dfill_data_g2[7] ,
         bypass_dfill_data_g2[8] , bypass_dfill_data_g2[9] ,
         bypass_dfill_data_g2[10] , bypass_dfill_data_g2[11] ,
         bypass_dfill_data_g2[12] , bypass_dfill_data_g2[13] ,
         bypass_dfill_data_g2[14] , bypass_dfill_data_g2[15] ,
         bypass_dfill_data_g2[16] , bypass_dfill_data_g2[17] ,
         bypass_dfill_data_g2[18] , bypass_dfill_data_g2[19] ,
         bypass_dfill_data_g2[20] , bypass_dfill_data_g2[21] ,
         bypass_dfill_data_g2[22] , bypass_dfill_data_g2[23] ,
         bypass_dfill_data_g2[24] , bypass_dfill_data_g2[25] ,
         bypass_dfill_data_g2[26] , bypass_dfill_data_g2[27] ,
         bypass_dfill_data_g2[28] , bypass_dfill_data_g2[29] ,
         bypass_dfill_data_g2[30] , bypass_dfill_data_g2[31] ,
         bypass_dfill_data_g2[32] , bypass_dfill_data_g2[33] ,
         bypass_dfill_data_g2[34] , bypass_dfill_data_g2[35] ,
         bypass_dfill_data_g2[36] , bypass_dfill_data_g2[37] ,
         bypass_dfill_data_g2[38] , bypass_dfill_data_g2[39] ,
         bypass_dfill_data_g2[40] , bypass_dfill_data_g2[41] ,
         bypass_dfill_data_g2[42] , bypass_dfill_data_g2[43] ,
         bypass_dfill_data_g2[44] , bypass_dfill_data_g2[45] ,
         bypass_dfill_data_g2[46] , bypass_dfill_data_g2[47] ,
         bypass_dfill_data_g2[48] , bypass_dfill_data_g2[49] ,
         bypass_dfill_data_g2[50] , bypass_dfill_data_g2[51] ,
         bypass_dfill_data_g2[52] , bypass_dfill_data_g2[53] ,
         bypass_dfill_data_g2[54] , bypass_dfill_data_g2[55] ,
         bypass_dfill_data_g2[56] , bypass_dfill_data_g2[57] ,
         bypass_dfill_data_g2[58] , bypass_dfill_data_g2[59] ,
         bypass_dfill_data_g2[60] , bypass_dfill_data_g2[61] ,
         bypass_dfill_data_g2[62] , bypass_dfill_data_g2[63] ,
         bypass_dfill_data_g[63] , bypass_dfill_data_g[62] ,
         bypass_dfill_data_g[61] , bypass_dfill_data_g[60] ,
         bypass_dfill_data_g[59] , bypass_dfill_data_g[58] ,
         bypass_dfill_data_g[57] , bypass_dfill_data_g[56] ,
         bypass_dfill_data_g[55] , bypass_dfill_data_g[54] ,
         bypass_dfill_data_g[53] , bypass_dfill_data_g[52] ,
         bypass_dfill_data_g[51] , bypass_dfill_data_g[50] ,
         bypass_dfill_data_g[49] , bypass_dfill_data_g[48] ,
         bypass_dfill_data_g[47] , bypass_dfill_data_g[46] ,
         bypass_dfill_data_g[45] , bypass_dfill_data_g[44] ,
         bypass_dfill_data_g[43] , bypass_dfill_data_g[42] ,
         bypass_dfill_data_g[41] , bypass_dfill_data_g[40] ,
         bypass_dfill_data_g[39] , bypass_dfill_data_g[38] ,
         bypass_dfill_data_g[37] , bypass_dfill_data_g[36] ,
         bypass_dfill_data_g[35] , bypass_dfill_data_g[34] ,
         bypass_dfill_data_g[33] , bypass_dfill_data_g[32] ,
         bypass_dfill_data_g[31] , bypass_dfill_data_g[30] ,
         bypass_dfill_data_g[29] , bypass_dfill_data_g[28] ,
         bypass_dfill_data_g[27] , bypass_dfill_data_g[26] ,
         bypass_dfill_data_g[25] , bypass_dfill_data_g[24] ,
         bypass_dfill_data_g[23] , bypass_dfill_data_g[22] ,
         bypass_dfill_data_g[21] , bypass_dfill_data_g[20] ,
         bypass_dfill_data_g[19] , bypass_dfill_data_g[18] ,
         bypass_dfill_data_g[17] , bypass_dfill_data_g[16] ,
         bypass_dfill_data_g[15] , bypass_dfill_data_g[14] ,
         bypass_dfill_data_g[13] , bypass_dfill_data_g[12] ,
         bypass_dfill_data_g[11] , bypass_dfill_data_g[10] ,
         bypass_dfill_data_g[9] , bypass_dfill_data_g[8] ,
         bypass_dfill_data_g[7] , bypass_dfill_data_g[6] ,
         bypass_dfill_data_g[5] , bypass_dfill_data_g[4] ,
         bypass_dfill_data_g[3] , bypass_dfill_data_g[2] ,
         bypass_dfill_data_g[1] , bypass_dfill_data_g[0] ,
         bypass_sehold_clk , ecc_error_data_m[63] , ecc_error_data_m[62] ,
         ecc_error_data_m[61] , ecc_error_data_m[60] ,
         ecc_error_data_m[59] , ecc_error_data_m[58] ,
         ecc_error_data_m[57] , ecc_error_data_m[56] ,
         ecc_error_data_m[55] , ecc_error_data_m[54] ,
         ecc_error_data_m[53] , ecc_error_data_m[52] ,
         ecc_error_data_m[51] , ecc_error_data_m[50] ,
         ecc_error_data_m[49] , ecc_error_data_m[48] ,
         ecc_error_data_m[47] , ecc_error_data_m[46] ,
         ecc_error_data_m[45] , ecc_error_data_m[44] ,
         ecc_error_data_m[43] , ecc_error_data_m[42] ,
         ecc_error_data_m[41] , ecc_error_data_m[40] ,
         ecc_error_data_m[39] , ecc_error_data_m[38] ,
         ecc_error_data_m[37] , ecc_error_data_m[36] ,
         ecc_error_data_m[35] , ecc_error_data_m[34] ,
         ecc_error_data_m[33] , ecc_error_data_m[32] ,
         ecc_error_data_m[31] , ecc_error_data_m[30] ,
         ecc_error_data_m[29] , ecc_error_data_m[28] ,
         ecc_error_data_m[27] , ecc_error_data_m[26] ,
         ecc_error_data_m[25] , ecc_error_data_m[24] ,
         ecc_error_data_m[23] , ecc_error_data_m[22] ,
         ecc_error_data_m[21] , ecc_error_data_m[20] ,
         ecc_error_data_m[19] , ecc_error_data_m[18] ,
         ecc_error_data_m[17] , ecc_error_data_m[16] ,
         ecc_error_data_m[15] , ecc_error_data_m[14] ,
         ecc_error_data_m[13] , ecc_error_data_m[12] ,
         ecc_error_data_m[11] , ecc_error_data_m[10] , ecc_error_data_m[9] ,
         ecc_error_data_m[8] , ecc_error_data_m[7] , ecc_error_data_m[6] ,
         ecc_error_data_m[5] , ecc_error_data_m[4] , ecc_error_data_m[3] ,
         ecc_error_data_m[2] , ecc_error_data_m[1] , ecc_error_data_m[0] ,
         ecc_ecc_datain_m[63] , ecc_ecc_datain_m[62] ,
         ecc_ecc_datain_m[61] , ecc_ecc_datain_m[60] ,
         ecc_ecc_datain_m[59] , ecc_ecc_datain_m[58] ,
         ecc_ecc_datain_m[57] , ecc_ecc_datain_m[56] ,
         ecc_ecc_datain_m[55] , ecc_ecc_datain_m[54] ,
         ecc_ecc_datain_m[53] , ecc_ecc_datain_m[52] ,
         ecc_ecc_datain_m[51] , ecc_ecc_datain_m[50] ,
         ecc_ecc_datain_m[49] , ecc_ecc_datain_m[48] ,
         ecc_ecc_datain_m[47] , ecc_ecc_datain_m[46] ,
         ecc_ecc_datain_m[45] , ecc_ecc_datain_m[44] ,
         ecc_ecc_datain_m[43] , ecc_ecc_datain_m[42] ,
         ecc_ecc_datain_m[41] , ecc_ecc_datain_m[40] ,
         ecc_ecc_datain_m[39] , ecc_ecc_datain_m[38] ,
         ecc_ecc_datain_m[37] , ecc_ecc_datain_m[36] ,
         ecc_ecc_datain_m[35] , ecc_ecc_datain_m[34] ,
         ecc_ecc_datain_m[33] , ecc_ecc_datain_m[32] ,
         ecc_ecc_datain_m[31] , ecc_ecc_datain_m[30] ,
         ecc_ecc_datain_m[29] , ecc_ecc_datain_m[28] ,
         ecc_ecc_datain_m[27] , ecc_ecc_datain_m[26] ,
         ecc_ecc_datain_m[25] , ecc_ecc_datain_m[24] ,
         ecc_ecc_datain_m[23] , ecc_ecc_datain_m[22] ,
         ecc_ecc_datain_m[21] , ecc_ecc_datain_m[20] ,
         ecc_ecc_datain_m[19] , ecc_ecc_datain_m[18] ,
         ecc_ecc_datain_m[17] , ecc_ecc_datain_m[16] ,
         ecc_ecc_datain_m[15] , ecc_ecc_datain_m[14] ,
         ecc_ecc_datain_m[13] , ecc_ecc_datain_m[12] ,
         ecc_ecc_datain_m[11] , ecc_ecc_datain_m[10] , ecc_ecc_datain_m[9] ,
         ecc_ecc_datain_m[8] , ecc_ecc_datain_m[7] , ecc_ecc_datain_m[6] ,
         ecc_ecc_datain_m[5] , ecc_ecc_datain_m[4] , ecc_ecc_datain_m[3] ,
         ecc_ecc_datain_m[2] , ecc_ecc_datain_m[1] , ecc_ecc_datain_m[0] ,
         ecc_err_m[6] , ecc_err_m[5] , ecc_err_m[4] , ecc_err_m[3] ,
         ecc_err_m[2] , ecc_err_m[1] , ecc_err_m[0] ,
         ecc_exu_lsu_rs3_data_m[63] , ecc_exu_lsu_rs3_data_m[62] ,
         ecc_exu_lsu_rs3_data_m[61] , ecc_exu_lsu_rs3_data_m[60] ,
         ecc_exu_lsu_rs3_data_m[59] , ecc_exu_lsu_rs3_data_m[58] ,
         ecc_exu_lsu_rs3_data_m[57] , ecc_exu_lsu_rs3_data_m[56] ,
         ecc_exu_lsu_rs3_data_m[55] , ecc_exu_lsu_rs3_data_m[54] ,
         ecc_exu_lsu_rs3_data_m[53] , ecc_exu_lsu_rs3_data_m[52] ,
         ecc_exu_lsu_rs3_data_m[51] , ecc_exu_lsu_rs3_data_m[50] ,
         ecc_exu_lsu_rs3_data_m[49] , ecc_exu_lsu_rs3_data_m[48] ,
         ecc_exu_lsu_rs3_data_m[47] , ecc_exu_lsu_rs3_data_m[46] ,
         ecc_exu_lsu_rs3_data_m[45] , ecc_exu_lsu_rs3_data_m[44] ,
         ecc_exu_lsu_rs3_data_m[43] , ecc_exu_lsu_rs3_data_m[42] ,
         ecc_exu_lsu_rs3_data_m[41] , ecc_exu_lsu_rs3_data_m[40] ,
         ecc_exu_lsu_rs3_data_m[39] , ecc_exu_lsu_rs3_data_m[38] ,
         ecc_exu_lsu_rs3_data_m[37] , ecc_exu_lsu_rs3_data_m[36] ,
         ecc_exu_lsu_rs3_data_m[35] , ecc_exu_lsu_rs3_data_m[34] ,
         ecc_exu_lsu_rs3_data_m[33] , ecc_exu_lsu_rs3_data_m[32] ,
         ecc_exu_lsu_rs3_data_m[31] , ecc_exu_lsu_rs3_data_m[30] ,
         ecc_exu_lsu_rs3_data_m[29] , ecc_exu_lsu_rs3_data_m[28] ,
         ecc_exu_lsu_rs3_data_m[27] , ecc_exu_lsu_rs3_data_m[26] ,
         ecc_exu_lsu_rs3_data_m[25] , ecc_exu_lsu_rs3_data_m[24] ,
         ecc_exu_lsu_rs3_data_m[23] , ecc_exu_lsu_rs3_data_m[22] ,
         ecc_exu_lsu_rs3_data_m[21] , ecc_exu_lsu_rs3_data_m[20] ,
         ecc_exu_lsu_rs3_data_m[19] , ecc_exu_lsu_rs3_data_m[18] ,
         ecc_exu_lsu_rs3_data_m[17] , ecc_exu_lsu_rs3_data_m[16] ,
         ecc_exu_lsu_rs3_data_m[15] , ecc_exu_lsu_rs3_data_m[14] ,
         ecc_exu_lsu_rs3_data_m[13] , ecc_exu_lsu_rs3_data_m[12] ,
         ecc_exu_lsu_rs3_data_m[11] , ecc_exu_lsu_rs3_data_m[10] ,
         ecc_exu_lsu_rs3_data_m[9] , ecc_exu_lsu_rs3_data_m[8] ,
         ecc_exu_lsu_rs3_data_m[7] , ecc_exu_lsu_rs3_data_m[6] ,
         ecc_exu_lsu_rs3_data_m[5] , ecc_exu_lsu_rs3_data_m[4] ,
         ecc_exu_lsu_rs3_data_m[3] , ecc_exu_lsu_rs3_data_m[2] ,
         ecc_exu_lsu_rs3_data_m[1] , ecc_exu_lsu_rs3_data_m[0] ,
         ecc_byp_alu_rs2_data_m[63] , ecc_byp_alu_rs2_data_m[62] ,
         ecc_byp_alu_rs2_data_m[61] , ecc_byp_alu_rs2_data_m[60] ,
         ecc_byp_alu_rs2_data_m[59] , ecc_byp_alu_rs2_data_m[58] ,
         ecc_byp_alu_rs2_data_m[57] , ecc_byp_alu_rs2_data_m[56] ,
         ecc_byp_alu_rs2_data_m[55] , ecc_byp_alu_rs2_data_m[54] ,
         ecc_byp_alu_rs2_data_m[53] , ecc_byp_alu_rs2_data_m[52] ,
         ecc_byp_alu_rs2_data_m[51] , ecc_byp_alu_rs2_data_m[50] ,
         ecc_byp_alu_rs2_data_m[49] , ecc_byp_alu_rs2_data_m[48] ,
         ecc_byp_alu_rs2_data_m[47] , ecc_byp_alu_rs2_data_m[46] ,
         ecc_byp_alu_rs2_data_m[45] , ecc_byp_alu_rs2_data_m[44] ,
         ecc_byp_alu_rs2_data_m[43] , ecc_byp_alu_rs2_data_m[42] ,
         ecc_byp_alu_rs2_data_m[41] , ecc_byp_alu_rs2_data_m[40] ,
         ecc_byp_alu_rs2_data_m[39] , ecc_byp_alu_rs2_data_m[38] ,
         ecc_byp_alu_rs2_data_m[37] , ecc_byp_alu_rs2_data_m[36] ,
         ecc_byp_alu_rs2_data_m[35] , ecc_byp_alu_rs2_data_m[34] ,
         ecc_byp_alu_rs2_data_m[33] , ecc_byp_alu_rs2_data_m[32] ,
         ecc_byp_alu_rs2_data_m[31] , ecc_byp_alu_rs2_data_m[30] ,
         ecc_byp_alu_rs2_data_m[29] , ecc_byp_alu_rs2_data_m[28] ,
         ecc_byp_alu_rs2_data_m[27] , ecc_byp_alu_rs2_data_m[26] ,
         ecc_byp_alu_rs2_data_m[25] , ecc_byp_alu_rs2_data_m[24] ,
         ecc_byp_alu_rs2_data_m[23] , ecc_byp_alu_rs2_data_m[22] ,
         ecc_byp_alu_rs2_data_m[21] , ecc_byp_alu_rs2_data_m[20] ,
         ecc_byp_alu_rs2_data_m[19] , ecc_byp_alu_rs2_data_m[18] ,
         ecc_byp_alu_rs2_data_m[17] , ecc_byp_alu_rs2_data_m[16] ,
         ecc_byp_alu_rs2_data_m[15] , ecc_byp_alu_rs2_data_m[14] ,
         ecc_byp_alu_rs2_data_m[13] , ecc_byp_alu_rs2_data_m[12] ,
         ecc_byp_alu_rs2_data_m[11] , ecc_byp_alu_rs2_data_m[10] ,
         ecc_byp_alu_rs2_data_m[9] , ecc_byp_alu_rs2_data_m[8] ,
         ecc_byp_alu_rs2_data_m[7] , ecc_byp_alu_rs2_data_m[6] ,
         ecc_byp_alu_rs2_data_m[5] , ecc_byp_alu_rs2_data_m[4] ,
         ecc_byp_alu_rs2_data_m[3] , ecc_byp_alu_rs2_data_m[2] ,
         ecc_byp_alu_rs2_data_m[1] , ecc_byp_alu_rs2_data_m[0] ,
         ecc_byp_ecc_rcc_data_m[63] , ecc_byp_ecc_rcc_data_m[62] ,
         ecc_byp_ecc_rcc_data_m[61] , ecc_byp_ecc_rcc_data_m[60] ,
         ecc_byp_ecc_rcc_data_m[59] , ecc_byp_ecc_rcc_data_m[58] ,
         ecc_byp_ecc_rcc_data_m[57] , ecc_byp_ecc_rcc_data_m[56] ,
         ecc_byp_ecc_rcc_data_m[55] , ecc_byp_ecc_rcc_data_m[54] ,
         ecc_byp_ecc_rcc_data_m[53] , ecc_byp_ecc_rcc_data_m[52] ,
         ecc_byp_ecc_rcc_data_m[51] , ecc_byp_ecc_rcc_data_m[50] ,
         ecc_byp_ecc_rcc_data_m[49] , ecc_byp_ecc_rcc_data_m[48] ,
         ecc_byp_ecc_rcc_data_m[47] , ecc_byp_ecc_rcc_data_m[46] ,
         ecc_byp_ecc_rcc_data_m[45] , ecc_byp_ecc_rcc_data_m[44] ,
         ecc_byp_ecc_rcc_data_m[43] , ecc_byp_ecc_rcc_data_m[42] ,
         ecc_byp_ecc_rcc_data_m[41] , ecc_byp_ecc_rcc_data_m[40] ,
         ecc_byp_ecc_rcc_data_m[39] , ecc_byp_ecc_rcc_data_m[38] ,
         ecc_byp_ecc_rcc_data_m[37] , ecc_byp_ecc_rcc_data_m[36] ,
         ecc_byp_ecc_rcc_data_m[35] , ecc_byp_ecc_rcc_data_m[34] ,
         ecc_byp_ecc_rcc_data_m[33] , ecc_byp_ecc_rcc_data_m[32] ,
         ecc_byp_ecc_rcc_data_m[31] , ecc_byp_ecc_rcc_data_m[30] ,
         ecc_byp_ecc_rcc_data_m[29] , ecc_byp_ecc_rcc_data_m[28] ,
         ecc_byp_ecc_rcc_data_m[27] , ecc_byp_ecc_rcc_data_m[26] ,
         ecc_byp_ecc_rcc_data_m[25] , ecc_byp_ecc_rcc_data_m[24] ,
         ecc_byp_ecc_rcc_data_m[23] , ecc_byp_ecc_rcc_data_m[22] ,
         ecc_byp_ecc_rcc_data_m[21] , ecc_byp_ecc_rcc_data_m[20] ,
         ecc_byp_ecc_rcc_data_m[19] , ecc_byp_ecc_rcc_data_m[18] ,
         ecc_byp_ecc_rcc_data_m[17] , ecc_byp_ecc_rcc_data_m[16] ,
         ecc_byp_ecc_rcc_data_m[15] , ecc_byp_ecc_rcc_data_m[14] ,
         ecc_byp_ecc_rcc_data_m[13] , ecc_byp_ecc_rcc_data_m[12] ,
         ecc_byp_ecc_rcc_data_m[11] , ecc_byp_ecc_rcc_data_m[10] ,
         ecc_byp_ecc_rcc_data_m[9] , ecc_byp_ecc_rcc_data_m[8] ,
         ecc_byp_ecc_rcc_data_m[7] , ecc_byp_ecc_rcc_data_m[6] ,
         ecc_byp_ecc_rcc_data_m[5] , ecc_byp_ecc_rcc_data_m[4] ,
         ecc_byp_ecc_rcc_data_m[3] , ecc_byp_ecc_rcc_data_m[2] ,
         ecc_byp_ecc_rcc_data_m[1] , ecc_byp_ecc_rcc_data_m[0] ,
         ecc_rs3_err_m[0] , ecc_rs3_err_m[1] , ecc_rs3_err_m[2] ,
         ecc_rs3_err_m[3] , ecc_rs3_err_m[4] , ecc_rs3_err_m[5] ,
         ecc_rs3_err_m[6] , ecc_rs2_err_m[0] , ecc_rs2_err_m[1] ,
         ecc_rs2_err_m[2] , ecc_rs2_err_m[3] , ecc_rs2_err_m[4] ,
         ecc_rs2_err_m[5] , ecc_rs2_err_m[6] , ecc_rs1_err_m[0] ,
         ecc_rs1_err_m[1] , ecc_rs1_err_m[2] , ecc_rs1_err_m[3] ,
         ecc_rs1_err_m[4] , ecc_rs1_err_m[5] , ecc_rs1_err_m[6] ,
         ecc_rs3_err_e[6] , ecc_rs3_err_e[5] , ecc_rs3_err_e[4] ,
         ecc_rs3_err_e[3] , ecc_rs3_err_e[2] , ecc_rs3_err_e[1] ,
         ecc_rs3_err_e[0] , ecc_rs2_err_e[6] , ecc_rs2_err_e[5] ,
         ecc_rs2_err_e[4] , ecc_rs2_err_e[3] , ecc_rs2_err_e[2] ,
         ecc_rs2_err_e[1] , ecc_rs2_err_e[0] , ecc_rs1_err_e[6] ,
         ecc_rs1_err_e[5] , ecc_rs1_err_e[4] , ecc_rs1_err_e[3] ,
         ecc_rs1_err_e[2] , ecc_rs1_err_e[1] , ecc_rs1_err_e[0] ,
         ecc_rs3_ecc_e[7] , ecc_rs3_ecc_e[6] , ecc_rs3_ecc_e[5] ,
         ecc_rs3_ecc_e[4] , ecc_rs3_ecc_e[3] , ecc_rs3_ecc_e[2] ,
         ecc_rs3_ecc_e[1] , ecc_rs3_ecc_e[0] , ecc_rs2_ecc_e[7] ,
         ecc_rs2_ecc_e[6] , ecc_rs2_ecc_e[5] , ecc_rs2_ecc_e[4] ,
         ecc_rs2_ecc_e[3] , ecc_rs2_ecc_e[2] , ecc_rs2_ecc_e[1] ,
         ecc_rs2_ecc_e[0] , ecc_rs1_ecc_e[7] , ecc_rs1_ecc_e[6] ,
         ecc_rs1_ecc_e[5] , ecc_rs1_ecc_e[4] , ecc_rs1_ecc_e[3] ,
         ecc_rs1_ecc_e[2] , ecc_rs1_ecc_e[1] , ecc_rs1_ecc_e[0] ,
         ecl_n145 , ecl_n144 , ecl_n143 , ecl_n142 , ecl_n141 ,
         ecl_n140 , ecl_n139 , ecl_n138 , ecl_n137 , ecl_n136 ,
         ecl_n135 , ecl_n134 , ecl_n133 , ecl_n132 , ecl_n131 ,
         ecl_n130 , ecl_n129 , ecl_n127 , ecl_n125 , ecl_n124 ,
         ecl_n123 , ecl_n122 , ecl_n121 , ecl_n120 , ecl_n119 ,
         ecl_n118 , ecl_n117 , ecl_n116 , ecl_n115 , ecl_n114 ,
         ecl_n113 , ecl_n112 , ecl_n111 , ecl_n110 , ecl_n109 ,
         ecl_n108 , ecl_n107 , ecl_n106 , ecl_n105 , ecl_n104 ,
         ecl_n103 , ecl_n102 , ecl_n101 , ecl_n100 , ecl_n99 , ecl_n98 ,
         ecl_n97 , ecl_n96 , ecl_n95 , ecl_n94 , ecl_n93 , ecl_n92 ,
         ecl_n91 , ecl_n90 , ecl_n89 , ecl_n88 , ecl_n87 , ecl_n86 ,
         ecl_n85 , ecl_n84 , ecl_n83 , ecl_n82 , ecl_n81 , ecl_n80 ,
         ecl_n79 , ecl_n78 , ecl_n77 , ecl_n76 , ecl_n75 , ecl_n74 ,
         ecl_n73 , ecl_n72 , ecl_n71 , ecl_n70 , ecl_n69 , ecl_n68 ,
         ecl_n67 , ecl_n66 , ecl_n65 , ecl_n64 , ecl_n63 , ecl_n62 ,
         ecl_n61 , ecl_n60 , ecl_n59 , ecl_n58 , ecl_n57 , ecl_n56 ,
         ecl_n55 , ecl_n54 , ecl_n53 , ecl_n52 , ecl_n51 , ecl_n50 ,
         ecl_n49 , ecl_n48 , ecl_n47 , ecl_n46 , ecl_n45 , ecl_n44 ,
         ecl_n43 , ecl_mdqctl_divcntl_muldone , ecl_ecl_div_signed_div ,
         ecl_mdqctl_divcntl_reset_div , ecl_ld_thr_match_dg2 ,
         ecl_ld_thr_match_dg , ecl_eccctl_wb_rd_m[4] ,
         ecl_eccctl_wb_rd_m[3] , ecl_eccctl_wb_rd_m[2] ,
         ecl_eccctl_wb_rd_m[1] , ecl_eccctl_wb_rd_m[0] ,
         ecl_mdqctl_wb_yreg_shift_g , ecl_mdqctl_wb_yreg_wen_g ,
         ecl_mdqctl_wb_mulsetcc_g , ecl_mdqctl_wb_divsetcc_g ,
         ecl_mdqctl_wb_multhr_g[1] , ecl_mdqctl_wb_multhr_g[0] ,
         ecl_mdqctl_wb_mulrd_g[4] , ecl_mdqctl_wb_mulrd_g[3] ,
         ecl_mdqctl_wb_mulrd_g[2] , ecl_mdqctl_wb_mulrd_g[1] ,
         ecl_mdqctl_wb_mulrd_g[0] , ecl_mdqctl_wb_divthr_g[1] ,
         ecl_mdqctl_wb_divthr_g[0] , ecl_mdqctl_wb_divrd_g[4] ,
         ecl_mdqctl_wb_divrd_g[3] , ecl_mdqctl_wb_divrd_g[2] ,
         ecl_mdqctl_wb_divrd_g[1] , ecl_mdqctl_wb_divrd_g[0] ,
         ecl_divcntl_wb_req_g , ecl_wb_byplog_wen_g2 ,
         ecl_wb_byplog_rd_g2[0] , ecl_wb_byplog_rd_g2[1] ,
         ecl_wb_byplog_rd_g2[2] , ecl_wb_byplog_rd_g2[3] ,
         ecl_wb_byplog_rd_g2[4] , ecl_wb_byplog_tid_w2[0] ,
         ecl_wb_byplog_tid_w2[1] , ecl_wb_byplog_rd_w2[0] ,
         ecl_wb_byplog_rd_w2[1] , ecl_wb_byplog_rd_w2[2] ,
         ecl_wb_byplog_rd_w2[3] , ecl_wb_byplog_rd_w2[4] , ecl_bypass_w ,
         ecl_wb_eccctl_spec_wen_next , ecl_bypass_m , ecl_wb_e ,
         ecl_divcntl_ccr_cc_w2[7] , ecl_divcntl_ccr_cc_w2[6] ,
         ecl_divcntl_ccr_cc_w2[3] , ecl_divcntl_ccr_cc_w2[2] ,
         ecl_divcntl_ccr_cc_w2[1] , ecl_divcntl_ccr_cc_w2[0] ,
         ecl_wb_ccr_setcc_g , ecl_wb_ccr_wrccr_w , ecl_thr_match_de ,
         ecl_thr_match_dm , ecl_fill_trap_m , ecl_div_zero_m ,
         ecl_early_ttype_vld_m , ecl_early_ttype_m[8] ,
         ecl_early_ttype_m[7] , ecl_early_ttype_m[6] ,
         ecl_early_ttype_m[5] , ecl_early_ttype_m[4] ,
         ecl_early_ttype_m[3] , ecl_early_ttype_m[2] ,
         ecl_early_ttype_m[1] , ecl_early_ttype_m[0] ,
         ecl_early2_ttype_e[5] , ecl_early2_ttype_e[4] ,
         ecl_early2_ttype_e[2] , ecl_pick_normal_ttype ,
         ecl_pick_not_aligned , ecl_early1_ttype_e[1] ,
         ecl_early1_ttype_e[2] , ecl_early1_ttype_e[3] ,
         ecl_early1_ttype_e[4] , ecl_early1_ttype_e[5] ,
         ecl_early_ttype_vld_e , ecl_std_e , ecl_std_d ,
         ecl_ecl_exu_kill_m , ecl_kill_rml_w , ecl_kill_rml_m ,
         ecl_flush_w1 , ecl_flush_w , ecl_part_early_flush_w ,
         ecl_tlu_priv_trap_w , ecl_part_early_flush_m , ecl_thr_match_mw1 ,
         ecl_inst_vld_w1 , ecl_ifu_tlu_flush_w , ecl_perr_store_next[3] ,
         ecl_perr_store_next[2] , ecl_perr_store_next[1] ,
         ecl_perr_store_next[0] , ecl_perr_store[0] , ecl_perr_store[1] ,
         ecl_perr_store[2] , ecl_perr_store[3] , ecl_ecl_irf_tid_w[0] ,
         ecl_ecl_irf_tid_w[1] , ecl_tid_w1[0] , ecl_tid_w1[1] ,
         ecl_tid_w[0] , ecl_tid_w[1] , ecl_tid_m[0] , ecl_tid_m[1] ,
         ecl_tid_e[0] , ecl_tid_e[1] , ecl_tid_d[0] , ecl_tid_d[1] ,
         ecl_ecl_irf_rd_w[0] , ecl_ecl_irf_rd_w[1] , ecl_ecl_irf_rd_w[2] ,
         ecl_ecl_irf_rd_w[3] , ecl_ecl_irf_rd_w[4] , ecl_rd_m[0] ,
         ecl_rd_m[1] , ecl_rd_m[2] , ecl_rd_m[3] , ecl_rd_m[4] ,
         ecl_real_rd_e[4] , ecl_rd_e[0] , ecl_rd_e[1] , ecl_rd_e[2] ,
         ecl_rd_e[3] , ecl_rd_e[4] , ecl_ifu_exu_range_check_other_e ,
         ecl_ifu_exu_range_check_jlret_m , ecl_ifu_exu_range_check_other_m ,
         ecl_alu_ecl_mem_addr_invalid_m_l , ecl_valid_range_check_jlret_e ,
         ecl_addr_mask_e , ecl_misalign_addr_e ,
         ecl_ifu_exu_range_check_jlret_e , ecl_alu_icc_e[3] ,
         ecl_alu_xcc_e[3] , ecl_alu_xcc_e[2] , ecl_adder_icc[0] ,
         ecl_adder_icc[1] , ecl_adder_xcc[1] , ecl_adder_xcc[0] ,
         ecl_restore_e , ecl_save_e , ecl_rs2_data_31_m ,
         ecl_muls_rs1_31_m_l , ecl_sub_e , ecl_next_yreg_data_31 ,
         ecl_muls_e , ecl_zero_rs2_d , ecl_thr_d[0] , ecl_thr_d[1] ,
         ecl_thr_d[2] , ecl_thr_d[3] , ecl_div_ecl_yreg_0_d , ecl_cc_e_1 ,
         ecl_cc_e_3 , ecl_cancel_rs3_ecc_e , ecl_read_tlusr_m ,
         ecl_read_tlusr_e , ecl_read_ffusr_e , ecl_read_yreg_e ,
         ecl_rs3_vld_e , ecl_rs3_vld_d , ecl_rs2_vld_e , ecl_rs1_vld_e ,
         ecl_ldxa_g , ecl_ialign_m , ecl_ialign_e , ecl_ifu_exu_tagop_e ,
         ecl_ifu_exu_tv_e , ecl_sel_sum_e , ecl_enshift_e ,
         ecl_shiftop_e_0 , ecl_shiftop_e[2] , ecl_shiftop_d[2] ,
         ecl_shiftop_d[1] , ecl_shiftop_d[0] , ecl_ifu_exu_aluop_e[0] ,
         ecl_ifu_exu_aluop_e[1] , ecl_ifu_exu_aluop_e[2] , ecl_ld_tid_g[0] ,
         ecl_ld_tid_g[1] , ecl_ld_rd_g[0] , ecl_ld_rd_g[1] ,
         ecl_ld_rd_g[2] , ecl_ld_rd_g[3] , ecl_ld_rd_g[4] ,
         ecl_ifu_exu_rs3_m[4] , ecl_ifu_exu_rs3_m[3] ,
         ecl_ifu_exu_rs3_m[2] , ecl_ifu_exu_rs3_m[1] ,
         ecl_ifu_exu_rs3_m[0] , ecl_ifu_exu_rs2_m[4] ,
         ecl_ifu_exu_rs2_m[3] , ecl_ifu_exu_rs2_m[2] ,
         ecl_ifu_exu_rs2_m[1] , ecl_ifu_exu_rs2_m[0] ,
         ecl_ifu_exu_rs1_m[4] , ecl_ifu_exu_rs1_m[3] ,
         ecl_ifu_exu_rs1_m[2] , ecl_ifu_exu_rs1_m[1] ,
         ecl_ifu_exu_rs1_m[0] , ecl_ifu_exu_rs3_e[4] ,
         ecl_ifu_exu_rs3_e[3] , ecl_ifu_exu_rs3_e[2] ,
         ecl_ifu_exu_rs3_e[1] , ecl_ifu_exu_rs3_e[0] ,
         ecl_ifu_exu_rs2_e[4] , ecl_ifu_exu_rs2_e[3] ,
         ecl_ifu_exu_rs2_e[2] , ecl_ifu_exu_rs2_e[1] ,
         ecl_ifu_exu_rs2_e[0] , ecl_ifu_exu_rs1_e[4] ,
         ecl_ifu_exu_rs1_e[3] , ecl_ifu_exu_rs1_e[2] ,
         ecl_ifu_exu_rs1_e[1] , ecl_ifu_exu_rs1_e[0] ,
         ecl_ifu_exu_rs3_d[0] , ecl_ifu_exu_rs3_d[1] ,
         ecl_ifu_exu_rs3_d[2] , ecl_ifu_exu_rs3_d[3] ,
         ecl_ifu_exu_rs3_d[4] , ecl_ifu_exu_rs2_d[0] ,
         ecl_ifu_exu_rs2_d[1] , ecl_ifu_exu_rs2_d[2] ,
         ecl_ifu_exu_rs2_d[3] , ecl_ifu_exu_rs2_d[4] ,
         ecl_ifu_exu_rs1_d[0] , ecl_ifu_exu_rs1_d[1] ,
         ecl_ifu_exu_rs1_d[2] , ecl_ifu_exu_rs1_d[3] ,
         ecl_ifu_exu_rs1_d[4] , ecl_ecl_reset_l , alu_n128 , alu_n127 ,
         alu_n126 , alu_n125 , alu_n124 , alu_n123 , alu_n122 ,
         alu_n121 , alu_n120 , alu_n119 , alu_n118 , alu_n117 ,
         alu_n116 , alu_n115 , alu_n114 , alu_n113 , alu_n112 ,
         alu_n111 , alu_n110 , alu_n109 , alu_n108 , alu_n107 ,
         alu_n106 , alu_n105 , alu_n104 , alu_n103 , alu_n102 ,
         alu_n101 , alu_n100 , alu_n99 , alu_n98 , alu_n97 , alu_n96 ,
         alu_n95 , alu_n94 , alu_n93 , alu_n92 , alu_n91 , alu_n90 ,
         alu_n89 , alu_n88 , alu_n87 , alu_n86 , alu_n85 , alu_n84 ,
         alu_n83 , alu_n82 , alu_n81 , alu_n80 , alu_n79 , alu_n78 ,
         alu_n77 , alu_n76 , alu_n75 , alu_n74 , alu_n73 , alu_n72 ,
         alu_n71 , alu_n70 , alu_n69 , alu_zcomp_in[63] ,
         alu_zcomp_in[62] , alu_zcomp_in[61] , alu_zcomp_in[60] ,
         alu_zcomp_in[59] , alu_zcomp_in[58] , alu_zcomp_in[57] ,
         alu_zcomp_in[56] , alu_zcomp_in[55] , alu_zcomp_in[54] ,
         alu_zcomp_in[53] , alu_zcomp_in[52] , alu_zcomp_in[51] ,
         alu_zcomp_in[50] , alu_zcomp_in[49] , alu_zcomp_in[48] ,
         alu_zcomp_in[47] , alu_zcomp_in[46] , alu_zcomp_in[45] ,
         alu_zcomp_in[44] , alu_zcomp_in[43] , alu_zcomp_in[42] ,
         alu_zcomp_in[41] , alu_zcomp_in[40] , alu_zcomp_in[39] ,
         alu_zcomp_in[38] , alu_zcomp_in[37] , alu_zcomp_in[36] ,
         alu_zcomp_in[35] , alu_zcomp_in[34] , alu_zcomp_in[33] ,
         alu_zcomp_in[32] , alu_zcomp_in[31] , alu_zcomp_in[30] ,
         alu_zcomp_in[29] , alu_zcomp_in[28] , alu_zcomp_in[27] ,
         alu_zcomp_in[26] , alu_zcomp_in[25] , alu_zcomp_in[24] ,
         alu_zcomp_in[23] , alu_zcomp_in[22] , alu_zcomp_in[21] ,
         alu_zcomp_in[20] , alu_zcomp_in[19] , alu_zcomp_in[18] ,
         alu_zcomp_in[17] , alu_zcomp_in[16] , alu_zcomp_in[15] ,
         alu_zcomp_in[14] , alu_zcomp_in[13] , alu_zcomp_in[12] ,
         alu_zcomp_in[11] , alu_zcomp_in[10] , alu_zcomp_in[9] ,
         alu_zcomp_in[8] , alu_zcomp_in[7] , alu_zcomp_in[6] ,
         alu_zcomp_in[5] , alu_zcomp_in[4] , alu_zcomp_in[3] ,
         alu_zcomp_in[2] , alu_zcomp_in[1] , alu_zcomp_in[0] ,
         alu_logic_out_0 , alu_logic_out_1 , alu_logic_out_2 ,
         alu_logic_out_3 , alu_logic_out_4 , alu_logic_out_5 ,
         alu_logic_out_6 , alu_logic_out_7 , alu_logic_out_8 ,
         alu_logic_out_9 , alu_logic_out_10 , alu_logic_out_11 ,
         alu_logic_out_12 , alu_logic_out_13 , alu_logic_out_14 ,
         alu_logic_out_15 , alu_logic_out_16 , alu_logic_out_17 ,
         alu_logic_out_18 , alu_logic_out_19 , alu_logic_out_20 ,
         alu_logic_out_21 , alu_logic_out_22 , alu_logic_out_23 ,
         alu_logic_out_24 , alu_logic_out_25 , alu_logic_out_26 ,
         alu_logic_out_27 , alu_logic_out_28 , alu_logic_out_29 ,
         alu_logic_out_30 , alu_logic_out[32] , alu_logic_out[33] ,
         alu_logic_out[34] , alu_logic_out[35] , alu_logic_out[36] ,
         alu_logic_out[37] , alu_logic_out[38] , alu_logic_out[39] ,
         alu_logic_out[40] , alu_logic_out[41] , alu_logic_out[42] ,
         alu_logic_out[43] , alu_logic_out[44] , alu_logic_out[45] ,
         alu_logic_out[46] , alu_logic_out[47] , alu_logic_out[48] ,
         alu_logic_out[49] , alu_logic_out[50] , alu_logic_out[51] ,
         alu_logic_out[52] , alu_logic_out[53] , alu_logic_out[54] ,
         alu_logic_out[55] , alu_logic_out[56] , alu_logic_out[57] ,
         alu_logic_out[58] , alu_logic_out[59] , alu_logic_out[60] ,
         alu_logic_out[61] , alu_logic_out[62] , alu_invert_e ,
         alu_spr_out[63] , alu_spr_out[62] , alu_spr_out[61] ,
         alu_spr_out[60] , alu_spr_out[59] , alu_spr_out[58] ,
         alu_spr_out[57] , alu_spr_out[56] , alu_spr_out[55] ,
         alu_spr_out[54] , alu_spr_out[53] , alu_spr_out[52] ,
         alu_spr_out[51] , alu_spr_out[50] , alu_spr_out[49] ,
         alu_spr_out[48] , alu_spr_out[47] , alu_spr_out[46] ,
         alu_spr_out[45] , alu_spr_out[44] , alu_spr_out[43] ,
         alu_spr_out[42] , alu_spr_out[41] , alu_spr_out[40] ,
         alu_spr_out[39] , alu_spr_out[38] , alu_spr_out[37] ,
         alu_spr_out[36] , alu_spr_out[35] , alu_spr_out[34] ,
         alu_spr_out[33] , alu_spr_out[32] , alu_spr_out[31] ,
         alu_spr_out[30] , alu_spr_out[29] , alu_spr_out[28] ,
         alu_spr_out[27] , alu_spr_out[26] , alu_spr_out[25] ,
         alu_spr_out[24] , alu_spr_out[23] , alu_spr_out[22] ,
         alu_spr_out[21] , alu_spr_out[20] , alu_spr_out[19] ,
         alu_spr_out[18] , alu_spr_out[17] , alu_spr_out[16] ,
         alu_spr_out[15] , alu_spr_out[14] , alu_spr_out[13] ,
         alu_spr_out[12] , alu_spr_out[11] , alu_spr_out[10] ,
         alu_spr_out[9] , alu_spr_out[8] , alu_spr_out[7] ,
         alu_spr_out[6] , alu_spr_out[5] , alu_spr_out[4] ,
         alu_spr_out[3] , alu_spr_out[2] , alu_spr_out[1] ,
         alu_spr_out[0] , alu_adder_out[48] , alu_adder_out[49] ,
         alu_adder_out[50] , alu_adder_out[51] , alu_adder_out[52] ,
         alu_adder_out[53] , alu_adder_out[54] , alu_adder_out[55] ,
         alu_adder_out[56] , alu_adder_out[57] , alu_adder_out[58] ,
         alu_adder_out[59] , alu_adder_out[60] , alu_adder_out[61] ,
         alu_adder_out[62] , alu_va_e[63] , alu_va_e[62] , alu_va_e[61] ,
         alu_va_e[60] , alu_va_e[59] , alu_va_e[58] , alu_va_e[57] ,
         alu_va_e[56] , alu_va_e[55] , alu_va_e[54] , alu_va_e[53] ,
         alu_va_e[52] , alu_va_e[51] , alu_va_e[50] , alu_va_e[49] ,
         alu_va_e[48] , shft_n5 , shft_lshift4_b1[8] , shft_lshift4_b1[9] ,
         shft_lshift4_b1[10] , shft_lshift4_b1[11] , shft_lshift4_b1[12] ,
         shft_lshift4_b1[13] , shft_lshift4_b1[14] , shft_lshift4_b1[15] ,
         shft_lshift4_b1[16] , shft_lshift4_b1[17] , shft_lshift4_b1[18] ,
         shft_lshift4_b1[19] , shft_lshift4_b1[20] , shft_lshift4_b1[21] ,
         shft_lshift4_b1[22] , shft_lshift4_b1[23] , shft_lshift4_b1[24] ,
         shft_lshift4_b1[25] , shft_lshift4_b1[26] , shft_lshift4_b1[27] ,
         shft_lshift4_b1[28] , shft_lshift4_b1[29] , shft_lshift4_b1[30] ,
         shft_lshift4_b1[31] , shft_lshift4_b1[32] , shft_lshift4_b1[33] ,
         shft_lshift4_b1[34] , shft_lshift4_b1[35] , shft_lshift4_b1[36] ,
         shft_lshift4_b1[37] , shft_lshift4_b1[38] , shft_lshift4_b1[39] ,
         shft_lshift4_b1[40] , shft_lshift4_b1[41] , shft_lshift4_b1[42] ,
         shft_lshift4_b1[43] , shft_lshift4_b1[44] , shft_lshift4_b1[45] ,
         shft_lshift4_b1[46] , shft_lshift4_b1[47] , shft_lshift4_b1[48] ,
         shft_lshift4_b1[49] , shft_lshift4_b1[50] , shft_lshift4_b1[51] ,
         shft_lshift4_b1[52] , shft_lshift4_b1[53] , shft_lshift4_b1[54] ,
         shft_lshift4_b1[55] , shft_lshift4_b1[56] , shft_lshift4_b1[57] ,
         shft_lshift4_b1[58] , shft_lshift4_b1[59] , shft_lshift4_b1[60] ,
         shft_lshift4_b1[61] , shft_lshift4_b1[62] , shft_lshift4_b1[63] ,
         shft_lshift16_b1[32] , shft_lshift16_b1[33] ,
         shft_lshift16_b1[34] , shft_lshift16_b1[35] ,
         shft_lshift16_b1[36] , shft_lshift16_b1[37] ,
         shft_lshift16_b1[38] , shft_lshift16_b1[39] ,
         shft_lshift16_b1[40] , shft_lshift16_b1[41] ,
         shft_lshift16_b1[42] , shft_lshift16_b1[43] ,
         shft_lshift16_b1[44] , shft_lshift16_b1[45] ,
         shft_lshift16_b1[46] , shft_lshift16_b1[47] ,
         shft_lshift16_b1[48] , shft_lshift16_b1[49] ,
         shft_lshift16_b1[50] , shft_lshift16_b1[51] ,
         shft_lshift16_b1[52] , shft_lshift16_b1[53] ,
         shft_lshift16_b1[54] , shft_lshift16_b1[55] ,
         shft_lshift16_b1[56] , shft_lshift16_b1[57] ,
         shft_lshift16_b1[58] , shft_lshift16_b1[59] ,
         shft_lshift16_b1[60] , shft_lshift16_b1[61] ,
         shft_lshift16_b1[62] , shft_lshift16_b1[63] ,
         shft_shifter_input_b1[32] , shft_shifter_input_b1[33] ,
         shft_shifter_input_b1[34] , shft_shifter_input_b1[35] ,
         shft_shifter_input_b1[36] , shft_shifter_input_b1[37] ,
         shft_shifter_input_b1[38] , shft_shifter_input_b1[39] ,
         shft_shifter_input_b1[40] , shft_shifter_input_b1[41] ,
         shft_shifter_input_b1[42] , shft_shifter_input_b1[43] ,
         shft_shifter_input_b1[44] , shft_shifter_input_b1[45] ,
         shft_shifter_input_b1[46] , shft_shifter_input_b1[47] ,
         shft_shifter_input_b1[48] , shft_shifter_input_b1[49] ,
         shft_shifter_input_b1[50] , shft_shifter_input_b1[51] ,
         shft_shifter_input_b1[52] , shft_shifter_input_b1[53] ,
         shft_shifter_input_b1[54] , shft_shifter_input_b1[55] ,
         shft_shifter_input_b1[56] , shft_shifter_input_b1[57] ,
         shft_shifter_input_b1[58] , shft_shifter_input_b1[59] ,
         shft_shifter_input_b1[60] , shft_shifter_input_b1[61] ,
         shft_shifter_input_b1[62] , shft_shifter_input_b1[63] ,
         shft_rshift4_b1[0] , shft_rshift4_b1[1] , shft_rshift4_b1[2] ,
         shft_rshift4_b1[3] , shft_rshift4_b1[4] , shft_rshift4_b1[5] ,
         shft_rshift4_b1[6] , shft_rshift4_b1[7] , shft_rshift4_b1[8] ,
         shft_rshift4_b1[9] , shft_rshift4_b1[10] , shft_rshift4_b1[11] ,
         shft_rshift4_b1[12] , shft_rshift4_b1[13] , shft_rshift4_b1[14] ,
         shft_rshift4_b1[15] , shft_rshift4_b1[16] , shft_rshift4_b1[17] ,
         shft_rshift4_b1[18] , shft_rshift4_b1[19] , shft_rshift4_b1[20] ,
         shft_rshift4_b1[21] , shft_rshift4_b1[22] , shft_rshift4_b1[23] ,
         shft_rshift4_b1[24] , shft_rshift4_b1[25] , shft_rshift4_b1[26] ,
         shft_rshift4_b1[27] , shft_rshift4_b1[28] , shft_rshift4_b1[29] ,
         shft_rshift4_b1[30] , shft_rshift4_b1[31] , shft_rshift4_b1[32] ,
         shft_rshift4_b1[33] , shft_rshift4_b1[34] , shft_rshift4_b1[35] ,
         shft_rshift4_b1[36] , shft_rshift4_b1[37] , shft_rshift4_b1[38] ,
         shft_rshift4_b1[39] , shft_rshift4_b1[40] , shft_rshift4_b1[41] ,
         shft_rshift4_b1[42] , shft_rshift4_b1[43] , shft_rshift4_b1[44] ,
         shft_rshift4_b1[45] , shft_rshift4_b1[46] , shft_rshift4_b1[47] ,
         shft_rshift4_b1[48] , shft_rshift4_b1[49] , shft_rshift4_b1[50] ,
         shft_rshift4_b1[51] , shft_rshift4_b1[52] , shft_rshift4_b1[53] ,
         shft_rshift4_b1[54] , shft_rshift4_b1[55] , shft_rshift4_b1[56] ,
         shft_rshift4_b1[57] , shft_rshift4_b1[58] , shft_rshift4_b1[59] ,
         shft_rshift4_b1[60] , shft_rshift4_b1[61] , shft_rshift4_b1[62] ,
         shft_rshift4_b1[63] , shft_rshift16_b1[0] , shft_rshift16_b1[1] ,
         shft_rshift16_b1[2] , shft_rshift16_b1[3] , shft_rshift16_b1[4] ,
         shft_rshift16_b1[5] , shft_rshift16_b1[6] , shft_rshift16_b1[7] ,
         shft_rshift16_b1[8] , shft_rshift16_b1[9] , shft_rshift16_b1[10] ,
         shft_rshift16_b1[11] , shft_rshift16_b1[12] ,
         shft_rshift16_b1[13] , shft_rshift16_b1[14] ,
         shft_rshift16_b1[15] , shft_rshift16_b1[16] ,
         shft_rshift16_b1[17] , shft_rshift16_b1[18] ,
         shft_rshift16_b1[19] , shft_rshift16_b1[20] ,
         shft_rshift16_b1[21] , shft_rshift16_b1[22] ,
         shft_rshift16_b1[23] , shft_rshift16_b1[24] ,
         shft_rshift16_b1[25] , shft_rshift16_b1[26] ,
         shft_rshift16_b1[27] , shft_rshift16_b1[28] ,
         shft_rshift16_b1[29] , shft_rshift16_b1[30] ,
         shft_rshift16_b1[31] , shft_rshift16_b1[32] ,
         shft_rshift16_b1[33] , shft_rshift16_b1[34] ,
         shft_rshift16_b1[35] , shft_rshift16_b1[36] ,
         shft_rshift16_b1[37] , shft_rshift16_b1[38] ,
         shft_rshift16_b1[39] , shft_rshift16_b1[40] ,
         shft_rshift16_b1[41] , shft_rshift16_b1[42] ,
         shft_rshift16_b1[43] , shft_rshift16_b1[44] ,
         shft_rshift16_b1[45] , shft_rshift16_b1[46] ,
         shft_rshift16_b1[47] , shft_rshift16_b1[48] ,
         shft_rshift16_b1[49] , shft_rshift16_b1[50] ,
         shft_rshift16_b1[51] , shft_rshift16_b1[52] ,
         shft_rshift16_b1[53] , shft_rshift16_b1[54] ,
         shft_rshift16_b1[55] , shft_rshift16_b1[56] ,
         shft_rshift16_b1[57] , shft_rshift16_b1[58] ,
         shft_rshift16_b1[59] , shft_rshift16_b1[60] ,
         shft_rshift16_b1[61] , shft_rshift16_b1[62] ,
         shft_rshift16_b1[63] , shft_rshifterinput_b1[0] ,
         shft_rshifterinput_b1[1] , shft_rshifterinput_b1[2] ,
         shft_rshifterinput_b1[3] , shft_rshifterinput_b1[4] ,
         shft_rshifterinput_b1[5] , shft_rshifterinput_b1[6] ,
         shft_rshifterinput_b1[7] , shft_rshifterinput_b1[8] ,
         shft_rshifterinput_b1[9] , shft_rshifterinput_b1[10] ,
         shft_rshifterinput_b1[11] , shft_rshifterinput_b1[12] ,
         shft_rshifterinput_b1[13] , shft_rshifterinput_b1[14] ,
         shft_rshifterinput_b1[15] , shft_rshifterinput_b1[16] ,
         shft_rshifterinput_b1[17] , shft_rshifterinput_b1[18] ,
         shft_rshifterinput_b1[19] , shft_rshifterinput_b1[20] ,
         shft_rshifterinput_b1[21] , shft_rshifterinput_b1[22] ,
         shft_rshifterinput_b1[23] , shft_rshifterinput_b1[24] ,
         shft_rshifterinput_b1[25] , shft_rshifterinput_b1[26] ,
         shft_rshifterinput_b1[27] , shft_rshifterinput_b1[28] ,
         shft_rshifterinput_b1[29] , shft_rshifterinput_b1[30] ,
         shft_rshifterinput_b1[31] , shft_rshifterinput_b1[32] ,
         shft_rshifterinput_b1[33] , shft_rshifterinput_b1[34] ,
         shft_rshifterinput_b1[35] , shft_rshifterinput_b1[36] ,
         shft_rshifterinput_b1[37] , shft_rshifterinput_b1[38] ,
         shft_rshifterinput_b1[39] , shft_rshifterinput_b1[40] ,
         shft_rshifterinput_b1[41] , shft_rshifterinput_b1[42] ,
         shft_rshifterinput_b1[43] , shft_rshifterinput_b1[44] ,
         shft_rshifterinput_b1[45] , shft_rshifterinput_b1[46] ,
         shft_rshifterinput_b1[47] , shft_rshifterinput_b1[48] ,
         shft_rshifterinput_b1[49] , shft_rshifterinput_b1[50] ,
         shft_rshifterinput_b1[51] , shft_rshifterinput_b1[52] ,
         shft_rshifterinput_b1[53] , shft_rshifterinput_b1[54] ,
         shft_rshifterinput_b1[55] , shft_rshifterinput_b1[56] ,
         shft_rshifterinput_b1[57] , shft_rshifterinput_b1[58] ,
         shft_rshifterinput_b1[59] , shft_rshifterinput_b1[60] ,
         shft_rshifterinput_b1[61] , shft_rshifterinput_b1[62] ,
         shft_rshifterinput_b1[63] , shft_rshift1[63] , shft_rshift1[62] ,
         shft_rshift1[61] , shft_rshift1[60] , shft_rshift1[59] ,
         shft_rshift1[58] , shft_rshift1[57] , shft_rshift1[56] ,
         shft_rshift1[55] , shft_rshift1[54] , shft_rshift1[53] ,
         shft_rshift1[52] , shft_rshift1[51] , shft_rshift1[50] ,
         shft_rshift1[49] , shft_rshift1[48] , shft_rshift1[47] ,
         shft_rshift1[46] , shft_rshift1[45] , shft_rshift1[44] ,
         shft_rshift1[43] , shft_rshift1[42] , shft_rshift1[41] ,
         shft_rshift1[40] , shft_rshift1[39] , shft_rshift1[38] ,
         shft_rshift1[37] , shft_rshift1[36] , shft_rshift1[35] ,
         shft_rshift1[34] , shft_rshift1[33] , shft_rshift1[32] ,
         shft_rshift1[31] , shft_rshift1[30] , shft_rshift1[29] ,
         shft_rshift1[28] , shft_rshift1[27] , shft_rshift1[26] ,
         shft_rshift1[25] , shft_rshift1[24] , shft_rshift1[23] ,
         shft_rshift1[22] , shft_rshift1[21] , shft_rshift1[20] ,
         shft_rshift1[19] , shft_rshift1[18] , shft_rshift1[17] ,
         shft_rshift1[16] , shft_rshift1[15] , shft_rshift1[14] ,
         shft_rshift1[13] , shft_rshift1[12] , shft_rshift1[11] ,
         shft_rshift1[10] , shft_rshift1[9] , shft_rshift1[8] ,
         shft_rshift1[7] , shft_rshift1[6] , shft_rshift1[5] ,
         shft_rshift1[4] , shft_rshift1[3] , shft_rshift1[2] ,
         shft_rshift1[1] , shft_rshift1[0] , shft_lshift1[63] ,
         shft_lshift1[62] , shft_lshift1[61] , shft_lshift1[60] ,
         shft_lshift1[59] , shft_lshift1[58] , shft_lshift1[57] ,
         shft_lshift1[56] , shft_lshift1[55] , shft_lshift1[54] ,
         shft_lshift1[53] , shft_lshift1[52] , shft_lshift1[51] ,
         shft_lshift1[50] , shft_lshift1[49] , shft_lshift1[48] ,
         shft_lshift1[47] , shft_lshift1[46] , shft_lshift1[45] ,
         shft_lshift1[44] , shft_lshift1[43] , shft_lshift1[42] ,
         shft_lshift1[41] , shft_lshift1[40] , shft_lshift1[39] ,
         shft_lshift1[38] , shft_lshift1[37] , shft_lshift1[36] ,
         shft_lshift1[35] , shft_lshift1[34] , shft_lshift1[33] ,
         shft_lshift1[32] , shft_lshift1[31] , shft_lshift1[30] ,
         shft_lshift1[29] , shft_lshift1[28] , shft_lshift1[27] ,
         shft_lshift1[26] , shft_lshift1[25] , shft_lshift1[24] ,
         shft_lshift1[23] , shft_lshift1[22] , shft_lshift1[21] ,
         shft_lshift1[20] , shft_lshift1[19] , shft_lshift1[18] ,
         shft_lshift1[17] , shft_lshift1[16] , shft_lshift1[15] ,
         shft_lshift1[14] , shft_lshift1[13] , shft_lshift1[12] ,
         shft_lshift1[11] , shft_lshift1[10] , shft_lshift1[9] ,
         shft_lshift1[8] , shft_lshift1[7] , shft_lshift1[6] ,
         shft_lshift1[5] , shft_lshift1[4] , shft_lshift1[3] ,
         shft_lshift1[2] , shft_shift16_e[0] , shft_shift16_e[1] ,
         shft_shift16_e[2] , shft_shift16_e[3] , div_n96 , div_n95 ,
         div_n94 , div_n93 , div_n92 , div_n91 , div_n90 , div_n89 ,
         div_n88 , div_n87 , div_n86 , div_n85 , div_n84 , div_n83 ,
         div_n82 , div_n81 , div_n80 , div_n79 , div_n78 , div_n77 ,
         div_n76 , div_n75 , div_n74 , div_n73 , div_n72 , div_n71 ,
         div_n70 , div_n69 , div_n68 , div_n67 , div_n66 , div_n65 ,
         div_n64 , div_n63 , div_n62 , div_n61 , div_n60 , div_n59 ,
         div_n58 , div_n57 , div_n56 , div_n55 , div_n54 , div_n53 ,
         div_n52 , div_n51 , div_n50 , div_n49 , div_n48 , div_n47 ,
         div_n46 , div_n45 , div_n44 , div_n43 , div_n42 , div_n41 ,
         div_n40 , div_n39 , div_n38 , div_n37 , div_mul_result_next[63] ,
         div_mul_result_next[62] , div_mul_result_next[61] ,
         div_mul_result_next[60] , div_mul_result_next[59] ,
         div_mul_result_next[58] , div_mul_result_next[57] ,
         div_mul_result_next[56] , div_mul_result_next[55] ,
         div_mul_result_next[54] , div_mul_result_next[53] ,
         div_mul_result_next[52] , div_mul_result_next[51] ,
         div_mul_result_next[50] , div_mul_result_next[49] ,
         div_mul_result_next[48] , div_mul_result_next[47] ,
         div_mul_result_next[46] , div_mul_result_next[45] ,
         div_mul_result_next[44] , div_mul_result_next[43] ,
         div_mul_result_next[42] , div_mul_result_next[41] ,
         div_mul_result_next[40] , div_mul_result_next[39] ,
         div_mul_result_next[38] , div_mul_result_next[37] ,
         div_mul_result_next[36] , div_mul_result_next[35] ,
         div_mul_result_next[34] , div_mul_result_next[33] ,
         div_mul_result_next[32] , div_mul_result_next[31] ,
         div_mul_result_next[30] , div_mul_result_next[29] ,
         div_mul_result_next[28] , div_mul_result_next[27] ,
         div_mul_result_next[26] , div_mul_result_next[25] ,
         div_mul_result_next[24] , div_mul_result_next[23] ,
         div_mul_result_next[22] , div_mul_result_next[21] ,
         div_mul_result_next[20] , div_mul_result_next[19] ,
         div_mul_result_next[18] , div_mul_result_next[17] ,
         div_mul_result_next[16] , div_mul_result_next[15] ,
         div_mul_result_next[14] , div_mul_result_next[13] ,
         div_mul_result_next[12] , div_mul_result_next[11] ,
         div_mul_result_next[10] , div_mul_result_next[9] ,
         div_mul_result_next[8] , div_mul_result_next[7] ,
         div_mul_result_next[6] , div_mul_result_next[5] ,
         div_mul_result_next[4] , div_mul_result_next[3] ,
         div_mul_result_next[2] , div_mul_result_next[1] ,
         div_mul_result_next[0] , div_next_mul_data[127] ,
         div_next_mul_data[126] , div_next_mul_data[125] ,
         div_next_mul_data[124] , div_next_mul_data[123] ,
         div_next_mul_data[122] , div_next_mul_data[121] ,
         div_next_mul_data[120] , div_next_mul_data[119] ,
         div_next_mul_data[118] , div_next_mul_data[117] ,
         div_next_mul_data[116] , div_next_mul_data[115] ,
         div_next_mul_data[114] , div_next_mul_data[113] ,
         div_next_mul_data[112] , div_next_mul_data[111] ,
         div_next_mul_data[110] , div_next_mul_data[109] ,
         div_next_mul_data[108] , div_next_mul_data[107] ,
         div_next_mul_data[106] , div_next_mul_data[105] ,
         div_next_mul_data[104] , div_next_mul_data[103] ,
         div_next_mul_data[102] , div_next_mul_data[101] ,
         div_next_mul_data[100] , div_next_mul_data[99] ,
         div_next_mul_data[98] , div_next_mul_data[97] ,
         div_next_mul_data[96] , div_next_mul_data[95] ,
         div_next_mul_data[94] , div_next_mul_data[93] ,
         div_next_mul_data[92] , div_next_mul_data[91] ,
         div_next_mul_data[90] , div_next_mul_data[89] ,
         div_next_mul_data[88] , div_next_mul_data[87] ,
         div_next_mul_data[86] , div_next_mul_data[85] ,
         div_next_mul_data[84] , div_next_mul_data[83] ,
         div_next_mul_data[82] , div_next_mul_data[81] ,
         div_next_mul_data[80] , div_next_mul_data[79] ,
         div_next_mul_data[78] , div_next_mul_data[77] ,
         div_next_mul_data[76] , div_next_mul_data[75] ,
         div_next_mul_data[74] , div_next_mul_data[73] ,
         div_next_mul_data[72] , div_next_mul_data[71] ,
         div_next_mul_data[70] , div_next_mul_data[69] ,
         div_next_mul_data[68] , div_next_mul_data[67] ,
         div_next_mul_data[66] , div_next_mul_data[65] ,
         div_next_mul_data[64] , div_next_mul_data[63] ,
         div_next_mul_data[62] , div_next_mul_data[61] ,
         div_next_mul_data[60] , div_next_mul_data[59] ,
         div_next_mul_data[58] , div_next_mul_data[57] ,
         div_next_mul_data[56] , div_next_mul_data[55] ,
         div_next_mul_data[54] , div_next_mul_data[53] ,
         div_next_mul_data[52] , div_next_mul_data[51] ,
         div_next_mul_data[50] , div_next_mul_data[49] ,
         div_next_mul_data[48] , div_next_mul_data[47] ,
         div_next_mul_data[46] , div_next_mul_data[45] ,
         div_next_mul_data[44] , div_next_mul_data[43] ,
         div_next_mul_data[42] , div_next_mul_data[41] ,
         div_next_mul_data[40] , div_next_mul_data[39] ,
         div_next_mul_data[38] , div_next_mul_data[37] ,
         div_next_mul_data[36] , div_next_mul_data[35] ,
         div_next_mul_data[34] , div_next_mul_data[33] ,
         div_next_mul_data[32] , div_next_mul_data[31] ,
         div_next_mul_data[30] , div_next_mul_data[29] ,
         div_next_mul_data[28] , div_next_mul_data[27] ,
         div_next_mul_data[26] , div_next_mul_data[25] ,
         div_next_mul_data[24] , div_next_mul_data[23] ,
         div_next_mul_data[22] , div_next_mul_data[21] ,
         div_next_mul_data[20] , div_next_mul_data[19] ,
         div_next_mul_data[18] , div_next_mul_data[17] ,
         div_next_mul_data[16] , div_next_mul_data[15] ,
         div_next_mul_data[14] , div_next_mul_data[13] ,
         div_next_mul_data[12] , div_next_mul_data[11] ,
         div_next_mul_data[10] , div_next_mul_data[9] ,
         div_next_mul_data[8] , div_next_mul_data[7] ,
         div_next_mul_data[6] , div_next_mul_data[5] ,
         div_next_mul_data[4] , div_next_mul_data[3] ,
         div_next_mul_data[2] , div_next_mul_data[1] ,
         div_next_mul_data[0] , div_z_in[63] , div_z_in[62] ,
         div_z_in[61] , div_z_in[60] , div_z_in[59] , div_z_in[58] ,
         div_z_in[57] , div_z_in[56] , div_z_in[55] , div_z_in[54] ,
         div_z_in[53] , div_z_in[52] , div_z_in[51] , div_z_in[50] ,
         div_z_in[49] , div_z_in[48] , div_z_in[47] , div_z_in[46] ,
         div_z_in[45] , div_z_in[44] , div_z_in[43] , div_z_in[42] ,
         div_z_in[41] , div_z_in[40] , div_z_in[39] , div_z_in[38] ,
         div_z_in[37] , div_z_in[36] , div_z_in[35] , div_z_in[34] ,
         div_z_in[33] , div_z_in[32] , div_z_in[31] , div_z_in[30] ,
         div_z_in[29] , div_z_in[28] , div_z_in[27] , div_z_in[26] ,
         div_z_in[25] , div_z_in[24] , div_z_in[23] , div_z_in[22] ,
         div_z_in[21] , div_z_in[20] , div_z_in[19] , div_z_in[18] ,
         div_z_in[17] , div_z_in[16] , div_z_in[15] , div_z_in[14] ,
         div_z_in[13] , div_z_in[12] , div_z_in[11] , div_z_in[10] ,
         div_z_in[9] , div_z_in[8] , div_z_in[7] , div_z_in[6] ,
         div_z_in[5] , div_z_in[4] , div_z_in[3] , div_z_in[2] ,
         div_z_in[1] , div_z_in[0] , div_spr_out[63] , div_spr_out[62] ,
         div_spr_out[61] , div_spr_out[60] , div_spr_out[59] ,
         div_spr_out[58] , div_spr_out[57] , div_spr_out[56] ,
         div_spr_out[55] , div_spr_out[54] , div_spr_out[53] ,
         div_spr_out[52] , div_spr_out[51] , div_spr_out[50] ,
         div_spr_out[49] , div_spr_out[48] , div_spr_out[47] ,
         div_spr_out[46] , div_spr_out[45] , div_spr_out[44] ,
         div_spr_out[43] , div_spr_out[42] , div_spr_out[41] ,
         div_spr_out[40] , div_spr_out[39] , div_spr_out[38] ,
         div_spr_out[37] , div_spr_out[36] , div_spr_out[35] ,
         div_spr_out[34] , div_spr_out[33] , div_spr_out[32] ,
         div_spr_out[31] , div_spr_out[30] , div_spr_out[29] ,
         div_spr_out[28] , div_spr_out[27] , div_spr_out[26] ,
         div_spr_out[25] , div_spr_out[24] , div_spr_out[23] ,
         div_spr_out[22] , div_spr_out[21] , div_spr_out[20] ,
         div_spr_out[19] , div_spr_out[18] , div_spr_out[17] ,
         div_spr_out[16] , div_spr_out[15] , div_spr_out[14] ,
         div_spr_out[13] , div_spr_out[12] , div_spr_out[11] ,
         div_spr_out[10] , div_spr_out[9] , div_spr_out[8] ,
         div_spr_out[7] , div_spr_out[6] , div_spr_out[5] ,
         div_spr_out[4] , div_spr_out[3] , div_spr_out[2] ,
         div_spr_out[1] , div_spr_out[0] , div_adder_out_0 ,
         div_adder_out_1 , div_adder_out_2 , div_adder_out_3 ,
         div_adder_out_4 , div_adder_out_5 , div_adder_out_6 ,
         div_adder_out_7 , div_adder_out_8 , div_adder_out_9 ,
         div_adder_out_10 , div_adder_out_11 , div_adder_out_12 ,
         div_adder_out_13 , div_adder_out_14 , div_adder_out_15 ,
         div_adder_out_16 , div_adder_out_17 , div_adder_out_18 ,
         div_adder_out_19 , div_adder_out_20 , div_adder_out_21 ,
         div_adder_out_22 , div_adder_out_23 , div_adder_out_24 ,
         div_adder_out_25 , div_adder_out_26 , div_adder_out_27 ,
         div_adder_out_28 , div_adder_out_29 , div_adder_out_30 ,
         div_adder_out[63] , div_adder_out[62] , div_adder_out[61] ,
         div_adder_out[60] , div_adder_out[59] , div_adder_out[58] ,
         div_adder_out[57] , div_adder_out[56] , div_adder_out[55] ,
         div_adder_out[54] , div_adder_out[53] , div_adder_out[52] ,
         div_adder_out[51] , div_adder_out[50] , div_adder_out[49] ,
         div_adder_out[48] , div_adder_out[47] , div_adder_out[46] ,
         div_adder_out[45] , div_adder_out[44] , div_adder_out[43] ,
         div_adder_out[42] , div_adder_out[41] , div_adder_out[40] ,
         div_adder_out[39] , div_adder_out[38] , div_adder_out[37] ,
         div_adder_out[36] , div_adder_out[35] , div_adder_out[34] ,
         div_adder_out[33] , div_adder_out[32] , div_adderin2[0] ,
         div_adderin2[1] , div_adderin2[2] , div_adderin2[3] ,
         div_adderin2[4] , div_adderin2[5] , div_adderin2[6] ,
         div_adderin2[7] , div_adderin2[8] , div_adderin2[9] ,
         div_adderin2[10] , div_adderin2[11] , div_adderin2[12] ,
         div_adderin2[13] , div_adderin2[14] , div_adderin2[15] ,
         div_adderin2[16] , div_adderin2[17] , div_adderin2[18] ,
         div_adderin2[19] , div_adderin2[20] , div_adderin2[21] ,
         div_adderin2[22] , div_adderin2[23] , div_adderin2[24] ,
         div_adderin2[25] , div_adderin2[26] , div_adderin2[27] ,
         div_adderin2[28] , div_adderin2[29] , div_adderin2[30] ,
         div_adderin2[31] , div_adderin2[32] , div_adderin2[33] ,
         div_adderin2[34] , div_adderin2[35] , div_adderin2[36] ,
         div_adderin2[37] , div_adderin2[38] , div_adderin2[39] ,
         div_adderin2[40] , div_adderin2[41] , div_adderin2[42] ,
         div_adderin2[43] , div_adderin2[44] , div_adderin2[45] ,
         div_adderin2[46] , div_adderin2[47] , div_adderin2[48] ,
         div_adderin2[49] , div_adderin2[50] , div_adderin2[51] ,
         div_adderin2[52] , div_adderin2[53] , div_adderin2[54] ,
         div_adderin2[55] , div_adderin2[56] , div_adderin2[57] ,
         div_adderin2[58] , div_adderin2[59] , div_adderin2[60] ,
         div_adderin2[61] , div_adderin2[62] , div_adderin2[63] ,
         div_adderin1[0] , div_adderin1[1] , div_adderin1[2] ,
         div_adderin1[3] , div_adderin1[4] , div_adderin1[5] ,
         div_adderin1[6] , div_adderin1[7] , div_adderin1[8] ,
         div_adderin1[9] , div_adderin1[10] , div_adderin1[11] ,
         div_adderin1[12] , div_adderin1[13] , div_adderin1[14] ,
         div_adderin1[15] , div_adderin1[16] , div_adderin1[17] ,
         div_adderin1[18] , div_adderin1[19] , div_adderin1[20] ,
         div_adderin1[21] , div_adderin1[22] , div_adderin1[23] ,
         div_adderin1[24] , div_adderin1[25] , div_adderin1[26] ,
         div_adderin1[27] , div_adderin1[28] , div_adderin1[29] ,
         div_adderin1[30] , div_adderin1[31] , div_adderin1[32] ,
         div_adderin1[33] , div_adderin1[34] , div_adderin1[35] ,
         div_adderin1[36] , div_adderin1[37] , div_adderin1[38] ,
         div_adderin1[39] , div_adderin1[40] , div_adderin1[41] ,
         div_adderin1[42] , div_adderin1[43] , div_adderin1[44] ,
         div_adderin1[45] , div_adderin1[46] , div_adderin1[47] ,
         div_adderin1[48] , div_adderin1[49] , div_adderin1[50] ,
         div_adderin1[51] , div_adderin1[52] , div_adderin1[53] ,
         div_adderin1[54] , div_adderin1[55] , div_adderin1[56] ,
         div_adderin1[57] , div_adderin1[58] , div_adderin1[59] ,
         div_adderin1[60] , div_adderin1[61] , div_adderin1[62] ,
         div_adderin1[63] , div_x[0] , div_x[1] , div_x[2] , div_x[3] ,
         div_x[4] , div_x[5] , div_x[6] , div_x[7] , div_x[8] ,
         div_x[9] , div_x[10] , div_x[11] , div_x[12] , div_x[13] ,
         div_x[14] , div_x[15] , div_x[16] , div_x[17] , div_x[18] ,
         div_x[19] , div_x[20] , div_x[21] , div_x[22] , div_x[23] ,
         div_x[24] , div_x[25] , div_x[26] , div_x[27] , div_x[28] ,
         div_x[29] , div_x[30] , div_x[31] , div_x[32] , div_x[33] ,
         div_x[34] , div_x[35] , div_x[36] , div_x[37] , div_x[38] ,
         div_x[39] , div_x[40] , div_x[41] , div_x[42] , div_x[43] ,
         div_x[44] , div_x[45] , div_x[46] , div_x[47] , div_x[48] ,
         div_x[49] , div_x[50] , div_x[51] , div_x[52] , div_x[53] ,
         div_x[54] , div_x[55] , div_x[56] , div_x[57] , div_x[58] ,
         div_x[59] , div_x[60] , div_x[61] , div_x[62] , div_xin[0] ,
         div_xin[1] , div_xin[2] , div_xin[3] , div_xin[4] , div_xin[5] ,
         div_xin[6] , div_xin[7] , div_xin[8] , div_xin[9] , div_xin[10] ,
         div_xin[11] , div_xin[12] , div_xin[13] , div_xin[14] ,
         div_xin[15] , div_xin[16] , div_xin[17] , div_xin[18] ,
         div_xin[19] , div_xin[20] , div_xin[21] , div_xin[22] ,
         div_xin[23] , div_xin[24] , div_xin[25] , div_xin[26] ,
         div_xin[27] , div_xin[28] , div_xin[29] , div_xin[30] ,
         div_xin[31] , div_xin[32] , div_xin[33] , div_xin[34] ,
         div_xin[35] , div_xin[36] , div_xin[37] , div_xin[38] ,
         div_xin[39] , div_xin[40] , div_xin[41] , div_xin[42] ,
         div_xin[43] , div_xin[44] , div_xin[45] , div_xin[46] ,
         div_xin[47] , div_xin[48] , div_xin[49] , div_xin[50] ,
         div_xin[51] , div_xin[52] , div_xin[53] , div_xin[54] ,
         div_xin[55] , div_xin[56] , div_xin[57] , div_xin[58] ,
         div_xin[59] , div_xin[60] , div_xin[61] , div_xin[62] ,
         div_xin[63] , div_dnext[127] , div_dnext[126] , div_dnext[125] ,
         div_dnext[124] , div_dnext[123] , div_dnext[122] ,
         div_dnext[121] , div_dnext[120] , div_dnext[119] ,
         div_dnext[118] , div_dnext[117] , div_dnext[116] ,
         div_dnext[115] , div_dnext[114] , div_dnext[113] ,
         div_dnext[112] , div_dnext[111] , div_dnext[110] ,
         div_dnext[109] , div_dnext[108] , div_dnext[107] ,
         div_dnext[106] , div_dnext[105] , div_dnext[104] ,
         div_dnext[103] , div_dnext[102] , div_dnext[101] ,
         div_dnext[100] , div_dnext[99] , div_dnext[98] , div_dnext[97] ,
         div_dnext[96] , div_dnext[95] , div_dnext[94] , div_dnext[93] ,
         div_dnext[92] , div_dnext[91] , div_dnext[90] , div_dnext[89] ,
         div_dnext[88] , div_dnext[87] , div_dnext[86] , div_dnext[85] ,
         div_dnext[84] , div_dnext[83] , div_dnext[82] , div_dnext[81] ,
         div_dnext[80] , div_dnext[79] , div_dnext[78] , div_dnext[77] ,
         div_dnext[76] , div_dnext[75] , div_dnext[74] , div_dnext[73] ,
         div_dnext[72] , div_dnext[71] , div_dnext[70] , div_dnext[69] ,
         div_dnext[68] , div_dnext[67] , div_dnext[66] , div_dnext[65] ,
         div_dnext[64] , div_dnext[63] , div_dnext[62] , div_dnext[61] ,
         div_dnext[60] , div_dnext[59] , div_dnext[58] , div_dnext[57] ,
         div_dnext[56] , div_dnext[55] , div_dnext[54] , div_dnext[53] ,
         div_dnext[52] , div_dnext[51] , div_dnext[50] , div_dnext[49] ,
         div_dnext[48] , div_dnext[47] , div_dnext[46] , div_dnext[45] ,
         div_dnext[44] , div_dnext[43] , div_dnext[42] , div_dnext[41] ,
         div_dnext[40] , div_dnext[39] , div_dnext[38] , div_dnext[37] ,
         div_dnext[36] , div_dnext[35] , div_dnext[34] , div_dnext[33] ,
         div_dnext[32] , div_dnext[31] , div_dnext[30] , div_dnext[29] ,
         div_dnext[28] , div_dnext[27] , div_dnext[26] , div_dnext[25] ,
         div_dnext[24] , div_dnext[23] , div_dnext[22] , div_dnext[21] ,
         div_dnext[20] , div_dnext[19] , div_dnext[18] , div_dnext[17] ,
         div_dnext[16] , div_dnext[15] , div_dnext[14] , div_dnext[13] ,
         div_dnext[12] , div_dnext[11] , div_dnext[10] , div_dnext[9] ,
         div_dnext[8] , div_dnext[7] , div_dnext[6] , div_dnext[5] ,
         div_dnext[4] , div_dnext[3] , div_dnext[2] , div_dnext[1] ,
         div_dnext[0] , div_din[94] , div_din[93] , div_din[92] ,
         div_din[91] , div_din[90] , div_din[89] , div_din[88] ,
         div_din[87] , div_din[86] , div_din[85] , div_din[84] ,
         div_din[83] , div_din[82] , div_din[81] , div_din[80] ,
         div_din[79] , div_din[78] , div_din[77] , div_din[76] ,
         div_din[75] , div_din[74] , div_din[73] , div_din[72] ,
         div_din[71] , div_din[70] , div_din[69] , div_din[68] ,
         div_din[67] , div_din[66] , div_din[65] , div_din[64] ,
         div_din[63] , div_out64[63] , div_out64[62] , div_out64[61] ,
         div_out64[60] , div_out64[59] , div_out64[58] , div_out64[57] ,
         div_out64[56] , div_out64[55] , div_out64[54] , div_out64[53] ,
         div_out64[52] , div_out64[51] , div_out64[50] , div_out64[49] ,
         div_out64[48] , div_out64[47] , div_out64[46] , div_out64[45] ,
         div_out64[44] , div_out64[43] , div_out64[42] , div_out64[41] ,
         div_out64[40] , div_out64[39] , div_out64[38] , div_out64[37] ,
         div_out64[36] , div_out64[35] , div_out64[34] , div_out64[33] ,
         div_out64[32] , div_out64[31] , div_out64[30] , div_out64[29] ,
         div_out64[28] , div_out64[27] , div_out64[26] , div_out64[25] ,
         div_out64[24] , div_out64[23] , div_out64[22] , div_out64[21] ,
         div_out64[20] , div_out64[19] , div_out64[18] , div_out64[17] ,
         div_out64[16] , div_out64[15] , div_out64[14] , div_out64[13] ,
         div_out64[12] , div_out64[11] , div_out64[10] , div_out64[9] ,
         div_out64[8] , div_out64[7] , div_out64[6] , div_out64[5] ,
         div_out64[4] , div_out64[3] , div_out64[2] , div_out64[1] ,
         div_out64[0] , div_neg32[30] , div_neg32[29] , div_neg32[28] ,
         div_neg32[27] , div_neg32[26] , div_neg32[25] , div_neg32[24] ,
         div_neg32[23] , div_neg32[22] , div_neg32[21] , div_neg32[20] ,
         div_neg32[19] , div_neg32[18] , div_neg32[17] , div_neg32[16] ,
         div_neg32[15] , div_neg32[14] , div_neg32[13] , div_neg32[12] ,
         div_neg32[11] , div_neg32[10] , div_neg32[9] , div_neg32[8] ,
         div_neg32[7] , div_neg32[6] , div_neg32[5] , div_neg32[4] ,
         div_neg32[3] , div_neg32[2] , div_neg32[1] , div_neg32[0] ,
         div_pos32[30] , div_pos32[29] , div_pos32[28] , div_pos32[27] ,
         div_pos32[26] , div_pos32[25] , div_pos32[24] , div_pos32[23] ,
         div_pos32[22] , div_pos32[21] , div_pos32[20] , div_pos32[19] ,
         div_pos32[18] , div_pos32[17] , div_pos32[16] , div_pos32[15] ,
         div_pos32[14] , div_pos32[13] , div_pos32[12] , div_pos32[11] ,
         div_pos32[10] , div_pos32[9] , div_pos32[8] , div_pos32[7] ,
         div_pos32[6] , div_pos32[5] , div_pos32[4] , div_pos32[3] ,
         div_pos32[2] , div_pos32[1] , div_pos32[0] , div_u32[31] ,
         div_u32[30] , div_u32[29] , div_u32[28] , div_u32[27] ,
         div_u32[26] , div_u32[25] , div_u32[24] , div_u32[23] ,
         div_u32[22] , div_u32[21] , div_u32[20] , div_u32[19] ,
         div_u32[18] , div_u32[17] , div_u32[16] , div_u32[15] ,
         div_u32[14] , div_u32[13] , div_u32[12] , div_u32[11] ,
         div_u32[10] , div_u32[9] , div_u32[8] , div_u32[7] , div_u32[6] ,
         div_u32[5] , div_u32[4] , div_u32[3] , div_u32[2] , div_u32[1] ,
         div_u32[0] , div_curr_q[0] , div_curr_q[1] , div_curr_q[2] ,
         div_curr_q[3] , div_curr_q[4] , div_curr_q[5] , div_curr_q[6] ,
         div_curr_q[7] , div_curr_q[8] , div_curr_q[9] , div_curr_q[10] ,
         div_curr_q[11] , div_curr_q[12] , div_curr_q[13] ,
         div_curr_q[14] , div_curr_q[15] , div_curr_q[16] ,
         div_curr_q[17] , div_curr_q[18] , div_curr_q[19] ,
         div_curr_q[20] , div_curr_q[21] , div_curr_q[22] ,
         div_curr_q[23] , div_curr_q[24] , div_curr_q[25] ,
         div_curr_q[26] , div_curr_q[27] , div_curr_q[28] ,
         div_curr_q[29] , div_curr_q[30] , div_curr_q[31] ,
         div_curr_q[32] , div_curr_q[33] , div_curr_q[34] ,
         div_curr_q[35] , div_curr_q[36] , div_curr_q[37] ,
         div_curr_q[38] , div_curr_q[39] , div_curr_q[40] ,
         div_curr_q[41] , div_curr_q[42] , div_curr_q[43] ,
         div_curr_q[44] , div_curr_q[45] , div_curr_q[46] ,
         div_curr_q[47] , div_curr_q[48] , div_curr_q[49] ,
         div_curr_q[50] , div_curr_q[51] , div_curr_q[52] ,
         div_curr_q[53] , div_curr_q[54] , div_curr_q[55] ,
         div_curr_q[56] , div_curr_q[57] , div_curr_q[58] ,
         div_curr_q[59] , div_curr_q[60] , div_curr_q[61] ,
         div_curr_q[62] , div_gencc_in_0 , div_gencc_in_1 ,
         div_gencc_in_2 , div_gencc_in_3 , div_gencc_in_4 ,
         div_gencc_in_5 , div_gencc_in_6 , div_gencc_in_7 ,
         div_gencc_in_8 , div_gencc_in_9 , div_gencc_in_10 ,
         div_gencc_in_11 , div_gencc_in_12 , div_gencc_in_13 ,
         div_gencc_in_14 , div_gencc_in_15 , div_gencc_in_16 ,
         div_gencc_in_17 , div_gencc_in_18 , div_gencc_in_19 ,
         div_gencc_in_20 , div_gencc_in_21 , div_gencc_in_22 ,
         div_gencc_in_23 , div_gencc_in_24 , div_gencc_in_25 ,
         div_gencc_in_26 , div_gencc_in_27 , div_gencc_in_28 ,
         div_gencc_in_29 , div_gencc_in_30 , div_gencc_in[32] ,
         div_gencc_in[33] , div_gencc_in[34] , div_gencc_in[35] ,
         div_gencc_in[36] , div_gencc_in[37] , div_gencc_in[38] ,
         div_gencc_in[39] , div_gencc_in[40] , div_gencc_in[41] ,
         div_gencc_in[42] , div_gencc_in[43] , div_gencc_in[44] ,
         div_gencc_in[45] , div_gencc_in[46] , div_gencc_in[47] ,
         div_gencc_in[48] , div_gencc_in[49] , div_gencc_in[50] ,
         div_gencc_in[51] , div_gencc_in[52] , div_gencc_in[53] ,
         div_gencc_in[54] , div_gencc_in[55] , div_gencc_in[56] ,
         div_gencc_in[57] , div_gencc_in[58] , div_gencc_in[59] ,
         div_gencc_in[60] , div_gencc_in[61] , div_gencc_in[62] ,
         div_gencc_in[63] , div_mul_result[0] , div_mul_result[1] ,
         div_mul_result[2] , div_mul_result[3] , div_mul_result[4] ,
         div_mul_result[5] , div_mul_result[6] , div_mul_result[7] ,
         div_mul_result[8] , div_mul_result[9] , div_mul_result[10] ,
         div_mul_result[11] , div_mul_result[12] , div_mul_result[13] ,
         div_mul_result[14] , div_mul_result[15] , div_mul_result[16] ,
         div_mul_result[17] , div_mul_result[18] , div_mul_result[19] ,
         div_mul_result[20] , div_mul_result[21] , div_mul_result[22] ,
         div_mul_result[23] , div_mul_result[24] , div_mul_result[25] ,
         div_mul_result[26] , div_mul_result[27] , div_mul_result[28] ,
         div_mul_result[29] , div_mul_result[30] , div_mul_result[31] ,
         div_mul_result[32] , div_mul_result[33] , div_mul_result[34] ,
         div_mul_result[35] , div_mul_result[36] , div_mul_result[37] ,
         div_mul_result[38] , div_mul_result[39] , div_mul_result[40] ,
         div_mul_result[41] , div_mul_result[42] , div_mul_result[43] ,
         div_mul_result[44] , div_mul_result[45] , div_mul_result[46] ,
         div_mul_result[47] , div_mul_result[48] , div_mul_result[49] ,
         div_mul_result[50] , div_mul_result[51] , div_mul_result[52] ,
         div_mul_result[53] , div_mul_result[54] , div_mul_result[55] ,
         div_mul_result[56] , div_mul_result[57] , div_mul_result[58] ,
         div_mul_result[59] , div_mul_result[60] , div_mul_result[61] ,
         div_mul_result[62] , div_mul_result[63] , div_d[0] , div_d[1] ,
         div_d[2] , div_d[3] , div_d[4] , div_d[5] , div_d[6] ,
         div_d[7] , div_d[8] , div_d[9] , div_d[10] , div_d[11] ,
         div_d[12] , div_d[13] , div_d[14] , div_d[15] , div_d[16] ,
         div_d[17] , div_d[18] , div_d[19] , div_d[20] , div_d[21] ,
         div_d[22] , div_d[23] , div_d[24] , div_d[25] , div_d[26] ,
         div_d[27] , div_d[28] , div_d[29] , div_d[30] , div_d[31] ,
         div_d[32] , div_d[33] , div_d[34] , div_d[35] , div_d[36] ,
         div_d[37] , div_d[38] , div_d[39] , div_d[40] , div_d[41] ,
         div_d[42] , div_d[43] , div_d[44] , div_d[45] , div_d[46] ,
         div_d[47] , div_d[48] , div_d[49] , div_d[50] , div_d[51] ,
         div_d[52] , div_d[53] , div_d[54] , div_d[55] , div_d[56] ,
         div_d[57] , div_d[58] , div_d[59] , div_d[60] , div_d[61] ,
         div_d_63 , div_dividend[62] , div_dividend[61] ,
         div_dividend[60] , div_dividend[59] , div_dividend[58] ,
         div_dividend[57] , div_dividend[56] , div_dividend[55] ,
         div_dividend[54] , div_dividend[53] , div_dividend[52] ,
         div_dividend[51] , div_dividend[50] , div_dividend[49] ,
         div_dividend[48] , div_dividend[47] , div_dividend[46] ,
         div_dividend[45] , div_dividend[44] , div_dividend[43] ,
         div_dividend[42] , div_dividend[41] , div_dividend[40] ,
         div_dividend[39] , div_dividend[38] , div_dividend[37] ,
         div_dividend[36] , div_dividend[35] , div_dividend[34] ,
         div_dividend[33] , div_dividend[32] , div_input_data_e[64] ,
         div_input_data_e[65] , div_input_data_e[66] ,
         div_input_data_e[67] , div_input_data_e[68] ,
         div_input_data_e[69] , div_input_data_e[70] ,
         div_input_data_e[71] , div_input_data_e[72] ,
         div_input_data_e[73] , div_input_data_e[74] ,
         div_input_data_e[75] , div_input_data_e[76] ,
         div_input_data_e[77] , div_input_data_e[78] ,
         div_input_data_e[79] , div_input_data_e[80] ,
         div_input_data_e[81] , div_input_data_e[82] ,
         div_input_data_e[83] , div_input_data_e[84] ,
         div_input_data_e[85] , div_input_data_e[86] ,
         div_input_data_e[87] , div_input_data_e[88] ,
         div_input_data_e[89] , div_input_data_e[90] ,
         div_input_data_e[91] , div_input_data_e[92] ,
         div_input_data_e[93] , div_input_data_e[94] ,
         div_input_data_e[95] , div_input_data_e[96] ,
         div_input_data_e[97] , div_input_data_e[98] ,
         div_input_data_e[99] , div_input_data_e[100] ,
         div_input_data_e[101] , div_input_data_e[102] ,
         div_input_data_e[103] , div_input_data_e[104] ,
         div_input_data_e[105] , div_input_data_e[106] ,
         div_input_data_e[107] , div_input_data_e[108] ,
         div_input_data_e[109] , div_input_data_e[110] ,
         div_input_data_e[111] , div_input_data_e[112] ,
         div_input_data_e[113] , div_input_data_e[114] ,
         div_input_data_e[115] , div_input_data_e[116] ,
         div_input_data_e[117] , div_input_data_e[118] ,
         div_input_data_e[119] , div_input_data_e[120] ,
         div_input_data_e[121] , div_input_data_e[122] ,
         div_input_data_e[123] , div_input_data_e[124] ,
         div_input_data_e[125] , div_input_data_e[126] ,
         div_input_data_e[127] , rml_n131 , rml_n130 , rml_n128 ,
         rml_n127 , rml_n126 , rml_n125 , rml_n124 , rml_n123 ,
         rml_n122 , rml_n121 , rml_n120 , rml_n119 , rml_n118 ,
         rml_n117 , rml_n116 , rml_n115 , rml_n114 , rml_n113 ,
         rml_n112 , rml_n111 , rml_n110 , rml_n109 , rml_n108 ,
         rml_n107 , rml_n106 , rml_n105 , rml_n104 , rml_n103 ,
         rml_n102 , rml_n101 , rml_n100 , rml_n99 , rml_n98 , rml_n97 ,
         rml_n95 , rml_n94 , rml_n93 , rml_n92 , rml_n91 , rml_n90 ,
         rml_n89 , rml_n88 , rml_n87 , rml_n86 , rml_n85 , rml_n84 ,
         rml_n83 , rml_n82 , rml_n81 , rml_n80 , rml_n79 , rml_n78 ,
         rml_n77 , rml_n76 , rml_n75 , rml_n74 , rml_n73 , rml_n72 ,
         rml_n71 , rml_n70 , rml_n69 , rml_n68 , rml_n67 , rml_n66 ,
         rml_n65 , rml_n64 , rml_n63 , rml_n62 , rml_n61 , rml_n60 ,
         rml_n59 , rml_n58 , rml_n57 , rml_n56 , rml_n55 , rml_n54 ,
         rml_n53 , rml_n52 , rml_n51 , rml_n50 , rml_n49 , rml_n48 ,
         rml_n47 , rml_n46 , rml_n45 , rml_n44 , rml_n43 , rml_n42 ,
         rml_n41 , rml_n40 , rml_n39 , rml_n38 , rml_n37 , rml_n36 ,
         rml_n35 , rml_agp_thr3_next[1] , rml_agp_thr3_next[0] ,
         rml_agp_thr2_next[1] , rml_agp_thr2_next[0] ,
         rml_agp_thr1_next[1] , rml_agp_thr1_next[0] , rml_new_agp[0] ,
         rml_new_agp[1] , rml_agp_thr0_next[1] , rml_agp_thr0_next[0] ,
         rml_agp_wen_thr3_w , rml_agp_wen_thr2_w , rml_agp_wen_thr1_w ,
         rml_agp_wen_thr0_w , rml_agp_thr3[0] , rml_agp_thr3[1] ,
         rml_agp_thr2[0] , rml_agp_thr2[1] , rml_agp_thr1[0] ,
         rml_agp_thr1[1] , rml_agp_thr0[0] , rml_agp_thr0[1] ,
         rml_agp_thr[0] , rml_agp_thr[1] , rml_agp_thr[2] ,
         rml_agp_thr[3] , rml_wstate_wen_w , rml_cleanwin_wen_w ,
         rml_next_cleanwin_w[2] , rml_next_cleanwin_w[1] ,
         rml_next_cleanwin_w[0] , rml_rml_cleanwin_wen_w ,
         rml_next_cleanwin_m[2] , rml_next_cleanwin_m[1] ,
         rml_next_cleanwin_m[0] , rml_cleanwin_wen_m ,
         rml_next_cleanwin_e[2] , rml_next_cleanwin_e[1] ,
         rml_next_cleanwin_e[0] , rml_rml_next_cleanwin_e[2] ,
         rml_rml_next_cleanwin_e[1] , rml_otherwin_wen_w ,
         rml_next_otherwin_w[2] , rml_next_otherwin_w[1] ,
         rml_next_otherwin_w[0] , rml_rml_otherwin_wen_w ,
         rml_next_otherwin_m[2] , rml_next_otherwin_m[1] ,
         rml_next_otherwin_m[0] , rml_otherwin_wen_m ,
         rml_next_otherwin_e[2] , rml_next_otherwin_e[1] ,
         rml_next_otherwin_e[0] , rml_rml_next_otherwin_e[2] ,
         rml_rml_next_otherwin_e[1] , rml_rml_ecl_otherwin_e[0] ,
         rml_rml_ecl_otherwin_e[1] , rml_rml_ecl_otherwin_e[2] ,
         rml_canrestore_wen_w , rml_next_canrestore_w[2] ,
         rml_next_canrestore_w[1] , rml_next_canrestore_w[0] ,
         rml_rml_canrestore_wen_w , rml_next_canrestore_m[2] ,
         rml_next_canrestore_m[1] , rml_next_canrestore_m[0] ,
         rml_canrestore_wen_m , rml_next_canrestore_e[2] ,
         rml_next_canrestore_e[1] , rml_next_canrestore_e[0] ,
         rml_canrestore_inc_e , rml_rml_next_canrestore_e[2] ,
         rml_rml_next_canrestore_e[1] , rml_canrestore_wen_e ,
         rml_cansave_wen_w , rml_next_cansave_w[2] , rml_next_cansave_w[1] ,
         rml_next_cansave_w[0] , rml_rml_cansave_wen_w ,
         rml_next_cansave_m[2] , rml_next_cansave_m[1] ,
         rml_next_cansave_m[0] , rml_cansave_wen_m , rml_next_cansave_e[2] ,
         rml_next_cansave_e[1] , rml_next_cansave_e[0] , rml_cansave_inc_e ,
         rml_rml_next_cansave_e[2] , rml_rml_next_cansave_e[1] ,
         rml_cansave_wen_e , rml_oddwin_m[3] , rml_oddwin_m[2] ,
         rml_oddwin_m[1] , rml_oddwin_m[0] , rml_oddwin_w[3] ,
         rml_oddwin_w[2] , rml_oddwin_w[1] , rml_oddwin_w[0] ,
         rml_full_swap_e , rml_cwp_wen_w , rml_cwp_wen_nokill_w ,
         rml_next_cwp_noreset_w[2] , rml_next_cwp_noreset_w[1] ,
         rml_next_cwp_noreset_w[0] , rml_next_cwp_m[0] , rml_next_cwp_m[1] ,
         rml_next_cwp_m[2] , rml_rml_cwp_wen_m , rml_next_cwp_e[0] ,
         rml_next_cwp_e[1] , rml_next_cwp_e[2] , rml_rml_next_cwp_e[2] ,
         rml_rml_next_cwp_e[1] , rml_cwp_wen_e , rml_spill_cwp_e[2] ,
         rml_spill_cwp_e[1] , rml_spill_cwp_e[0] , rml_rml_ecl_cwp_e[0] ,
         rml_rml_ecl_cwp_e[1] , rml_rml_ecl_cwp_e[2] , rml_kill_restore_w ,
         rml_kill_restore_m , rml_did_restore_w , rml_did_restore_m ,
         rml_swap_locals_ins , rml_swap_e , rml_rml_ecl_other_d ,
         rml_rml_ecl_kill_e , rml_rml_ecl_cleanwin_e[0] ,
         rml_rml_ecl_cleanwin_e[1] , rml_rml_ecl_cleanwin_e[2] ,
         rml_spill_m , rml_rml_ecl_cansave_e[0] , rml_rml_ecl_cansave_e[1] ,
         rml_rml_ecl_cansave_e[2] , rml_rml_ecl_canrestore_e[0] ,
         rml_rml_ecl_canrestore_e[1] , rml_rml_ecl_canrestore_e[2] ,
         rml_win_trap_m , rml_win_trap_e , rml_exu_tlu_spill_e ,
         rml_rml_kill_w , rml_win_trap_w , rml_restore_e , rml_save_m ,
         rml_save_e , rml_thr_d[3] , rml_tid_e[0] , rml_tid_e[1] ,
         rml_tid_d[0] , rml_tid_d[1] , rml_rml_reset_l ,
         bypass_irf_write_clkbuf_n1 , bypass_irf_write_clkbuf_clken ,
         bypass_irf_write_clkbuf_N1 , bypass_irf_write_clkbuf_tmb_l ,
         bypass_dfill_data_mux_n129 , bypass_dfill_data_mux_n128 ,
         bypass_dfill_data_mux_n127 , bypass_dfill_data_mux_n126 ,
         bypass_dfill_data_mux_n125 , bypass_dfill_data_mux_n124 ,
         bypass_dfill_data_mux_n123 , bypass_dfill_data_mux_n122 ,
         bypass_dfill_data_mux_n121 , bypass_dfill_data_mux_n120 ,
         bypass_dfill_data_mux_n119 , bypass_dfill_data_mux_n118 ,
         bypass_dfill_data_mux_n117 , bypass_dfill_data_mux_n116 ,
         bypass_dfill_data_mux_n115 , bypass_dfill_data_mux_n114 ,
         bypass_dfill_data_mux_n113 , bypass_dfill_data_mux_n112 ,
         bypass_dfill_data_mux_n111 , bypass_dfill_data_mux_n110 ,
         bypass_dfill_data_mux_n109 , bypass_dfill_data_mux_n108 ,
         bypass_dfill_data_mux_n107 , bypass_dfill_data_mux_n106 ,
         bypass_dfill_data_mux_n105 , bypass_dfill_data_mux_n104 ,
         bypass_dfill_data_mux_n103 , bypass_dfill_data_mux_n102 ,
         bypass_dfill_data_mux_n101 , bypass_dfill_data_mux_n100 ,
         bypass_dfill_data_mux_n99 , bypass_dfill_data_mux_n98 ,
         bypass_dfill_data_mux_n97 , bypass_dfill_data_mux_n96 ,
         bypass_dfill_data_mux_n95 , bypass_dfill_data_mux_n94 ,
         bypass_dfill_data_mux_n93 , bypass_dfill_data_mux_n92 ,
         bypass_dfill_data_mux_n91 , bypass_dfill_data_mux_n90 ,
         bypass_dfill_data_mux_n89 , bypass_dfill_data_mux_n88 ,
         bypass_dfill_data_mux_n87 , bypass_dfill_data_mux_n86 ,
         bypass_dfill_data_mux_n85 , bypass_dfill_data_mux_n84 ,
         bypass_dfill_data_mux_n83 , bypass_dfill_data_mux_n82 ,
         bypass_dfill_data_mux_n81 , bypass_dfill_data_mux_n80 ,
         bypass_dfill_data_mux_n79 , bypass_dfill_data_mux_n78 ,
         bypass_dfill_data_mux_n77 , bypass_dfill_data_mux_n76 ,
         bypass_dfill_data_mux_n75 , bypass_dfill_data_mux_n74 ,
         bypass_dfill_data_mux_n73 , bypass_dfill_data_mux_n72 ,
         bypass_dfill_data_mux_n71 , bypass_dfill_data_mux_n70 ,
         bypass_dfill_data_mux_n69 , bypass_dfill_data_mux_n68 ,
         bypass_dfill_data_mux_n67 , bypass_dfill_data_mux_n66 ,
         bypass_dfill_data_mux_n65 , bypass_dfill_data_mux_n64 ,
         bypass_dfill_data_mux_n63 , bypass_dfill_data_mux_n62 ,
         bypass_dfill_data_mux_n61 , bypass_dfill_data_mux_n60 ,
         bypass_dfill_data_mux_n59 , bypass_dfill_data_mux_n58 ,
         bypass_dfill_data_mux_n57 , bypass_dfill_data_mux_n56 ,
         bypass_dfill_data_mux_n55 , bypass_dfill_data_mux_n54 ,
         bypass_dfill_data_mux_n53 , bypass_dfill_data_mux_n52 ,
         bypass_dfill_data_mux_n51 , bypass_dfill_data_mux_n50 ,
         bypass_dfill_data_mux_n49 , bypass_dfill_data_mux_n48 ,
         bypass_dfill_data_mux_n47 , bypass_dfill_data_mux_n46 ,
         bypass_dfill_data_mux_n45 , bypass_dfill_data_mux_n44 ,
         bypass_dfill_data_mux_n43 , bypass_dfill_data_mux_n42 ,
         bypass_dfill_data_mux_n41 , bypass_dfill_data_mux_n40 ,
         bypass_dfill_data_mux_n39 , bypass_dfill_data_mux_n38 ,
         bypass_dfill_data_mux_n37 , bypass_dfill_data_mux_n36 ,
         bypass_dfill_data_mux_n35 , bypass_dfill_data_mux_n34 ,
         bypass_dfill_data_mux_n33 , bypass_dfill_data_mux_n32 ,
         bypass_dfill_data_mux_n31 , bypass_dfill_data_mux_n30 ,
         bypass_dfill_data_mux_n29 , bypass_dfill_data_mux_n28 ,
         bypass_dfill_data_mux_n27 , bypass_dfill_data_mux_n26 ,
         bypass_dfill_data_mux_n25 , bypass_dfill_data_mux_n24 ,
         bypass_dfill_data_mux_n23 , bypass_dfill_data_mux_n22 ,
         bypass_dfill_data_mux_n21 , bypass_dfill_data_mux_n20 ,
         bypass_dfill_data_mux_n19 , bypass_dfill_data_mux_n18 ,
         bypass_dfill_data_mux_n17 , bypass_dfill_data_mux_n16 ,
         bypass_dfill_data_mux_n15 , bypass_dfill_data_mux_n14 ,
         bypass_dfill_data_mux_n13 , bypass_dfill_data_mux_n12 ,
         bypass_dfill_data_mux_n11 , bypass_dfill_data_mux_n10 ,
         bypass_dfill_data_mux_n9 , bypass_dfill_data_mux_n8 ,
         bypass_dfill_data_mux_n7 , bypass_dfill_data_mux_n6 ,
         bypass_dfill_data_mux_n5 , bypass_dfill_data_mux_n4 ,
         bypass_dfill_data_mux_n3 , bypass_dfill_data_mux_n2 ,
         bypass_dfill_data_dff_n129 , bypass_dfill_data_dff_n127 ,
         bypass_dfill_data_dff_n125 , bypass_dfill_data_dff_n123 ,
         bypass_dfill_data_dff_n121 , bypass_dfill_data_dff_n119 ,
         bypass_dfill_data_dff_n117 , bypass_dfill_data_dff_n115 ,
         bypass_dfill_data_dff_n113 , bypass_dfill_data_dff_n111 ,
         bypass_dfill_data_dff_n109 , bypass_dfill_data_dff_n107 ,
         bypass_dfill_data_dff_n105 , bypass_dfill_data_dff_n103 ,
         bypass_dfill_data_dff_n101 , bypass_dfill_data_dff_n99 ,
         bypass_dfill_data_dff_n97 , bypass_dfill_data_dff_n95 ,
         bypass_dfill_data_dff_n93 , bypass_dfill_data_dff_n91 ,
         bypass_dfill_data_dff_n89 , bypass_dfill_data_dff_n87 ,
         bypass_dfill_data_dff_n85 , bypass_dfill_data_dff_n83 ,
         bypass_dfill_data_dff_n81 , bypass_dfill_data_dff_n79 ,
         bypass_dfill_data_dff_n77 , bypass_dfill_data_dff_n75 ,
         bypass_dfill_data_dff_n73 , bypass_dfill_data_dff_n71 ,
         bypass_dfill_data_dff_n69 , bypass_dfill_data_dff_n67 ,
         bypass_dfill_data_dff_n65 , bypass_dfill_data_dff_n63 ,
         bypass_dfill_data_dff_n61 , bypass_dfill_data_dff_n59 ,
         bypass_dfill_data_dff_n57 , bypass_dfill_data_dff_n55 ,
         bypass_dfill_data_dff_n53 , bypass_dfill_data_dff_n51 ,
         bypass_dfill_data_dff_n49 , bypass_dfill_data_dff_n47 ,
         bypass_dfill_data_dff_n45 , bypass_dfill_data_dff_n43 ,
         bypass_dfill_data_dff_n41 , bypass_dfill_data_dff_n39 ,
         bypass_dfill_data_dff_n37 , bypass_dfill_data_dff_n35 ,
         bypass_dfill_data_dff_n33 , bypass_dfill_data_dff_n31 ,
         bypass_dfill_data_dff_n29 , bypass_dfill_data_dff_n27 ,
         bypass_dfill_data_dff_n25 , bypass_dfill_data_dff_n23 ,
         bypass_dfill_data_dff_n21 , bypass_dfill_data_dff_n19 ,
         bypass_dfill_data_dff_n17 , bypass_dfill_data_dff_n15 ,
         bypass_dfill_data_dff_n13 , bypass_dfill_data_dff_n11 ,
         bypass_dfill_data_dff_n9 , bypass_dfill_data_dff_n7 ,
         bypass_dfill_data_dff_n5 , bypass_dfill_data_dff_n3 ,
         bypass_dfill_data_dff_n1 , bypass_ifu_exu_sr_mux_n384 ,
         bypass_ifu_exu_sr_mux_n383 , bypass_ifu_exu_sr_mux_n382 ,
         bypass_ifu_exu_sr_mux_n381 , bypass_ifu_exu_sr_mux_n380 ,
         bypass_ifu_exu_sr_mux_n379 , bypass_ifu_exu_sr_mux_n378 ,
         bypass_ifu_exu_sr_mux_n376 , bypass_ifu_exu_sr_mux_n375 ,
         bypass_ifu_exu_sr_mux_n374 , bypass_ifu_exu_sr_mux_n372 ,
         bypass_ifu_exu_sr_mux_n370 , bypass_ifu_exu_sr_mux_n369 ,
         bypass_ifu_exu_sr_mux_n368 , bypass_ifu_exu_sr_mux_n366 ,
         bypass_ifu_exu_sr_mux_n364 , bypass_ifu_exu_sr_mux_n363 ,
         bypass_ifu_exu_sr_mux_n362 , bypass_ifu_exu_sr_mux_n360 ,
         bypass_ifu_exu_sr_mux_n358 , bypass_ifu_exu_sr_mux_n357 ,
         bypass_ifu_exu_sr_mux_n356 , bypass_ifu_exu_sr_mux_n354 ,
         bypass_ifu_exu_sr_mux_n352 , bypass_ifu_exu_sr_mux_n351 ,
         bypass_ifu_exu_sr_mux_n350 , bypass_ifu_exu_sr_mux_n348 ,
         bypass_ifu_exu_sr_mux_n346 , bypass_ifu_exu_sr_mux_n345 ,
         bypass_ifu_exu_sr_mux_n344 , bypass_ifu_exu_sr_mux_n342 ,
         bypass_ifu_exu_sr_mux_n340 , bypass_ifu_exu_sr_mux_n339 ,
         bypass_ifu_exu_sr_mux_n338 , bypass_ifu_exu_sr_mux_n336 ,
         bypass_ifu_exu_sr_mux_n334 , bypass_ifu_exu_sr_mux_n333 ,
         bypass_ifu_exu_sr_mux_n332 , bypass_ifu_exu_sr_mux_n330 ,
         bypass_ifu_exu_sr_mux_n328 , bypass_ifu_exu_sr_mux_n327 ,
         bypass_ifu_exu_sr_mux_n326 , bypass_ifu_exu_sr_mux_n324 ,
         bypass_ifu_exu_sr_mux_n322 , bypass_ifu_exu_sr_mux_n321 ,
         bypass_ifu_exu_sr_mux_n320 , bypass_ifu_exu_sr_mux_n318 ,
         bypass_ifu_exu_sr_mux_n317 , bypass_ifu_exu_sr_mux_n316 ,
         bypass_ifu_exu_sr_mux_n315 , bypass_ifu_exu_sr_mux_n314 ,
         bypass_ifu_exu_sr_mux_n313 , bypass_ifu_exu_sr_mux_n312 ,
         bypass_ifu_exu_sr_mux_n310 , bypass_ifu_exu_sr_mux_n309 ,
         bypass_ifu_exu_sr_mux_n308 , bypass_ifu_exu_sr_mux_n306 ,
         bypass_ifu_exu_sr_mux_n304 , bypass_ifu_exu_sr_mux_n303 ,
         bypass_ifu_exu_sr_mux_n302 , bypass_ifu_exu_sr_mux_n300 ,
         bypass_ifu_exu_sr_mux_n298 , bypass_ifu_exu_sr_mux_n297 ,
         bypass_ifu_exu_sr_mux_n296 , bypass_ifu_exu_sr_mux_n294 ,
         bypass_ifu_exu_sr_mux_n292 , bypass_ifu_exu_sr_mux_n291 ,
         bypass_ifu_exu_sr_mux_n290 , bypass_ifu_exu_sr_mux_n288 ,
         bypass_ifu_exu_sr_mux_n286 , bypass_ifu_exu_sr_mux_n285 ,
         bypass_ifu_exu_sr_mux_n284 , bypass_ifu_exu_sr_mux_n282 ,
         bypass_ifu_exu_sr_mux_n280 , bypass_ifu_exu_sr_mux_n279 ,
         bypass_ifu_exu_sr_mux_n278 , bypass_ifu_exu_sr_mux_n276 ,
         bypass_ifu_exu_sr_mux_n274 , bypass_ifu_exu_sr_mux_n273 ,
         bypass_ifu_exu_sr_mux_n272 , bypass_ifu_exu_sr_mux_n270 ,
         bypass_ifu_exu_sr_mux_n268 , bypass_ifu_exu_sr_mux_n267 ,
         bypass_ifu_exu_sr_mux_n266 , bypass_ifu_exu_sr_mux_n264 ,
         bypass_ifu_exu_sr_mux_n262 , bypass_ifu_exu_sr_mux_n261 ,
         bypass_ifu_exu_sr_mux_n260 , bypass_ifu_exu_sr_mux_n258 ,
         bypass_ifu_exu_sr_mux_n256 , bypass_ifu_exu_sr_mux_n255 ,
         bypass_ifu_exu_sr_mux_n254 , bypass_ifu_exu_sr_mux_n252 ,
         bypass_ifu_exu_sr_mux_n251 , bypass_ifu_exu_sr_mux_n250 ,
         bypass_ifu_exu_sr_mux_n249 , bypass_ifu_exu_sr_mux_n248 ,
         bypass_ifu_exu_sr_mux_n247 , bypass_ifu_exu_sr_mux_n246 ,
         bypass_ifu_exu_sr_mux_n244 , bypass_ifu_exu_sr_mux_n243 ,
         bypass_ifu_exu_sr_mux_n242 , bypass_ifu_exu_sr_mux_n240 ,
         bypass_ifu_exu_sr_mux_n238 , bypass_ifu_exu_sr_mux_n237 ,
         bypass_ifu_exu_sr_mux_n236 , bypass_ifu_exu_sr_mux_n232 ,
         bypass_ifu_exu_sr_mux_n231 , bypass_ifu_exu_sr_mux_n230 ,
         bypass_ifu_exu_sr_mux_n226 , bypass_ifu_exu_sr_mux_n225 ,
         bypass_ifu_exu_sr_mux_n224 , bypass_ifu_exu_sr_mux_n220 ,
         bypass_ifu_exu_sr_mux_n219 , bypass_ifu_exu_sr_mux_n218 ,
         bypass_ifu_exu_sr_mux_n214 , bypass_ifu_exu_sr_mux_n213 ,
         bypass_ifu_exu_sr_mux_n212 , bypass_ifu_exu_sr_mux_n208 ,
         bypass_ifu_exu_sr_mux_n207 , bypass_ifu_exu_sr_mux_n206 ,
         bypass_ifu_exu_sr_mux_n202 , bypass_ifu_exu_sr_mux_n201 ,
         bypass_ifu_exu_sr_mux_n200 , bypass_ifu_exu_sr_mux_n196 ,
         bypass_ifu_exu_sr_mux_n195 , bypass_ifu_exu_sr_mux_n194 ,
         bypass_ifu_exu_sr_mux_n190 , bypass_ifu_exu_sr_mux_n189 ,
         bypass_ifu_exu_sr_mux_n188 , bypass_ifu_exu_sr_mux_n186 ,
         bypass_ifu_exu_sr_mux_n185 , bypass_ifu_exu_sr_mux_n184 ,
         bypass_ifu_exu_sr_mux_n183 , bypass_ifu_exu_sr_mux_n182 ,
         bypass_ifu_exu_sr_mux_n181 , bypass_ifu_exu_sr_mux_n178 ,
         bypass_ifu_exu_sr_mux_n177 , bypass_ifu_exu_sr_mux_n176 ,
         bypass_ifu_exu_sr_mux_n172 , bypass_ifu_exu_sr_mux_n171 ,
         bypass_ifu_exu_sr_mux_n170 , bypass_ifu_exu_sr_mux_n166 ,
         bypass_ifu_exu_sr_mux_n165 , bypass_ifu_exu_sr_mux_n164 ,
         bypass_ifu_exu_sr_mux_n160 , bypass_ifu_exu_sr_mux_n159 ,
         bypass_ifu_exu_sr_mux_n158 , bypass_ifu_exu_sr_mux_n154 ,
         bypass_ifu_exu_sr_mux_n153 , bypass_ifu_exu_sr_mux_n152 ,
         bypass_ifu_exu_sr_mux_n148 , bypass_ifu_exu_sr_mux_n147 ,
         bypass_ifu_exu_sr_mux_n146 , bypass_ifu_exu_sr_mux_n142 ,
         bypass_ifu_exu_sr_mux_n141 , bypass_ifu_exu_sr_mux_n140 ,
         bypass_ifu_exu_sr_mux_n136 , bypass_ifu_exu_sr_mux_n135 ,
         bypass_ifu_exu_sr_mux_n134 , bypass_ifu_exu_sr_mux_n130 ,
         bypass_ifu_exu_sr_mux_n129 , bypass_ifu_exu_sr_mux_n128 ,
         bypass_ifu_exu_sr_mux_n124 , bypass_ifu_exu_sr_mux_n123 ,
         bypass_ifu_exu_sr_mux_n122 , bypass_ifu_exu_sr_mux_n120 ,
         bypass_ifu_exu_sr_mux_n119 , bypass_ifu_exu_sr_mux_n118 ,
         bypass_ifu_exu_sr_mux_n117 , bypass_ifu_exu_sr_mux_n116 ,
         bypass_ifu_exu_sr_mux_n115 , bypass_ifu_exu_sr_mux_n112 ,
         bypass_ifu_exu_sr_mux_n111 , bypass_ifu_exu_sr_mux_n110 ,
         bypass_ifu_exu_sr_mux_n106 , bypass_ifu_exu_sr_mux_n105 ,
         bypass_ifu_exu_sr_mux_n104 , bypass_ifu_exu_sr_mux_n100 ,
         bypass_ifu_exu_sr_mux_n99 , bypass_ifu_exu_sr_mux_n98 ,
         bypass_ifu_exu_sr_mux_n94 , bypass_ifu_exu_sr_mux_n93 ,
         bypass_ifu_exu_sr_mux_n92 , bypass_ifu_exu_sr_mux_n88 ,
         bypass_ifu_exu_sr_mux_n87 , bypass_ifu_exu_sr_mux_n86 ,
         bypass_ifu_exu_sr_mux_n82 , bypass_ifu_exu_sr_mux_n81 ,
         bypass_ifu_exu_sr_mux_n80 , bypass_ifu_exu_sr_mux_n76 ,
         bypass_ifu_exu_sr_mux_n75 , bypass_ifu_exu_sr_mux_n74 ,
         bypass_ifu_exu_sr_mux_n70 , bypass_ifu_exu_sr_mux_n69 ,
         bypass_ifu_exu_sr_mux_n68 , bypass_ifu_exu_sr_mux_n64 ,
         bypass_ifu_exu_sr_mux_n63 , bypass_ifu_exu_sr_mux_n62 ,
         bypass_ifu_exu_sr_mux_n58 , bypass_ifu_exu_sr_mux_n57 ,
         bypass_ifu_exu_sr_mux_n56 , bypass_ifu_exu_sr_mux_n54 ,
         bypass_ifu_exu_sr_mux_n53 , bypass_ifu_exu_sr_mux_n52 ,
         bypass_ifu_exu_sr_mux_n51 , bypass_ifu_exu_sr_mux_n50 ,
         bypass_ifu_exu_sr_mux_n49 , bypass_ifu_exu_sr_mux_n46 ,
         bypass_ifu_exu_sr_mux_n45 , bypass_ifu_exu_sr_mux_n44 ,
         bypass_ifu_exu_sr_mux_n40 , bypass_ifu_exu_sr_mux_n39 ,
         bypass_ifu_exu_sr_mux_n38 , bypass_ifu_exu_sr_mux_n34 ,
         bypass_ifu_exu_sr_mux_n33 , bypass_ifu_exu_sr_mux_n32 ,
         bypass_ifu_exu_sr_mux_n28 , bypass_ifu_exu_sr_mux_n27 ,
         bypass_ifu_exu_sr_mux_n26 , bypass_ifu_exu_sr_mux_n24 ,
         bypass_ifu_exu_sr_mux_n23 , bypass_ifu_exu_sr_mux_n22 ,
         bypass_ifu_exu_sr_mux_n21 , bypass_ifu_exu_sr_mux_n20 ,
         bypass_ifu_exu_sr_mux_n19 , bypass_ifu_exu_sr_mux_n18 ,
         bypass_ifu_exu_sr_mux_n17 , bypass_ifu_exu_sr_mux_n16 ,
         bypass_ifu_exu_sr_mux_n15 , bypass_ifu_exu_sr_mux_n14 ,
         bypass_ifu_exu_sr_mux_n13 , bypass_ifu_exu_sr_mux_n12 ,
         bypass_ifu_exu_sr_mux_n10 , bypass_ifu_exu_sr_mux_n9 ,
         bypass_ifu_exu_sr_mux_n8 , bypass_ifu_exu_sr_mux_n6 ,
         bypass_ifu_exu_sr_mux_n4 , bypass_ifu_exu_sr_mux_n3 ,
         bypass_ifu_exu_sr_mux_n2 , bypass_sr_out_mux_n256 ,
         bypass_sr_out_mux_n255 , bypass_sr_out_mux_n254 ,
         bypass_sr_out_mux_n253 , bypass_sr_out_mux_n252 ,
         bypass_sr_out_mux_n251 , bypass_sr_out_mux_n250 ,
         bypass_sr_out_mux_n249 , bypass_sr_out_mux_n248 ,
         bypass_sr_out_mux_n247 , bypass_sr_out_mux_n246 ,
         bypass_sr_out_mux_n245 , bypass_sr_out_mux_n244 ,
         bypass_sr_out_mux_n243 , bypass_sr_out_mux_n242 ,
         bypass_sr_out_mux_n241 , bypass_sr_out_mux_n240 ,
         bypass_sr_out_mux_n239 , bypass_sr_out_mux_n238 ,
         bypass_sr_out_mux_n237 , bypass_sr_out_mux_n236 ,
         bypass_sr_out_mux_n235 , bypass_sr_out_mux_n234 ,
         bypass_sr_out_mux_n233 , bypass_sr_out_mux_n232 ,
         bypass_sr_out_mux_n231 , bypass_sr_out_mux_n230 ,
         bypass_sr_out_mux_n229 , bypass_sr_out_mux_n228 ,
         bypass_sr_out_mux_n227 , bypass_sr_out_mux_n226 ,
         bypass_sr_out_mux_n225 , bypass_sr_out_mux_n224 ,
         bypass_sr_out_mux_n223 , bypass_sr_out_mux_n222 ,
         bypass_sr_out_mux_n221 , bypass_sr_out_mux_n220 ,
         bypass_sr_out_mux_n219 , bypass_sr_out_mux_n218 ,
         bypass_sr_out_mux_n217 , bypass_sr_out_mux_n216 ,
         bypass_sr_out_mux_n215 , bypass_sr_out_mux_n214 ,
         bypass_sr_out_mux_n213 , bypass_sr_out_mux_n212 ,
         bypass_sr_out_mux_n211 , bypass_sr_out_mux_n210 ,
         bypass_sr_out_mux_n209 , bypass_sr_out_mux_n208 ,
         bypass_sr_out_mux_n207 , bypass_sr_out_mux_n206 ,
         bypass_sr_out_mux_n205 , bypass_sr_out_mux_n204 ,
         bypass_sr_out_mux_n203 , bypass_sr_out_mux_n202 ,
         bypass_sr_out_mux_n201 , bypass_sr_out_mux_n200 ,
         bypass_sr_out_mux_n199 , bypass_sr_out_mux_n198 ,
         bypass_sr_out_mux_n197 , bypass_sr_out_mux_n196 ,
         bypass_sr_out_mux_n195 , bypass_sr_out_mux_n194 ,
         bypass_sr_out_mux_n193 , bypass_sr_out_mux_n192 ,
         bypass_sr_out_mux_n191 , bypass_sr_out_mux_n190 ,
         bypass_sr_out_mux_n189 , bypass_sr_out_mux_n188 ,
         bypass_sr_out_mux_n187 , bypass_sr_out_mux_n186 ,
         bypass_sr_out_mux_n185 , bypass_sr_out_mux_n184 ,
         bypass_sr_out_mux_n183 , bypass_sr_out_mux_n182 ,
         bypass_sr_out_mux_n181 , bypass_sr_out_mux_n180 ,
         bypass_sr_out_mux_n179 , bypass_sr_out_mux_n178 ,
         bypass_sr_out_mux_n177 , bypass_sr_out_mux_n176 ,
         bypass_sr_out_mux_n175 , bypass_sr_out_mux_n174 ,
         bypass_sr_out_mux_n173 , bypass_sr_out_mux_n172 ,
         bypass_sr_out_mux_n171 , bypass_sr_out_mux_n170 ,
         bypass_sr_out_mux_n169 , bypass_sr_out_mux_n168 ,
         bypass_sr_out_mux_n167 , bypass_sr_out_mux_n166 ,
         bypass_sr_out_mux_n165 , bypass_sr_out_mux_n164 ,
         bypass_sr_out_mux_n163 , bypass_sr_out_mux_n162 ,
         bypass_sr_out_mux_n161 , bypass_sr_out_mux_n160 ,
         bypass_sr_out_mux_n159 , bypass_sr_out_mux_n158 ,
         bypass_sr_out_mux_n157 , bypass_sr_out_mux_n156 ,
         bypass_sr_out_mux_n155 , bypass_sr_out_mux_n154 ,
         bypass_sr_out_mux_n153 , bypass_sr_out_mux_n152 ,
         bypass_sr_out_mux_n151 , bypass_sr_out_mux_n150 ,
         bypass_sr_out_mux_n149 , bypass_sr_out_mux_n148 ,
         bypass_sr_out_mux_n147 , bypass_sr_out_mux_n146 ,
         bypass_sr_out_mux_n145 , bypass_sr_out_mux_n144 ,
         bypass_sr_out_mux_n143 , bypass_sr_out_mux_n142 ,
         bypass_sr_out_mux_n141 , bypass_sr_out_mux_n140 ,
         bypass_sr_out_mux_n139 , bypass_sr_out_mux_n138 ,
         bypass_sr_out_mux_n137 , bypass_sr_out_mux_n136 ,
         bypass_sr_out_mux_n135 , bypass_sr_out_mux_n134 ,
         bypass_sr_out_mux_n133 , bypass_sr_out_mux_n132 ,
         bypass_sr_out_mux_n131 , bypass_sr_out_mux_n130 ,
         bypass_sr_out_mux_n129 , bypass_sr_out_mux_n128 ,
         bypass_sr_out_mux_n127 , bypass_sr_out_mux_n126 ,
         bypass_sr_out_mux_n125 , bypass_sr_out_mux_n124 ,
         bypass_sr_out_mux_n123 , bypass_sr_out_mux_n122 ,
         bypass_sr_out_mux_n121 , bypass_sr_out_mux_n120 ,
         bypass_sr_out_mux_n119 , bypass_sr_out_mux_n118 ,
         bypass_sr_out_mux_n117 , bypass_sr_out_mux_n116 ,
         bypass_sr_out_mux_n115 , bypass_sr_out_mux_n114 ,
         bypass_sr_out_mux_n113 , bypass_sr_out_mux_n112 ,
         bypass_sr_out_mux_n111 , bypass_sr_out_mux_n110 ,
         bypass_sr_out_mux_n109 , bypass_sr_out_mux_n108 ,
         bypass_sr_out_mux_n107 , bypass_sr_out_mux_n106 ,
         bypass_sr_out_mux_n105 , bypass_sr_out_mux_n104 ,
         bypass_sr_out_mux_n103 , bypass_sr_out_mux_n102 ,
         bypass_sr_out_mux_n101 , bypass_sr_out_mux_n100 ,
         bypass_sr_out_mux_n99 , bypass_sr_out_mux_n98 ,
         bypass_sr_out_mux_n97 , bypass_sr_out_mux_n96 ,
         bypass_sr_out_mux_n95 , bypass_sr_out_mux_n94 ,
         bypass_sr_out_mux_n93 , bypass_sr_out_mux_n92 ,
         bypass_sr_out_mux_n91 , bypass_sr_out_mux_n90 ,
         bypass_sr_out_mux_n89 , bypass_sr_out_mux_n88 ,
         bypass_sr_out_mux_n87 , bypass_sr_out_mux_n86 ,
         bypass_sr_out_mux_n85 , bypass_sr_out_mux_n84 ,
         bypass_sr_out_mux_n83 , bypass_sr_out_mux_n82 ,
         bypass_sr_out_mux_n81 , bypass_sr_out_mux_n80 ,
         bypass_sr_out_mux_n79 , bypass_sr_out_mux_n78 ,
         bypass_sr_out_mux_n77 , bypass_sr_out_mux_n76 ,
         bypass_sr_out_mux_n75 , bypass_sr_out_mux_n74 ,
         bypass_sr_out_mux_n73 , bypass_sr_out_mux_n72 ,
         bypass_sr_out_mux_n71 , bypass_sr_out_mux_n70 ,
         bypass_sr_out_mux_n69 , bypass_sr_out_mux_n68 ,
         bypass_sr_out_mux_n67 , bypass_sr_out_mux_n66 ,
         bypass_sr_out_mux_n65 , bypass_sr_out_mux_n64 ,
         bypass_sr_out_mux_n63 , bypass_sr_out_mux_n62 ,
         bypass_sr_out_mux_n61 , bypass_sr_out_mux_n60 ,
         bypass_sr_out_mux_n59 , bypass_sr_out_mux_n58 ,
         bypass_sr_out_mux_n57 , bypass_sr_out_mux_n56 ,
         bypass_sr_out_mux_n55 , bypass_sr_out_mux_n54 ,
         bypass_sr_out_mux_n53 , bypass_sr_out_mux_n52 ,
         bypass_sr_out_mux_n51 , bypass_sr_out_mux_n50 ,
         bypass_sr_out_mux_n49 , bypass_sr_out_mux_n48 ,
         bypass_sr_out_mux_n47 , bypass_sr_out_mux_n46 ,
         bypass_sr_out_mux_n45 , bypass_sr_out_mux_n44 ,
         bypass_sr_out_mux_n43 , bypass_sr_out_mux_n42 ,
         bypass_sr_out_mux_n41 , bypass_sr_out_mux_n40 ,
         bypass_sr_out_mux_n39 , bypass_sr_out_mux_n38 ,
         bypass_sr_out_mux_n37 , bypass_sr_out_mux_n36 ,
         bypass_sr_out_mux_n35 , bypass_sr_out_mux_n34 ,
         bypass_sr_out_mux_n33 , bypass_sr_out_mux_n32 ,
         bypass_sr_out_mux_n31 , bypass_sr_out_mux_n30 ,
         bypass_sr_out_mux_n29 , bypass_sr_out_mux_n28 ,
         bypass_sr_out_mux_n27 , bypass_sr_out_mux_n26 ,
         bypass_sr_out_mux_n25 , bypass_sr_out_mux_n24 ,
         bypass_sr_out_mux_n23 , bypass_sr_out_mux_n22 ,
         bypass_sr_out_mux_n21 , bypass_sr_out_mux_n20 ,
         bypass_sr_out_mux_n19 , bypass_sr_out_mux_n18 ,
         bypass_sr_out_mux_n17 , bypass_sr_out_mux_n16 ,
         bypass_sr_out_mux_n15 , bypass_sr_out_mux_n14 ,
         bypass_sr_out_mux_n13 , bypass_sr_out_mux_n12 ,
         bypass_sr_out_mux_n11 , bypass_sr_out_mux_n10 ,
         bypass_sr_out_mux_n9 , bypass_sr_out_mux_n8 ,
         bypass_sr_out_mux_n7 , bypass_sr_out_mux_n6 ,
         bypass_sr_out_mux_n5 , bypass_sr_out_mux_n4 ,
         bypass_sr_out_mux_n3 , bypass_sr_out_mux_n2 ,
         bypass_sr_out_mux_n1 , bypass_rs3h_data_dff_n65 ,
         bypass_rs3h_data_dff_n63 , bypass_rs3h_data_dff_n61 ,
         bypass_rs3h_data_dff_n59 , bypass_rs3h_data_dff_n57 ,
         bypass_rs3h_data_dff_n55 , bypass_rs3h_data_dff_n53 ,
         bypass_rs3h_data_dff_n51 , bypass_rs3h_data_dff_n49 ,
         bypass_rs3h_data_dff_n47 , bypass_rs3h_data_dff_n45 ,
         bypass_rs3h_data_dff_n43 , bypass_rs3h_data_dff_n41 ,
         bypass_rs3h_data_dff_n39 , bypass_rs3h_data_dff_n37 ,
         bypass_rs3h_data_dff_n35 , bypass_rs3h_data_dff_n33 ,
         bypass_rs3h_data_dff_n31 , bypass_rs3h_data_dff_n29 ,
         bypass_rs3h_data_dff_n27 , bypass_rs3h_data_dff_n25 ,
         bypass_rs3h_data_dff_n23 , bypass_rs3h_data_dff_n21 ,
         bypass_rs3h_data_dff_n19 , bypass_rs3h_data_dff_n17 ,
         bypass_rs3h_data_dff_n15 , bypass_rs3h_data_dff_n13 ,
         bypass_rs3h_data_dff_n11 , bypass_rs3h_data_dff_n9 ,
         bypass_rs3h_data_dff_n7 , bypass_rs3h_data_dff_n5 ,
         bypass_rs3h_data_dff_n3 , bypass_rs3h_data_dff_n1 ,
         bypass_rs3h_w2_mux_n128 , bypass_rs3h_w2_mux_n127 ,
         bypass_rs3h_w2_mux_n126 , bypass_rs3h_w2_mux_n125 ,
         bypass_rs3h_w2_mux_n124 , bypass_rs3h_w2_mux_n123 ,
         bypass_rs3h_w2_mux_n122 , bypass_rs3h_w2_mux_n121 ,
         bypass_rs3h_w2_mux_n120 , bypass_rs3h_w2_mux_n119 ,
         bypass_rs3h_w2_mux_n118 , bypass_rs3h_w2_mux_n117 ,
         bypass_rs3h_w2_mux_n116 , bypass_rs3h_w2_mux_n115 ,
         bypass_rs3h_w2_mux_n114 , bypass_rs3h_w2_mux_n113 ,
         bypass_rs3h_w2_mux_n112 , bypass_rs3h_w2_mux_n111 ,
         bypass_rs3h_w2_mux_n110 , bypass_rs3h_w2_mux_n109 ,
         bypass_rs3h_w2_mux_n108 , bypass_rs3h_w2_mux_n107 ,
         bypass_rs3h_w2_mux_n106 , bypass_rs3h_w2_mux_n105 ,
         bypass_rs3h_w2_mux_n104 , bypass_rs3h_w2_mux_n103 ,
         bypass_rs3h_w2_mux_n102 , bypass_rs3h_w2_mux_n101 ,
         bypass_rs3h_w2_mux_n100 , bypass_rs3h_w2_mux_n99 ,
         bypass_rs3h_w2_mux_n98 , bypass_rs3h_w2_mux_n97 ,
         bypass_rs3h_w2_mux_n96 , bypass_rs3h_w2_mux_n95 ,
         bypass_rs3h_w2_mux_n94 , bypass_rs3h_w2_mux_n93 ,
         bypass_rs3h_w2_mux_n92 , bypass_rs3h_w2_mux_n91 ,
         bypass_rs3h_w2_mux_n90 , bypass_rs3h_w2_mux_n89 ,
         bypass_rs3h_w2_mux_n88 , bypass_rs3h_w2_mux_n87 ,
         bypass_rs3h_w2_mux_n86 , bypass_rs3h_w2_mux_n85 ,
         bypass_rs3h_w2_mux_n84 , bypass_rs3h_w2_mux_n83 ,
         bypass_rs3h_w2_mux_n82 , bypass_rs3h_w2_mux_n81 ,
         bypass_rs3h_w2_mux_n80 , bypass_rs3h_w2_mux_n79 ,
         bypass_rs3h_w2_mux_n78 , bypass_rs3h_w2_mux_n77 ,
         bypass_rs3h_w2_mux_n76 , bypass_rs3h_w2_mux_n75 ,
         bypass_rs3h_w2_mux_n74 , bypass_rs3h_w2_mux_n73 ,
         bypass_rs3h_w2_mux_n72 , bypass_rs3h_w2_mux_n71 ,
         bypass_rs3h_w2_mux_n70 , bypass_rs3h_w2_mux_n69 ,
         bypass_rs3h_w2_mux_n68 , bypass_rs3h_w2_mux_n67 ,
         bypass_rs3h_w2_mux_n66 , bypass_rs3h_w2_mux_n65 ,
         bypass_rs3h_w2_mux_n64 , bypass_rs3h_w2_mux_n63 ,
         bypass_rs3h_w2_mux_n62 , bypass_rs3h_w2_mux_n61 ,
         bypass_rs3h_w2_mux_n60 , bypass_rs3h_w2_mux_n59 ,
         bypass_rs3h_w2_mux_n58 , bypass_rs3h_w2_mux_n57 ,
         bypass_rs3h_w2_mux_n56 , bypass_rs3h_w2_mux_n55 ,
         bypass_rs3h_w2_mux_n54 , bypass_rs3h_w2_mux_n53 ,
         bypass_rs3h_w2_mux_n52 , bypass_rs3h_w2_mux_n51 ,
         bypass_rs3h_w2_mux_n50 , bypass_rs3h_w2_mux_n49 ,
         bypass_rs3h_w2_mux_n48 , bypass_rs3h_w2_mux_n47 ,
         bypass_rs3h_w2_mux_n46 , bypass_rs3h_w2_mux_n45 ,
         bypass_rs3h_w2_mux_n44 , bypass_rs3h_w2_mux_n43 ,
         bypass_rs3h_w2_mux_n42 , bypass_rs3h_w2_mux_n41 ,
         bypass_rs3h_w2_mux_n40 , bypass_rs3h_w2_mux_n39 ,
         bypass_rs3h_w2_mux_n38 , bypass_rs3h_w2_mux_n37 ,
         bypass_rs3h_w2_mux_n36 , bypass_rs3h_w2_mux_n35 ,
         bypass_rs3h_w2_mux_n34 , bypass_rs3h_w2_mux_n33 ,
         bypass_rs3h_w2_mux_n32 , bypass_rs3h_w2_mux_n31 ,
         bypass_rs3h_w2_mux_n30 , bypass_rs3h_w2_mux_n29 ,
         bypass_rs3h_w2_mux_n28 , bypass_rs3h_w2_mux_n27 ,
         bypass_rs3h_w2_mux_n26 , bypass_rs3h_w2_mux_n25 ,
         bypass_rs3h_w2_mux_n24 , bypass_rs3h_w2_mux_n23 ,
         bypass_rs3h_w2_mux_n22 , bypass_rs3h_w2_mux_n21 ,
         bypass_rs3h_w2_mux_n20 , bypass_rs3h_w2_mux_n19 ,
         bypass_rs3h_w2_mux_n18 , bypass_rs3h_w2_mux_n17 ,
         bypass_rs3h_w2_mux_n16 , bypass_rs3h_w2_mux_n15 ,
         bypass_rs3h_w2_mux_n14 , bypass_rs3h_w2_mux_n13 ,
         bypass_rs3h_w2_mux_n12 , bypass_rs3h_w2_mux_n11 ,
         bypass_rs3h_w2_mux_n10 , bypass_rs3h_w2_mux_n9 ,
         bypass_rs3h_w2_mux_n8 , bypass_rs3h_w2_mux_n7 ,
         bypass_rs3h_w2_mux_n6 , bypass_rs3h_w2_mux_n5 ,
         bypass_rs3h_w2_mux_n4 , bypass_rs3h_w2_mux_n3 ,
         bypass_rs3h_w2_mux_n2 , bypass_rs3h_w2_mux_n1 ,
         bypass_mux_rs3h_data_1_n192 , bypass_mux_rs3h_data_1_n191 ,
         bypass_mux_rs3h_data_1_n190 , bypass_mux_rs3h_data_1_n187 ,
         bypass_mux_rs3h_data_1_n186 , bypass_mux_rs3h_data_1_n185 ,
         bypass_mux_rs3h_data_1_n184 , bypass_mux_rs3h_data_1_n181 ,
         bypass_mux_rs3h_data_1_n180 , bypass_mux_rs3h_data_1_n179 ,
         bypass_mux_rs3h_data_1_n178 , bypass_mux_rs3h_data_1_n175 ,
         bypass_mux_rs3h_data_1_n174 , bypass_mux_rs3h_data_1_n173 ,
         bypass_mux_rs3h_data_1_n172 , bypass_mux_rs3h_data_1_n169 ,
         bypass_mux_rs3h_data_1_n168 , bypass_mux_rs3h_data_1_n167 ,
         bypass_mux_rs3h_data_1_n166 , bypass_mux_rs3h_data_1_n163 ,
         bypass_mux_rs3h_data_1_n162 , bypass_mux_rs3h_data_1_n161 ,
         bypass_mux_rs3h_data_1_n160 , bypass_mux_rs3h_data_1_n157 ,
         bypass_mux_rs3h_data_1_n156 , bypass_mux_rs3h_data_1_n155 ,
         bypass_mux_rs3h_data_1_n154 , bypass_mux_rs3h_data_1_n151 ,
         bypass_mux_rs3h_data_1_n150 , bypass_mux_rs3h_data_1_n149 ,
         bypass_mux_rs3h_data_1_n148 , bypass_mux_rs3h_data_1_n145 ,
         bypass_mux_rs3h_data_1_n144 , bypass_mux_rs3h_data_1_n143 ,
         bypass_mux_rs3h_data_1_n142 , bypass_mux_rs3h_data_1_n139 ,
         bypass_mux_rs3h_data_1_n138 , bypass_mux_rs3h_data_1_n137 ,
         bypass_mux_rs3h_data_1_n136 , bypass_mux_rs3h_data_1_n133 ,
         bypass_mux_rs3h_data_1_n132 , bypass_mux_rs3h_data_1_n131 ,
         bypass_mux_rs3h_data_1_n130 , bypass_mux_rs3h_data_1_n127 ,
         bypass_mux_rs3h_data_1_n126 , bypass_mux_rs3h_data_1_n125 ,
         bypass_mux_rs3h_data_1_n124 , bypass_mux_rs3h_data_1_n121 ,
         bypass_mux_rs3h_data_1_n120 , bypass_mux_rs3h_data_1_n119 ,
         bypass_mux_rs3h_data_1_n118 , bypass_mux_rs3h_data_1_n115 ,
         bypass_mux_rs3h_data_1_n114 , bypass_mux_rs3h_data_1_n113 ,
         bypass_mux_rs3h_data_1_n112 , bypass_mux_rs3h_data_1_n109 ,
         bypass_mux_rs3h_data_1_n108 , bypass_mux_rs3h_data_1_n107 ,
         bypass_mux_rs3h_data_1_n106 , bypass_mux_rs3h_data_1_n103 ,
         bypass_mux_rs3h_data_1_n102 , bypass_mux_rs3h_data_1_n101 ,
         bypass_mux_rs3h_data_1_n100 , bypass_mux_rs3h_data_1_n97 ,
         bypass_mux_rs3h_data_1_n96 , bypass_mux_rs3h_data_1_n95 ,
         bypass_mux_rs3h_data_1_n94 , bypass_mux_rs3h_data_1_n91 ,
         bypass_mux_rs3h_data_1_n90 , bypass_mux_rs3h_data_1_n89 ,
         bypass_mux_rs3h_data_1_n88 , bypass_mux_rs3h_data_1_n85 ,
         bypass_mux_rs3h_data_1_n84 , bypass_mux_rs3h_data_1_n83 ,
         bypass_mux_rs3h_data_1_n82 , bypass_mux_rs3h_data_1_n79 ,
         bypass_mux_rs3h_data_1_n78 , bypass_mux_rs3h_data_1_n77 ,
         bypass_mux_rs3h_data_1_n76 , bypass_mux_rs3h_data_1_n73 ,
         bypass_mux_rs3h_data_1_n72 , bypass_mux_rs3h_data_1_n71 ,
         bypass_mux_rs3h_data_1_n70 , bypass_mux_rs3h_data_1_n67 ,
         bypass_mux_rs3h_data_1_n66 , bypass_mux_rs3h_data_1_n65 ,
         bypass_mux_rs3h_data_1_n64 , bypass_mux_rs3h_data_1_n61 ,
         bypass_mux_rs3h_data_1_n60 , bypass_mux_rs3h_data_1_n59 ,
         bypass_mux_rs3h_data_1_n58 , bypass_mux_rs3h_data_1_n55 ,
         bypass_mux_rs3h_data_1_n54 , bypass_mux_rs3h_data_1_n53 ,
         bypass_mux_rs3h_data_1_n52 , bypass_mux_rs3h_data_1_n49 ,
         bypass_mux_rs3h_data_1_n48 , bypass_mux_rs3h_data_1_n47 ,
         bypass_mux_rs3h_data_1_n46 , bypass_mux_rs3h_data_1_n43 ,
         bypass_mux_rs3h_data_1_n42 , bypass_mux_rs3h_data_1_n41 ,
         bypass_mux_rs3h_data_1_n40 , bypass_mux_rs3h_data_1_n37 ,
         bypass_mux_rs3h_data_1_n36 , bypass_mux_rs3h_data_1_n35 ,
         bypass_mux_rs3h_data_1_n34 , bypass_mux_rs3h_data_1_n31 ,
         bypass_mux_rs3h_data_1_n30 , bypass_mux_rs3h_data_1_n29 ,
         bypass_mux_rs3h_data_1_n28 , bypass_mux_rs3h_data_1_n25 ,
         bypass_mux_rs3h_data_1_n24 , bypass_mux_rs3h_data_1_n23 ,
         bypass_mux_rs3h_data_1_n22 , bypass_mux_rs3h_data_1_n19 ,
         bypass_mux_rs3h_data_1_n18 , bypass_mux_rs3h_data_1_n17 ,
         bypass_mux_rs3h_data_1_n16 , bypass_mux_rs3h_data_1_n13 ,
         bypass_mux_rs3h_data_1_n12 , bypass_mux_rs3h_data_1_n11 ,
         bypass_mux_rs3h_data_1_n10 , bypass_mux_rs3h_data_1_n7 ,
         bypass_mux_rs3h_data_1_n6 , bypass_mux_rs3h_data_1_n5 ,
         bypass_mux_rs3h_data_1_n4 , bypass_mux_rs3h_data_1_n1 ,
         bypass_w1_eccgen_n127 , bypass_w1_eccgen_n126 ,
         bypass_w1_eccgen_n125 , bypass_w1_eccgen_n124 ,
         bypass_w1_eccgen_n123 , bypass_w1_eccgen_n122 ,
         bypass_w1_eccgen_n121 , bypass_w1_eccgen_n120 ,
         bypass_w1_eccgen_n119 , bypass_w1_eccgen_n118 ,
         bypass_w1_eccgen_n117 , bypass_w1_eccgen_n116 ,
         bypass_w1_eccgen_n115 , bypass_w1_eccgen_n114 ,
         bypass_w1_eccgen_n113 , bypass_w1_eccgen_n112 ,
         bypass_w1_eccgen_n111 , bypass_w1_eccgen_n110 ,
         bypass_w1_eccgen_n109 , bypass_w1_eccgen_n108 ,
         bypass_w1_eccgen_n107 , bypass_w1_eccgen_n106 ,
         bypass_w1_eccgen_n105 , bypass_w1_eccgen_n104 ,
         bypass_w1_eccgen_n103 , bypass_w1_eccgen_n102 ,
         bypass_w1_eccgen_n101 , bypass_w1_eccgen_n100 ,
         bypass_w1_eccgen_n99 , bypass_w1_eccgen_n98 ,
         bypass_w1_eccgen_n97 , bypass_w1_eccgen_n96 ,
         bypass_w1_eccgen_n95 , bypass_w1_eccgen_n94 ,
         bypass_w1_eccgen_n93 , bypass_w1_eccgen_n92 ,
         bypass_w1_eccgen_n91 , bypass_w1_eccgen_n90 ,
         bypass_w1_eccgen_n89 , bypass_w1_eccgen_n88 ,
         bypass_w1_eccgen_n87 , bypass_w1_eccgen_n86 ,
         bypass_w1_eccgen_n85 , bypass_w1_eccgen_n84 ,
         bypass_w1_eccgen_n83 , bypass_w1_eccgen_n82 ,
         bypass_w1_eccgen_n81 , bypass_w1_eccgen_n80 ,
         bypass_w1_eccgen_n79 , bypass_w1_eccgen_n78 ,
         bypass_w1_eccgen_n77 , bypass_w1_eccgen_n76 ,
         bypass_w1_eccgen_n75 , bypass_w1_eccgen_n74 ,
         bypass_w1_eccgen_n73 , bypass_w1_eccgen_n72 ,
         bypass_w1_eccgen_n71 , bypass_w1_eccgen_n70 ,
         bypass_w1_eccgen_n69 , bypass_w1_eccgen_n68 ,
         bypass_w1_eccgen_n67 , bypass_w1_eccgen_n66 ,
         bypass_w1_eccgen_n65 , bypass_w1_eccgen_n64 ,
         bypass_w1_eccgen_n63 , bypass_w1_eccgen_n62 ,
         bypass_w1_eccgen_n61 , bypass_w1_eccgen_n60 ,
         bypass_w1_eccgen_n59 , bypass_w1_eccgen_n58 ,
         bypass_w1_eccgen_n57 , bypass_w1_eccgen_n56 ,
         bypass_w1_eccgen_n55 , bypass_w1_eccgen_n54 ,
         bypass_w1_eccgen_n53 , bypass_w1_eccgen_n52 ,
         bypass_w1_eccgen_n51 , bypass_w1_eccgen_n50 ,
         bypass_w1_eccgen_n49 , bypass_w1_eccgen_n48 ,
         bypass_w1_eccgen_n47 , bypass_w1_eccgen_n46 ,
         bypass_w1_eccgen_n45 , bypass_w1_eccgen_n44 ,
         bypass_w1_eccgen_n43 , bypass_w1_eccgen_n42 ,
         bypass_w1_eccgen_n41 , bypass_w1_eccgen_n40 ,
         bypass_w1_eccgen_n39 , bypass_w1_eccgen_n38 ,
         bypass_w1_eccgen_n37 , bypass_w1_eccgen_n36 ,
         bypass_w1_eccgen_n35 , bypass_w1_eccgen_n34 ,
         bypass_w1_eccgen_n33 , bypass_w1_eccgen_n32 ,
         bypass_w1_eccgen_n31 , bypass_w1_eccgen_n30 ,
         bypass_w1_eccgen_n29 , bypass_w1_eccgen_n28 ,
         bypass_w1_eccgen_n27 , bypass_w1_eccgen_n26 ,
         bypass_w1_eccgen_n25 , bypass_w1_eccgen_n24 ,
         bypass_w1_eccgen_n23 , bypass_w1_eccgen_n22 ,
         bypass_w1_eccgen_n21 , bypass_w1_eccgen_n20 ,
         bypass_w1_eccgen_n19 , bypass_w1_eccgen_n18 ,
         bypass_w1_eccgen_n17 , bypass_w1_eccgen_n16 ,
         bypass_w1_eccgen_n15 , bypass_w1_eccgen_n14 ,
         bypass_w1_eccgen_n13 , bypass_w1_eccgen_n12 ,
         bypass_w1_eccgen_n11 , bypass_w1_eccgen_n10 , bypass_w1_eccgen_n9 ,
         bypass_w1_eccgen_n8 , bypass_w1_eccgen_n7 , bypass_w1_eccgen_n6 ,
         bypass_w1_eccgen_n5 , bypass_w1_eccgen_n4 , bypass_w1_eccgen_n3 ,
         bypass_w1_eccgen_n2 , bypass_w1_eccgen_n1 ,
         bypass_w1_eccgen_p7_g[0] , bypass_w1_eccgen_p7_g[1] ,
         bypass_w1_eccgen_p7_g[2] , bypass_w1_eccgen_p7_g[3] ,
         bypass_w1_eccgen_p7_g[4] , bypass_w1_eccgen_p7_g[5] ,
         bypass_w1_eccgen_p7_g[6] , bypass_w1_eccgen_p7_g[7] ,
         bypass_w1_eccgen_p7_w[7] , bypass_w1_eccgen_p7_w[6] ,
         bypass_w1_eccgen_p7_w[5] , bypass_w1_eccgen_p7_w[4] ,
         bypass_w1_eccgen_p7_w[3] , bypass_w1_eccgen_p7_w[2] ,
         bypass_w1_eccgen_p7_w[1] , bypass_w1_eccgen_p7_w[0] ,
         bypass_w1_eccgen_p6_g[1] , bypass_w1_eccgen_p6_g[0] ,
         bypass_w1_eccgen_p6_w[1] , bypass_w1_eccgen_p6_w[0] ,
         bypass_w1_eccgen_p5_g[1] , bypass_w1_eccgen_p5_g[0] ,
         bypass_w1_eccgen_p5_w[1] , bypass_w1_eccgen_p5_w[0] ,
         bypass_w1_eccgen_p4_g[3] , bypass_w1_eccgen_p4_g[2] ,
         bypass_w1_eccgen_p4_g[1] , bypass_w1_eccgen_p4_g[0] ,
         bypass_w1_eccgen_p4_w[0] , bypass_w1_eccgen_p4_w[1] ,
         bypass_w1_eccgen_p4_w[2] , bypass_w1_eccgen_p4_w[3] ,
         bypass_w1_eccgen_p3_g[0] , bypass_w1_eccgen_p3_g[1] ,
         bypass_w1_eccgen_p3_g[2] , bypass_w1_eccgen_p3_g[3] ,
         bypass_w1_eccgen_p3_g[4] , bypass_w1_eccgen_p3_g[5] ,
         bypass_w1_eccgen_p3_g[6] , bypass_w1_eccgen_p3_g[7] ,
         bypass_w1_eccgen_p3_w[7] , bypass_w1_eccgen_p3_w[6] ,
         bypass_w1_eccgen_p3_w[5] , bypass_w1_eccgen_p3_w[4] ,
         bypass_w1_eccgen_p3_w[3] , bypass_w1_eccgen_p3_w[2] ,
         bypass_w1_eccgen_p3_w[1] , bypass_w1_eccgen_p3_w[0] ,
         bypass_w1_eccgen_p2_g[7] , bypass_w1_eccgen_p2_g[6] ,
         bypass_w1_eccgen_p2_g[5] , bypass_w1_eccgen_p2_g[4] ,
         bypass_w1_eccgen_p2_g[3] , bypass_w1_eccgen_p2_g[2] ,
         bypass_w1_eccgen_p2_g[1] , bypass_w1_eccgen_p2_g[0] ,
         bypass_w1_eccgen_p2_w[7] , bypass_w1_eccgen_p2_w[6] ,
         bypass_w1_eccgen_p2_w[5] , bypass_w1_eccgen_p2_w[4] ,
         bypass_w1_eccgen_p2_w[3] , bypass_w1_eccgen_p2_w[2] ,
         bypass_w1_eccgen_p2_w[1] , bypass_w1_eccgen_p2_w[0] ,
         bypass_w1_eccgen_p1_g[7] , bypass_w1_eccgen_p1_g[6] ,
         bypass_w1_eccgen_p1_g[5] , bypass_w1_eccgen_p1_g[4] ,
         bypass_w1_eccgen_p1_g[3] , bypass_w1_eccgen_p1_g[2] ,
         bypass_w1_eccgen_p1_g[1] , bypass_w1_eccgen_p1_g[0] ,
         bypass_w1_eccgen_p1_w[7] , bypass_w1_eccgen_p1_w[6] ,
         bypass_w1_eccgen_p1_w[5] , bypass_w1_eccgen_p1_w[4] ,
         bypass_w1_eccgen_p1_w[3] , bypass_w1_eccgen_p1_w[2] ,
         bypass_w1_eccgen_p1_w[1] , bypass_w1_eccgen_p1_w[0] ,
         bypass_w1_eccgen_p0_g[7] , bypass_w1_eccgen_p0_g[6] ,
         bypass_w1_eccgen_p0_g[5] , bypass_w1_eccgen_p0_g[4] ,
         bypass_w1_eccgen_p0_g[3] , bypass_w1_eccgen_p0_g[2] ,
         bypass_w1_eccgen_p0_g[1] , bypass_w1_eccgen_p0_g[0] ,
         bypass_w1_eccgen_p0_w[7] , bypass_w1_eccgen_p0_w[6] ,
         bypass_w1_eccgen_p0_w[5] , bypass_w1_eccgen_p0_w[4] ,
         bypass_w1_eccgen_p0_w[3] , bypass_w1_eccgen_p0_w[2] ,
         bypass_w1_eccgen_p0_w[1] , bypass_w1_eccgen_p0_w[0] ,
         bypass_w1_eccgen_msk_w4 , bypass_w1_eccgen_msk_w5 ,
         ecc_rs1_ecc_d2e_n17 , ecc_rs1_ecc_d2e_n15 , ecc_rs1_ecc_d2e_n13 ,
         ecc_rs1_ecc_d2e_n11 , ecc_rs1_ecc_d2e_n9 , ecc_rs1_ecc_d2e_n7 ,
         ecc_rs1_ecc_d2e_n5 , ecc_rs1_ecc_d2e_n3 , ecc_rs1_ecc_d2e_n1 ,
         ecc_chk_rs1_n138 , ecc_chk_rs1_n137 , ecc_chk_rs1_n136 ,
         ecc_chk_rs1_n135 , ecc_chk_rs1_n134 , ecc_chk_rs1_n133 ,
         ecc_chk_rs1_n132 , ecc_chk_rs1_n131 , ecc_chk_rs1_n130 ,
         ecc_chk_rs1_n129 , ecc_chk_rs1_n128 , ecc_chk_rs1_n127 ,
         ecc_chk_rs1_n126 , ecc_chk_rs1_n125 , ecc_chk_rs1_n124 ,
         ecc_chk_rs1_n123 , ecc_chk_rs1_n122 , ecc_chk_rs1_n121 ,
         ecc_chk_rs1_n120 , ecc_chk_rs1_n119 , ecc_chk_rs1_n118 ,
         ecc_chk_rs1_n117 , ecc_chk_rs1_n116 , ecc_chk_rs1_n115 ,
         ecc_chk_rs1_n114 , ecc_chk_rs1_n113 , ecc_chk_rs1_n112 ,
         ecc_chk_rs1_n111 , ecc_chk_rs1_n110 , ecc_chk_rs1_n109 ,
         ecc_chk_rs1_n108 , ecc_chk_rs1_n107 , ecc_chk_rs1_n106 ,
         ecc_chk_rs1_n105 , ecc_chk_rs1_n104 , ecc_chk_rs1_n103 ,
         ecc_chk_rs1_n102 , ecc_chk_rs1_n101 , ecc_chk_rs1_n100 ,
         ecc_chk_rs1_n99 , ecc_chk_rs1_n98 , ecc_chk_rs1_n97 ,
         ecc_chk_rs1_n96 , ecc_chk_rs1_n95 , ecc_chk_rs1_n94 ,
         ecc_chk_rs1_n93 , ecc_chk_rs1_n92 , ecc_chk_rs1_n91 ,
         ecc_chk_rs1_n90 , ecc_chk_rs1_n89 , ecc_chk_rs1_n88 ,
         ecc_chk_rs1_n87 , ecc_chk_rs1_n86 , ecc_chk_rs1_n85 ,
         ecc_chk_rs1_n84 , ecc_chk_rs1_n83 , ecc_chk_rs1_n82 ,
         ecc_chk_rs1_n81 , ecc_chk_rs1_n80 , ecc_chk_rs1_n79 ,
         ecc_chk_rs1_n78 , ecc_chk_rs1_n77 , ecc_chk_rs1_n76 ,
         ecc_chk_rs1_n75 , ecc_chk_rs1_n74 , ecc_chk_rs1_n73 ,
         ecc_chk_rs1_n72 , ecc_chk_rs1_n71 , ecc_chk_rs1_n70 ,
         ecc_chk_rs1_n69 , ecc_chk_rs1_n68 , ecc_chk_rs1_n67 ,
         ecc_chk_rs1_n66 , ecc_chk_rs1_n65 , ecc_chk_rs1_n64 ,
         ecc_chk_rs1_n63 , ecc_chk_rs1_n62 , ecc_chk_rs1_n61 ,
         ecc_chk_rs1_n60 , ecc_chk_rs1_n59 , ecc_chk_rs1_n58 ,
         ecc_chk_rs1_n57 , ecc_chk_rs1_n56 , ecc_chk_rs1_n55 ,
         ecc_chk_rs1_n54 , ecc_chk_rs1_n53 , ecc_chk_rs1_n52 ,
         ecc_chk_rs1_n51 , ecc_chk_rs1_n50 , ecc_chk_rs1_n49 ,
         ecc_chk_rs1_n48 , ecc_chk_rs1_n47 , ecc_chk_rs1_n46 ,
         ecc_chk_rs1_n45 , ecc_chk_rs1_n44 , ecc_chk_rs1_n43 ,
         ecc_chk_rs1_n42 , ecc_chk_rs1_n41 , ecc_chk_rs1_n40 ,
         ecc_chk_rs1_n39 , ecc_chk_rs1_n38 , ecc_chk_rs1_n37 ,
         ecc_chk_rs1_n36 , ecc_chk_rs1_n35 , ecc_chk_rs1_n34 ,
         ecc_chk_rs1_n33 , ecc_chk_rs1_n32 , ecc_chk_rs1_n31 ,
         ecc_chk_rs1_n30 , ecc_chk_rs1_n29 , ecc_chk_rs1_n28 ,
         ecc_chk_rs1_n27 , ecc_chk_rs1_n26 , ecc_chk_rs1_n25 ,
         ecc_chk_rs1_n24 , ecc_chk_rs1_n23 , ecc_chk_rs1_n22 ,
         ecc_chk_rs1_n21 , ecc_chk_rs1_n20 , ecc_chk_rs1_n19 ,
         ecc_chk_rs1_n18 , ecc_chk_rs1_n17 , ecc_chk_rs1_n16 ,
         ecc_chk_rs1_n15 , ecc_chk_rs1_n14 , ecc_chk_rs1_n13 ,
         ecc_chk_rs1_n12 , ecc_chk_rs1_n11 , ecc_chk_rs1_n10 ,
         ecc_chk_rs1_n9 , ecc_chk_rs1_n8 , ecc_chk_rs1_n7 ,
         ecc_chk_rs1_n6 , ecc_chk_rs1_n5 , ecc_chk_rs1_n3 ,
         ecc_chk_rs1_n2 , ecc_chk_rs1_parity , ecc_rs1_err_e2m_n15 ,
         ecc_rs1_err_e2m_n13 , ecc_rs1_err_e2m_n11 , ecc_rs1_err_e2m_n9 ,
         ecc_rs1_err_e2m_n7 , ecc_rs1_err_e2m_n5 , ecc_rs1_err_e2m_n3 ,
         ecc_rs1_err_e2m_n1 , ecc_syn_mux_n28 , ecc_syn_mux_n27 ,
         ecc_syn_mux_n26 , ecc_syn_mux_n25 , ecc_syn_mux_n24 ,
         ecc_syn_mux_n23 , ecc_syn_mux_n22 , ecc_syn_mux_n21 ,
         ecc_syn_mux_n20 , ecc_syn_mux_n19 , ecc_syn_mux_n18 ,
         ecc_syn_mux_n17 , ecc_syn_mux_n16 , ecc_syn_mux_n15 ,
         ecc_syn_mux_n14 , ecc_syn_mux_n13 , ecc_syn_mux_n12 ,
         ecc_syn_mux_n11 , ecc_syn_mux_n10 , ecc_syn_mux_n9 ,
         ecc_syn_mux_n8 , ecc_syn_mux_n7 , ecc_syn_mux_n6 ,
         ecc_syn_mux_n5 , ecc_syn_mux_n4 , ecc_syn_mux_n3 ,
         ecc_syn_mux_n2 , ecc_syn_mux_n1 , ecc_decode_n49 ,
         ecc_decode_n48 , ecc_decode_n47 , ecc_decode_n46 ,
         ecc_decode_n45 , ecc_decode_n44 , ecc_decode_n43 ,
         ecc_decode_n42 , ecc_decode_n41 , ecc_decode_n40 ,
         ecc_decode_n39 , ecc_decode_n38 , ecc_decode_n37 ,
         ecc_decode_n36 , ecc_decode_n35 , ecc_decode_n34 ,
         ecc_decode_n33 , ecc_decode_n32 , ecc_decode_n31 ,
         ecc_decode_n30 , ecc_decode_n29 , ecc_decode_n28 ,
         ecc_decode_n27 , ecc_decode_n26 , ecc_decode_n25 ,
         ecc_decode_n24 , ecc_decode_n23 , ecc_decode_n22 ,
         ecc_decode_n21 , ecc_decode_n20 , ecc_decode_n19 ,
         ecc_decode_n18 , ecc_decode_n17 , ecc_decode_n16 ,
         ecc_decode_n15 , ecl_dff_rs1_s2d_n11 , ecl_dff_rs1_s2d_n9 ,
         ecl_dff_rs1_s2d_n7 , ecl_dff_rs1_s2d_n5 , ecl_dff_rs1_s2d_n3 ,
         ecl_dff_rs1_s2d_n1 , ecl_dff_ld_tid_m2g_n5 ,
         ecl_dff_ld_tid_m2g_n3 , ecl_dff_ld_tid_m2g_n1 ,
         ecl_dff_aluop_d2e_n7 , ecl_dff_aluop_d2e_n5 ,
         ecl_dff_aluop_d2e_n3 , ecl_dff_aluop_d2e_n1 ,
         ecl_dff_enshift_d2e_n3 , ecl_yreg0_mux_n6 , ecl_yreg0_mux_n5 ,
         ecl_yreg0_mux_n4 , ecl_yreg0_mux_n3 , ecl_yreg0_mux_n2 ,
         ecl_yreg0_mux_n1 , ecl_perr_dff_n9 , ecl_perr_dff_n7 ,
         ecl_perr_dff_n5 , ecl_perr_dff_n3 , ecl_perr_dff_n2 ,
         ecl_ttype_mux_n36 , ecl_ttype_mux_n35 , ecl_ttype_mux_n33 ,
         ecl_ttype_mux_n31 , ecl_ttype_mux_n29 , ecl_ttype_mux_n28 ,
         ecl_ttype_mux_n27 , ecl_ttype_mux_n25 , ecl_ttype_mux_n24 ,
         ecl_ttype_mux_n23 , ecl_ttype_mux_n21 , ecl_ttype_mux_n20 ,
         ecl_ttype_mux_n19 , ecl_ttype_mux_n17 , ecl_ttype_mux_n16 ,
         ecl_ttype_mux_n15 , ecl_ttype_mux_n13 , ecl_ttype_mux_n12 ,
         ecl_ttype_mux_n11 , ecl_ttype_mux_n9 , ecl_ttype_mux_n7 ,
         ecl_ttype_mux_n5 , ecl_ttype_e2m_n19 , ecl_ttype_e2m_n17 ,
         ecl_ttype_e2m_n15 , ecl_ttype_e2m_n13 , ecl_ttype_e2m_n11 ,
         ecl_ttype_e2m_n9 , ecl_ttype_e2m_n7 , ecl_ttype_e2m_n5 ,
         ecl_ttype_e2m_n3 , ecl_ttype_e2m_n1 , ecl_ccr_n54 , ecl_ccr_n53 ,
         ecl_ccr_n52 , ecl_ccr_n51 , ecl_ccr_n50 , ecl_ccr_n49 ,
         ecl_ccr_n48 , ecl_ccr_n47 , ecl_ccr_n46 , ecl_ccr_n45 ,
         ecl_ccr_n44 , ecl_ccr_n43 , ecl_ccr_n42 , ecl_ccr_n41 ,
         ecl_ccr_n40 , ecl_ccr_n39 , ecl_ccr_n38 , ecl_ccr_n37 ,
         ecl_ccr_n36 , ecl_ccr_n35 , ecl_ccr_n34 , ecl_ccr_n33 ,
         ecl_ccr_n32 , ecl_ccr_n31 , ecl_ccr_n30 , ecl_ccr_n29 ,
         ecl_ccr_n28 , ecl_ccr_n27 , ecl_ccr_n26 , ecl_ccr_n25 ,
         ecl_ccr_n24 , ecl_ccr_n23 , ecl_ccr_n22 , ecl_ccr_n21 ,
         ecl_ccr_n20 , ecl_ccr_n19 , ecl_ccr_n18 , ecl_ccr_n17 ,
         ecl_ccr_n16 , ecl_ccr_n15 , ecl_ccr_n14 , ecl_ccr_n13 ,
         ecl_ccr_n12 , ecl_ccr_use_cc_w , ecl_ccr_partial_cc_d[7] ,
         ecl_ccr_partial_cc_d[6] , ecl_ccr_partial_cc_d[5] ,
         ecl_ccr_partial_cc_d[4] , ecl_ccr_partial_cc_d[3] ,
         ecl_ccr_partial_cc_d[2] , ecl_ccr_partial_cc_d[1] ,
         ecl_ccr_partial_cc_d[0] , ecl_ccr_ccr_d[7] , ecl_ccr_ccr_d[6] ,
         ecl_ccr_ccr_d[5] , ecl_ccr_ccr_d[4] , ecl_ccr_ccr_d[3] ,
         ecl_ccr_ccr_d[2] , ecl_ccr_ccr_d[1] , ecl_ccr_ccr_d[0] ,
         ecl_ccr_ccrin_thr3[7] , ecl_ccr_ccrin_thr3[6] ,
         ecl_ccr_ccrin_thr3[5] , ecl_ccr_ccrin_thr3[4] ,
         ecl_ccr_ccrin_thr3[3] , ecl_ccr_ccrin_thr3[2] ,
         ecl_ccr_ccrin_thr3[1] , ecl_ccr_ccrin_thr3[0] ,
         ecl_ccr_ccrin_thr2[7] , ecl_ccr_ccrin_thr2[6] ,
         ecl_ccr_ccrin_thr2[5] , ecl_ccr_ccrin_thr2[4] ,
         ecl_ccr_ccrin_thr2[3] , ecl_ccr_ccrin_thr2[2] ,
         ecl_ccr_ccrin_thr2[1] , ecl_ccr_ccrin_thr2[0] ,
         ecl_ccr_ccrin_thr1[7] , ecl_ccr_ccrin_thr1[6] ,
         ecl_ccr_ccrin_thr1[5] , ecl_ccr_ccrin_thr1[4] ,
         ecl_ccr_ccrin_thr1[3] , ecl_ccr_ccrin_thr1[2] ,
         ecl_ccr_ccrin_thr1[1] , ecl_ccr_ccrin_thr1[0] ,
         ecl_ccr_ccrin_thr0[7] , ecl_ccr_ccrin_thr0[6] ,
         ecl_ccr_ccrin_thr0[5] , ecl_ccr_ccrin_thr0[4] ,
         ecl_ccr_ccrin_thr0[3] , ecl_ccr_ccrin_thr0[2] ,
         ecl_ccr_ccrin_thr0[1] , ecl_ccr_ccrin_thr0[0] ,
         ecl_ccr_wen_thr3_w , ecl_ccr_wen_thr2_w , ecl_ccr_wen_thr1_w ,
         ecl_ccr_wen_thr0_w , ecl_ccr_thr_w2[0] , ecl_ccr_thr_w2[1] ,
         ecl_ccr_setcc_w2 , ecl_ccr_exu_ifu_cc_w[0] ,
         ecl_ccr_exu_ifu_cc_w[1] , ecl_ccr_exu_ifu_cc_w[2] ,
         ecl_ccr_exu_ifu_cc_w[3] , ecl_ccr_exu_ifu_cc_w[4] ,
         ecl_ccr_exu_ifu_cc_w[5] , ecl_ccr_exu_ifu_cc_w[6] ,
         ecl_ccr_exu_ifu_cc_w[7] , ecl_ccr_setcc_w , ecl_ccr_alu_cc_w[0] ,
         ecl_ccr_alu_cc_w[1] , ecl_ccr_alu_cc_w[2] , ecl_ccr_alu_cc_w[3] ,
         ecl_ccr_alu_cc_w[4] , ecl_ccr_alu_cc_w[5] , ecl_ccr_alu_cc_w[6] ,
         ecl_ccr_alu_cc_w[7] , ecl_ccr_ccr_m[7] , ecl_ccr_ccr_m[6] ,
         ecl_ccr_ccr_m[5] , ecl_ccr_ccr_m[4] , ecl_ccr_ccr_m[3] ,
         ecl_ccr_ccr_m[2] , ecl_ccr_ccr_m[1] , ecl_ccr_ccr_m[0] ,
         ecl_ccr_valid_setcc_m , ecl_ccr_setcc_m , ecl_ccr_alu_cc_m[0] ,
         ecl_ccr_alu_cc_m[1] , ecl_ccr_alu_cc_m[2] , ecl_ccr_alu_cc_m[3] ,
         ecl_ccr_alu_cc_m[4] , ecl_ccr_alu_cc_m[5] , ecl_ccr_alu_cc_m[6] ,
         ecl_ccr_alu_cc_m[7] , ecl_ccr_valid_setcc_e , ecl_ccr_setcc_e ,
         ecl_writeback_n200 , ecl_writeback_n199 , ecl_writeback_n198 ,
         ecl_writeback_n197 , ecl_writeback_n196 , ecl_writeback_n195 ,
         ecl_writeback_n194 , ecl_writeback_n193 , ecl_writeback_n192 ,
         ecl_writeback_n191 , ecl_writeback_n190 , ecl_writeback_n189 ,
         ecl_writeback_n188 , ecl_writeback_n187 , ecl_writeback_n186 ,
         ecl_writeback_n185 , ecl_writeback_n184 , ecl_writeback_n183 ,
         ecl_writeback_n182 , ecl_writeback_n181 , ecl_writeback_n180 ,
         ecl_writeback_n179 , ecl_writeback_n178 , ecl_writeback_n177 ,
         ecl_writeback_n176 , ecl_writeback_n175 , ecl_writeback_n174 ,
         ecl_writeback_n173 , ecl_writeback_n172 , ecl_writeback_n171 ,
         ecl_writeback_n170 , ecl_writeback_n169 , ecl_writeback_n168 ,
         ecl_writeback_n167 , ecl_writeback_n166 , ecl_writeback_n165 ,
         ecl_writeback_n164 , ecl_writeback_n162 , ecl_writeback_n161 ,
         ecl_writeback_n160 , ecl_writeback_n159 , ecl_writeback_n158 ,
         ecl_writeback_n157 , ecl_writeback_n156 , ecl_writeback_n155 ,
         ecl_writeback_n154 , ecl_writeback_n153 , ecl_writeback_n152 ,
         ecl_writeback_n151 , ecl_writeback_n150 , ecl_writeback_n149 ,
         ecl_writeback_n148 , ecl_writeback_n147 , ecl_writeback_n146 ,
         ecl_writeback_n145 , ecl_writeback_n144 , ecl_writeback_n143 ,
         ecl_writeback_n142 , ecl_writeback_n141 , ecl_writeback_n140 ,
         ecl_writeback_n139 , ecl_writeback_n138 , ecl_writeback_n137 ,
         ecl_writeback_n136 , ecl_writeback_n135 , ecl_writeback_n134 ,
         ecl_writeback_n133 , ecl_writeback_n132 , ecl_writeback_n131 ,
         ecl_writeback_n130 , ecl_writeback_n129 , ecl_writeback_n128 ,
         ecl_writeback_n127 , ecl_writeback_n126 , ecl_writeback_n125 ,
         ecl_writeback_n124 , ecl_writeback_n123 , ecl_writeback_n122 ,
         ecl_writeback_n121 , ecl_writeback_n120 , ecl_writeback_n119 ,
         ecl_writeback_n118 , ecl_writeback_n117 , ecl_writeback_n116 ,
         ecl_writeback_n115 , ecl_writeback_n114 , ecl_writeback_n113 ,
         ecl_writeback_n112 , ecl_writeback_n111 , ecl_writeback_n110 ,
         ecl_writeback_n109 , ecl_writeback_n108 , ecl_writeback_n107 ,
         ecl_writeback_n106 , ecl_writeback_n105 , ecl_writeback_n104 ,
         ecl_writeback_n103 , ecl_writeback_n102 , ecl_writeback_n101 ,
         ecl_writeback_n100 , ecl_writeback_n99 , ecl_writeback_n98 ,
         ecl_writeback_n97 , ecl_writeback_n96 , ecl_writeback_n94 ,
         ecl_writeback_n93 , ecl_writeback_n92 , ecl_writeback_n91 ,
         ecl_writeback_n90 , ecl_writeback_n89 , ecl_writeback_n88 ,
         ecl_writeback_n86 , ecl_writeback_n85 , ecl_writeback_n84 ,
         ecl_writeback_n83 , ecl_writeback_n82 , ecl_writeback_n81 ,
         ecl_writeback_n80 , ecl_writeback_n79 , ecl_writeback_n78 ,
         ecl_writeback_n77 , ecl_writeback_n76 , ecl_writeback_n75 ,
         ecl_writeback_n74 , ecl_writeback_n73 , ecl_writeback_n72 ,
         ecl_writeback_n71 , ecl_writeback_n70 , ecl_writeback_n69 ,
         ecl_writeback_n68 , ecl_writeback_n67 , ecl_writeback_n66 ,
         ecl_writeback_n65 , ecl_writeback_n64 , ecl_writeback_n63 ,
         ecl_writeback_n62 , ecl_writeback_n61 , ecl_writeback_n60 ,
         ecl_writeback_n59 , ecl_writeback_n58 , ecl_writeback_n57 ,
         ecl_writeback_n56 , ecl_writeback_n55 , ecl_writeback_n54 ,
         ecl_writeback_n53 , ecl_writeback_n52 , ecl_writeback_n51 ,
         ecl_writeback_n50 , ecl_writeback_n49 , ecl_writeback_n48 ,
         ecl_writeback_n47 , ecl_writeback_n46 , ecl_writeback_n45 ,
         ecl_writeback_n44 , ecl_writeback_n43 , ecl_writeback_n19 ,
         ecl_writeback_short_longop_done_m ,
         ecl_writeback_short_longop_done_e ,
         ecl_writeback_restore_ready_next , ecl_writeback_restore_ready ,
         ecl_writeback_restore_w , ecl_writeback_vld_restore_e ,
         ecl_writeback_return_e , ecl_writeback_rdpr_mux2_out[5] ,
         ecl_writeback_rdpr_mux2_out[4] , ecl_writeback_rdpr_mux2_out[3] ,
         ecl_writeback_rdpr_mux2_out[2] , ecl_writeback_rdpr_mux2_out[1] ,
         ecl_writeback_rdpr_mux2_out[0] , ecl_writeback_sel_wstate_d ,
         ecl_writeback_sel_cwp_d , ecl_writeback_rdpr_mux1_out[2] ,
         ecl_writeback_rdpr_mux1_out[1] , ecl_writeback_rdpr_mux1_out[0] ,
         ecl_writeback_sel_cansave_d , ecl_writeback_sel_cleanwin_d ,
         ecl_writeback_sraddr_m[6] , ecl_writeback_sraddr_m[5] ,
         ecl_writeback_sraddr_m[4] , ecl_writeback_sraddr_m[3] ,
         ecl_writeback_sraddr_m[2] , ecl_writeback_sraddr_m[1] ,
         ecl_writeback_sraddr_m[0] , ecl_writeback_yreg_wen_w1 ,
         ecl_writeback_yreg_wen_w , ecl_writeback_wrsr_w ,
         ecl_writeback_sraddr_w[0] , ecl_writeback_sraddr_w[1] ,
         ecl_writeback_sraddr_w[2] , ecl_writeback_sraddr_w[3] ,
         ecl_writeback_sraddr_w[4] , ecl_writeback_sraddr_w[5] ,
         ecl_writeback_sraddr_w[6] , ecl_writeback_sraddr_e[0] ,
         ecl_writeback_sraddr_e[1] , ecl_writeback_sraddr_e[2] ,
         ecl_writeback_sraddr_e[3] , ecl_writeback_sraddr_e[4] ,
         ecl_writeback_sraddr_e[5] , ecl_writeback_sraddr_e[6] ,
         ecl_writeback_wb_w , ecl_writeback_valid_m ,
         ecl_writeback_valid_e , ecl_writeback_inst_vld_noflush_wen_w ,
         ecl_writeback_inst_vld_noflush_wen_m ,
         ecl_writeback_wen_no_inst_vld_w , ecl_writeback_wen_no_inst_vld_m ,
         ecl_writeback_setcc_g , ecl_writeback_restore_tid[0] ,
         ecl_writeback_restore_tid[1] , ecl_writeback_restore_rd[0] ,
         ecl_writeback_restore_rd[1] , ecl_writeback_restore_rd[2] ,
         ecl_writeback_restore_rd[3] , ecl_writeback_restore_rd[4] ,
         ecl_writeback_ecl_irf_wen_g , ecl_writeback_ecl_sel_div_g ,
         ecl_writeback_ecl_sel_mul_g , ecl_writeback_wrsr_m ,
         ecl_writeback_dfill_tid_g2[0] , ecl_writeback_dfill_tid_g2[1] ,
         ecl_writeback_ld_g , ecl_eccctl_n35 , ecl_eccctl_n34 ,
         ecl_eccctl_n33 , ecl_eccctl_n32 , ecl_eccctl_n31 ,
         ecl_eccctl_n30 , ecl_eccctl_n29 , ecl_eccctl_n28 ,
         ecl_eccctl_n27 , ecl_eccctl_n26 , ecl_eccctl_n25 ,
         ecl_eccctl_n24 , ecl_eccctl_n23 , ecl_eccctl_n22 ,
         ecl_eccctl_n21 , ecl_eccctl_n20 , ecl_eccctl_n19 ,
         ecl_eccctl_n18 , ecl_eccctl_n17 , ecl_eccctl_n16 ,
         ecl_eccctl_n15 , ecl_eccctl_n14 , ecl_eccctl_inj_irferr_m ,
         ecl_eccctl_cwp_e[2] , ecl_eccctl_cwp_e[1] , ecl_eccctl_cwp_e[0] ,
         ecl_eccctl_rs2_ce_m , ecl_eccctl_rs3_ue_m , ecl_eccctl_rs2_ue_m ,
         ecl_eccctl_rs1_ce_m , ecl_eccctl_rs1_ue_m , ecl_eccctl_sel_rs3_m ,
         ecl_eccctl_sel_rs2_m , ecl_eccctl_sel_rs1_m ,
         ecl_eccctl_sel_rs2_e , ecl_eccctl_cwp_m[2] , ecl_eccctl_cwp_m[1] ,
         ecl_eccctl_cwp_m[0] , ecl_eccctl_gl_m[1] , ecl_eccctl_gl_m[0] ,
         ecl_eccctl_nceen_m , ecl_eccctl_flag_ecc_ce_e ,
         ecl_eccctl_flag_ecc_ue_e , ecl_eccctl_rs3_sel_rf_e ,
         ecl_eccctl_rs2_sel_rf_e , ecl_eccctl_rs1_sel_rf_e ,
         ecl_byplog_rs1_n50 , ecl_byplog_rs1_n49 , ecl_byplog_rs1_n48 ,
         ecl_byplog_rs1_n47 , ecl_byplog_rs1_n46 , ecl_byplog_rs1_n45 ,
         ecl_byplog_rs1_n44 , ecl_byplog_rs1_n43 , ecl_byplog_rs1_n42 ,
         ecl_byplog_rs1_n41 , ecl_byplog_rs1_n40 , ecl_byplog_rs1_n39 ,
         ecl_byplog_rs1_n38 , ecl_byplog_rs1_n37 , ecl_byplog_rs1_n36 ,
         ecl_byplog_rs1_n35 , ecl_byplog_rs1_n34 , ecl_byplog_rs1_n33 ,
         ecl_byplog_rs1_n32 , ecl_byplog_rs1_n31 , ecl_byplog_rs1_n30 ,
         ecl_byplog_rs1_n29 , ecl_byplog_rs1_n28 , ecl_byplog_rs1_n27 ,
         ecl_byplog_rs1_n26 , ecl_byplog_rs1_n25 , ecl_byplog_rs1_n24 ,
         ecl_byplog_rs1_n23 , ecl_byplog_rs1_n22 , ecl_byplog_rs1_n21 ,
         ecl_byplog_rs1_n20 , ecl_byplog_rs1_n19 , ecl_byplog_rs1_n18 ,
         ecl_byplog_rs1_n17 , ecl_byplog_rs1_n16 , ecl_byplog_rs1_n15 ,
         ecl_byplog_rs1_n14 , ecl_byplog_rs1_N3 , ecl_byplog_rs1_N2 ,
         ecl_byplog_rs1_N1 , ecl_byplog_rs1_N0 , ecl_byplog_rs1_match_w2 ,
         ecl_byplog_rs1_match_w , ecl_byplog_rs2_n51 , ecl_byplog_rs2_n50 ,
         ecl_byplog_rs2_n49 , ecl_byplog_rs2_n48 , ecl_byplog_rs2_n47 ,
         ecl_byplog_rs2_n46 , ecl_byplog_rs2_n44 , ecl_byplog_rs2_n42 ,
         ecl_byplog_rs2_n41 , ecl_byplog_rs2_n40 , ecl_byplog_rs2_n39 ,
         ecl_byplog_rs2_n38 , ecl_byplog_rs2_n37 , ecl_byplog_rs2_n36 ,
         ecl_byplog_rs2_n35 , ecl_byplog_rs2_n34 , ecl_byplog_rs2_n33 ,
         ecl_byplog_rs2_n32 , ecl_byplog_rs2_n31 , ecl_byplog_rs2_n30 ,
         ecl_byplog_rs2_n29 , ecl_byplog_rs2_n27 , ecl_byplog_rs2_n26 ,
         ecl_byplog_rs2_n25 , ecl_byplog_rs2_n24 , ecl_byplog_rs2_n23 ,
         ecl_byplog_rs2_n22 , ecl_byplog_rs2_n21 , ecl_byplog_rs2_n20 ,
         ecl_byplog_rs2_n19 , ecl_byplog_rs2_n18 , ecl_byplog_rs2_n17 ,
         ecl_byplog_rs2_n16 , ecl_byplog_rs2_n15 , ecl_byplog_rs2_n14 ,
         ecl_byplog_rs2_n13 , ecl_byplog_rs2_n12 , ecl_byplog_rs2_N3 ,
         ecl_byplog_rs2_N2 , ecl_byplog_rs2_N1 , ecl_byplog_rs2_N0 ,
         ecl_byplog_rs2_match_w2 , ecl_byplog_rs2_match_w ,
         ecl_divcntl_n89 , ecl_divcntl_n88 , ecl_divcntl_n87 ,
         ecl_divcntl_n86 , ecl_divcntl_n85 , ecl_divcntl_n84 ,
         ecl_divcntl_n83 , ecl_divcntl_n82 , ecl_divcntl_n81 ,
         ecl_divcntl_n80 , ecl_divcntl_n79 , ecl_divcntl_n78 ,
         ecl_divcntl_n77 , ecl_divcntl_n76 , ecl_divcntl_n75 ,
         ecl_divcntl_n74 , ecl_divcntl_n73 , ecl_divcntl_n72 ,
         ecl_divcntl_n71 , ecl_divcntl_n70 , ecl_divcntl_n69 ,
         ecl_divcntl_n68 , ecl_divcntl_n67 , ecl_divcntl_n66 ,
         ecl_divcntl_n65 , ecl_divcntl_n64 , ecl_divcntl_n63 ,
         ecl_divcntl_n62 , ecl_divcntl_n61 , ecl_divcntl_n60 ,
         ecl_divcntl_n59 , ecl_divcntl_n58 , ecl_divcntl_n57 ,
         ecl_divcntl_n56 , ecl_divcntl_n55 , ecl_divcntl_n54 ,
         ecl_divcntl_n53 , ecl_divcntl_n52 , ecl_divcntl_n51 ,
         ecl_divcntl_n50 , ecl_divcntl_n49 , ecl_divcntl_n48 ,
         ecl_divcntl_n47 , ecl_divcntl_n46 , ecl_divcntl_n45 ,
         ecl_divcntl_n44 , ecl_divcntl_n43 , ecl_divcntl_n42 ,
         ecl_divcntl_n41 , ecl_divcntl_n40 , ecl_divcntl_n39 ,
         ecl_divcntl_n38 , ecl_divcntl_n37 , ecl_divcntl_n36 ,
         ecl_divcntl_n35 , ecl_divcntl_n34 , ecl_divcntl_n33 ,
         ecl_divcntl_n32 , ecl_divcntl_n31 , ecl_divcntl_n30 ,
         ecl_divcntl_n29 , ecl_divcntl_n28 , ecl_divcntl_n27 ,
         ecl_divcntl_n26 , ecl_divcntl_n25 , ecl_divcntl_n24 ,
         ecl_divcntl_n23 , ecl_divcntl_N56 , ecl_divcntl_muls_v ,
         ecl_divcntl_next_muls_v , ecl_divcntl_div_adder_out_31_w ,
         ecl_divcntl_rs2_data_31_w , ecl_divcntl_muls_rs1_data_31_w ,
         ecl_divcntl_muls_c , ecl_divcntl_next_muls_c ,
         ecl_divcntl_low32_nonzero_d1 , ecl_divcntl_sel_div_d1 ,
         ecl_divcntl_gencc_in_31_d1 , ecl_divcntl_upper32_equal_d1 ,
         ecl_divcntl_gencc_in_msb_l_d1 , ecl_divcntl_inputs_neg_q ,
         ecl_divcntl_inputs_neg_d , ecl_divcntl_last_cin_next ,
         ecl_divcntl_zero_rem_q , ecl_divcntl_last_cin ,
         ecl_divcntl_sub_next , ecl_divcntl_sub_next_nocout[1] ,
         ecl_divcntl_sub_next_nocout[0] , ecl_divcntl_firstlast_sub ,
         ecl_divcntl_q_next , ecl_divcntl_q_next_nocout[1] ,
         ecl_divcntl_q_next_nocout[0] , ecl_divcntl_subtract ,
         ecl_divcntl_cntr[5] , ecl_divcntl_cntr[4] , ecl_divcntl_cntr[3] ,
         ecl_divcntl_cntr[2] , ecl_divcntl_cntr[1] , ecl_divcntl_cntr[0] ,
         ecl_divcntl_next_state[5] , ecl_divcntl_next_state[4] ,
         ecl_divcntl_next_state[3] , ecl_divcntl_next_state[2] ,
         ecl_divcntl_next_state[1] , ecl_divcntl_next_state[0] ,
         ecl_divcntl_div_state_0 , ecl_divcntl_div_state_1 ,
         ecl_divcntl_div_state[3] , ecl_divcntl_div_state[4] ,
         ecl_divcntl_div_state[5] , ecl_mdqctl_n63 , ecl_mdqctl_n62 ,
         ecl_mdqctl_n61 , ecl_mdqctl_n60 , ecl_mdqctl_n59 ,
         ecl_mdqctl_n56 , ecl_mdqctl_n55 , ecl_mdqctl_n54 ,
         ecl_mdqctl_n52 , ecl_mdqctl_n51 , ecl_mdqctl_n50 ,
         ecl_mdqctl_n49 , ecl_mdqctl_n48 , ecl_mdqctl_n47 ,
         ecl_mdqctl_n46 , ecl_mdqctl_n45 , ecl_mdqctl_n44 ,
         ecl_mdqctl_n43 , ecl_mdqctl_n42 , ecl_mdqctl_n41 ,
         ecl_mdqctl_n40 , ecl_mdqctl_n39 , ecl_mdqctl_n38 ,
         ecl_mdqctl_n37 , ecl_mdqctl_n36 , ecl_mdqctl_n35 ,
         ecl_mdqctl_n34 , ecl_mdqctl_n33 , ecl_mdqctl_n32 ,
         ecl_mdqctl_n31 , ecl_mdqctl_n30 , ecl_mdqctl_n29 ,
         ecl_mdqctl_n28 , ecl_mdqctl_n27 , ecl_mdqctl_n26 ,
         ecl_mdqctl_n25 , ecl_mdqctl_n24 , ecl_mdqctl_n23 ,
         ecl_mdqctl_n22 , ecl_mdqctl_n21 , ecl_mdqctl_n20 ,
         ecl_mdqctl_n19 , ecl_mdqctl_n18 , ecl_mdqctl_n17 ,
         ecl_mdqctl_n16 , ecl_mdqctl_n15 , ecl_mdqctl_n14 ,
         ecl_mdqctl_n13 , ecl_mdqctl_n12 , ecl_mdqctl_next_mul_done ,
         ecl_mdqctl_mul_done_c3 , ecl_mdqctl_mul_done_c2 ,
         ecl_mdqctl_mul_done_valid_c1 , ecl_mdqctl_mul_done_c1 ,
         ecl_mdqctl_mul_done_valid_c0 , ecl_mdqctl_mul_done_c0 ,
         ecl_mdqctl_mul_done_ack , ecl_mdqctl_mul_ready_next ,
         ecl_mdqctl_mul_data_next[9] , ecl_mdqctl_mul_data_next[8] ,
         ecl_mdqctl_mul_data_next[7] , ecl_mdqctl_mul_data_next[6] ,
         ecl_mdqctl_mul_data_next[5] , ecl_mdqctl_mul_data_next[4] ,
         ecl_mdqctl_mul_data_next[3] , ecl_mdqctl_mul_data_next[2] ,
         ecl_mdqctl_mul_data_next[1] , ecl_mdqctl_mul_data_next[0] ,
         ecl_mdqctl_mul_data[8] , ecl_mdqctl_mul_data[9] ,
         ecl_mdqctl_ismul_w , ecl_mdqctl_ismul_m_valid ,
         ecl_mdqctl_ismul_m , ecl_mdqctl_ismul_e ,
         ecl_mdqctl_isdiv_m_valid , ecl_mdqctl_isdiv_e_valid ,
         ecl_mdqctl_isdiv_m , ecl_mdqctl_div_zero_unqual_m ,
         ecl_mdqctl_isdiv_w , ecl_mdqctl_div_zero_e ,
         ecl_mdqctl_div_data_7 , ecl_mdqctl_div_data[11] ,
         ecl_mdqctl_curr_div_vld , ecl_mdqctl_div_data_next[11] ,
         ecl_mdqctl_div_data_next[10] , ecl_mdqctl_div_data_next[9] ,
         ecl_mdqctl_div_data_next[8] , ecl_mdqctl_div_data_next[7] ,
         ecl_mdqctl_div_data_next[6] , ecl_mdqctl_div_data_next[5] ,
         ecl_mdqctl_div_data_next[4] , ecl_mdqctl_div_data_next[3] ,
         ecl_mdqctl_div_data_next[2] , ecl_mdqctl_div_data_next[1] ,
         ecl_mdqctl_div_data_next[0] , ecl_mdqctl_new_div_vld ,
         alu_regzcmp_high_nonzero , alu_regzcmp_low_nonzero ,
         alu_addsub_cout64_e , alu_addsub_rs2_data_0 ,
         alu_addsub_rs2_data_1 , alu_addsub_rs2_data_2 ,
         alu_addsub_rs2_data_3 , alu_addsub_rs2_data_4 ,
         alu_addsub_rs2_data_5 , alu_addsub_rs2_data_6 ,
         alu_addsub_rs2_data_7 , alu_addsub_rs2_data_8 ,
         alu_addsub_rs2_data_9 , alu_addsub_rs2_data_10 ,
         alu_addsub_rs2_data_11 , alu_addsub_rs2_data_12 ,
         alu_addsub_rs2_data_13 , alu_addsub_rs2_data_14 ,
         alu_addsub_rs2_data_15 , alu_addsub_rs2_data_16 ,
         alu_addsub_rs2_data_17 , alu_addsub_rs2_data_18 ,
         alu_addsub_rs2_data_19 , alu_addsub_rs2_data_20 ,
         alu_addsub_rs2_data_21 , alu_addsub_rs2_data_22 ,
         alu_addsub_rs2_data_23 , alu_addsub_rs2_data_24 ,
         alu_addsub_rs2_data_25 , alu_addsub_rs2_data_26 ,
         alu_addsub_rs2_data_27 , alu_addsub_rs2_data_28 ,
         alu_addsub_rs2_data_29 , alu_addsub_rs2_data_30 ,
         alu_addsub_rs2_data[32] , alu_addsub_rs2_data[33] ,
         alu_addsub_rs2_data[34] , alu_addsub_rs2_data[35] ,
         alu_addsub_rs2_data[36] , alu_addsub_rs2_data[37] ,
         alu_addsub_rs2_data[38] , alu_addsub_rs2_data[39] ,
         alu_addsub_rs2_data[40] , alu_addsub_rs2_data[41] ,
         alu_addsub_rs2_data[42] , alu_addsub_rs2_data[43] ,
         alu_addsub_rs2_data[44] , alu_addsub_rs2_data[45] ,
         alu_addsub_rs2_data[46] , alu_addsub_rs2_data[47] ,
         alu_addsub_rs2_data[48] , alu_addsub_rs2_data[49] ,
         alu_addsub_rs2_data[50] , alu_addsub_rs2_data[51] ,
         alu_addsub_rs2_data[52] , alu_addsub_rs2_data[53] ,
         alu_addsub_rs2_data[54] , alu_addsub_rs2_data[55] ,
         alu_addsub_rs2_data[56] , alu_addsub_rs2_data[57] ,
         alu_addsub_rs2_data[58] , alu_addsub_rs2_data[59] ,
         alu_addsub_rs2_data[60] , alu_addsub_rs2_data[61] ,
         alu_addsub_rs2_data[62] , alu_addsub_subtract_e[63] ,
         alu_addsub_subtract_e[62] , alu_addsub_subtract_e[61] ,
         alu_addsub_subtract_e[60] , alu_addsub_subtract_e[59] ,
         alu_addsub_subtract_e[58] , alu_addsub_subtract_e[57] ,
         alu_addsub_subtract_e[56] , alu_addsub_subtract_e[55] ,
         alu_addsub_subtract_e[54] , alu_addsub_subtract_e[53] ,
         alu_addsub_subtract_e[52] , alu_addsub_subtract_e[51] ,
         alu_addsub_subtract_e[50] , alu_addsub_subtract_e[49] ,
         alu_addsub_subtract_e[48] , alu_addsub_subtract_e[47] ,
         alu_addsub_subtract_e[46] , alu_addsub_subtract_e[45] ,
         alu_addsub_subtract_e[44] , alu_addsub_subtract_e[43] ,
         alu_addsub_subtract_e[42] , alu_addsub_subtract_e[41] ,
         alu_addsub_subtract_e[40] , alu_addsub_subtract_e[39] ,
         alu_addsub_subtract_e[38] , alu_addsub_subtract_e[37] ,
         alu_addsub_subtract_e[36] , alu_addsub_subtract_e[35] ,
         alu_addsub_subtract_e[34] , alu_addsub_subtract_e[33] ,
         alu_addsub_subtract_e[32] , alu_addsub_subtract_e[31] ,
         alu_addsub_subtract_e[30] , alu_addsub_subtract_e[29] ,
         alu_addsub_subtract_e[28] , alu_addsub_subtract_e[27] ,
         alu_addsub_subtract_e[26] , alu_addsub_subtract_e[25] ,
         alu_addsub_subtract_e[24] , alu_addsub_subtract_e[23] ,
         alu_addsub_subtract_e[22] , alu_addsub_subtract_e[21] ,
         alu_addsub_subtract_e[20] , alu_addsub_subtract_e[19] ,
         alu_addsub_subtract_e[18] , alu_addsub_subtract_e[17] ,
         alu_addsub_subtract_e[16] , alu_addsub_subtract_e[15] ,
         alu_addsub_subtract_e[14] , alu_addsub_subtract_e[13] ,
         alu_addsub_subtract_e[12] , alu_addsub_subtract_e[11] ,
         alu_addsub_subtract_e[10] , alu_addsub_subtract_e[9] ,
         alu_addsub_subtract_e[8] , alu_addsub_subtract_e[7] ,
         alu_addsub_subtract_e[6] , alu_addsub_subtract_e[5] ,
         alu_addsub_subtract_e[4] , alu_addsub_subtract_e[3] ,
         alu_addsub_subtract_e[2] , alu_addsub_subtract_e[1] ,
         alu_addsub_subtract_e[0] , alu_logic_n160 , alu_logic_n159 ,
         alu_logic_n158 , alu_logic_n157 , alu_logic_n156 ,
         alu_logic_n155 , alu_logic_n154 , alu_logic_n153 ,
         alu_logic_n152 , alu_logic_n151 , alu_logic_n150 ,
         alu_logic_n149 , alu_logic_n148 , alu_logic_n147 ,
         alu_logic_n146 , alu_logic_n145 , alu_logic_n144 ,
         alu_logic_n143 , alu_logic_n142 , alu_logic_n141 ,
         alu_logic_n140 , alu_logic_n139 , alu_logic_n138 ,
         alu_logic_n137 , alu_logic_n136 , alu_logic_n135 ,
         alu_logic_n134 , alu_logic_n133 , alu_logic_n132 ,
         alu_logic_n131 , alu_logic_n130 , alu_logic_n129 ,
         alu_logic_n128 , alu_logic_n127 , alu_logic_n126 ,
         alu_logic_n125 , alu_logic_n124 , alu_logic_n123 ,
         alu_logic_n122 , alu_logic_n121 , alu_logic_n120 ,
         alu_logic_n119 , alu_logic_n118 , alu_logic_n117 ,
         alu_logic_n116 , alu_logic_n115 , alu_logic_n114 ,
         alu_logic_n113 , alu_logic_n112 , alu_logic_n111 ,
         alu_logic_n110 , alu_logic_n109 , alu_logic_n108 ,
         alu_logic_n107 , alu_logic_n106 , alu_logic_n105 ,
         alu_logic_n104 , alu_logic_n103 , alu_logic_n102 ,
         alu_logic_n101 , alu_logic_n100 , alu_logic_n99 , alu_logic_n98 ,
         alu_logic_n97 , alu_logic_n96 , alu_logic_n95 , alu_logic_n94 ,
         alu_logic_n93 , alu_logic_n92 , alu_logic_n91 , alu_logic_n90 ,
         alu_logic_n89 , alu_logic_n88 , alu_logic_n87 , alu_logic_n86 ,
         alu_logic_n85 , alu_logic_n84 , alu_logic_n83 , alu_logic_n82 ,
         alu_logic_n81 , alu_logic_n80 , alu_logic_n79 , alu_logic_n78 ,
         alu_logic_n77 , alu_logic_n76 , alu_logic_n75 , alu_logic_n74 ,
         alu_logic_n73 , alu_logic_n72 , alu_logic_n71 , alu_logic_n70 ,
         alu_logic_n69 , alu_logic_n68 , alu_logic_n67 , alu_logic_n66 ,
         alu_logic_n65 , alu_logic_n64 , alu_logic_n63 , alu_logic_n62 ,
         alu_logic_n61 , alu_logic_n60 , alu_logic_n59 , alu_logic_n58 ,
         alu_logic_n57 , alu_logic_n56 , alu_logic_n55 , alu_logic_n54 ,
         alu_logic_n53 , alu_logic_n52 , alu_logic_n51 , alu_logic_n50 ,
         alu_logic_n49 , alu_logic_n48 , alu_logic_n47 , alu_logic_n46 ,
         alu_logic_n45 , alu_logic_n44 , alu_logic_n43 , alu_logic_n42 ,
         alu_logic_n41 , alu_logic_n40 , alu_logic_n39 , alu_logic_n38 ,
         alu_logic_n37 , alu_logic_n36 , alu_logic_n35 , alu_logic_n34 ,
         alu_logic_n33 , alu_logic_rs1_data_bf1[0] ,
         alu_logic_rs1_data_bf1[1] , alu_logic_rs1_data_bf1[2] ,
         alu_logic_rs1_data_bf1[3] , alu_logic_rs1_data_bf1[4] ,
         alu_logic_rs1_data_bf1[5] , alu_logic_rs1_data_bf1[6] ,
         alu_logic_rs1_data_bf1[7] , alu_logic_rs1_data_bf1[8] ,
         alu_logic_rs1_data_bf1[9] , alu_logic_rs1_data_bf1[10] ,
         alu_logic_rs1_data_bf1[11] , alu_logic_rs1_data_bf1[12] ,
         alu_logic_rs1_data_bf1[13] , alu_logic_rs1_data_bf1[14] ,
         alu_logic_rs1_data_bf1[15] , alu_logic_rs1_data_bf1[16] ,
         alu_logic_rs1_data_bf1[17] , alu_logic_rs1_data_bf1[18] ,
         alu_logic_rs1_data_bf1[19] , alu_logic_rs1_data_bf1[20] ,
         alu_logic_rs1_data_bf1[21] , alu_logic_rs1_data_bf1[22] ,
         alu_logic_rs1_data_bf1[23] , alu_logic_rs1_data_bf1[24] ,
         alu_logic_rs1_data_bf1[25] , alu_logic_rs1_data_bf1[26] ,
         alu_logic_rs1_data_bf1[27] , alu_logic_rs1_data_bf1[28] ,
         alu_logic_rs1_data_bf1[29] , alu_logic_rs1_data_bf1[30] ,
         alu_logic_rs1_data_bf1[31] , alu_logic_rs1_data_bf1[32] ,
         alu_logic_rs1_data_bf1[33] , alu_logic_rs1_data_bf1[34] ,
         alu_logic_rs1_data_bf1[35] , alu_logic_rs1_data_bf1[36] ,
         alu_logic_rs1_data_bf1[37] , alu_logic_rs1_data_bf1[38] ,
         alu_logic_rs1_data_bf1[39] , alu_logic_rs1_data_bf1[40] ,
         alu_logic_rs1_data_bf1[41] , alu_logic_rs1_data_bf1[42] ,
         alu_logic_rs1_data_bf1[43] , alu_logic_rs1_data_bf1[44] ,
         alu_logic_rs1_data_bf1[45] , alu_logic_rs1_data_bf1[46] ,
         alu_logic_rs1_data_bf1[47] , alu_logic_rs1_data_bf1[48] ,
         alu_logic_rs1_data_bf1[49] , alu_logic_rs1_data_bf1[50] ,
         alu_logic_rs1_data_bf1[51] , alu_logic_rs1_data_bf1[52] ,
         alu_logic_rs1_data_bf1[53] , alu_logic_rs1_data_bf1[54] ,
         alu_logic_rs1_data_bf1[55] , alu_logic_rs1_data_bf1[56] ,
         alu_logic_rs1_data_bf1[57] , alu_logic_rs1_data_bf1[58] ,
         alu_logic_rs1_data_bf1[59] , alu_logic_rs1_data_bf1[60] ,
         alu_logic_rs1_data_bf1[61] , alu_logic_rs1_data_bf1[62] ,
         alu_logic_rs1_data_bf1[63] , alu_logic_mov_data[63] ,
         alu_logic_mov_data[62] , alu_logic_mov_data[61] ,
         alu_logic_mov_data[60] , alu_logic_mov_data[59] ,
         alu_logic_mov_data[58] , alu_logic_mov_data[57] ,
         alu_logic_mov_data[56] , alu_logic_mov_data[55] ,
         alu_logic_mov_data[54] , alu_logic_mov_data[53] ,
         alu_logic_mov_data[52] , alu_logic_mov_data[51] ,
         alu_logic_mov_data[50] , alu_logic_mov_data[49] ,
         alu_logic_mov_data[48] , alu_logic_mov_data[47] ,
         alu_logic_mov_data[46] , alu_logic_mov_data[45] ,
         alu_logic_mov_data[44] , alu_logic_mov_data[43] ,
         alu_logic_mov_data[42] , alu_logic_mov_data[41] ,
         alu_logic_mov_data[40] , alu_logic_mov_data[39] ,
         alu_logic_mov_data[38] , alu_logic_mov_data[37] ,
         alu_logic_mov_data[36] , alu_logic_mov_data[35] ,
         alu_logic_mov_data[34] , alu_logic_mov_data[33] ,
         alu_logic_mov_data[32] , alu_logic_result_xor[63] ,
         alu_logic_result_xor[62] , alu_logic_result_xor[61] ,
         alu_logic_result_xor[60] , alu_logic_result_xor[59] ,
         alu_logic_result_xor[58] , alu_logic_result_xor[57] ,
         alu_logic_result_xor[56] , alu_logic_result_xor[55] ,
         alu_logic_result_xor[54] , alu_logic_result_xor[53] ,
         alu_logic_result_xor[52] , alu_logic_result_xor[51] ,
         alu_logic_result_xor[50] , alu_logic_result_xor[49] ,
         alu_logic_result_xor[48] , alu_logic_result_xor[47] ,
         alu_logic_result_xor[46] , alu_logic_result_xor[45] ,
         alu_logic_result_xor[44] , alu_logic_result_xor[43] ,
         alu_logic_result_xor[42] , alu_logic_result_xor[41] ,
         alu_logic_result_xor[40] , alu_logic_result_xor[39] ,
         alu_logic_result_xor[38] , alu_logic_result_xor[37] ,
         alu_logic_result_xor[36] , alu_logic_result_xor[35] ,
         alu_logic_result_xor[34] , alu_logic_result_xor[33] ,
         alu_logic_result_xor[32] , alu_logic_result_xor[31] ,
         alu_logic_result_xor[30] , alu_logic_result_xor[29] ,
         alu_logic_result_xor[28] , alu_logic_result_xor[27] ,
         alu_logic_result_xor[26] , alu_logic_result_xor[25] ,
         alu_logic_result_xor[24] , alu_logic_result_xor[23] ,
         alu_logic_result_xor[22] , alu_logic_result_xor[21] ,
         alu_logic_result_xor[20] , alu_logic_result_xor[19] ,
         alu_logic_result_xor[18] , alu_logic_result_xor[17] ,
         alu_logic_result_xor[16] , alu_logic_result_xor[15] ,
         alu_logic_result_xor[14] , alu_logic_result_xor[13] ,
         alu_logic_result_xor[12] , alu_logic_result_xor[11] ,
         alu_logic_result_xor[10] , alu_logic_result_xor[9] ,
         alu_logic_result_xor[8] , alu_logic_result_xor[7] ,
         alu_logic_result_xor[6] , alu_logic_result_xor[5] ,
         alu_logic_result_xor[4] , alu_logic_result_xor[3] ,
         alu_logic_result_xor[2] , alu_logic_result_xor[1] ,
         alu_logic_result_xor[0] , alu_logic_result_or[63] ,
         alu_logic_result_or[62] , alu_logic_result_or[61] ,
         alu_logic_result_or[60] , alu_logic_result_or[59] ,
         alu_logic_result_or[58] , alu_logic_result_or[57] ,
         alu_logic_result_or[56] , alu_logic_result_or[55] ,
         alu_logic_result_or[54] , alu_logic_result_or[53] ,
         alu_logic_result_or[52] , alu_logic_result_or[51] ,
         alu_logic_result_or[50] , alu_logic_result_or[49] ,
         alu_logic_result_or[48] , alu_logic_result_or[47] ,
         alu_logic_result_or[46] , alu_logic_result_or[45] ,
         alu_logic_result_or[44] , alu_logic_result_or[43] ,
         alu_logic_result_or[42] , alu_logic_result_or[41] ,
         alu_logic_result_or[40] , alu_logic_result_or[39] ,
         alu_logic_result_or[38] , alu_logic_result_or[37] ,
         alu_logic_result_or[36] , alu_logic_result_or[35] ,
         alu_logic_result_or[34] , alu_logic_result_or[33] ,
         alu_logic_result_or[32] , alu_logic_result_or[31] ,
         alu_logic_result_or[30] , alu_logic_result_or[29] ,
         alu_logic_result_or[28] , alu_logic_result_or[27] ,
         alu_logic_result_or[26] , alu_logic_result_or[25] ,
         alu_logic_result_or[24] , alu_logic_result_or[23] ,
         alu_logic_result_or[22] , alu_logic_result_or[21] ,
         alu_logic_result_or[20] , alu_logic_result_or[19] ,
         alu_logic_result_or[18] , alu_logic_result_or[17] ,
         alu_logic_result_or[16] , alu_logic_result_or[15] ,
         alu_logic_result_or[14] , alu_logic_result_or[13] ,
         alu_logic_result_or[12] , alu_logic_result_or[11] ,
         alu_logic_result_or[10] , alu_logic_result_or[9] ,
         alu_logic_result_or[8] , alu_logic_result_or[7] ,
         alu_logic_result_or[6] , alu_logic_result_or[5] ,
         alu_logic_result_or[4] , alu_logic_result_or[3] ,
         alu_logic_result_or[2] , alu_logic_result_or[1] ,
         alu_logic_result_or[0] , alu_logic_result_and[63] ,
         alu_logic_result_and[62] , alu_logic_result_and[61] ,
         alu_logic_result_and[60] , alu_logic_result_and[59] ,
         alu_logic_result_and[58] , alu_logic_result_and[57] ,
         alu_logic_result_and[56] , alu_logic_result_and[55] ,
         alu_logic_result_and[54] , alu_logic_result_and[53] ,
         alu_logic_result_and[52] , alu_logic_result_and[51] ,
         alu_logic_result_and[50] , alu_logic_result_and[49] ,
         alu_logic_result_and[48] , alu_logic_result_and[47] ,
         alu_logic_result_and[46] , alu_logic_result_and[45] ,
         alu_logic_result_and[44] , alu_logic_result_and[43] ,
         alu_logic_result_and[42] , alu_logic_result_and[41] ,
         alu_logic_result_and[40] , alu_logic_result_and[39] ,
         alu_logic_result_and[38] , alu_logic_result_and[37] ,
         alu_logic_result_and[36] , alu_logic_result_and[35] ,
         alu_logic_result_and[34] , alu_logic_result_and[33] ,
         alu_logic_result_and[32] , alu_logic_result_and[31] ,
         alu_logic_result_and[30] , alu_logic_result_and[29] ,
         alu_logic_result_and[28] , alu_logic_result_and[27] ,
         alu_logic_result_and[26] , alu_logic_result_and[25] ,
         alu_logic_result_and[24] , alu_logic_result_and[23] ,
         alu_logic_result_and[22] , alu_logic_result_and[21] ,
         alu_logic_result_and[20] , alu_logic_result_and[19] ,
         alu_logic_result_and[18] , alu_logic_result_and[17] ,
         alu_logic_result_and[16] , alu_logic_result_and[15] ,
         alu_logic_result_and[14] , alu_logic_result_and[13] ,
         alu_logic_result_and[12] , alu_logic_result_and[11] ,
         alu_logic_result_and[10] , alu_logic_result_and[9] ,
         alu_logic_result_and[8] , alu_logic_result_and[7] ,
         alu_logic_result_and[6] , alu_logic_result_and[5] ,
         alu_logic_result_and[4] , alu_logic_result_and[3] ,
         alu_logic_result_and[2] , alu_logic_result_and[1] ,
         alu_logic_result_and[0] , alu_chk_mem_addr_n30 ,
         alu_chk_mem_addr_n29 , alu_chk_mem_addr_n28 ,
         alu_chk_mem_addr_n27 , alu_chk_mem_addr_n26 ,
         alu_chk_mem_addr_n25 , alu_chk_mem_addr_n24 ,
         alu_chk_mem_addr_n23 , alu_chk_mem_addr_n22 ,
         alu_chk_mem_addr_n21 , alu_chk_mem_addr_n20 ,
         alu_chk_mem_addr_n19 , alu_chk_mem_addr_n18 ,
         alu_chk_mem_addr_n17 , alu_chk_mem_addr_n16 ,
         alu_chk_mem_addr_n15 , alu_chk_mem_addr_n14 ,
         alu_chk_mem_addr_n13 , alu_chk_mem_addr_n12 ,
         alu_chk_mem_addr_n11 , alu_chk_mem_addr_n10 , alu_chk_mem_addr_n9 ,
         alu_chk_mem_addr_n8 , alu_chk_mem_addr_n7 , alu_chk_mem_addr_n6 ,
         alu_chk_mem_addr_n5 , alu_chk_mem_addr_n4 , alu_chk_mem_addr_n3 ,
         alu_chk_mem_addr_n2 , alu_chk_mem_addr_n1 ,
         shft_mux_rshift_extend_n65 , shft_mux_rshift_extend_n64 ,
         shft_mux_rshift_extend_n63 , shft_mux_rshift_extend_n62 ,
         shft_mux_rshift_extend_n61 , shft_mux_rshift_extend_n60 ,
         shft_mux_rshift_extend_n59 , shft_mux_rshift_extend_n58 ,
         shft_mux_rshift_extend_n57 , shft_mux_rshift_extend_n56 ,
         shft_mux_rshift_extend_n55 , shft_mux_rshift_extend_n54 ,
         shft_mux_rshift_extend_n53 , shft_mux_rshift_extend_n52 ,
         shft_mux_rshift_extend_n51 , shft_mux_rshift_extend_n49 ,
         shft_mux_rshift_extend_n47 , shft_mux_rshift_extend_n45 ,
         shft_mux_rshift_extend_n43 , shft_mux_rshift_extend_n42 ,
         shft_mux_rshift_extend_n41 , shft_mux_rshift_extend_n39 ,
         shft_mux_rshift_extend_n37 , shft_mux_rshift_extend_n35 ,
         shft_mux_rshift_extend_n33 , shft_mux_rshift_extend_n31 ,
         shft_mux_rshift_extend_n30 , shft_mux_rshift_extend_n29 ,
         shft_mux_rshift_extend_n27 , shft_mux_rshift_extend_n25 ,
         shft_mux_rshift_extend_n24 , shft_mux_rshift_extend_n23 ,
         shft_mux_rshift_extend_n22 , shft_mux_rshift_extend_n21 ,
         shft_mux_rshift_extend_n20 , shft_mux_rshift_extend_n19 ,
         shft_mux_rshift_extend_n18 , shft_mux_rshift_extend_n17 ,
         shft_mux_rshift_extend_n16 , shft_mux_rshift_extend_n15 ,
         shft_mux_rshift_extend_n14 , shft_mux_rshift_extend_n13 ,
         shft_mux_rshift_extend_n12 , shft_mux_rshift_extend_n11 ,
         shft_mux_rshift_extend_n10 , shft_mux_rshift_extend_n9 ,
         shft_mux_rshift_extend_n8 , shft_mux_rshift_extend_n7 ,
         shft_mux_rshift_extend_n6 , shft_mux_rshift_extend_n5 ,
         shft_mux_rshift_extend_n4 , shft_mux_rshift_extend_n3 ,
         shft_mux_rshift_extend_n2 , div_u32eql_notequal ,
         div_u32eql_inxor[31] , div_u32eql_inxor[30] ,
         div_u32eql_inxor[29] , div_u32eql_inxor[28] ,
         div_u32eql_inxor[27] , div_u32eql_inxor[26] ,
         div_u32eql_inxor[25] , div_u32eql_inxor[24] ,
         div_u32eql_inxor[23] , div_u32eql_inxor[22] ,
         div_u32eql_inxor[21] , div_u32eql_inxor[20] ,
         div_u32eql_inxor[19] , div_u32eql_inxor[18] ,
         div_u32eql_inxor[17] , div_u32eql_inxor[16] ,
         div_u32eql_inxor[15] , div_u32eql_inxor[14] ,
         div_u32eql_inxor[13] , div_u32eql_inxor[12] ,
         div_u32eql_inxor[11] , div_u32eql_inxor[9] , div_u32eql_inxor[8] ,
         div_u32eql_inxor[7] , div_u32eql_inxor[6] , div_u32eql_inxor[5] ,
         div_u32eql_inxor[4] , div_u32eql_inxor[3] , div_u32eql_inxor[2] ,
         div_u32eql_inxor[1] , div_low32or_n30 , div_low32or_n29 ,
         div_low32or_n28 , div_low32or_n27 , div_low32or_n26 ,
         div_low32or_n25 , div_low32or_n24 , div_low32or_n23 ,
         div_low32or_n22 , div_low32or_n21 , div_low32or_n20 ,
         div_low32or_n19 , div_low32or_n18 , div_low32or_n17 ,
         div_low32or_n16 , div_low32or_n15 , div_low32or_n14 ,
         div_low32or_n13 , div_low32or_n12 , div_low32or_n11 ,
         div_low32or_n10 , div_low32or_n9 , div_low32or_n8 ,
         div_low32or_n7 , div_low32or_n6 , div_low32or_n5 ,
         div_low32or_n4 , div_low32or_n3 , div_low32or_n2 ,
         div_low32or_n1 , div_d_mux_n512 , div_d_mux_n511 ,
         div_d_mux_n510 , div_d_mux_n509 , div_d_mux_n508 ,
         div_d_mux_n507 , div_d_mux_n505 , div_d_mux_n504 ,
         div_d_mux_n503 , div_d_mux_n501 , div_d_mux_n500 ,
         div_d_mux_n499 , div_d_mux_n497 , div_d_mux_n496 ,
         div_d_mux_n495 , div_d_mux_n493 , div_d_mux_n492 ,
         div_d_mux_n491 , div_d_mux_n489 , div_d_mux_n488 ,
         div_d_mux_n487 , div_d_mux_n485 , div_d_mux_n484 ,
         div_d_mux_n483 , div_d_mux_n481 , div_d_mux_n480 ,
         div_d_mux_n479 , div_d_mux_n477 , div_d_mux_n476 ,
         div_d_mux_n475 , div_d_mux_n473 , div_d_mux_n472 ,
         div_d_mux_n471 , div_d_mux_n469 , div_d_mux_n468 ,
         div_d_mux_n467 , div_d_mux_n466 , div_d_mux_n465 ,
         div_d_mux_n464 , div_d_mux_n463 , div_d_mux_n461 ,
         div_d_mux_n460 , div_d_mux_n459 , div_d_mux_n457 ,
         div_d_mux_n456 , div_d_mux_n455 , div_d_mux_n453 ,
         div_d_mux_n452 , div_d_mux_n451 , div_d_mux_n449 ,
         div_d_mux_n448 , div_d_mux_n447 , div_d_mux_n445 ,
         div_d_mux_n444 , div_d_mux_n443 , div_d_mux_n441 ,
         div_d_mux_n440 , div_d_mux_n439 , div_d_mux_n437 ,
         div_d_mux_n436 , div_d_mux_n435 , div_d_mux_n433 ,
         div_d_mux_n432 , div_d_mux_n431 , div_d_mux_n429 ,
         div_d_mux_n428 , div_d_mux_n427 , div_d_mux_n425 ,
         div_d_mux_n424 , div_d_mux_n423 , div_d_mux_n422 ,
         div_d_mux_n421 , div_d_mux_n420 , div_d_mux_n419 ,
         div_d_mux_n417 , div_d_mux_n416 , div_d_mux_n415 ,
         div_d_mux_n413 , div_d_mux_n412 , div_d_mux_n411 ,
         div_d_mux_n409 , div_d_mux_n408 , div_d_mux_n407 ,
         div_d_mux_n405 , div_d_mux_n404 , div_d_mux_n403 ,
         div_d_mux_n401 , div_d_mux_n400 , div_d_mux_n399 ,
         div_d_mux_n397 , div_d_mux_n396 , div_d_mux_n395 ,
         div_d_mux_n393 , div_d_mux_n392 , div_d_mux_n391 ,
         div_d_mux_n389 , div_d_mux_n388 , div_d_mux_n387 ,
         div_d_mux_n386 , div_d_mux_n385 , div_d_mux_n384 ,
         div_d_mux_n383 , div_d_mux_n382 , div_d_mux_n381 ,
         div_d_mux_n380 , div_d_mux_n379 , div_d_mux_n378 ,
         div_d_mux_n377 , div_d_mux_n376 , div_d_mux_n375 ,
         div_d_mux_n374 , div_d_mux_n373 , div_d_mux_n372 ,
         div_d_mux_n371 , div_d_mux_n370 , div_d_mux_n369 ,
         div_d_mux_n368 , div_d_mux_n367 , div_d_mux_n366 ,
         div_d_mux_n365 , div_d_mux_n364 , div_d_mux_n363 ,
         div_d_mux_n362 , div_d_mux_n361 , div_d_mux_n360 ,
         div_d_mux_n359 , div_d_mux_n358 , div_d_mux_n357 ,
         div_d_mux_n356 , div_d_mux_n355 , div_d_mux_n354 ,
         div_d_mux_n353 , div_d_mux_n352 , div_d_mux_n351 ,
         div_d_mux_n350 , div_d_mux_n349 , div_d_mux_n348 ,
         div_d_mux_n347 , div_d_mux_n346 , div_d_mux_n345 ,
         div_d_mux_n344 , div_d_mux_n343 , div_d_mux_n342 ,
         div_d_mux_n341 , div_d_mux_n340 , div_d_mux_n339 ,
         div_d_mux_n338 , div_d_mux_n337 , div_d_mux_n336 ,
         div_d_mux_n335 , div_d_mux_n334 , div_d_mux_n333 ,
         div_d_mux_n332 , div_d_mux_n331 , div_d_mux_n330 ,
         div_d_mux_n329 , div_d_mux_n328 , div_d_mux_n327 ,
         div_d_mux_n326 , div_d_mux_n325 , div_d_mux_n324 ,
         div_d_mux_n323 , div_d_mux_n322 , div_d_mux_n321 ,
         div_d_mux_n320 , div_d_mux_n319 , div_d_mux_n318 ,
         div_d_mux_n317 , div_d_mux_n316 , div_d_mux_n315 ,
         div_d_mux_n314 , div_d_mux_n313 , div_d_mux_n312 ,
         div_d_mux_n311 , div_d_mux_n310 , div_d_mux_n309 ,
         div_d_mux_n308 , div_d_mux_n307 , div_d_mux_n306 ,
         div_d_mux_n305 , div_d_mux_n304 , div_d_mux_n303 ,
         div_d_mux_n302 , div_d_mux_n301 , div_d_mux_n300 ,
         div_d_mux_n299 , div_d_mux_n298 , div_d_mux_n297 ,
         div_d_mux_n296 , div_d_mux_n295 , div_d_mux_n294 ,
         div_d_mux_n293 , div_d_mux_n292 , div_d_mux_n291 ,
         div_d_mux_n290 , div_d_mux_n289 , div_d_mux_n288 ,
         div_d_mux_n287 , div_d_mux_n286 , div_d_mux_n285 ,
         div_d_mux_n284 , div_d_mux_n283 , div_d_mux_n282 ,
         div_d_mux_n281 , div_d_mux_n280 , div_d_mux_n279 ,
         div_d_mux_n278 , div_d_mux_n277 , div_d_mux_n276 ,
         div_d_mux_n275 , div_d_mux_n274 , div_d_mux_n273 ,
         div_d_mux_n272 , div_d_mux_n271 , div_d_mux_n270 ,
         div_d_mux_n269 , div_d_mux_n268 , div_d_mux_n267 ,
         div_d_mux_n266 , div_d_mux_n265 , div_d_mux_n264 ,
         div_d_mux_n263 , div_d_mux_n262 , div_d_mux_n261 ,
         div_d_mux_n260 , div_d_mux_n259 , div_d_mux_n258 ,
         div_d_mux_n257 , div_d_mux_n256 , div_d_mux_n255 ,
         div_d_mux_n254 , div_d_mux_n253 , div_d_mux_n252 ,
         div_d_mux_n251 , div_d_mux_n250 , div_d_mux_n249 ,
         div_d_mux_n248 , div_d_mux_n247 , div_d_mux_n246 ,
         div_d_mux_n245 , div_d_mux_n244 , div_d_mux_n243 ,
         div_d_mux_n242 , div_d_mux_n241 , div_d_mux_n240 ,
         div_d_mux_n239 , div_d_mux_n238 , div_d_mux_n237 ,
         div_d_mux_n236 , div_d_mux_n235 , div_d_mux_n234 ,
         div_d_mux_n233 , div_d_mux_n232 , div_d_mux_n231 ,
         div_d_mux_n230 , div_d_mux_n229 , div_d_mux_n228 ,
         div_d_mux_n227 , div_d_mux_n226 , div_d_mux_n225 ,
         div_d_mux_n224 , div_d_mux_n223 , div_d_mux_n222 ,
         div_d_mux_n221 , div_d_mux_n220 , div_d_mux_n219 ,
         div_d_mux_n218 , div_d_mux_n217 , div_d_mux_n216 ,
         div_d_mux_n215 , div_d_mux_n214 , div_d_mux_n213 ,
         div_d_mux_n212 , div_d_mux_n211 , div_d_mux_n210 ,
         div_d_mux_n209 , div_d_mux_n208 , div_d_mux_n207 ,
         div_d_mux_n206 , div_d_mux_n205 , div_d_mux_n204 ,
         div_d_mux_n203 , div_d_mux_n202 , div_d_mux_n201 ,
         div_d_mux_n200 , div_d_mux_n199 , div_d_mux_n198 ,
         div_d_mux_n197 , div_d_mux_n196 , div_d_mux_n195 ,
         div_d_mux_n194 , div_d_mux_n193 , div_d_mux_n192 ,
         div_d_mux_n191 , div_d_mux_n190 , div_d_mux_n189 ,
         div_d_mux_n188 , div_d_mux_n187 , div_d_mux_n186 ,
         div_d_mux_n185 , div_d_mux_n184 , div_d_mux_n183 ,
         div_d_mux_n182 , div_d_mux_n181 , div_d_mux_n180 ,
         div_d_mux_n179 , div_d_mux_n178 , div_d_mux_n177 ,
         div_d_mux_n176 , div_d_mux_n175 , div_d_mux_n174 ,
         div_d_mux_n173 , div_d_mux_n172 , div_d_mux_n171 ,
         div_d_mux_n170 , div_d_mux_n169 , div_d_mux_n168 ,
         div_d_mux_n167 , div_d_mux_n166 , div_d_mux_n165 ,
         div_d_mux_n164 , div_d_mux_n163 , div_d_mux_n162 ,
         div_d_mux_n161 , div_d_mux_n160 , div_d_mux_n159 ,
         div_d_mux_n158 , div_d_mux_n157 , div_d_mux_n156 ,
         div_d_mux_n155 , div_d_mux_n154 , div_d_mux_n153 ,
         div_d_mux_n152 , div_d_mux_n151 , div_d_mux_n150 ,
         div_d_mux_n149 , div_d_mux_n148 , div_d_mux_n147 ,
         div_d_mux_n146 , div_d_mux_n145 , div_d_mux_n144 ,
         div_d_mux_n143 , div_d_mux_n142 , div_d_mux_n141 ,
         div_d_mux_n140 , div_d_mux_n139 , div_d_mux_n138 ,
         div_d_mux_n137 , div_d_mux_n136 , div_d_mux_n135 ,
         div_d_mux_n134 , div_d_mux_n133 , div_d_mux_n132 ,
         div_d_mux_n131 , div_d_mux_n130 , div_d_mux_n129 ,
         div_d_mux_n128 , div_d_mux_n127 , div_d_mux_n126 ,
         div_d_mux_n125 , div_d_mux_n124 , div_d_mux_n123 ,
         div_d_mux_n122 , div_d_mux_n121 , div_d_mux_n120 ,
         div_d_mux_n119 , div_d_mux_n118 , div_d_mux_n117 ,
         div_d_mux_n116 , div_d_mux_n115 , div_d_mux_n114 ,
         div_d_mux_n113 , div_d_mux_n112 , div_d_mux_n111 ,
         div_d_mux_n110 , div_d_mux_n109 , div_d_mux_n108 ,
         div_d_mux_n107 , div_d_mux_n106 , div_d_mux_n105 ,
         div_d_mux_n104 , div_d_mux_n103 , div_d_mux_n102 ,
         div_d_mux_n101 , div_d_mux_n100 , div_d_mux_n99 , div_d_mux_n98 ,
         div_d_mux_n97 , div_d_mux_n96 , div_d_mux_n95 , div_d_mux_n94 ,
         div_d_mux_n93 , div_d_mux_n92 , div_d_mux_n91 , div_d_mux_n90 ,
         div_d_mux_n89 , div_d_mux_n88 , div_d_mux_n87 , div_d_mux_n86 ,
         div_d_mux_n85 , div_d_mux_n84 , div_d_mux_n83 , div_d_mux_n82 ,
         div_d_mux_n81 , div_d_mux_n80 , div_d_mux_n79 , div_d_mux_n78 ,
         div_d_mux_n77 , div_d_mux_n76 , div_d_mux_n75 , div_d_mux_n74 ,
         div_d_mux_n73 , div_d_mux_n72 , div_d_mux_n71 , div_d_mux_n70 ,
         div_d_mux_n69 , div_d_mux_n68 , div_d_mux_n67 , div_d_mux_n66 ,
         div_d_mux_n65 , div_d_mux_n64 , div_d_mux_n63 , div_d_mux_n62 ,
         div_d_mux_n61 , div_d_mux_n60 , div_d_mux_n59 , div_d_mux_n58 ,
         div_d_mux_n57 , div_d_mux_n56 , div_d_mux_n55 , div_d_mux_n54 ,
         div_d_mux_n53 , div_d_mux_n52 , div_d_mux_n51 , div_d_mux_n50 ,
         div_d_mux_n49 , div_d_mux_n48 , div_d_mux_n47 , div_d_mux_n46 ,
         div_d_mux_n45 , div_d_mux_n44 , div_d_mux_n43 , div_d_mux_n42 ,
         div_d_mux_n41 , div_d_mux_n40 , div_d_mux_n39 , div_d_mux_n38 ,
         div_d_mux_n37 , div_d_mux_n36 , div_d_mux_n35 , div_d_mux_n34 ,
         div_d_mux_n33 , div_d_mux_n32 , div_d_mux_n31 , div_d_mux_n30 ,
         div_d_mux_n29 , div_d_mux_n28 , div_d_mux_n27 , div_d_mux_n26 ,
         div_d_mux_n25 , div_d_mux_n24 , div_d_mux_n23 , div_d_mux_n21 ,
         div_d_mux_n20 , div_d_mux_n19 , div_d_mux_n17 , div_d_mux_n16 ,
         div_d_mux_n15 , div_d_mux_n13 , div_d_mux_n12 , div_d_mux_n11 ,
         div_d_mux_n9 , div_d_mux_n8 , div_d_mux_n7 , div_d_mux_n5 ,
         div_d_mux_n4 , div_d_mux_n3 , div_d_mux_n2 , div_d_mux_n1 ,
         div_d_dff_n257 , div_d_dff_n255 , div_d_dff_n253 ,
         div_d_dff_n251 , div_d_dff_n249 , div_d_dff_n247 ,
         div_d_dff_n245 , div_d_dff_n243 , div_d_dff_n241 ,
         div_d_dff_n239 , div_d_dff_n237 , div_d_dff_n235 ,
         div_d_dff_n233 , div_d_dff_n231 , div_d_dff_n229 ,
         div_d_dff_n227 , div_d_dff_n225 , div_d_dff_n223 ,
         div_d_dff_n221 , div_d_dff_n219 , div_d_dff_n217 ,
         div_d_dff_n215 , div_d_dff_n213 , div_d_dff_n211 ,
         div_d_dff_n209 , div_d_dff_n207 , div_d_dff_n205 ,
         div_d_dff_n203 , div_d_dff_n201 , div_d_dff_n199 ,
         div_d_dff_n197 , div_d_dff_n195 , div_d_dff_n193 ,
         div_d_dff_n191 , div_d_dff_n189 , div_d_dff_n187 ,
         div_d_dff_n185 , div_d_dff_n183 , div_d_dff_n181 ,
         div_d_dff_n179 , div_d_dff_n177 , div_d_dff_n175 ,
         div_d_dff_n173 , div_d_dff_n171 , div_d_dff_n169 ,
         div_d_dff_n167 , div_d_dff_n165 , div_d_dff_n163 ,
         div_d_dff_n161 , div_d_dff_n159 , div_d_dff_n157 ,
         div_d_dff_n155 , div_d_dff_n153 , div_d_dff_n151 ,
         div_d_dff_n149 , div_d_dff_n147 , div_d_dff_n145 ,
         div_d_dff_n143 , div_d_dff_n141 , div_d_dff_n139 ,
         div_d_dff_n137 , div_d_dff_n135 , div_d_dff_n133 ,
         div_d_dff_n131 , div_d_dff_n129 , div_d_dff_n127 ,
         div_d_dff_n125 , div_d_dff_n123 , div_d_dff_n121 ,
         div_d_dff_n119 , div_d_dff_n117 , div_d_dff_n115 ,
         div_d_dff_n113 , div_d_dff_n111 , div_d_dff_n109 ,
         div_d_dff_n107 , div_d_dff_n105 , div_d_dff_n103 ,
         div_d_dff_n101 , div_d_dff_n99 , div_d_dff_n97 , div_d_dff_n95 ,
         div_d_dff_n93 , div_d_dff_n91 , div_d_dff_n89 , div_d_dff_n87 ,
         div_d_dff_n85 , div_d_dff_n83 , div_d_dff_n81 , div_d_dff_n79 ,
         div_d_dff_n77 , div_d_dff_n75 , div_d_dff_n73 , div_d_dff_n71 ,
         div_d_dff_n69 , div_d_dff_n67 , div_d_dff_n65 , div_d_dff_n63 ,
         div_d_dff_n61 , div_d_dff_n59 , div_d_dff_n57 , div_d_dff_n55 ,
         div_d_dff_n53 , div_d_dff_n51 , div_d_dff_n49 , div_d_dff_n47 ,
         div_d_dff_n45 , div_d_dff_n43 , div_d_dff_n41 , div_d_dff_n39 ,
         div_d_dff_n37 , div_d_dff_n35 , div_d_dff_n33 , div_d_dff_n31 ,
         div_d_dff_n29 , div_d_dff_n27 , div_d_dff_n25 , div_d_dff_n23 ,
         div_d_dff_n21 , div_d_dff_n19 , div_d_dff_n17 , div_d_dff_n15 ,
         div_d_dff_n13 , div_d_dff_n11 , div_d_dff_n9 , div_d_dff_n7 ,
         div_d_dff_n5 , div_d_dff_n3 , div_d_dff_n1 , div_spr_n127 ,
         div_spr_n126 , div_spr_n125 , div_spr_n124 , div_spr_n123 ,
         div_spr_n122 , div_spr_n121 , div_spr_n120 , div_spr_n119 ,
         div_spr_n118 , div_spr_n117 , div_spr_n116 , div_spr_n115 ,
         div_spr_n114 , div_spr_n113 , div_spr_n112 , div_spr_n111 ,
         div_spr_n110 , div_spr_n109 , div_spr_n108 , div_spr_n107 ,
         div_spr_n106 , div_spr_n105 , div_spr_n104 , div_spr_n103 ,
         div_spr_n102 , div_spr_n101 , div_spr_n100 , div_spr_n99 ,
         div_spr_n98 , div_spr_n97 , div_spr_n96 , div_spr_n95 ,
         div_spr_n94 , div_spr_n93 , div_spr_n92 , div_spr_n91 ,
         div_spr_n90 , div_spr_n89 , div_spr_n88 , div_spr_n87 ,
         div_spr_n86 , div_spr_n85 , div_spr_n84 , div_spr_n83 ,
         div_spr_n82 , div_spr_n81 , div_spr_n80 , div_spr_n79 ,
         div_spr_n78 , div_spr_n77 , div_spr_n76 , div_spr_n75 ,
         div_spr_n74 , div_spr_n73 , div_spr_n72 , div_spr_n71 ,
         div_spr_n70 , div_spr_n69 , div_spr_n68 , div_spr_n67 ,
         div_spr_n66 , div_spr_n65 , div_spr_n64 , div_spr_n63 ,
         div_spr_n62 , div_spr_n61 , div_spr_n60 , div_spr_n59 ,
         div_spr_n58 , div_spr_n57 , div_spr_n56 , div_spr_n55 ,
         div_spr_n54 , div_spr_n53 , div_spr_n52 , div_spr_n51 ,
         div_spr_n50 , div_spr_n49 , div_spr_n48 , div_spr_n47 ,
         div_spr_n46 , div_spr_n45 , div_spr_n44 , div_spr_n43 ,
         div_spr_n42 , div_spr_n41 , div_spr_n40 , div_spr_n39 ,
         div_spr_n38 , div_spr_n37 , div_spr_n36 , div_spr_n35 ,
         div_spr_n34 , div_spr_n33 , div_spr_n32 , div_spr_n31 ,
         div_spr_n30 , div_spr_n29 , div_spr_n28 , div_spr_n27 ,
         div_spr_n26 , div_spr_n25 , div_spr_n24 , div_spr_n23 ,
         div_spr_n22 , div_spr_n21 , div_spr_n20 , div_spr_n19 ,
         div_spr_n18 , div_spr_n17 , div_spr_n16 , div_spr_n15 ,
         div_spr_n14 , div_spr_n13 , div_spr_n12 , div_spr_n11 ,
         div_spr_n10 , div_spr_n9 , div_spr_n8 , div_spr_n7 , div_spr_n6 ,
         div_spr_n5 , div_spr_n4 , div_spr_n3 , div_spr_n2 , div_spr_n1 ,
         div_yreg_next_yreg_thr3[31] , div_yreg_next_yreg_thr3[30] ,
         div_yreg_next_yreg_thr3[29] , div_yreg_next_yreg_thr3[28] ,
         div_yreg_next_yreg_thr3[27] , div_yreg_next_yreg_thr3[26] ,
         div_yreg_next_yreg_thr3[25] , div_yreg_next_yreg_thr3[24] ,
         div_yreg_next_yreg_thr3[23] , div_yreg_next_yreg_thr3[22] ,
         div_yreg_next_yreg_thr3[21] , div_yreg_next_yreg_thr3[20] ,
         div_yreg_next_yreg_thr3[19] , div_yreg_next_yreg_thr3[18] ,
         div_yreg_next_yreg_thr3[17] , div_yreg_next_yreg_thr3[16] ,
         div_yreg_next_yreg_thr3[15] , div_yreg_next_yreg_thr3[14] ,
         div_yreg_next_yreg_thr3[13] , div_yreg_next_yreg_thr3[12] ,
         div_yreg_next_yreg_thr3[11] , div_yreg_next_yreg_thr3[10] ,
         div_yreg_next_yreg_thr3[9] , div_yreg_next_yreg_thr3[8] ,
         div_yreg_next_yreg_thr3[7] , div_yreg_next_yreg_thr3[6] ,
         div_yreg_next_yreg_thr3[5] , div_yreg_next_yreg_thr3[4] ,
         div_yreg_next_yreg_thr3[3] , div_yreg_next_yreg_thr3[2] ,
         div_yreg_next_yreg_thr3[1] , div_yreg_next_yreg_thr3[0] ,
         div_yreg_next_yreg_thr2[31] , div_yreg_next_yreg_thr2[30] ,
         div_yreg_next_yreg_thr2[29] , div_yreg_next_yreg_thr2[28] ,
         div_yreg_next_yreg_thr2[27] , div_yreg_next_yreg_thr2[26] ,
         div_yreg_next_yreg_thr2[25] , div_yreg_next_yreg_thr2[24] ,
         div_yreg_next_yreg_thr2[23] , div_yreg_next_yreg_thr2[22] ,
         div_yreg_next_yreg_thr2[21] , div_yreg_next_yreg_thr2[20] ,
         div_yreg_next_yreg_thr2[19] , div_yreg_next_yreg_thr2[18] ,
         div_yreg_next_yreg_thr2[17] , div_yreg_next_yreg_thr2[16] ,
         div_yreg_next_yreg_thr2[15] , div_yreg_next_yreg_thr2[14] ,
         div_yreg_next_yreg_thr2[13] , div_yreg_next_yreg_thr2[12] ,
         div_yreg_next_yreg_thr2[11] , div_yreg_next_yreg_thr2[10] ,
         div_yreg_next_yreg_thr2[9] , div_yreg_next_yreg_thr2[8] ,
         div_yreg_next_yreg_thr2[7] , div_yreg_next_yreg_thr2[6] ,
         div_yreg_next_yreg_thr2[5] , div_yreg_next_yreg_thr2[4] ,
         div_yreg_next_yreg_thr2[3] , div_yreg_next_yreg_thr2[2] ,
         div_yreg_next_yreg_thr2[1] , div_yreg_next_yreg_thr2[0] ,
         div_yreg_next_yreg_thr1[31] , div_yreg_next_yreg_thr1[30] ,
         div_yreg_next_yreg_thr1[29] , div_yreg_next_yreg_thr1[28] ,
         div_yreg_next_yreg_thr1[27] , div_yreg_next_yreg_thr1[26] ,
         div_yreg_next_yreg_thr1[25] , div_yreg_next_yreg_thr1[24] ,
         div_yreg_next_yreg_thr1[23] , div_yreg_next_yreg_thr1[22] ,
         div_yreg_next_yreg_thr1[21] , div_yreg_next_yreg_thr1[20] ,
         div_yreg_next_yreg_thr1[19] , div_yreg_next_yreg_thr1[18] ,
         div_yreg_next_yreg_thr1[17] , div_yreg_next_yreg_thr1[16] ,
         div_yreg_next_yreg_thr1[15] , div_yreg_next_yreg_thr1[14] ,
         div_yreg_next_yreg_thr1[13] , div_yreg_next_yreg_thr1[12] ,
         div_yreg_next_yreg_thr1[11] , div_yreg_next_yreg_thr1[10] ,
         div_yreg_next_yreg_thr1[9] , div_yreg_next_yreg_thr1[8] ,
         div_yreg_next_yreg_thr1[7] , div_yreg_next_yreg_thr1[6] ,
         div_yreg_next_yreg_thr1[5] , div_yreg_next_yreg_thr1[4] ,
         div_yreg_next_yreg_thr1[3] , div_yreg_next_yreg_thr1[2] ,
         div_yreg_next_yreg_thr1[1] , div_yreg_next_yreg_thr1[0] ,
         div_yreg_next_yreg_thr0[31] , div_yreg_next_yreg_thr0[30] ,
         div_yreg_next_yreg_thr0[29] , div_yreg_next_yreg_thr0[28] ,
         div_yreg_next_yreg_thr0[27] , div_yreg_next_yreg_thr0[26] ,
         div_yreg_next_yreg_thr0[25] , div_yreg_next_yreg_thr0[24] ,
         div_yreg_next_yreg_thr0[23] , div_yreg_next_yreg_thr0[22] ,
         div_yreg_next_yreg_thr0[21] , div_yreg_next_yreg_thr0[20] ,
         div_yreg_next_yreg_thr0[19] , div_yreg_next_yreg_thr0[18] ,
         div_yreg_next_yreg_thr0[17] , div_yreg_next_yreg_thr0[16] ,
         div_yreg_next_yreg_thr0[15] , div_yreg_next_yreg_thr0[14] ,
         div_yreg_next_yreg_thr0[13] , div_yreg_next_yreg_thr0[12] ,
         div_yreg_next_yreg_thr0[11] , div_yreg_next_yreg_thr0[10] ,
         div_yreg_next_yreg_thr0[9] , div_yreg_next_yreg_thr0[8] ,
         div_yreg_next_yreg_thr0[7] , div_yreg_next_yreg_thr0[6] ,
         div_yreg_next_yreg_thr0[5] , div_yreg_next_yreg_thr0[4] ,
         div_yreg_next_yreg_thr0[3] , div_yreg_next_yreg_thr0[2] ,
         div_yreg_next_yreg_thr0[1] , div_yreg_next_yreg_thr0[0] ,
         div_yreg_yreg_data_w1[0] , div_yreg_yreg_data_w1[1] ,
         div_yreg_yreg_data_w1[2] , div_yreg_yreg_data_w1[3] ,
         div_yreg_yreg_data_w1[4] , div_yreg_yreg_data_w1[5] ,
         div_yreg_yreg_data_w1[6] , div_yreg_yreg_data_w1[7] ,
         div_yreg_yreg_data_w1[8] , div_yreg_yreg_data_w1[9] ,
         div_yreg_yreg_data_w1[10] , div_yreg_yreg_data_w1[11] ,
         div_yreg_yreg_data_w1[12] , div_yreg_yreg_data_w1[13] ,
         div_yreg_yreg_data_w1[14] , div_yreg_yreg_data_w1[15] ,
         div_yreg_yreg_data_w1[16] , div_yreg_yreg_data_w1[17] ,
         div_yreg_yreg_data_w1[18] , div_yreg_yreg_data_w1[19] ,
         div_yreg_yreg_data_w1[20] , div_yreg_yreg_data_w1[21] ,
         div_yreg_yreg_data_w1[22] , div_yreg_yreg_data_w1[23] ,
         div_yreg_yreg_data_w1[24] , div_yreg_yreg_data_w1[25] ,
         div_yreg_yreg_data_w1[26] , div_yreg_yreg_data_w1[27] ,
         div_yreg_yreg_data_w1[28] , div_yreg_yreg_data_w1[29] ,
         div_yreg_yreg_data_w1[30] , div_yreg_yreg_data_w1[31] ,
         div_yreg_div_ecl_yreg_0[0] , div_yreg_div_ecl_yreg_0[1] ,
         div_yreg_div_ecl_yreg_0[2] , div_yreg_div_ecl_yreg_0[3] ,
         div_yreg_yreg_thr0[1] , div_yreg_yreg_thr0[2] ,
         div_yreg_yreg_thr0[3] , div_yreg_yreg_thr0[4] ,
         div_yreg_yreg_thr0[5] , div_yreg_yreg_thr0[6] ,
         div_yreg_yreg_thr0[7] , div_yreg_yreg_thr0[8] ,
         div_yreg_yreg_thr0[9] , div_yreg_yreg_thr0[10] ,
         div_yreg_yreg_thr0[11] , div_yreg_yreg_thr0[12] ,
         div_yreg_yreg_thr0[13] , div_yreg_yreg_thr0[14] ,
         div_yreg_yreg_thr0[15] , div_yreg_yreg_thr0[16] ,
         div_yreg_yreg_thr0[17] , div_yreg_yreg_thr0[18] ,
         div_yreg_yreg_thr0[19] , div_yreg_yreg_thr0[20] ,
         div_yreg_yreg_thr0[21] , div_yreg_yreg_thr0[22] ,
         div_yreg_yreg_thr0[23] , div_yreg_yreg_thr0[24] ,
         div_yreg_yreg_thr0[25] , div_yreg_yreg_thr0[26] ,
         div_yreg_yreg_thr0[27] , div_yreg_yreg_thr0[28] ,
         div_yreg_yreg_thr0[29] , div_yreg_yreg_thr0[30] ,
         div_yreg_yreg_thr0[31] , div_yreg_yreg_thr1[1] ,
         div_yreg_yreg_thr1[2] , div_yreg_yreg_thr1[3] ,
         div_yreg_yreg_thr1[4] , div_yreg_yreg_thr1[5] ,
         div_yreg_yreg_thr1[6] , div_yreg_yreg_thr1[7] ,
         div_yreg_yreg_thr1[8] , div_yreg_yreg_thr1[9] ,
         div_yreg_yreg_thr1[10] , div_yreg_yreg_thr1[11] ,
         div_yreg_yreg_thr1[12] , div_yreg_yreg_thr1[13] ,
         div_yreg_yreg_thr1[14] , div_yreg_yreg_thr1[15] ,
         div_yreg_yreg_thr1[16] , div_yreg_yreg_thr1[17] ,
         div_yreg_yreg_thr1[18] , div_yreg_yreg_thr1[19] ,
         div_yreg_yreg_thr1[20] , div_yreg_yreg_thr1[21] ,
         div_yreg_yreg_thr1[22] , div_yreg_yreg_thr1[23] ,
         div_yreg_yreg_thr1[24] , div_yreg_yreg_thr1[25] ,
         div_yreg_yreg_thr1[26] , div_yreg_yreg_thr1[27] ,
         div_yreg_yreg_thr1[28] , div_yreg_yreg_thr1[29] ,
         div_yreg_yreg_thr1[30] , div_yreg_yreg_thr1[31] ,
         div_yreg_yreg_thr2[1] , div_yreg_yreg_thr2[2] ,
         div_yreg_yreg_thr2[3] , div_yreg_yreg_thr2[4] ,
         div_yreg_yreg_thr2[5] , div_yreg_yreg_thr2[6] ,
         div_yreg_yreg_thr2[7] , div_yreg_yreg_thr2[8] ,
         div_yreg_yreg_thr2[9] , div_yreg_yreg_thr2[10] ,
         div_yreg_yreg_thr2[11] , div_yreg_yreg_thr2[12] ,
         div_yreg_yreg_thr2[13] , div_yreg_yreg_thr2[14] ,
         div_yreg_yreg_thr2[15] , div_yreg_yreg_thr2[16] ,
         div_yreg_yreg_thr2[17] , div_yreg_yreg_thr2[18] ,
         div_yreg_yreg_thr2[19] , div_yreg_yreg_thr2[20] ,
         div_yreg_yreg_thr2[21] , div_yreg_yreg_thr2[22] ,
         div_yreg_yreg_thr2[23] , div_yreg_yreg_thr2[24] ,
         div_yreg_yreg_thr2[25] , div_yreg_yreg_thr2[26] ,
         div_yreg_yreg_thr2[27] , div_yreg_yreg_thr2[28] ,
         div_yreg_yreg_thr2[29] , div_yreg_yreg_thr2[30] ,
         div_yreg_yreg_thr2[31] , div_yreg_yreg_thr3[1] ,
         div_yreg_yreg_thr3[2] , div_yreg_yreg_thr3[3] ,
         div_yreg_yreg_thr3[4] , div_yreg_yreg_thr3[5] ,
         div_yreg_yreg_thr3[6] , div_yreg_yreg_thr3[7] ,
         div_yreg_yreg_thr3[8] , div_yreg_yreg_thr3[9] ,
         div_yreg_yreg_thr3[10] , div_yreg_yreg_thr3[11] ,
         div_yreg_yreg_thr3[12] , div_yreg_yreg_thr3[13] ,
         div_yreg_yreg_thr3[14] , div_yreg_yreg_thr3[15] ,
         div_yreg_yreg_thr3[16] , div_yreg_yreg_thr3[17] ,
         div_yreg_yreg_thr3[18] , div_yreg_yreg_thr3[19] ,
         div_yreg_yreg_thr3[20] , div_yreg_yreg_thr3[21] ,
         div_yreg_yreg_thr3[22] , div_yreg_yreg_thr3[23] ,
         div_yreg_yreg_thr3[24] , div_yreg_yreg_thr3[25] ,
         div_yreg_yreg_thr3[26] , div_yreg_yreg_thr3[27] ,
         div_yreg_yreg_thr3[28] , div_yreg_yreg_thr3[29] ,
         div_yreg_yreg_thr3[30] , div_yreg_yreg_thr3[31] ,
         rml_wtype_mux_n12 , rml_wtype_mux_n11 , rml_wtype_mux_n10 ,
         rml_wtype_mux_n9 , rml_wtype_mux_n8 , rml_wtype_mux_n7 ,
         rml_wtype_mux_n5 , rml_wtype_mux_n4 , rml_wtype_mux_n3 ,
         rml_cwp_inc_n6 , rml_cwp_inc_n5 , rml_cwp_inc_n4 ,
         rml_cwp_inc_n3 , rml_cwp_inc_n2 , rml_next_cwp_mux_n12 ,
         rml_next_cwp_mux_n11 , rml_next_cwp_mux_n10 , rml_next_cwp_mux_n9 ,
         rml_next_cwp_mux_n8 , rml_next_cwp_mux_n7 , rml_next_cwp_mux_n6 ,
         rml_next_cwp_mux_n5 , rml_next_cwp_mux_n4 , rml_next_cwp_mux_n3 ,
         rml_next_cwp_mux_n2 , rml_next_cwp_mux_n1 , rml_oddwin_dff_n9 ,
         rml_oddwin_dff_n7 , rml_oddwin_dff_n5 , rml_oddwin_dff_n3 ,
         rml_oddwin_dff_n1 , rml_cwp_n104 , rml_cwp_n103 , rml_cwp_n102 ,
         rml_cwp_n101 , rml_cwp_n100 , rml_cwp_n99 , rml_cwp_n98 ,
         rml_cwp_n97 , rml_cwp_n96 , rml_cwp_n95 , rml_cwp_n94 ,
         rml_cwp_n93 , rml_cwp_n92 , rml_cwp_n91 , rml_cwp_n90 ,
         rml_cwp_n89 , rml_cwp_n88 , rml_cwp_n87 , rml_cwp_n86 ,
         rml_cwp_n85 , rml_cwp_n84 , rml_cwp_n83 , rml_cwp_n82 ,
         rml_cwp_n81 , rml_cwp_n80 , rml_cwp_n79 , rml_cwp_n78 ,
         rml_cwp_n77 , rml_cwp_n76 , rml_cwp_n75 , rml_cwp_n74 ,
         rml_cwp_n73 , rml_cwp_n72 , rml_cwp_n71 , rml_cwp_n70 ,
         rml_cwp_n69 , rml_cwp_n68 , rml_cwp_n67 , rml_cwp_n66 ,
         rml_cwp_n65 , rml_cwp_n64 , rml_cwp_n63 , rml_cwp_n62 ,
         rml_cwp_n61 , rml_cwp_n60 , rml_cwp_n59 , rml_cwp_n58 ,
         rml_cwp_n57 , rml_cwp_n56 , rml_cwp_n55 , rml_cwp_n54 ,
         rml_cwp_n53 , rml_cwp_n52 , rml_cwp_n51 , rml_cwp_n50 ,
         rml_cwp_n49 , rml_cwp_n48 , rml_cwp_n47 , rml_cwp_n46 ,
         rml_cwp_n45 , rml_cwp_n44 , rml_cwp_n43 , rml_cwp_n42 ,
         rml_cwp_n41 , rml_cwp_n40 , rml_cwp_n39 , rml_cwp_n38 ,
         rml_cwp_n37 , rml_cwp_n36 , rml_cwp_n35 , rml_cwp_n34 ,
         rml_cwp_n33 , rml_cwp_n32 , rml_cwp_n31 , rml_cwp_n30 ,
         rml_cwp_n29 , rml_cwp_n28 , rml_cwp_n27 , rml_cwp_n26 ,
         rml_cwp_n25 , rml_cwp_N99 , rml_cwp_cwp_fastcmplt_w ,
         rml_cwp_cwp_fastcmplt_m , rml_cwp_cwp_cmplt_next ,
         rml_cwp_swap_done_next_cycle[3] , rml_cwp_swap_done_next_cycle[2] ,
         rml_cwp_swap_done_next_cycle[1] , rml_cwp_swap_done_next_cycle[0] ,
         rml_cwp_spill_wtype_next[2] , rml_cwp_spill_wtype_next[1] ,
         rml_cwp_spill_wtype_next[0] , rml_cwp_just_swapped ,
         rml_cwp_swapping , rml_cwp_swap_state[1] , rml_cwp_swap_state[0] ,
         rml_cwp_swap_sel[3] , rml_cwp_swap_sel[2] , rml_cwp_swap_sel[1] ,
         rml_cwp_swap_sel[0] , rml_cwp_next_swap_thr[3] ,
         rml_cwp_next_swap_thr[2] , rml_cwp_next_swap_thr[1] ,
         rml_cwp_next_swap_thr[0] , rml_cwp_swap_req_vec[3] ,
         rml_cwp_swap_req_vec[2] , rml_cwp_swap_req_vec[1] ,
         rml_cwp_swap_req_vec[0] , rml_cwp_swap_slot3_state[1] ,
         rml_cwp_swap_slot2_state[1] , rml_cwp_swap_slot1_state[1] ,
         rml_cwp_swap_slot0_state[1] , rml_cwp_swap_slot3_state_valid[0] ,
         rml_cwp_swap_slot3_state_valid[1] , rml_cwp_next_slot3_state[1] ,
         rml_cwp_next_slot3_state[0] , rml_cwp_swap_slot2_state_valid[0] ,
         rml_cwp_swap_slot2_state_valid[1] , rml_cwp_next_slot2_state[1] ,
         rml_cwp_next_slot2_state[0] , rml_cwp_swap_slot1_state_valid[0] ,
         rml_cwp_swap_slot1_state_valid[1] , rml_cwp_next_slot1_state[1] ,
         rml_cwp_next_slot1_state[0] , rml_cwp_swap_slot0_state_valid[0] ,
         rml_cwp_swap_slot0_state_valid[1] , rml_cwp_next_slot0_state[1] ,
         rml_cwp_next_slot0_state[0] , rml_cwp_swap_slot3_data[0] ,
         rml_cwp_swap_slot3_data[1] , rml_cwp_swap_slot3_data[2] ,
         rml_cwp_swap_slot3_data[3] , rml_cwp_swap_slot3_data[4] ,
         rml_cwp_swap_slot3_data[5] , rml_cwp_swap_slot3_data[6] ,
         rml_cwp_swap_slot3_data[7] , rml_cwp_swap_slot3_data[8] ,
         rml_cwp_swap_slot3_data[9] , rml_cwp_swap_slot3_data[10] ,
         rml_cwp_swap_slot3_data[11] , rml_cwp_swap_slot3_data[12] ,
         rml_cwp_next_slot3_data[12] , rml_cwp_next_slot3_data[11] ,
         rml_cwp_next_slot3_data[10] , rml_cwp_next_slot3_data[9] ,
         rml_cwp_next_slot3_data[8] , rml_cwp_next_slot3_data[7] ,
         rml_cwp_next_slot3_data[6] , rml_cwp_next_slot3_data[5] ,
         rml_cwp_next_slot3_data[4] , rml_cwp_next_slot3_data[3] ,
         rml_cwp_next_slot3_data[2] , rml_cwp_next_slot3_data[1] ,
         rml_cwp_next_slot3_data[0] , rml_cwp_swap_slot2_data[0] ,
         rml_cwp_swap_slot2_data[1] , rml_cwp_swap_slot2_data[2] ,
         rml_cwp_swap_slot2_data[3] , rml_cwp_swap_slot2_data[4] ,
         rml_cwp_swap_slot2_data[5] , rml_cwp_swap_slot2_data[6] ,
         rml_cwp_swap_slot2_data[7] , rml_cwp_swap_slot2_data[8] ,
         rml_cwp_swap_slot2_data[9] , rml_cwp_swap_slot2_data[10] ,
         rml_cwp_swap_slot2_data[11] , rml_cwp_swap_slot2_data[12] ,
         rml_cwp_next_slot2_data[12] , rml_cwp_next_slot2_data[11] ,
         rml_cwp_next_slot2_data[10] , rml_cwp_next_slot2_data[9] ,
         rml_cwp_next_slot2_data[8] , rml_cwp_next_slot2_data[7] ,
         rml_cwp_next_slot2_data[6] , rml_cwp_next_slot2_data[5] ,
         rml_cwp_next_slot2_data[4] , rml_cwp_next_slot2_data[3] ,
         rml_cwp_next_slot2_data[2] , rml_cwp_next_slot2_data[1] ,
         rml_cwp_next_slot2_data[0] , rml_cwp_swap_slot1_data[0] ,
         rml_cwp_swap_slot1_data[1] , rml_cwp_swap_slot1_data[2] ,
         rml_cwp_swap_slot1_data[3] , rml_cwp_swap_slot1_data[4] ,
         rml_cwp_swap_slot1_data[5] , rml_cwp_swap_slot1_data[6] ,
         rml_cwp_swap_slot1_data[7] , rml_cwp_swap_slot1_data[8] ,
         rml_cwp_swap_slot1_data[9] , rml_cwp_swap_slot1_data[10] ,
         rml_cwp_swap_slot1_data[11] , rml_cwp_swap_slot1_data[12] ,
         rml_cwp_next_slot1_data[12] , rml_cwp_next_slot1_data[11] ,
         rml_cwp_next_slot1_data[10] , rml_cwp_next_slot1_data[9] ,
         rml_cwp_next_slot1_data[8] , rml_cwp_next_slot1_data[7] ,
         rml_cwp_next_slot1_data[6] , rml_cwp_next_slot1_data[5] ,
         rml_cwp_next_slot1_data[4] , rml_cwp_next_slot1_data[3] ,
         rml_cwp_next_slot1_data[2] , rml_cwp_next_slot1_data[1] ,
         rml_cwp_next_slot1_data[0] , rml_cwp_swap_slot0_data[0] ,
         rml_cwp_swap_slot0_data[1] , rml_cwp_swap_slot0_data[2] ,
         rml_cwp_swap_slot0_data[3] , rml_cwp_swap_slot0_data[4] ,
         rml_cwp_swap_slot0_data[5] , rml_cwp_swap_slot0_data[6] ,
         rml_cwp_swap_slot0_data[7] , rml_cwp_swap_slot0_data[8] ,
         rml_cwp_swap_slot0_data[9] , rml_cwp_swap_slot0_data[10] ,
         rml_cwp_swap_slot0_data[11] , rml_cwp_swap_slot0_data[12] ,
         rml_cwp_next_slot0_data[12] , rml_cwp_next_slot0_data[11] ,
         rml_cwp_next_slot0_data[10] , rml_cwp_next_slot0_data[9] ,
         rml_cwp_next_slot0_data[8] , rml_cwp_next_slot0_data[7] ,
         rml_cwp_next_slot0_data[6] , rml_cwp_next_slot0_data[5] ,
         rml_cwp_next_slot0_data[4] , rml_cwp_next_slot0_data[3] ,
         rml_cwp_next_slot0_data[2] , rml_cwp_next_slot0_data[1] ,
         rml_cwp_next_slot0_data[0] , rml_cwp_swap_next_state[3] ,
         rml_cwp_swap_next_state[2] , rml_cwp_swap_next_state[1] ,
         rml_cwp_swap_next_state[0] , rml_cwp_swap_keep_state[3] ,
         rml_cwp_swap_keep_state[2] , rml_cwp_swap_keep_state[1] ,
         rml_cwp_swap_keep_state[0] , rml_cwp_swap_sel_tlu[0] ,
         rml_cwp_cwpccr_update_w , rml_cwp_tlu_swap_data[12] ,
         rml_cwp_full_swap_w , rml_cwp_full_swap_m ,
         rml_cwp_tlu_exu_cwp_w[0] , rml_cwp_tlu_exu_cwp_w[1] ,
         rml_cwp_tlu_exu_cwp_w[2] , rml_cwp_cwp_thr0_next[2] ,
         rml_cwp_cwp_thr0_next[1] , rml_cwp_cwp_thr1_next[2] ,
         rml_cwp_cwp_thr1_next[1] , rml_cwp_cwp_thr2_next[2] ,
         rml_cwp_cwp_thr2_next[1] , rml_cwp_cwp_thr3_next[2] ,
         rml_cwp_cwp_thr3_next[1] , rml_cwp_cwp_wen_tlu_w[3] ,
         rml_cwp_cwp_wen_tlu_w[2] , rml_cwp_cwp_wen_tlu_w[1] ,
         rml_cwp_cwp_wen_tlu_w[0] , rml_cwp_valid_tlu_swap_w ,
         rml_cwp_spill_next , rml_cwp_swap_thr[0] , rml_cwp_swap_thr[1] ,
         rml_cwp_swap_thr[2] , rml_cwp_swap_thr[3] ,
         rml_cwp_trap_old_cwp_m[2] , rml_cwp_trap_old_cwp_m[1] ,
         rml_cwp_trap_old_cwp_m[0] , rml_cwp_old_cwp_w[0] ,
         rml_cwp_old_cwp_w[1] , rml_cwp_old_cwp_w[2] ,
         rml_cwp_new_swap_cwp[0] , rml_cwp_new_swap_cwp[1] ,
         rml_cwp_new_swap_cwp[2] , rml_cwp_swap_data[6] ,
         rml_cwp_swap_data[7] , rml_cwp_swap_data[8] ,
         rml_cwp_swap_data_12 , rml_cwp_old_swap_cwp[2] ,
         rml_cwp_old_swap_cwp[1] , rml_cwp_old_swap_cwp[0] ,
         rml_cwp_swap_tid[0] , rml_cwp_swap_tid[1] , rml_cwp_thr_e[0] ,
         rml_cwp_thr_e[2] , rml_cwp_thr_e[3] , rml_next_cansave_mux_n7 ,
         rml_next_cansave_mux_n6 , rml_next_cansave_mux_n5 ,
         rml_next_cansave_mux_n4 , rml_next_cansave_mux_n3 ,
         rml_next_cansave_mux_n2 , rml_cansave_reg_n8 , rml_cansave_reg_n7 ,
         rml_cansave_reg_n6 , rml_cansave_reg_n5 ,
         rml_cansave_reg_data_thr3_next[2] ,
         rml_cansave_reg_data_thr3_next[1] ,
         rml_cansave_reg_data_thr3_next[0] ,
         rml_cansave_reg_data_thr2_next[2] ,
         rml_cansave_reg_data_thr2_next[1] ,
         rml_cansave_reg_data_thr2_next[0] ,
         rml_cansave_reg_data_thr1_next[2] ,
         rml_cansave_reg_data_thr1_next[1] ,
         rml_cansave_reg_data_thr1_next[0] ,
         rml_cansave_reg_data_thr0_next[2] ,
         rml_cansave_reg_data_thr0_next[1] ,
         rml_cansave_reg_data_thr0_next[0] , rml_cansave_reg_data_thr3[0] ,
         rml_cansave_reg_data_thr3[1] , rml_cansave_reg_data_thr3[2] ,
         rml_cansave_reg_data_thr2[0] , rml_cansave_reg_data_thr2[1] ,
         rml_cansave_reg_data_thr2[2] , rml_cansave_reg_data_thr1[0] ,
         rml_cansave_reg_data_thr1[1] , rml_cansave_reg_data_thr1[2] ,
         rml_cansave_reg_data_thr0[0] , rml_cansave_reg_data_thr0[1] ,
         rml_cansave_reg_data_thr0[2] , rml_mux_agp_out1_n12 ,
         rml_mux_agp_out1_n11 , rml_mux_agp_out1_n10 , rml_mux_agp_out1_n9 ,
         rml_mux_agp_out1_n8 , rml_mux_agp_out1_n7 , rml_mux_agp_out1_n6 ,
         rml_mux_agp_out1_n5 , rml_mux_agp_out1_n4 , rml_mux_agp_out1_n3 ,
         rml_mux_agp_out1_n2 , rml_mux_agp_out1_n1 , rml_agp_next0_mux_n5 ,
         rml_agp_next0_mux_n4 , rml_agp_next0_mux_n3 ,
         rml_agp_next0_mux_n2 , ecl_ccr_mux_ccr_m_n17 ,
         ecl_ccr_mux_ccr_m_n16 , ecl_ccr_mux_ccr_m_n15 ,
         ecl_ccr_mux_ccr_m_n14 , ecl_ccr_mux_ccr_m_n13 ,
         ecl_ccr_mux_ccr_m_n12 , ecl_ccr_mux_ccr_m_n11 ,
         ecl_ccr_mux_ccr_m_n10 , ecl_ccr_mux_ccr_m_n9 ,
         ecl_ccr_mux_ccr_m_n8 , ecl_ccr_mux_ccr_m_n7 ,
         ecl_ccr_mux_ccr_m_n6 , ecl_ccr_mux_ccr_m_n5 ,
         ecl_ccr_mux_ccr_m_n4 , ecl_ccr_mux_ccr_m_n3 ,
         ecl_ccr_mux_ccr_m_n2 , ecl_ccr_mux_ccrin0_n32 ,
         ecl_ccr_mux_ccrin0_n31 , ecl_ccr_mux_ccrin0_n30 ,
         ecl_ccr_mux_ccrin0_n29 , ecl_ccr_mux_ccrin0_n28 ,
         ecl_ccr_mux_ccrin0_n27 , ecl_ccr_mux_ccrin0_n26 ,
         ecl_ccr_mux_ccrin0_n25 , ecl_ccr_mux_ccrin0_n24 ,
         ecl_ccr_mux_ccrin0_n23 , ecl_ccr_mux_ccrin0_n22 ,
         ecl_ccr_mux_ccrin0_n21 , ecl_ccr_mux_ccrin0_n20 ,
         ecl_ccr_mux_ccrin0_n19 , ecl_ccr_mux_ccrin0_n18 ,
         ecl_ccr_mux_ccrin0_n17 , ecl_ccr_mux_ccrin0_n16 ,
         ecl_ccr_mux_ccrin0_n14 , ecl_ccr_mux_ccrin0_n12 ,
         ecl_ccr_mux_ccrin0_n10 , ecl_ccr_mux_ccrin0_n8 ,
         ecl_ccr_mux_ccrin0_n7 , ecl_ccr_mux_ccrin0_n6 ,
         ecl_ccr_mux_ccrin0_n5 , ecl_ccr_mux_ccrin0_n4 ,
         ecl_ccr_mux_ccrin0_n3 , ecl_ccr_mux_ccrin0_n2 ,
         ecl_ccr_mux_ccrin0_n1 , ecl_ccr_mux_ccrin0_sel2 ,
         ecl_ccr_mux_ccr_out_n48 , ecl_ccr_mux_ccr_out_n47 ,
         ecl_ccr_mux_ccr_out_n46 , ecl_ccr_mux_ccr_out_n45 ,
         ecl_ccr_mux_ccr_out_n44 , ecl_ccr_mux_ccr_out_n43 ,
         ecl_ccr_mux_ccr_out_n42 , ecl_ccr_mux_ccr_out_n41 ,
         ecl_ccr_mux_ccr_out_n40 , ecl_ccr_mux_ccr_out_n39 ,
         ecl_ccr_mux_ccr_out_n38 , ecl_ccr_mux_ccr_out_n37 ,
         ecl_ccr_mux_ccr_out_n36 , ecl_ccr_mux_ccr_out_n35 ,
         ecl_ccr_mux_ccr_out_n34 , ecl_ccr_mux_ccr_out_n33 ,
         ecl_ccr_mux_ccr_out_n32 , ecl_ccr_mux_ccr_out_n31 ,
         ecl_ccr_mux_ccr_out_n30 , ecl_ccr_mux_ccr_out_n29 ,
         ecl_ccr_mux_ccr_out_n28 , ecl_ccr_mux_ccr_out_n27 ,
         ecl_ccr_mux_ccr_out_n26 , ecl_ccr_mux_ccr_out_n25 ,
         ecl_ccr_mux_ccr_out_n24 , ecl_ccr_mux_ccr_out_n23 ,
         ecl_ccr_mux_ccr_out_n22 , ecl_ccr_mux_ccr_out_n21 ,
         ecl_ccr_mux_ccr_out_n20 , ecl_ccr_mux_ccr_out_n19 ,
         ecl_ccr_mux_ccr_out_n18 , ecl_ccr_mux_ccr_out_n17 ,
         ecl_ccr_mux_ccr_out_n16 , ecl_ccr_mux_ccr_out_n15 ,
         ecl_ccr_mux_ccr_out_n14 , ecl_ccr_mux_ccr_out_n13 ,
         ecl_ccr_mux_ccr_out_n12 , ecl_ccr_mux_ccr_out_n11 ,
         ecl_ccr_mux_ccr_out_n10 , ecl_ccr_mux_ccr_out_n9 ,
         ecl_ccr_mux_ccr_out_n8 , ecl_ccr_mux_ccr_out_n7 ,
         ecl_ccr_mux_ccr_out_n6 , ecl_ccr_mux_ccr_out_n5 ,
         ecl_ccr_mux_ccr_out_n4 , ecl_ccr_mux_ccr_out_n3 ,
         ecl_ccr_mux_ccr_out_n2 , ecl_ccr_mux_ccr_out_n1 ,
         ecl_writeback_rd_g_mux_n30 , ecl_writeback_rd_g_mux_n29 ,
         ecl_writeback_rd_g_mux_n28 , ecl_writeback_rd_g_mux_n27 ,
         ecl_writeback_rd_g_mux_n26 , ecl_writeback_rd_g_mux_n25 ,
         ecl_writeback_rd_g_mux_n24 , ecl_writeback_rd_g_mux_n23 ,
         ecl_writeback_rd_g_mux_n22 , ecl_writeback_rd_g_mux_n21 ,
         ecl_writeback_rd_g_mux_n20 , ecl_writeback_rd_g_mux_n19 ,
         ecl_writeback_rd_g_mux_n18 , ecl_writeback_rd_g_mux_n17 ,
         ecl_writeback_rd_g_mux_n16 , ecl_writeback_rd_g_mux_n15 ,
         ecl_writeback_rd_g_mux_n14 , ecl_writeback_rd_g_mux_n13 ,
         ecl_writeback_rd_g_mux_n12 , ecl_writeback_rd_g_mux_n11 ,
         ecl_writeback_rd_g_mux_n10 , ecl_writeback_rd_g_mux_n9 ,
         ecl_writeback_rd_g_mux_n8 , ecl_writeback_rd_g_mux_n7 ,
         ecl_writeback_rd_g_mux_n6 , ecl_writeback_rd_g_mux_n5 ,
         ecl_writeback_rd_g_mux_n4 , ecl_writeback_rd_g_mux_n3 ,
         ecl_writeback_rd_g_mux_n2 , ecl_writeback_rd_g_mux_n1 ,
         ecl_writeback_setcc_g_mux_n3 , ecl_writeback_setcc_g_mux_n2 ,
         ecl_writeback_dff_wb_m2w_n2 , ecl_writeback_rdpr_mux1_n18 ,
         ecl_writeback_rdpr_mux1_n17 , ecl_writeback_rdpr_mux1_n16 ,
         ecl_writeback_rdpr_mux1_n15 , ecl_writeback_rdpr_mux1_n14 ,
         ecl_writeback_rdpr_mux1_n13 , ecl_writeback_rdpr_mux1_n12 ,
         ecl_writeback_rdpr_mux1_n11 , ecl_writeback_rdpr_mux1_n10 ,
         ecl_writeback_rdpr_mux1_n9 , ecl_writeback_rdpr_mux1_n8 ,
         ecl_writeback_rdpr_mux1_n7 , ecl_writeback_rdpr_mux1_n6 ,
         ecl_writeback_rdpr_mux1_n5 , ecl_writeback_rdpr_mux1_n4 ,
         ecl_writeback_rdpr_mux1_n3 , ecl_writeback_rdpr_mux1_n2 ,
         ecl_writeback_rdpr_mux1_n1 , ecl_writeback_restore_tid_dff_n15 ,
         ecl_writeback_restore_tid_dff_n14 ,
         ecl_writeback_restore_tid_dff_n13 ,
         ecl_writeback_restore_tid_dff_n10 ,
         ecl_writeback_restore_tid_dff_n9 ,
         ecl_writeback_restore_tid_dff_n8 ,
         ecl_writeback_restore_tid_dff_n6 ,
         ecl_writeback_restore_tid_dff_n4 ,
         ecl_writeback_restore_tid_dff_n3 ,
         ecl_writeback_restore_tid_dff_n2 ,
         ecl_writeback_restore_rd_dff_n27 ,
         ecl_writeback_restore_rd_dff_n26 ,
         ecl_writeback_restore_rd_dff_n25 ,
         ecl_writeback_restore_rd_dff_n24 ,
         ecl_writeback_restore_rd_dff_n23 ,
         ecl_writeback_restore_rd_dff_n22 ,
         ecl_writeback_restore_rd_dff_n20 ,
         ecl_writeback_restore_rd_dff_n18 ,
         ecl_writeback_restore_rd_dff_n16 ,
         ecl_writeback_restore_rd_dff_n14 ,
         ecl_writeback_restore_rd_dff_n12 ,
         ecl_writeback_restore_rd_dff_n10 , ecl_writeback_restore_rd_dff_n8 ,
         ecl_writeback_restore_rd_dff_n6 , ecl_writeback_restore_rd_dff_n5 ,
         ecl_writeback_restore_rd_dff_n3 , ecl_writeback_restore_rd_dff_n2 ,
         ecl_eccctl_ecc_rd_mux_n20 , ecl_eccctl_ecc_rd_mux_n19 ,
         ecl_eccctl_ecc_rd_mux_n18 , ecl_eccctl_ecc_rd_mux_n17 ,
         ecl_eccctl_ecc_rd_mux_n16 , ecl_eccctl_ecc_rd_mux_n15 ,
         ecl_eccctl_ecc_rd_mux_n14 , ecl_eccctl_ecc_rd_mux_n13 ,
         ecl_eccctl_ecc_rd_mux_n12 , ecl_eccctl_ecc_rd_mux_n11 ,
         ecl_eccctl_ecc_rd_mux_n10 , ecl_eccctl_ecc_rd_mux_n9 ,
         ecl_eccctl_ecc_rd_mux_n8 , ecl_eccctl_ecc_rd_mux_n7 ,
         ecl_eccctl_ecc_rd_mux_n6 , ecl_eccctl_ecc_rd_mux_n5 ,
         ecl_eccctl_ecc_rd_mux_n4 , ecl_eccctl_ecc_rd_mux_n3 ,
         ecl_eccctl_ecc_rd_mux_n2 , ecl_eccctl_ecc_rd_mux_n1 ,
         ecl_eccctl_ecc_synd7_mux_n4 , ecl_eccctl_ecc_synd7_mux_n3 ,
         ecl_eccctl_ecc_synd7_mux_n2 , ecl_eccctl_ecc_synd7_mux_n1 ,
         ecl_byplog_rs1_w_comp7_n12 , ecl_byplog_rs1_w_comp7_n11 ,
         ecl_byplog_rs1_w_comp7_n10 , ecl_byplog_rs1_w_comp7_n9 ,
         ecl_byplog_rs1_w_comp7_n8 , ecl_byplog_rs1_w_comp7_n7 ,
         ecl_byplog_rs1_w_comp7_n6 , ecl_byplog_rs1_w_comp7_n5 ,
         ecl_byplog_rs1_w_comp7_n4 , ecl_byplog_rs1_w_comp7_n3 ,
         ecl_byplog_rs1_w_comp7_n2 , ecl_byplog_rs1_w_comp7_n1 ,
         ecl_divcntl_divstate_dff_n13 , ecl_divcntl_divstate_dff_n11 ,
         ecl_divcntl_divstate_dff_n9 , ecl_divcntl_divstate_dff_n7 ,
         ecl_divcntl_divstate_dff_n5 , ecl_divcntl_divstate_dff_n3 ,
         ecl_divcntl_divstate_dff_n1 , ecl_divcntl_cnt6_n32 ,
         ecl_divcntl_cnt6_n31 , ecl_divcntl_cnt6_n30 ,
         ecl_divcntl_cnt6_n29 , ecl_divcntl_cnt6_n28 ,
         ecl_divcntl_cnt6_n27 , ecl_divcntl_cnt6_n26 ,
         ecl_divcntl_cnt6_n25 , ecl_divcntl_cnt6_n24 ,
         ecl_divcntl_cnt6_n23 , ecl_divcntl_cnt6_n22 ,
         ecl_divcntl_cnt6_n21 , ecl_divcntl_cnt6_n20 ,
         ecl_divcntl_cnt6_n19 , ecl_divcntl_cnt6_n18 ,
         ecl_divcntl_cnt6_n17 , ecl_divcntl_cnt6_n16 ,
         ecl_divcntl_cnt6_n15 , ecl_divcntl_cnt6_n14 ,
         ecl_divcntl_cnt6_n12 , ecl_divcntl_cnt6_n11 ,
         ecl_divcntl_cnt6_n10 , ecl_divcntl_cnt6_n9 ,
         ecl_divcntl_cnt6_next_cntr[5] , ecl_divcntl_cnt6_next_cntr[4] ,
         ecl_divcntl_cnt6_next_cntr[3] , ecl_divcntl_cnt6_next_cntr[2] ,
         ecl_divcntl_cnt6_next_cntr[1] , ecl_divcntl_qnext_cout_mux_n3 ,
         ecl_divcntl_qnext_cout_mux_n2 , ecl_divcntl_inputs_neg_dff_n9 ,
         ecl_divcntl_inputs_neg_dff_n8 , ecl_divcntl_inputs_neg_dff_n6 ,
         ecl_divcntl_inputs_neg_dff_n4 , ecl_divcntl_inputs_neg_dff_n3 ,
         ecl_mdqctl_div_data_mux_n25 , ecl_mdqctl_div_data_mux_n23 ,
         ecl_mdqctl_div_data_mux_n22 , ecl_mdqctl_div_data_mux_n21 ,
         ecl_mdqctl_div_data_mux_n20 , ecl_mdqctl_div_data_mux_n19 ,
         ecl_mdqctl_div_data_mux_n18 , ecl_mdqctl_div_data_mux_n17 ,
         ecl_mdqctl_div_data_mux_n16 , ecl_mdqctl_div_data_mux_n15 ,
         ecl_mdqctl_div_data_mux_n14 , ecl_mdqctl_div_data_mux_n13 ,
         ecl_mdqctl_div_data_mux_n12 , ecl_mdqctl_div_data_mux_n11 ,
         ecl_mdqctl_div_data_mux_n10 , ecl_mdqctl_div_data_mux_n9 ,
         ecl_mdqctl_div_data_mux_n8 , ecl_mdqctl_div_data_mux_n7 ,
         ecl_mdqctl_div_data_mux_n6 , ecl_mdqctl_div_data_mux_n5 ,
         ecl_mdqctl_div_data_mux_n4 , ecl_mdqctl_div_data_mux_n3 ,
         ecl_mdqctl_div_data_mux_n2 , ecl_mdqctl_div_data_dff_n25 ,
         ecl_mdqctl_div_data_dff_n23 , ecl_mdqctl_div_data_dff_n21 ,
         ecl_mdqctl_div_data_dff_n19 , ecl_mdqctl_div_data_dff_n17 ,
         ecl_mdqctl_div_data_dff_n15 , ecl_mdqctl_div_data_dff_n13 ,
         ecl_mdqctl_div_data_dff_n11 , ecl_mdqctl_div_data_dff_n9 ,
         ecl_mdqctl_div_data_dff_n7 , ecl_mdqctl_div_data_dff_n5 ,
         ecl_mdqctl_div_data_dff_n2 , ecl_mdqctl_mul_data_dff_n21 ,
         ecl_mdqctl_mul_data_dff_n19 , ecl_mdqctl_mul_data_dff_n17 ,
         ecl_mdqctl_mul_data_dff_n15 , ecl_mdqctl_mul_data_dff_n13 ,
         ecl_mdqctl_mul_data_dff_n11 , ecl_mdqctl_mul_data_dff_n9 ,
         ecl_mdqctl_mul_data_dff_n7 , ecl_mdqctl_mul_data_dff_n5 ,
         ecl_mdqctl_mul_data_dff_n3 , ecl_mdqctl_mul_data_dff_n1 ,
         rml_cwp_slot0_data_mux_n52 , rml_cwp_slot0_data_mux_n51 ,
         rml_cwp_slot0_data_mux_n50 , rml_cwp_slot0_data_mux_n49 ,
         rml_cwp_slot0_data_mux_n48 , rml_cwp_slot0_data_mux_n46 ,
         rml_cwp_slot0_data_mux_n44 , rml_cwp_slot0_data_mux_n42 ,
         rml_cwp_slot0_data_mux_n39 , rml_cwp_slot0_data_mux_n38 ,
         rml_cwp_slot0_data_mux_n36 , rml_cwp_slot0_data_mux_n35 ,
         rml_cwp_slot0_data_mux_n34 , rml_cwp_slot0_data_mux_n33 ,
         rml_cwp_slot0_data_mux_n32 , rml_cwp_slot0_data_mux_n31 ,
         rml_cwp_slot0_data_mux_n30 , rml_cwp_slot0_data_mux_n29 ,
         rml_cwp_slot0_data_mux_n28 , rml_cwp_slot0_data_mux_n27 ,
         rml_cwp_slot0_data_mux_n26 , rml_cwp_slot0_data_mux_n25 ,
         rml_cwp_slot0_data_mux_n24 , rml_cwp_slot0_data_mux_n23 ,
         rml_cwp_slot0_data_mux_n22 , rml_cwp_slot0_data_mux_n21 ,
         rml_cwp_slot0_data_mux_n20 , rml_cwp_slot0_data_mux_n19 ,
         rml_cwp_slot0_data_mux_n18 , rml_cwp_slot0_data_mux_n17 ,
         rml_cwp_slot0_data_mux_n16 , rml_cwp_slot0_data_mux_n14 ,
         rml_cwp_slot0_data_mux_n10 , rml_cwp_slot0_data_mux_n8 ,
         rml_cwp_slot0_data_mux_n6 , rml_cwp_slot0_data_mux_n4 ,
         rml_cwp_slot0_data_mux_n2 , rml_cwp_slot0_data_mux_sel2 ,
         rml_cwp_slot0_data_dff_n31 , rml_cwp_slot0_data_dff_n29 ,
         rml_cwp_slot0_data_dff_n27 , rml_cwp_slot0_data_dff_n25 ,
         rml_cwp_slot0_data_dff_n23 , rml_cwp_slot0_data_dff_n21 ,
         rml_cwp_slot0_data_dff_n19 , rml_cwp_slot0_data_dff_n17 ,
         rml_cwp_slot0_data_dff_n15 , rml_cwp_slot0_data_dff_n13 ,
         rml_cwp_slot0_data_dff_n11 , rml_cwp_slot0_data_dff_n9 ,
         rml_cwp_slot0_data_dff_n7 , rml_cwp_slot0_data_dff_n5 ,
         rml_cwp_slot0_data_dff_n2 , rml_cwp_cwp_output_queue_n38 ,
         rml_cwp_cwp_output_queue_n37 , rml_cwp_cwp_output_queue_n36 ,
         rml_cwp_cwp_output_queue_n35 , rml_cwp_cwp_output_queue_n34 ,
         rml_cwp_cwp_output_queue_n33 , rml_cwp_cwp_output_queue_n32 ,
         rml_cwp_cwp_output_queue_n31 , rml_cwp_cwp_output_queue_n30 ,
         rml_cwp_cwp_output_queue_n29 , rml_cwp_cwp_output_queue_n28 ,
         rml_cwp_cwp_output_queue_n27 , rml_cwp_cwp_output_queue_n26 ,
         rml_cwp_cwp_output_queue_n25 , rml_cwp_cwp_output_queue_n24 ,
         rml_cwp_cwp_output_queue_n23 , rml_cwp_cwp_output_queue_n22 ,
         rml_cwp_cwp_output_queue_n21 , rml_cwp_cwp_output_queue_n20 ,
         rml_cwp_cwp_output_queue_n19 , rml_cwp_cwp_output_queue_n18 ,
         rml_cwp_cwp_output_queue_n17 , rml_cwp_cwp_output_queue_n16 ,
         rml_cwp_cwp_output_queue_n15 , rml_cwp_cwp_output_queue_n14 ,
         rml_cwp_cwp_output_queue_n13 , rml_cwp_cwp_output_queue_n12 ,
         rml_cwp_cwp_output_queue_n11 , rml_cwp_cwp_output_queue_n10 ,
         rml_cwp_cwp_output_queue_pv[0] , rml_cwp_cwp_output_queue_pv[1] ,
         rml_cwp_cwp_output_queue_pv[2] , rml_cwp_cwp_output_queue_pv[3] ,
         rml_cwp_cwp_output_queue_next_pv[3] ,
         rml_cwp_cwp_output_queue_next_pv[2] ,
         rml_cwp_cwp_output_queue_next_pv[1] ,
         rml_cwp_cwp_output_queue_next_pv[0] , rml_cwp_cwp_output_mux_n90 ,
         rml_cwp_cwp_output_mux_n89 , rml_cwp_cwp_output_mux_n88 ,
         rml_cwp_cwp_output_mux_n87 , rml_cwp_cwp_output_mux_n86 ,
         rml_cwp_cwp_output_mux_n85 , rml_cwp_cwp_output_mux_n84 ,
         rml_cwp_cwp_output_mux_n83 , rml_cwp_cwp_output_mux_n82 ,
         rml_cwp_cwp_output_mux_n81 , rml_cwp_cwp_output_mux_n80 ,
         rml_cwp_cwp_output_mux_n79 , rml_cwp_cwp_output_mux_n78 ,
         rml_cwp_cwp_output_mux_n77 , rml_cwp_cwp_output_mux_n76 ,
         rml_cwp_cwp_output_mux_n75 , rml_cwp_cwp_output_mux_n74 ,
         rml_cwp_cwp_output_mux_n73 , rml_cwp_cwp_output_mux_n72 ,
         rml_cwp_cwp_output_mux_n71 , rml_cwp_cwp_output_mux_n70 ,
         rml_cwp_cwp_output_mux_n69 , rml_cwp_cwp_output_mux_n68 ,
         rml_cwp_cwp_output_mux_n67 , rml_cwp_cwp_output_mux_n66 ,
         rml_cwp_cwp_output_mux_n65 , rml_cwp_cwp_output_mux_n64 ,
         rml_cwp_cwp_output_mux_n63 , rml_cwp_cwp_output_mux_n62 ,
         rml_cwp_cwp_output_mux_n61 , rml_cwp_cwp_output_mux_n60 ,
         rml_cwp_cwp_output_mux_n59 , rml_cwp_cwp_output_mux_n58 ,
         rml_cwp_cwp_output_mux_n57 , rml_cwp_cwp_output_mux_n56 ,
         rml_cwp_cwp_output_mux_n55 , rml_cwp_cwp_output_mux_n54 ,
         rml_cwp_cwp_output_mux_n53 , rml_cwp_cwp_output_mux_n52 ,
         rml_cwp_cwp_output_mux_n51 , rml_cwp_cwp_output_mux_n50 ,
         rml_cwp_cwp_output_mux_n49 , rml_cwp_cwp_output_mux_n48 ,
         rml_cwp_cwp_output_mux_n47 , rml_cwp_cwp_output_mux_n46 ,
         rml_cwp_cwp_output_mux_n45 , rml_cwp_cwp_output_mux_n44 ,
         rml_cwp_cwp_output_mux_n43 , rml_cwp_cwp_output_mux_n42 ,
         rml_cwp_cwp_output_mux_n41 , rml_cwp_cwp_output_mux_n40 ,
         rml_cwp_cwp_output_mux_n39 , rml_cwp_cwp_output_mux_n38 ,
         rml_cwp_cwp_output_mux_n37 , rml_cwp_cwp_output_mux_n36 ,
         rml_cwp_cwp_output_mux_n35 , rml_cwp_cwp_output_mux_n34 ,
         rml_cwp_cwp_output_mux_n33 , rml_cwp_cwp_output_mux_n32 ,
         rml_cwp_cwp_output_mux_n31 , rml_cwp_cwp_output_mux_n30 ,
         rml_cwp_cwp_output_mux_n29 , rml_cwp_cwp_output_mux_n28 ,
         rml_cwp_cwp_output_mux_n27 , rml_cwp_cwp_output_mux_n26 ,
         rml_cwp_cwp_output_mux_n25 , rml_cwp_cwp_output_mux_n24 ,
         rml_cwp_cwp_output_mux_n23 , rml_cwp_cwp_output_mux_n22 ,
         rml_cwp_cwp_output_mux_n21 , rml_cwp_cwp_output_mux_n20 ,
         rml_cwp_cwp_output_mux_n19 , rml_cwp_cwp_output_mux_n18 ,
         rml_cwp_cwp_output_mux_n17 , rml_cwp_cwp_output_mux_n16 ,
         rml_cwp_cwp_output_mux_n15 , rml_cwp_cwp_output_mux_n14 ,
         rml_cwp_cwp_output_mux_n13 , rml_cwp_cwp_output_mux_n12 ,
         rml_cwp_cwp_output_mux_n11 , rml_cwp_cwp_output_mux_n10 ,
         rml_cwp_cwp_output_mux_n9 , rml_cwp_cwp_output_mux_n8 ,
         rml_cwp_cwp_output_mux_n7 , rml_cwp_cwp_output_mux_n6 ,
         rml_cwp_cwp_output_mux_n5 , rml_cwp_cwp_output_mux_n4 ,
         rml_cwp_cwp_output_mux_n3 , rml_cwp_cwp_output_mux_n2 ,
         rml_cwp_cwp_output_mux_n1 , bypass_mux_rs3_data_2_in1[0] ,
         bypass_mux_rs3_data_2_in1[1] , bypass_mux_rs3_data_2_in1[2] ,
         bypass_mux_rs3_data_2_in1[3] , bypass_mux_rs3_data_2_in1[4] ,
         bypass_mux_rs3_data_2_in1[5] , bypass_mux_rs3_data_2_in1[6] ,
         bypass_mux_rs3_data_2_in1[7] , bypass_mux_rs3_data_2_in1[8] ,
         bypass_mux_rs3_data_2_in1[9] , bypass_mux_rs3_data_2_in1[10] ,
         bypass_mux_rs3_data_2_in1[11] , bypass_mux_rs3_data_2_in1[12] ,
         bypass_mux_rs3_data_2_in1[13] , bypass_mux_rs3_data_2_in1[14] ,
         bypass_mux_rs3_data_2_in1[15] , bypass_mux_rs3_data_2_in1[16] ,
         bypass_mux_rs3_data_2_in1[17] , bypass_mux_rs3_data_2_in1[18] ,
         bypass_mux_rs3_data_2_in1[19] , bypass_mux_rs3_data_2_in1[20] ,
         bypass_mux_rs3_data_2_in1[21] , bypass_mux_rs3_data_2_in1[22] ,
         bypass_mux_rs3_data_2_in1[23] , bypass_mux_rs3_data_2_in1[24] ,
         bypass_mux_rs3_data_2_in1[25] , bypass_mux_rs3_data_2_in1[26] ,
         bypass_mux_rs3_data_2_in1[27] , bypass_mux_rs3_data_2_in1[28] ,
         bypass_mux_rs3_data_2_in1[29] , bypass_mux_rs3_data_2_in1[30] ,
         bypass_mux_rs3_data_2_in1[31] , bypass_mux_rs3_data_2_in1[32] ,
         bypass_mux_rs3_data_2_in1[33] , bypass_mux_rs3_data_2_in1[34] ,
         bypass_mux_rs3_data_2_in1[35] , bypass_mux_rs3_data_2_in1[36] ,
         bypass_mux_rs3_data_2_in1[37] , bypass_mux_rs3_data_2_in1[38] ,
         bypass_mux_rs3_data_2_in1[39] , bypass_mux_rs3_data_2_in1[40] ,
         bypass_mux_rs3_data_2_in1[41] , bypass_mux_rs3_data_2_in1[42] ,
         bypass_mux_rs3_data_2_in1[43] , bypass_mux_rs3_data_2_in1[44] ,
         bypass_mux_rs3_data_2_in1[45] , bypass_mux_rs3_data_2_in1[46] ,
         bypass_mux_rs3_data_2_in1[47] , bypass_mux_rs3_data_2_in1[48] ,
         bypass_mux_rs3_data_2_in1[49] , bypass_mux_rs3_data_2_in1[50] ,
         bypass_mux_rs3_data_2_in1[51] , bypass_mux_rs3_data_2_in1[52] ,
         bypass_mux_rs3_data_2_in1[53] , bypass_mux_rs3_data_2_in1[54] ,
         bypass_mux_rs3_data_2_in1[55] , bypass_mux_rs3_data_2_in1[56] ,
         bypass_mux_rs3_data_2_in1[57] , bypass_mux_rs3_data_2_in1[58] ,
         bypass_mux_rs3_data_2_in1[59] , bypass_mux_rs3_data_2_in1[60] ,
         bypass_mux_rs3_data_2_in1[61] , bypass_mux_rs3_data_2_in1[62] ,
         bypass_mux_rs3_data_2_in1[63] , bypass_mux_rs2_data_2_in1[0] ,
         bypass_mux_rs2_data_2_in1[1] , bypass_mux_rs2_data_2_in1[2] ,
         bypass_mux_rs2_data_2_in1[3] , bypass_mux_rs2_data_2_in1[4] ,
         bypass_mux_rs2_data_2_in1[5] , bypass_mux_rs2_data_2_in1[6] ,
         bypass_mux_rs2_data_2_in1[7] , bypass_mux_rs2_data_2_in1[8] ,
         bypass_mux_rs2_data_2_in1[9] , bypass_mux_rs2_data_2_in1[10] ,
         bypass_mux_rs2_data_2_in1[11] , bypass_mux_rs2_data_2_in1[12] ,
         bypass_mux_rs2_data_2_in1[13] , bypass_mux_rs2_data_2_in1[14] ,
         bypass_mux_rs2_data_2_in1[15] , bypass_mux_rs2_data_2_in1[16] ,
         bypass_mux_rs2_data_2_in1[17] , bypass_mux_rs2_data_2_in1[18] ,
         bypass_mux_rs2_data_2_in1[19] , bypass_mux_rs2_data_2_in1[20] ,
         bypass_mux_rs2_data_2_in1[21] , bypass_mux_rs2_data_2_in1[22] ,
         bypass_mux_rs2_data_2_in1[23] , bypass_mux_rs2_data_2_in1[24] ,
         bypass_mux_rs2_data_2_in1[25] , bypass_mux_rs2_data_2_in1[26] ,
         bypass_mux_rs2_data_2_in1[27] , bypass_mux_rs2_data_2_in1[28] ,
         bypass_mux_rs2_data_2_in1[29] , bypass_mux_rs2_data_2_in1[30] ,
         bypass_mux_rs2_data_2_in1[31] , bypass_mux_rs2_data_2_in1[32] ,
         bypass_mux_rs2_data_2_in1[33] , bypass_mux_rs2_data_2_in1[34] ,
         bypass_mux_rs2_data_2_in1[35] , bypass_mux_rs2_data_2_in1[36] ,
         bypass_mux_rs2_data_2_in1[37] , bypass_mux_rs2_data_2_in1[38] ,
         bypass_mux_rs2_data_2_in1[39] , bypass_mux_rs2_data_2_in1[40] ,
         bypass_mux_rs2_data_2_in1[41] , bypass_mux_rs2_data_2_in1[42] ,
         bypass_mux_rs2_data_2_in1[43] , bypass_mux_rs2_data_2_in1[44] ,
         bypass_mux_rs2_data_2_in1[45] , bypass_mux_rs2_data_2_in1[46] ,
         bypass_mux_rs2_data_2_in1[47] , bypass_mux_rs2_data_2_in1[48] ,
         bypass_mux_rs2_data_2_in1[49] , bypass_mux_rs2_data_2_in1[50] ,
         bypass_mux_rs2_data_2_in1[51] , bypass_mux_rs2_data_2_in1[52] ,
         bypass_mux_rs2_data_2_in1[53] , bypass_mux_rs2_data_2_in1[54] ,
         bypass_mux_rs2_data_2_in1[55] , bypass_mux_rs2_data_2_in1[56] ,
         bypass_mux_rs2_data_2_in1[57] , bypass_mux_rs2_data_2_in1[58] ,
         bypass_mux_rs2_data_2_in1[59] , bypass_mux_rs2_data_2_in1[60] ,
         bypass_mux_rs2_data_2_in1[61] , bypass_mux_rs2_data_2_in1[62] ,
         bypass_mux_rs2_data_2_in1[63] , bypass_mux_rcc_data_2_in1[0] ,
         bypass_mux_rcc_data_2_in1[1] , bypass_mux_rcc_data_2_in1[2] ,
         bypass_mux_rcc_data_2_in1[3] , bypass_mux_rcc_data_2_in1[4] ,
         bypass_mux_rcc_data_2_in1[5] , bypass_mux_rcc_data_2_in1[6] ,
         bypass_mux_rcc_data_2_in1[7] , bypass_mux_rcc_data_2_in1[8] ,
         bypass_mux_rcc_data_2_in1[9] , bypass_mux_rcc_data_2_in1[10] ,
         bypass_mux_rcc_data_2_in1[11] , bypass_mux_rcc_data_2_in1[12] ,
         bypass_mux_rcc_data_2_in1[13] , bypass_mux_rcc_data_2_in1[14] ,
         bypass_mux_rcc_data_2_in1[15] , bypass_mux_rcc_data_2_in1[16] ,
         bypass_mux_rcc_data_2_in1[17] , bypass_mux_rcc_data_2_in1[18] ,
         bypass_mux_rcc_data_2_in1[19] , bypass_mux_rcc_data_2_in1[20] ,
         bypass_mux_rcc_data_2_in1[21] , bypass_mux_rcc_data_2_in1[22] ,
         bypass_mux_rcc_data_2_in1[23] , bypass_mux_rcc_data_2_in1[24] ,
         bypass_mux_rcc_data_2_in1[25] , bypass_mux_rcc_data_2_in1[26] ,
         bypass_mux_rcc_data_2_in1[27] , bypass_mux_rcc_data_2_in1[28] ,
         bypass_mux_rcc_data_2_in1[29] , bypass_mux_rcc_data_2_in1[30] ,
         bypass_mux_rcc_data_2_in1[31] , bypass_mux_rcc_data_2_in1[32] ,
         bypass_mux_rcc_data_2_in1[33] , bypass_mux_rcc_data_2_in1[34] ,
         bypass_mux_rcc_data_2_in1[35] , bypass_mux_rcc_data_2_in1[36] ,
         bypass_mux_rcc_data_2_in1[37] , bypass_mux_rcc_data_2_in1[38] ,
         bypass_mux_rcc_data_2_in1[39] , bypass_mux_rcc_data_2_in1[40] ,
         bypass_mux_rcc_data_2_in1[41] , bypass_mux_rcc_data_2_in1[42] ,
         bypass_mux_rcc_data_2_in1[43] , bypass_mux_rcc_data_2_in1[44] ,
         bypass_mux_rcc_data_2_in1[45] , bypass_mux_rcc_data_2_in1[46] ,
         bypass_mux_rcc_data_2_in1[47] , bypass_mux_rcc_data_2_in1[48] ,
         bypass_mux_rcc_data_2_in1[49] , bypass_mux_rcc_data_2_in1[50] ,
         bypass_mux_rcc_data_2_in1[51] , bypass_mux_rcc_data_2_in1[52] ,
         bypass_mux_rcc_data_2_in1[53] , bypass_mux_rcc_data_2_in1[54] ,
         bypass_mux_rcc_data_2_in1[55] , bypass_mux_rcc_data_2_in1[56] ,
         bypass_mux_rcc_data_2_in1[57] , bypass_mux_rcc_data_2_in1[58] ,
         bypass_mux_rcc_data_2_in1[59] , bypass_mux_rcc_data_2_in1[60] ,
         bypass_mux_rcc_data_2_in1[61] , bypass_mux_rcc_data_2_in1[62] ,
         bypass_mux_rcc_data_2_in1[63] , bypass_mux_rs3h_data_2_in1[0] ,
         bypass_mux_rs3h_data_2_in1[1] , bypass_mux_rs3h_data_2_in1[2] ,
         bypass_mux_rs3h_data_2_in1[3] , bypass_mux_rs3h_data_2_in1[4] ,
         bypass_mux_rs3h_data_2_in1[5] , bypass_mux_rs3h_data_2_in1[6] ,
         bypass_mux_rs3h_data_2_in1[7] , bypass_mux_rs3h_data_2_in1[8] ,
         bypass_mux_rs3h_data_2_in1[9] , bypass_mux_rs3h_data_2_in1[10] ,
         bypass_mux_rs3h_data_2_in1[11] , bypass_mux_rs3h_data_2_in1[12] ,
         bypass_mux_rs3h_data_2_in1[13] , bypass_mux_rs3h_data_2_in1[14] ,
         bypass_mux_rs3h_data_2_in1[15] , bypass_mux_rs3h_data_2_in1[16] ,
         bypass_mux_rs3h_data_2_in1[17] , bypass_mux_rs3h_data_2_in1[18] ,
         bypass_mux_rs3h_data_2_in1[19] , bypass_mux_rs3h_data_2_in1[20] ,
         bypass_mux_rs3h_data_2_in1[21] , bypass_mux_rs3h_data_2_in1[22] ,
         bypass_mux_rs3h_data_2_in1[23] , bypass_mux_rs3h_data_2_in1[24] ,
         bypass_mux_rs3h_data_2_in1[25] , bypass_mux_rs3h_data_2_in1[26] ,
         bypass_mux_rs3h_data_2_in1[27] , bypass_mux_rs3h_data_2_in1[28] ,
         bypass_mux_rs3h_data_2_in1[29] , bypass_mux_rs3h_data_2_in1[30] ,
         bypass_mux_rs3h_data_2_in1[31] , bypass_w2_eccgen_p7_g[0] ,
         bypass_w2_eccgen_p7_g[1] , bypass_w2_eccgen_p7_g[2] ,
         bypass_w2_eccgen_p7_g[3] , bypass_w2_eccgen_p7_g[4] ,
         bypass_w2_eccgen_p7_g[5] , bypass_w2_eccgen_p7_g[6] ,
         bypass_w2_eccgen_p7_g[7] , bypass_w2_eccgen_p7_w[7] ,
         bypass_w2_eccgen_p7_w[6] , bypass_w2_eccgen_p7_w[5] ,
         bypass_w2_eccgen_p7_w[4] , bypass_w2_eccgen_p7_w[3] ,
         bypass_w2_eccgen_p7_w[2] , bypass_w2_eccgen_p7_w[1] ,
         bypass_w2_eccgen_p7_w[0] , bypass_w2_eccgen_p6_g[1] ,
         bypass_w2_eccgen_p6_g[0] , bypass_w2_eccgen_p6_w[1] ,
         bypass_w2_eccgen_p6_w[0] , bypass_w2_eccgen_p5_g[1] ,
         bypass_w2_eccgen_p5_g[0] , bypass_w2_eccgen_p5_w[1] ,
         bypass_w2_eccgen_p5_w[0] , bypass_w2_eccgen_p4_g[3] ,
         bypass_w2_eccgen_p4_g[2] , bypass_w2_eccgen_p4_g[1] ,
         bypass_w2_eccgen_p4_g[0] , bypass_w2_eccgen_p4_w[0] ,
         bypass_w2_eccgen_p4_w[1] , bypass_w2_eccgen_p4_w[2] ,
         bypass_w2_eccgen_p4_w[3] , bypass_w2_eccgen_p3_g[0] ,
         bypass_w2_eccgen_p3_g[1] , bypass_w2_eccgen_p3_g[2] ,
         bypass_w2_eccgen_p3_g[3] , bypass_w2_eccgen_p3_g[4] ,
         bypass_w2_eccgen_p3_g[5] , bypass_w2_eccgen_p3_g[6] ,
         bypass_w2_eccgen_p3_g[7] , bypass_w2_eccgen_p3_w[7] ,
         bypass_w2_eccgen_p3_w[6] , bypass_w2_eccgen_p3_w[5] ,
         bypass_w2_eccgen_p3_w[4] , bypass_w2_eccgen_p3_w[3] ,
         bypass_w2_eccgen_p3_w[2] , bypass_w2_eccgen_p3_w[1] ,
         bypass_w2_eccgen_p3_w[0] , bypass_w2_eccgen_p2_g[7] ,
         bypass_w2_eccgen_p2_g[6] , bypass_w2_eccgen_p2_g[5] ,
         bypass_w2_eccgen_p2_g[4] , bypass_w2_eccgen_p2_g[3] ,
         bypass_w2_eccgen_p2_g[2] , bypass_w2_eccgen_p2_g[1] ,
         bypass_w2_eccgen_p2_g[0] , bypass_w2_eccgen_p2_w[7] ,
         bypass_w2_eccgen_p2_w[6] , bypass_w2_eccgen_p2_w[5] ,
         bypass_w2_eccgen_p2_w[4] , bypass_w2_eccgen_p2_w[3] ,
         bypass_w2_eccgen_p2_w[2] , bypass_w2_eccgen_p2_w[1] ,
         bypass_w2_eccgen_p2_w[0] , bypass_w2_eccgen_p1_g[7] ,
         bypass_w2_eccgen_p1_g[6] , bypass_w2_eccgen_p1_g[5] ,
         bypass_w2_eccgen_p1_g[4] , bypass_w2_eccgen_p1_g[3] ,
         bypass_w2_eccgen_p1_g[2] , bypass_w2_eccgen_p1_g[1] ,
         bypass_w2_eccgen_p1_g[0] , bypass_w2_eccgen_p1_w[7] ,
         bypass_w2_eccgen_p1_w[6] , bypass_w2_eccgen_p1_w[5] ,
         bypass_w2_eccgen_p1_w[4] , bypass_w2_eccgen_p1_w[3] ,
         bypass_w2_eccgen_p1_w[2] , bypass_w2_eccgen_p1_w[1] ,
         bypass_w2_eccgen_p1_w[0] , bypass_w2_eccgen_p0_g[7] ,
         bypass_w2_eccgen_p0_g[6] , bypass_w2_eccgen_p0_g[5] ,
         bypass_w2_eccgen_p0_g[4] , bypass_w2_eccgen_p0_g[3] ,
         bypass_w2_eccgen_p0_g[2] , bypass_w2_eccgen_p0_g[1] ,
         bypass_w2_eccgen_p0_g[0] , bypass_w2_eccgen_p0_w[7] ,
         bypass_w2_eccgen_p0_w[6] , bypass_w2_eccgen_p0_w[5] ,
         bypass_w2_eccgen_p0_w[4] , bypass_w2_eccgen_p0_w[3] ,
         bypass_w2_eccgen_p0_w[2] , bypass_w2_eccgen_p0_w[1] ,
         bypass_w2_eccgen_p0_w[0] , bypass_w2_eccgen_msk_w4 ,
         bypass_w2_eccgen_msk_w5 , ecc_chk_rs3_parity , ecc_chk_rs2_parity ,
         ecl_eccctl_ecc_sel_rs3_dff_din[0] , ecl_ld_thr_match_sg_dff_din[0] ,
         ecl_ld_thr_match_sm_dff_din[0] , ecl_thr_match_se_dff_din[0] ,
         ecl_thr_match_sd_dff_din[0] , ecl_thr_match_ew_dff_din[0] ,
         ecl_c_used_dff_din[0] , ecl_dff_sel_sum_d2e_din[0] ,
         ecl_byplog_rs3h_N3 , ecl_byplog_rs3h_N2 , ecl_byplog_rs3h_N1 ,
         ecl_byplog_rs3h_N0 , ecl_byplog_rs3h_match_w2 ,
         ecl_byplog_rs3h_match_w , ecl_byplog_rs3_N3 , ecl_byplog_rs3_N2 ,
         ecl_byplog_rs3_N1 , ecl_byplog_rs3_N0 , ecl_byplog_rs3_match_w2 ,
         ecl_byplog_rs3_match_w , rml_lo_wstate_reg_data_thr3_next[2] ,
         rml_lo_wstate_reg_data_thr3_next[1] ,
         rml_lo_wstate_reg_data_thr3_next[0] ,
         rml_lo_wstate_reg_data_thr2_next[2] ,
         rml_lo_wstate_reg_data_thr2_next[1] ,
         rml_lo_wstate_reg_data_thr2_next[0] ,
         rml_lo_wstate_reg_data_thr1_next[2] ,
         rml_lo_wstate_reg_data_thr1_next[1] ,
         rml_lo_wstate_reg_data_thr1_next[0] ,
         rml_lo_wstate_reg_data_thr0_next[2] ,
         rml_lo_wstate_reg_data_thr0_next[1] ,
         rml_lo_wstate_reg_data_thr0_next[0] ,
         rml_lo_wstate_reg_data_thr3[0] , rml_lo_wstate_reg_data_thr3[1] ,
         rml_lo_wstate_reg_data_thr3[2] , rml_lo_wstate_reg_data_thr2[0] ,
         rml_lo_wstate_reg_data_thr2[1] , rml_lo_wstate_reg_data_thr2[2] ,
         rml_lo_wstate_reg_data_thr1[0] , rml_lo_wstate_reg_data_thr1[1] ,
         rml_lo_wstate_reg_data_thr1[2] , rml_lo_wstate_reg_data_thr0[0] ,
         rml_lo_wstate_reg_data_thr0[1] , rml_lo_wstate_reg_data_thr0[2] ,
         rml_hi_wstate_reg_data_thr3_next[2] ,
         rml_hi_wstate_reg_data_thr3_next[1] ,
         rml_hi_wstate_reg_data_thr3_next[0] ,
         rml_hi_wstate_reg_data_thr2_next[2] ,
         rml_hi_wstate_reg_data_thr2_next[1] ,
         rml_hi_wstate_reg_data_thr2_next[0] ,
         rml_hi_wstate_reg_data_thr1_next[2] ,
         rml_hi_wstate_reg_data_thr1_next[1] ,
         rml_hi_wstate_reg_data_thr1_next[0] ,
         rml_hi_wstate_reg_data_thr0_next[2] ,
         rml_hi_wstate_reg_data_thr0_next[1] ,
         rml_hi_wstate_reg_data_thr0_next[0] ,
         rml_hi_wstate_reg_data_thr3[0] , rml_hi_wstate_reg_data_thr3[1] ,
         rml_hi_wstate_reg_data_thr3[2] , rml_hi_wstate_reg_data_thr2[0] ,
         rml_hi_wstate_reg_data_thr2[1] , rml_hi_wstate_reg_data_thr2[2] ,
         rml_hi_wstate_reg_data_thr1[0] , rml_hi_wstate_reg_data_thr1[1] ,
         rml_hi_wstate_reg_data_thr1[2] , rml_hi_wstate_reg_data_thr0[0] ,
         rml_hi_wstate_reg_data_thr0[1] , rml_hi_wstate_reg_data_thr0[2] ,
         rml_cleanwin_reg_data_thr3_next[2] ,
         rml_cleanwin_reg_data_thr3_next[1] ,
         rml_cleanwin_reg_data_thr3_next[0] ,
         rml_cleanwin_reg_data_thr2_next[2] ,
         rml_cleanwin_reg_data_thr2_next[1] ,
         rml_cleanwin_reg_data_thr2_next[0] ,
         rml_cleanwin_reg_data_thr1_next[2] ,
         rml_cleanwin_reg_data_thr1_next[1] ,
         rml_cleanwin_reg_data_thr1_next[0] ,
         rml_cleanwin_reg_data_thr0_next[2] ,
         rml_cleanwin_reg_data_thr0_next[1] ,
         rml_cleanwin_reg_data_thr0_next[0] , rml_cleanwin_reg_data_thr3[0] ,
         rml_cleanwin_reg_data_thr3[1] , rml_cleanwin_reg_data_thr3[2] ,
         rml_cleanwin_reg_data_thr2[0] , rml_cleanwin_reg_data_thr2[1] ,
         rml_cleanwin_reg_data_thr2[2] , rml_cleanwin_reg_data_thr1[0] ,
         rml_cleanwin_reg_data_thr1[1] , rml_cleanwin_reg_data_thr1[2] ,
         rml_cleanwin_reg_data_thr0[0] , rml_cleanwin_reg_data_thr0[1] ,
         rml_cleanwin_reg_data_thr0[2] , rml_otherwin_reg_data_thr3_next[2] ,
         rml_otherwin_reg_data_thr3_next[1] ,
         rml_otherwin_reg_data_thr3_next[0] ,
         rml_otherwin_reg_data_thr2_next[2] ,
         rml_otherwin_reg_data_thr2_next[1] ,
         rml_otherwin_reg_data_thr2_next[0] ,
         rml_otherwin_reg_data_thr1_next[2] ,
         rml_otherwin_reg_data_thr1_next[1] ,
         rml_otherwin_reg_data_thr1_next[0] ,
         rml_otherwin_reg_data_thr0_next[2] ,
         rml_otherwin_reg_data_thr0_next[1] ,
         rml_otherwin_reg_data_thr0_next[0] , rml_otherwin_reg_data_thr3[0] ,
         rml_otherwin_reg_data_thr3[1] , rml_otherwin_reg_data_thr3[2] ,
         rml_otherwin_reg_data_thr2[0] , rml_otherwin_reg_data_thr2[1] ,
         rml_otherwin_reg_data_thr2[2] , rml_otherwin_reg_data_thr1[0] ,
         rml_otherwin_reg_data_thr1[1] , rml_otherwin_reg_data_thr1[2] ,
         rml_otherwin_reg_data_thr0[0] , rml_otherwin_reg_data_thr0[1] ,
         rml_otherwin_reg_data_thr0[2] ,
         rml_canrestore_reg_data_thr3_next[2] ,
         rml_canrestore_reg_data_thr3_next[1] ,
         rml_canrestore_reg_data_thr3_next[0] ,
         rml_canrestore_reg_data_thr2_next[2] ,
         rml_canrestore_reg_data_thr2_next[1] ,
         rml_canrestore_reg_data_thr2_next[0] ,
         rml_canrestore_reg_data_thr1_next[2] ,
         rml_canrestore_reg_data_thr1_next[1] ,
         rml_canrestore_reg_data_thr1_next[0] ,
         rml_canrestore_reg_data_thr0_next[2] ,
         rml_canrestore_reg_data_thr0_next[1] ,
         rml_canrestore_reg_data_thr0_next[0] ,
         rml_canrestore_reg_data_thr3[0] , rml_canrestore_reg_data_thr3[1] ,
         rml_canrestore_reg_data_thr3[2] , rml_canrestore_reg_data_thr2[0] ,
         rml_canrestore_reg_data_thr2[1] , rml_canrestore_reg_data_thr2[2] ,
         rml_canrestore_reg_data_thr1[0] , rml_canrestore_reg_data_thr1[1] ,
         rml_canrestore_reg_data_thr1[2] , rml_canrestore_reg_data_thr0[0] ,
         rml_canrestore_reg_data_thr0[1] , rml_canrestore_reg_data_thr0[2] ,
         ecl_divcntl_subnext_mux_in1[0] , ecl_ccr_mux_ccr_bypass1_sel0 ,
         ecl_ccr_mux_ccrin3_sel2 , ecl_ccr_mux_ccrin2_sel2 ,
         ecl_ccr_mux_ccrin1_sel2 , ecl_writeback_rdpr_mux2_sel3 ,
         rml_cwp_cwp_next3_mux_sel0 , rml_cwp_cwp_next2_mux_sel0 ,
         rml_cwp_cwp_next1_mux_sel0 , rml_cwp_cwp_next0_mux_sel0 , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15034, n15035,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15410, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
         n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936,
         n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
         n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952,
         n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960,
         n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
         n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
         n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
         n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
         n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000,
         n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008,
         n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
         n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024,
         n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032,
         n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
         n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
         n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
         n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064,
         n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072,
         n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080,
         n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
         n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096,
         n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
         n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
         n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120,
         n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
         n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136,
         n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144,
         n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152,
         n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
         n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168,
         n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
         n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184,
         n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192,
         n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
         n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208,
         n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216,
         n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224,
         n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
         n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240,
         n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
         n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256,
         n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264,
         n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
         n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280,
         n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288,
         n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296,
         n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
         n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
         n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320,
         n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328,
         n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
         n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
         n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352,
         n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360,
         n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368,
         n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
         n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
         n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392,
         n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400,
         n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
         n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
         n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424,
         n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432,
         n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440,
         n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
         n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456,
         n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464,
         n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472,
         n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
         n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
         n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496,
         n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504,
         n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512,
         n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
         n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528,
         n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536,
         n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544,
         n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
         n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
         n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568,
         n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
         n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
         n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592,
         n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600,
         n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608,
         n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616,
         n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
         n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
         n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640,
         n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
         n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656,
         n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664,
         n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672,
         n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680,
         n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688,
         n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
         n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
         n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712,
         n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
         n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728,
         n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736,
         n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744,
         n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752,
         n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760,
         n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
         n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
         n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
         n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
         n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800,
         n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808,
         n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816,
         n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824,
         n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832,
         n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
         n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
         n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856,
         n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
         n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872,
         n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880,
         n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888,
         n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896,
         n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904,
         n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
         n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
         n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928,
         n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
         n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944,
         n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952,
         n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960,
         n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968,
         n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976,
         n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
         n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
         n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000,
         n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
         n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016,
         n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024,
         n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032,
         n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040,
         n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
         n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
         n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
         n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072,
         n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
         n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088,
         n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096,
         n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104,
         n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112,
         n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120,
         n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
         n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
         n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144,
         n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
         n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160,
         n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168,
         n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176,
         n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
         n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192,
         n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
         n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
         n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216,
         n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
         n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232,
         n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240,
         n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
         n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256,
         n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264,
         n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
         n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
         n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288,
         n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
         n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304,
         n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
         n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320,
         n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328,
         n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336,
         n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
         n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
         n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360,
         n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
         n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
         n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384,
         n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392,
         n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400,
         n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408,
         n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
         n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
         n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432,
         n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
         n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448,
         n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456,
         n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464,
         n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472,
         n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480,
         n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
         n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
         n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
         n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,
         n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520,
         n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528,
         n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536,
         n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544,
         n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552,
         n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
         n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
         n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576,
         n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
         n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592,
         n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600,
         n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608,
         n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616,
         n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
         n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
         n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
         n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648,
         n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
         n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664,
         n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672,
         n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680,
         n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688,
         n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696,
         n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
         n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
         n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720,
         n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,
         n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736,
         n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744,
         n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752,
         n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760,
         n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768,
         n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
         n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
         n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792,
         n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
         n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808,
         n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816,
         n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824,
         n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832,
         n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840,
         n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
         n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
         n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864,
         n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
         n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880,
         n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888,
         n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896,
         n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904,
         n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,
         n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920,
         n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
         n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936,
         n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
         n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952,
         n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960,
         n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968,
         n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976,
         n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
         n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992,
         n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
         n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008,
         n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,
         n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024,
         n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032,
         n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040,
         n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048,
         n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,
         n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064,
         n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
         n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080,
         n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
         n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096,
         n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104,
         n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
         n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120,
         n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
         n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136,
         n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
         n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152,
         n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
         n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
         n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176,
         n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184,
         n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192,
         n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
         n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208,
         n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216,
         n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224,
         n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
         n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
         n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248,
         n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256,
         n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264,
         n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
         n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280,
         n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288,
         n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296,
         n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
         n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312,
         n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320,
         n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328,
         n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336,
         n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
         n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352,
         n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360,
         n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368,
         n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
         n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384,
         n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392,
         n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400,
         n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408,
         n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
         n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424,
         n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432,
         n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440,
         n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
         n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456,
         n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,
         n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472,
         n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480,
         n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488,
         n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496,
         n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504,
         n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512,
         n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
         n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528,
         n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536,
         n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544,
         n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
         n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560,
         n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568,
         n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576,
         n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584,
         n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
         n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600,
         n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608,
         n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616,
         n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624,
         n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632,
         n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640,
         n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648,
         n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656,
         n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
         n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672,
         n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,
         n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688,
         n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696,
         n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
         n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712,
         n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720,
         n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728,
         n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
         n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744,
         n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
         n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760,
         n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768,
         n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
         n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784,
         n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792,
         n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800,
         n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
         n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816,
         n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
         n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832,
         n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840,
         n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848,
         n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856,
         n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864,
         n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872,
         n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
         n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888,
         n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,
         n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904,
         n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
         n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,
         n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928,
         n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936,
         n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944,
         n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,
         n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960,
         n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968,
         n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976,
         n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984,
         n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992,
         n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000,
         n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008,
         n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016,
         n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,
         n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032,
         n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040,
         n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048,
         n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056,
         n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064,
         n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072,
         n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080,
         n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088,
         n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
         n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104,
         n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,
         n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120,
         n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128,
         n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136,
         n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144,
         n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152,
         n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160,
         n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
         n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176,
         n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184,
         n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192,
         n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200,
         n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
         n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216,
         n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224,
         n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232,
         n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
         n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
         n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256,
         n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264,
         n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272,
         n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
         n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288,
         n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296,
         n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304,
         n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,
         n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
         n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328,
         n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336,
         n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344,
         n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
         n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360,
         n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368,
         n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376,
         n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384,
         n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
         n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400,
         n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408,
         n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416,
         n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424,
         n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432,
         n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440,
         n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448,
         n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456,
         n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,
         n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472,
         n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480,
         n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488,
         n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496,
         n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504,
         n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512,
         n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520,
         n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528,
         n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,
         n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544,
         n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552,
         n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560,
         n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,
         n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576,
         n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584,
         n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592,
         n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600,
         n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,
         n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616,
         n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624,
         n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632,
         n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640,
         n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648,
         n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656,
         n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664,
         n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672,
         n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,
         n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688,
         n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696,
         n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704,
         n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712,
         n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720,
         n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728,
         n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736,
         n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744,
         n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752,
         n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760,
         n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768,
         n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776,
         n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,
         n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792,
         n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800,
         n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808,
         n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816,
         n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824,
         n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832,
         n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840,
         n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,
         n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856,
         n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864,
         n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872,
         n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880,
         n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888,
         n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896,
         n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904,
         n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912,
         n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
         n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928,
         n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936,
         n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,
         n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952,
         n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960,
         n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968,
         n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976,
         n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984,
         n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,
         n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000,
         n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008,
         n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
         n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024,
         n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,
         n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040,
         n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048,
         n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056,
         n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
         n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072,
         n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080,
         n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
         n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096,
         n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,
         n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112,
         n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120,
         n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128,
         n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
         n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144,
         n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152,
         n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160,
         n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168,
         n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176,
         n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184,
         n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192,
         n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200,
         n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
         n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216,
         n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224,
         n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232,
         n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240,
         n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248,
         n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256,
         n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264,
         n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272,
         n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280,
         n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288,
         n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296,
         n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
         n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312,
         n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320,
         n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328,
         n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336,
         n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344,
         n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352,
         n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360,
         n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368,
         n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376,
         n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384,
         n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392,
         n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400,
         n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408,
         n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
         n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
         n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432,
         n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440,
         n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448,
         n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456,
         n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464,
         n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472,
         n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480,
         n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488,
         n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,
         n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504,
         n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512,
         n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520,
         n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528,
         n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536,
         n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544,
         n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552,
         n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,
         n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568,
         n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576,
         n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584,
         n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592,
         n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600,
         n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608,
         n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616,
         n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624,
         n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,
         n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640,
         n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648,
         n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656,
         n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664,
         n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672,
         n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680,
         n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688,
         n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696,
         n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704,
         n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712,
         n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720,
         n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728,
         n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736,
         n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744,
         n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752,
         n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760,
         n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768,
         n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776,
         n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784,
         n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792,
         n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800,
         n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808,
         n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816,
         n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824,
         n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832,
         n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840,
         n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848,
         n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856,
         n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864,
         n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872,
         n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880,
         n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888,
         n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896,
         n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904,
         n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912,
         n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920,
         n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,
         n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936,
         n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944,
         n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952,
         n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960,
         n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968,
         n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,
         n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
         n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992,
         n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,
         n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008,
         n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016,
         n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024,
         n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032,
         n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040,
         n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
         n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,
         n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064,
         n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
         n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080,
         n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088,
         n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096,
         n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104,
         n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,
         n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120,
         n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,
         n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136,
         n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
         n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152,
         n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160,
         n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168,
         n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176,
         n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
         n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192,
         n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,
         n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208,
         n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
         n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224,
         n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232,
         n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240,
         n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248,
         n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,
         n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264,
         n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,
         n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280,
         n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
         n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296,
         n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304,
         n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312,
         n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
         n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328,
         n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336,
         n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,
         n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352,
         n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360,
         n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368,
         n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376,
         n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384,
         n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
         n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400,
         n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408,
         n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,
         n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
         n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432,
         n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440,
         n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448,
         n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456,
         n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464,
         n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472,
         n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480,
         n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
         n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
         n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504,
         n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512,
         n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520,
         n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
         n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536,
         n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544,
         n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552,
         n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,
         n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
         n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576,
         n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584,
         n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592,
         n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
         n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608,
         n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616,
         n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624,
         n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632,
         n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
         n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648,
         n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656,
         n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
         n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
         n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680,
         n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688,
         n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696,
         n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704,
         n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
         n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720,
         n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728,
         n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
         n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744,
         n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752,
         n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,
         n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768,
         n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776,
         n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
         n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792,
         n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800,
         n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
         n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816,
         n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824,
         n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
         n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840,
         n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848,
         n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
         n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864,
         n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
         n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880,
         n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888,
         n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896,
         n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
         n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912,
         n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920,
         n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
         n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936,
         n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,
         n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952,
         n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960,
         n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968,
         n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
         n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984,
         n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992,
         n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,
         n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008,
         n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016,
         n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024,
         n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,
         n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040,
         n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048,
         n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056,
         n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064,
         n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
         n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
         n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088,
         n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096,
         n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104,
         n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112,
         n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120,
         n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128,
         n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,
         n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
         n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152,
         n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160,
         n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168,
         n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176,
         n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184,
         n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192,
         n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200,
         n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,
         n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
         n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224,
         n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232,
         n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240,
         n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248,
         n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256,
         n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264,
         n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272,
         n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280,
         n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
         n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296,
         n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304,
         n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312,
         n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320,
         n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328,
         n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336,
         n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344,
         n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
         n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
         n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368,
         n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376,
         n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384,
         n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392,
         n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400,
         n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408,
         n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
         n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424,
         n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
         n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440,
         n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448,
         n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456,
         n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464,
         n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472,
         n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480,
         n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
         n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496,
         n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
         n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512,
         n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520,
         n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528,
         n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536,
         n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544,
         n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552,
         n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560,
         n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568,
         n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
         n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584,
         n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592,
         n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600,
         n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608,
         n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616,
         n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624,
         n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632,
         n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640,
         n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
         n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656,
         n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664,
         n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672,
         n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680,
         n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688,
         n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696,
         n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704,
         n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712,
         n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,
         n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728,
         n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736,
         n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744,
         n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752,
         n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760,
         n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768,
         n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776,
         n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784,
         n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
         n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800,
         n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808,
         n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816,
         n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
         n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832,
         n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840,
         n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848,
         n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856,
         n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,
         n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872,
         n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880,
         n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
         n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896,
         n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904,
         n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912,
         n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920,
         n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928,
         n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,
         n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944,
         n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952,
         n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
         n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
         n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976,
         n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984,
         n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992,
         n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000,
         n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
         n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016,
         n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024,
         n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032,
         n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,
         n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048,
         n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056,
         n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064,
         n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072,
         n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,
         n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088,
         n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096,
         n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104,
         n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,
         n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120,
         n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128,
         n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,
         n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144,
         n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
         n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160,
         n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168,
         n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176,
         n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
         n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192,
         n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200,
         n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208,
         n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216,
         n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224,
         n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232,
         n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240,
         n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,
         n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256,
         n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264,
         n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272,
         n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280,
         n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288,
         n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296,
         n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304,
         n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312,
         n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320,
         n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328,
         n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336,
         n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344,
         n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352,
         n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360,
         n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368,
         n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376,
         n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384,
         n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
         n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400,
         n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408,
         n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416,
         n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424,
         n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
         n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440,
         n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448,
         n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456,
         n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
         n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472,
         n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480,
         n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488,
         n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
         n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504,
         n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512,
         n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520,
         n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528,
         n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536,
         n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544,
         n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552,
         n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560,
         n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568,
         n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576,
         n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584,
         n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592,
         n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600,
         n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608,
         n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616,
         n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624,
         n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632,
         n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640,
         n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648,
         n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656,
         n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664,
         n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672,
         n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680,
         n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688,
         n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696,
         n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704,
         n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712,
         n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720,
         n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728,
         n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736,
         n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744,
         n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752,
         n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760,
         n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768,
         n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776,
         n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784,
         n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792,
         n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800,
         n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808,
         n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816,
         n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824,
         n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832,
         n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840,
         n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848,
         n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856,
         n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864,
         n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872,
         n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880,
         n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888,
         n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896,
         n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904,
         n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912,
         n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920,
         n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928,
         n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936,
         n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944,
         n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952,
         n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960,
         n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968,
         n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976,
         n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984,
         n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992,
         n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000,
         n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008,
         n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016,
         n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024,
         n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032,
         n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040,
         n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048,
         n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056,
         n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064,
         n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072,
         n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080,
         n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088,
         n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096,
         n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104,
         n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112,
         n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120,
         n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128,
         n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136,
         n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144,
         n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152,
         n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160,
         n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168,
         n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176,
         n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184,
         n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192,
         n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200,
         n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208,
         n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216,
         n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224,
         n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232,
         n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240,
         n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248,
         n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256,
         n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264,
         n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272,
         n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280,
         n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288,
         n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296,
         n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304,
         n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312,
         n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320,
         n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328,
         n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336,
         n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344,
         n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352,
         n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360,
         n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368,
         n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376,
         n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384,
         n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392,
         n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400,
         n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408,
         n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416,
         n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424,
         n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432,
         n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440,
         n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448,
         n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
         n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464,
         n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472,
         n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480,
         n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488,
         n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496,
         n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504,
         n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512,
         n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520,
         n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528,
         n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536,
         n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544,
         n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552,
         n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560,
         n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568,
         n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576,
         n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584,
         n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592,
         n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600,
         n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608,
         n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616,
         n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624,
         n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632,
         n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640,
         n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648,
         n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656,
         n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
         n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672,
         n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680,
         n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688,
         n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696,
         n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704,
         n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712,
         n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720,
         n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728,
         n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736,
         n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744,
         n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752,
         n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760,
         n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768,
         n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776,
         n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784,
         n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792,
         n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800,
         n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808,
         n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816,
         n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824,
         n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832,
         n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840,
         n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848,
         n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856,
         n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864,
         n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872,
         n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880,
         n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888,
         n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896,
         n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904,
         n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912,
         n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920,
         n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928,
         n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936,
         n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944,
         n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952,
         n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960,
         n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968,
         n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976,
         n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984,
         n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992,
         n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000,
         n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008,
         n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016,
         n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024,
         n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032,
         n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040,
         n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048,
         n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056,
         n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064,
         n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072,
         n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
         n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088,
         n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096,
         n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104,
         n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112,
         n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120,
         n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128,
         n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136,
         n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144,
         n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152,
         n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160,
         n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168,
         n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176,
         n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184,
         n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192,
         n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200,
         n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208,
         n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216,
         n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224,
         n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232,
         n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240,
         n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248,
         n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256,
         n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264,
         n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272,
         n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280,
         n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288,
         n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296,
         n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304,
         n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312,
         n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320,
         n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328,
         n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336,
         n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344,
         n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352,
         n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360,
         n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368,
         n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376,
         n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384,
         n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392,
         n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400,
         n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408,
         n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416,
         n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424,
         n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432,
         n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
         n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448,
         n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456,
         n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464,
         n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472,
         n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480,
         n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488,
         n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496,
         n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504,
         n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
         n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520,
         n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528,
         n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536,
         n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544,
         n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552,
         n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560,
         n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568,
         n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576,
         n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584,
         n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592,
         n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600,
         n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608,
         n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616,
         n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624,
         n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632,
         n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640,
         n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648,
         n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656,
         n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664,
         n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672,
         n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680,
         n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688,
         n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696,
         n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704,
         n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712,
         n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720,
         n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728,
         n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736,
         n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744,
         n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752,
         n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760,
         n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768,
         n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776,
         n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784,
         n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792,
         n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
         n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808,
         n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816,
         n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824,
         n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832,
         n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840,
         n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848,
         n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856,
         n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864,
         n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872,
         n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880,
         n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888,
         n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896,
         n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904,
         n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912,
         n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920,
         n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928,
         n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936,
         n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944,
         n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952,
         n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960,
         n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968,
         n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976,
         n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984,
         n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992,
         n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000,
         n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008,
         n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016,
         n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024,
         n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032,
         n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040,
         n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048,
         n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056,
         n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064,
         n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072,
         n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080,
         n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088,
         n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096,
         n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104,
         n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112,
         n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120,
         n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128,
         n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136,
         n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144,
         n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152,
         n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160,
         n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168,
         n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176,
         n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184,
         n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192,
         n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200,
         n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208,
         n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216,
         n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224,
         n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232,
         n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240,
         n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248,
         n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256,
         n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264,
         n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272,
         n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280,
         n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288,
         n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296,
         n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304,
         n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312,
         n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320,
         n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328,
         n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336,
         n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344,
         n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352,
         n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360,
         n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368,
         n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376,
         n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384,
         n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392,
         n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400,
         n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408,
         n30413, n30414, n30425, n30426, n30437, n30438, n30447, n30448,
         n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456,
         n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464,
         n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472,
         n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480,
         n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488,
         n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496,
         n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504,
         n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512,
         n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520,
         n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528,
         n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536,
         n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544,
         n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552,
         n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560,
         n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568,
         n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576,
         n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584,
         n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592,
         n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600,
         n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608,
         n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616,
         n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624,
         n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632,
         n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640,
         n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648,
         n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656,
         n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664,
         n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672,
         n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680,
         n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688,
         n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696,
         n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704,
         n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712,
         n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720,
         n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728,
         n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736,
         n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744,
         n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752,
         n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760,
         n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768,
         n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776,
         n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784,
         n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792,
         n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800,
         n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808,
         n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816,
         n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824,
         n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832,
         n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840,
         n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848,
         n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856,
         n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864,
         n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872,
         n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880,
         n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888,
         n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896,
         n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904,
         n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912,
         n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920,
         n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928,
         n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936,
         n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944,
         n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952,
         n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960,
         n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968,
         n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976,
         n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984,
         n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992,
         n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000,
         n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008,
         n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016,
         n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024,
         n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032,
         n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040,
         n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048,
         n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056,
         n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064,
         n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072,
         n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080,
         n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088,
         n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096,
         n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104,
         n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112,
         n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120,
         n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128,
         n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136,
         n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144,
         n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152,
         n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160,
         n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168,
         n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176,
         n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184,
         n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192,
         n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200,
         n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208,
         n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216,
         n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224,
         n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232,
         n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240,
         n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248,
         n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256,
         n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264,
         n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272,
         n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280,
         n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288,
         n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296,
         n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304,
         n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312,
         n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320,
         n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328,
         n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336,
         n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344,
         n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352,
         n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360,
         n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368,
         n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376,
         n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384,
         n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392,
         n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400,
         n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408,
         n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416,
         n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424,
         n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432,
         n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440,
         n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448,
         n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456,
         n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464,
         n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472,
         n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480,
         n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488,
         n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496,
         n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504,
         n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512,
         n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520,
         n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528,
         n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536,
         n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544,
         n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552,
         n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560,
         n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568,
         n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576,
         n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584,
         n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592,
         n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600,
         n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608,
         n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616,
         n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624,
         n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632,
         n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640,
         n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648,
         n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656,
         n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664,
         n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672,
         n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680,
         n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688,
         n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696,
         n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704;
  wire   [63:0] byp_alu_rcc_data_e;
  wire   [7:0] byp_ecc_rs1_synd_d;
  wire   [7:0] byp_ecc_rs2_synd_d;
  wire   [7:0] byp_ecc_rs3_synd_d;
  wire   [63:0] alu_byp_rd_data_e;
  wire   [63:0] div_byp_muldivout_g;
  wire   [63:0] ecc_byp_ecc_result_m;
  wire   [7:0] ecl_byp_ecc_mask_m_l;
  wire   [2:0] ecl_byp_3lsb_m;
  wire   [7:0] ecl_byp_eclpr_e;
  wire   [31:0] div_byp_yreg_e;
  wire   [3:0] ecl_div_yreg_wen_l;
  wire   [3:0] ecl_div_yreg_wen_w;
  wire   [3:0] ecl_shft_shift4_e;
  wire   [3:0] ecl_shft_shift1_e;
  wire   [3:0] ecl_div_thr_e;
  wire   [3:0] ecl_rml_thr_m;
  wire   [3:0] ecl_rml_thr_w;
  wire   [2:0] ecl_rml_xor_data_e;
  wire   [2:0] rml_ecl_canrestore_d;
  wire   [2:0] rml_ecl_cansave_d;
  wire   [2:0] rml_ecl_cleanwin_d;
  wire   [2:0] rml_ecl_cwp_d;
  wire   [1:0] rml_ecl_gl_e;
  wire   [2:0] rml_ecl_otherwin_d;
  wire   [3:0] rml_ecl_swap_done;
  wire   [5:0] rml_ecl_wstate_d;
  wire   [2:0] rml_ecl_wtype_e;
  wire   [63:0] shft_alu_shift_out_e;
  tri   [1:0] tlu_exu_agp_tid;
  tri   tlu_exu_agp_swap;
  tri   [1:0] tlu_exu_agp;
  tri   sehold;
  tri   se;
  tri   rclk;
  tri   [1:0] ifu_exu_tid_s2;
  tri   [4:0] ifu_exu_rs3_s;
  tri   [4:0] ifu_exu_rs2_s;
  tri   [4:0] ifu_exu_rs1_s;
  tri   ifu_exu_ren3_s;
  tri   ifu_exu_ren2_s;
  tri   ifu_exu_ren1_s;
  tri   arst_l;
  tri   mem_write_disable;
  tri   short_si0;
  tri   [1:0] rml_irf_old_e_cwp_e;
  tri   [1:0] rml_irf_new_e_cwp_e;
  tri   [71:0] irf_byp_rs1_data_d_l;
  tri   [71:0] irf_byp_rs2_data_d_l;
  tri   [71:0] irf_byp_rs3_data_d_l;
  tri   [31:0] irf_byp_rs3h_data_d_l;
  tri   ecl_irf_wen_w;
  tri   [4:0] ecl_irf_rd_m;
  tri   [4:0] ecl_irf_rd_g;
  tri   [71:0] byp_irf_rd_data_w;
  tri   [71:0] byp_irf_rd_data_w2;
  tri   [1:0] ecl_irf_tid_m;
  tri   [1:0] ecl_irf_tid_g;
  tri   [2:0] rml_irf_old_lo_cwp_e;
  tri   [2:0] rml_irf_new_lo_cwp_e;
  tri   rml_irf_swap_even_e;
  tri   rml_irf_swap_odd_e;
  tri   rml_irf_swap_local_e;
  tri   rml_irf_kill_restore_w;
  tri   [1:0] rml_irf_cwpswap_tid_e;
  tri   [1:0] rml_irf_old_agp;
  tri   ecl_wb_byplog_wen_w2 ;
  tri   short_scan0_1;
  assign exu_lsu_early_va_e[10] = exu_ifu_brpc_e[10];
  assign exu_lsu_early_va_e[9] = exu_ifu_brpc_e[9];
  assign exu_lsu_early_va_e[8] = exu_ifu_brpc_e[8];
  assign exu_lsu_early_va_e[7] = exu_ifu_brpc_e[7];
  assign exu_mmu_early_va_e[7] = exu_ifu_brpc_e[7];
  assign exu_lsu_early_va_e[6] = exu_ifu_brpc_e[6];
  assign exu_mmu_early_va_e[6] = exu_ifu_brpc_e[6];
  assign exu_lsu_early_va_e[5] = exu_ifu_brpc_e[5];
  assign exu_mmu_early_va_e[5] = exu_ifu_brpc_e[5];
  assign exu_lsu_early_va_e[4] = exu_ifu_brpc_e[4];
  assign exu_mmu_early_va_e[4] = exu_ifu_brpc_e[4];
  assign exu_lsu_early_va_e[3] = exu_ifu_brpc_e[3];
  assign exu_mmu_early_va_e[3] = exu_ifu_brpc_e[3];
  assign exu_mmu_early_va_e[2] = exu_ifu_brpc_e[2];
  assign exu_mmu_early_va_e[1] = exu_ifu_brpc_e[1];
  assign exu_mmu_early_va_e[0] = exu_ifu_brpc_e[0];
  assign short_so1 = 1'b0;
  assign short_so0 = 1'b0;
  assign so0 = 1'b0;

BUFX1 exu_exu_assign_1(.A(ifu_exu_kill_e), .Y(ecl_rml_kill_e));
BUFX1 exu_exu_assign_2(.A(ifu_exu_use_rsr_e_l), .Y(ecl_byp_sel_alu_e));
XOR2X1 exu_ecc_U67(.A(ecc_error_data_m[0]), .B(exu_n15186), .Y(ecc_byp_ecc_result_m[0]));
XOR2X1 exu_ecc_U66(.A(ecc_error_data_m[10]), .B(exu_n15185), .Y(ecc_byp_ecc_result_m[10]));
XOR2X1 exu_ecc_U65(.A(ecc_error_data_m[11]), .B(exu_n15184), .Y(ecc_byp_ecc_result_m[11]));
XOR2X1 exu_ecc_U64(.A(ecc_error_data_m[12]), .B(exu_n15183), .Y(ecc_byp_ecc_result_m[12]));
XOR2X1 exu_ecc_U63(.A(ecc_error_data_m[13]), .B(exu_n15182), .Y(ecc_byp_ecc_result_m[13]));
XOR2X1 exu_ecc_U62(.A(ecc_error_data_m[14]), .B(exu_n15181), .Y(ecc_byp_ecc_result_m[14]));
XOR2X1 exu_ecc_U61(.A(ecc_error_data_m[15]), .B(exu_n15180), .Y(ecc_byp_ecc_result_m[15]));
XOR2X1 exu_ecc_U60(.A(ecc_error_data_m[16]), .B(exu_n15179), .Y(ecc_byp_ecc_result_m[16]));
XOR2X1 exu_ecc_U59(.A(ecc_error_data_m[17]), .B(exu_n15178), .Y(ecc_byp_ecc_result_m[17]));
XOR2X1 exu_ecc_U58(.A(ecc_error_data_m[18]), .B(exu_n15177), .Y(ecc_byp_ecc_result_m[18]));
XOR2X1 exu_ecc_U57(.A(ecc_error_data_m[19]), .B(exu_n15176), .Y(ecc_byp_ecc_result_m[19]));
XOR2X1 exu_ecc_U56(.A(ecc_error_data_m[1]), .B(exu_n15175), .Y(ecc_byp_ecc_result_m[1]));
XOR2X1 exu_ecc_U55(.A(ecc_error_data_m[20]), .B(exu_n15174), .Y(ecc_byp_ecc_result_m[20]));
XOR2X1 exu_ecc_U54(.A(ecc_error_data_m[21]), .B(exu_n15173), .Y(ecc_byp_ecc_result_m[21]));
XOR2X1 exu_ecc_U53(.A(ecc_error_data_m[22]), .B(exu_n15172), .Y(ecc_byp_ecc_result_m[22]));
XOR2X1 exu_ecc_U52(.A(ecc_error_data_m[23]), .B(exu_n15171), .Y(ecc_byp_ecc_result_m[23]));
XOR2X1 exu_ecc_U51(.A(ecc_error_data_m[24]), .B(exu_n15170), .Y(ecc_byp_ecc_result_m[24]));
XOR2X1 exu_ecc_U50(.A(ecc_error_data_m[25]), .B(exu_n15169), .Y(ecc_byp_ecc_result_m[25]));
XOR2X1 exu_ecc_U49(.A(exu_n15116), .B(exu_n15168), .Y(ecc_byp_ecc_result_m[26]));
XOR2X1 exu_ecc_U48(.A(exu_n15115), .B(exu_n15167), .Y(ecc_byp_ecc_result_m[27]));
XOR2X1 exu_ecc_U47(.A(exu_n15114), .B(exu_n15166), .Y(ecc_byp_ecc_result_m[28]));
XOR2X1 exu_ecc_U46(.A(exu_n15113), .B(exu_n15165), .Y(ecc_byp_ecc_result_m[29]));
XOR2X1 exu_ecc_U45(.A(ecc_error_data_m[2]), .B(exu_n15164), .Y(ecc_byp_ecc_result_m[2]));
XOR2X1 exu_ecc_U44(.A(exu_n15112), .B(exu_n15163), .Y(ecc_byp_ecc_result_m[30]));
XOR2X1 exu_ecc_U43(.A(exu_n15111), .B(exu_n15162), .Y(ecc_byp_ecc_result_m[31]));
XOR2X1 exu_ecc_U42(.A(exu_n15110), .B(exu_n15161), .Y(ecc_byp_ecc_result_m[32]));
XOR2X1 exu_ecc_U41(.A(exu_n15109), .B(exu_n15160), .Y(ecc_byp_ecc_result_m[33]));
XOR2X1 exu_ecc_U40(.A(exu_n15108), .B(exu_n15159), .Y(ecc_byp_ecc_result_m[34]));
XOR2X1 exu_ecc_U39(.A(exu_n15107), .B(exu_n15158), .Y(ecc_byp_ecc_result_m[35]));
XOR2X1 exu_ecc_U38(.A(exu_n15106), .B(exu_n15157), .Y(ecc_byp_ecc_result_m[36]));
XOR2X1 exu_ecc_U37(.A(exu_n15105), .B(exu_n15156), .Y(ecc_byp_ecc_result_m[37]));
XOR2X1 exu_ecc_U36(.A(exu_n15104), .B(exu_n15155), .Y(ecc_byp_ecc_result_m[38]));
XOR2X1 exu_ecc_U35(.A(exu_n15103), .B(exu_n15154), .Y(ecc_byp_ecc_result_m[39]));
XOR2X1 exu_ecc_U34(.A(ecc_error_data_m[3]), .B(exu_n15153), .Y(ecc_byp_ecc_result_m[3]));
XOR2X1 exu_ecc_U33(.A(exu_n15102), .B(exu_n15152), .Y(ecc_byp_ecc_result_m[40]));
XOR2X1 exu_ecc_U32(.A(exu_n15101), .B(exu_n15151), .Y(ecc_byp_ecc_result_m[41]));
XOR2X1 exu_ecc_U31(.A(exu_n15100), .B(exu_n15150), .Y(ecc_byp_ecc_result_m[42]));
XOR2X1 exu_ecc_U30(.A(exu_n15099), .B(exu_n15149), .Y(ecc_byp_ecc_result_m[43]));
XOR2X1 exu_ecc_U29(.A(exu_n15098), .B(exu_n15148), .Y(ecc_byp_ecc_result_m[44]));
XOR2X1 exu_ecc_U28(.A(exu_n15097), .B(exu_n15147), .Y(ecc_byp_ecc_result_m[45]));
XOR2X1 exu_ecc_U27(.A(exu_n15096), .B(exu_n15146), .Y(ecc_byp_ecc_result_m[46]));
XOR2X1 exu_ecc_U26(.A(exu_n15095), .B(exu_n15145), .Y(ecc_byp_ecc_result_m[47]));
XOR2X1 exu_ecc_U25(.A(exu_n15094), .B(exu_n15144), .Y(ecc_byp_ecc_result_m[48]));
XOR2X1 exu_ecc_U24(.A(exu_n15093), .B(exu_n15143), .Y(ecc_byp_ecc_result_m[49]));
XOR2X1 exu_ecc_U23(.A(exu_n15092), .B(exu_n15142), .Y(ecc_byp_ecc_result_m[4]));
XOR2X1 exu_ecc_U22(.A(exu_n15091), .B(exu_n15141), .Y(ecc_byp_ecc_result_m[50]));
XOR2X1 exu_ecc_U21(.A(exu_n15090), .B(exu_n15140), .Y(ecc_byp_ecc_result_m[51]));
XOR2X1 exu_ecc_U20(.A(exu_n15089), .B(exu_n15139), .Y(ecc_byp_ecc_result_m[52]));
XOR2X1 exu_ecc_U19(.A(exu_n15088), .B(exu_n15138), .Y(ecc_byp_ecc_result_m[53]));
XOR2X1 exu_ecc_U18(.A(exu_n15087), .B(exu_n15137), .Y(ecc_byp_ecc_result_m[54]));
XOR2X1 exu_ecc_U17(.A(exu_n15086), .B(exu_n15136), .Y(ecc_byp_ecc_result_m[55]));
XOR2X1 exu_ecc_U16(.A(exu_n15085), .B(exu_n15135), .Y(ecc_byp_ecc_result_m[56]));
XOR2X1 exu_ecc_U15(.A(exu_n15084), .B(exu_n15134), .Y(ecc_byp_ecc_result_m[57]));
XOR2X1 exu_ecc_U14(.A(exu_n15083), .B(exu_n15133), .Y(ecc_byp_ecc_result_m[58]));
XOR2X1 exu_ecc_U13(.A(exu_n15082), .B(exu_n15132), .Y(ecc_byp_ecc_result_m[59]));
XOR2X1 exu_ecc_U12(.A(ecc_error_data_m[5]), .B(exu_n15131), .Y(ecc_byp_ecc_result_m[5]));
XOR2X1 exu_ecc_U11(.A(exu_n15081), .B(exu_n15130), .Y(ecc_byp_ecc_result_m[60]));
XOR2X1 exu_ecc_U10(.A(exu_n15080), .B(exu_n15129), .Y(ecc_byp_ecc_result_m[61]));
XOR2X1 exu_ecc_U9(.A(exu_n15079), .B(exu_n15128), .Y(ecc_byp_ecc_result_m[62]));
XOR2X1 exu_ecc_U8(.A(exu_n15078), .B(exu_n15127), .Y(ecc_byp_ecc_result_m[63]));
XOR2X1 exu_ecc_U7(.A(ecc_error_data_m[6]), .B(exu_n15126), .Y(ecc_byp_ecc_result_m[6]));
XOR2X1 exu_ecc_U6(.A(ecc_error_data_m[7]), .B(exu_n15125), .Y(ecc_byp_ecc_result_m[7]));
XOR2X1 exu_ecc_U5(.A(ecc_error_data_m[8]), .B(exu_n15124), .Y(ecc_byp_ecc_result_m[8]));
XOR2X1 exu_ecc_U4(.A(ecc_error_data_m[9]), .B(exu_n15123), .Y(ecc_byp_ecc_result_m[9]));
XOR2X1 exu_ecl_U252(.A(ecl_sub_e), .B(exu_n15795), .Y(ecl_n145));
XNOR2X1 exu_ecl_U244(.A(ecl_sub_e), .B(alu_addsub_cout64_e), .Y(ecl_n135));
XOR2X1 exu_ecl_U192(.A(div_input_data_e[64]), .B(alu_logic_rs1_data_bf1[0]), .Y(ecl_rml_xor_data_e[0]));
XOR2X1 exu_ecl_U191(.A(div_input_data_e[65]), .B(alu_logic_rs1_data_bf1[1]), .Y(ecl_rml_xor_data_e[1]));
XOR2X1 exu_ecl_U190(.A(div_input_data_e[66]), .B(alu_logic_rs1_data_bf1[2]), .Y(ecl_rml_xor_data_e[2]));
NOR2X1 exu_ecl_U181(.A(exu_tlu_ue_trap_m), .B(exu_n16403), .Y(exu_tlu_ttype_m[7]));
XOR2X1 exu_ecl_U177(.A(ecl_tid_w[1]), .B(ecl_tid_m[1]), .Y(ecl_n91));
XOR2X1 exu_ecl_U176(.A(exu_n16577), .B(ecl_tid_w[0]), .Y(ecl_n93));
XOR2X1 exu_ecl_U161(.A(lsu_exu_thr_m[1]), .B(ifu_exu_tid_s2[1]), .Y(ecl_n79));
XOR2X1 exu_ecl_U160(.A(lsu_exu_thr_m[0]), .B(ifu_exu_tid_s2[0]), .Y(ecl_n80));
XNOR2X1 exu_ecl_U155(.A(ifu_exu_invert_d), .B(exu_n15122), .Y(ecl_c_used_dff_din[0]));
XOR2X1 exu_ecl_U154(.A(ecl_tid_w[1]), .B(ecl_tid_e[1]), .Y(ecl_n74));
XOR2X1 exu_ecl_U153(.A(ecl_tid_w[0]), .B(ecl_tid_e[0]), .Y(ecl_n75));
XOR2X1 exu_ecl_U151(.A(ecl_tid_e[1]), .B(ifu_exu_tid_s2[1]), .Y(ecl_n72));
XOR2X1 exu_ecl_U150(.A(ecl_tid_e[0]), .B(ifu_exu_tid_s2[0]), .Y(ecl_n73));
XOR2X1 exu_ecl_U148(.A(ecl_tid_d[1]), .B(ifu_exu_tid_s2[1]), .Y(ecl_n70));
XOR2X1 exu_ecl_U147(.A(ecl_tid_d[0]), .B(ifu_exu_tid_s2[0]), .Y(ecl_n71));
XNOR2X1 exu_ecl_U145(.A(ecl_cc_e_3), .B(ecl_cc_e_1), .Y(ecl_div_muls_rs1_31_e_l));
XOR2X1 exu_ecl_U141(.A(ecl_ld_tid_g[1]), .B(ifu_exu_tid_s2[1]), .Y(ecl_n65));
XOR2X1 exu_ecl_U140(.A(ecl_ld_tid_g[0]), .B(ifu_exu_tid_s2[0]), .Y(ecl_n66));
XNOR2X1 exu_ecl_U112(.A(ecl_rd_e[4]), .B(exu_n15121), .Y(ecl_real_rd_e[4]));
XNOR2X1 exu_div_U290(.A(exu_n16591), .B(div_x[0]), .Y(div_adderin2[0]));
XNOR2X1 exu_div_U289(.A(exu_n16591), .B(div_x[10]), .Y(div_adderin2[10]));
XNOR2X1 exu_div_U288(.A(exu_n16591), .B(div_x[11]), .Y(div_adderin2[11]));
XNOR2X1 exu_div_U287(.A(exu_n16591), .B(div_x[12]), .Y(div_adderin2[12]));
XNOR2X1 exu_div_U286(.A(exu_n15987), .B(div_x[13]), .Y(div_adderin2[13]));
XNOR2X1 exu_div_U285(.A(exu_n16591), .B(div_x[14]), .Y(div_adderin2[14]));
XNOR2X1 exu_div_U284(.A(exu_n15987), .B(div_x[15]), .Y(div_adderin2[15]));
XNOR2X1 exu_div_U283(.A(exu_n16591), .B(div_x[16]), .Y(div_adderin2[16]));
XNOR2X1 exu_div_U282(.A(exu_n15987), .B(div_x[17]), .Y(div_adderin2[17]));
XNOR2X1 exu_div_U281(.A(exu_n16591), .B(div_x[18]), .Y(div_adderin2[18]));
XNOR2X1 exu_div_U280(.A(exu_n15987), .B(div_x[19]), .Y(div_adderin2[19]));
XNOR2X1 exu_div_U279(.A(exu_n16591), .B(div_x[1]), .Y(div_adderin2[1]));
XNOR2X1 exu_div_U278(.A(exu_n15987), .B(div_x[20]), .Y(div_adderin2[20]));
XNOR2X1 exu_div_U277(.A(exu_n16591), .B(div_x[21]), .Y(div_adderin2[21]));
XNOR2X1 exu_div_U276(.A(exu_n15987), .B(div_x[22]), .Y(div_adderin2[22]));
XNOR2X1 exu_div_U275(.A(exu_n16591), .B(div_x[23]), .Y(div_adderin2[23]));
XNOR2X1 exu_div_U274(.A(exu_n15987), .B(div_x[24]), .Y(div_adderin2[24]));
XNOR2X1 exu_div_U273(.A(exu_n15987), .B(div_x[25]), .Y(div_adderin2[25]));
XNOR2X1 exu_div_U272(.A(exu_n15987), .B(div_x[26]), .Y(div_adderin2[26]));
XNOR2X1 exu_div_U271(.A(exu_n15987), .B(div_x[27]), .Y(div_adderin2[27]));
XNOR2X1 exu_div_U270(.A(exu_n15987), .B(div_x[28]), .Y(div_adderin2[28]));
XNOR2X1 exu_div_U269(.A(exu_n15987), .B(div_x[29]), .Y(div_adderin2[29]));
XNOR2X1 exu_div_U268(.A(exu_n15987), .B(div_x[2]), .Y(div_adderin2[2]));
XNOR2X1 exu_div_U267(.A(exu_n15987), .B(div_x[30]), .Y(div_adderin2[30]));
XNOR2X1 exu_div_U266(.A(exu_n15987), .B(div_x[31]), .Y(div_adderin2[31]));
XNOR2X1 exu_div_U265(.A(exu_n15987), .B(div_x[32]), .Y(div_adderin2[32]));
XNOR2X1 exu_div_U264(.A(exu_n15987), .B(div_x[33]), .Y(div_adderin2[33]));
XNOR2X1 exu_div_U263(.A(exu_n15987), .B(div_x[34]), .Y(div_adderin2[34]));
XNOR2X1 exu_div_U262(.A(exu_n16591), .B(div_x[35]), .Y(div_adderin2[35]));
XNOR2X1 exu_div_U261(.A(exu_n16591), .B(div_x[36]), .Y(div_adderin2[36]));
XNOR2X1 exu_div_U260(.A(exu_n16591), .B(div_x[37]), .Y(div_adderin2[37]));
XNOR2X1 exu_div_U259(.A(exu_n16591), .B(div_x[38]), .Y(div_adderin2[38]));
XNOR2X1 exu_div_U258(.A(exu_n16591), .B(div_x[39]), .Y(div_adderin2[39]));
XNOR2X1 exu_div_U257(.A(exu_n16591), .B(div_x[3]), .Y(div_adderin2[3]));
XNOR2X1 exu_div_U256(.A(exu_n15987), .B(div_x[40]), .Y(div_adderin2[40]));
XNOR2X1 exu_div_U255(.A(exu_n16591), .B(div_x[41]), .Y(div_adderin2[41]));
XNOR2X1 exu_div_U254(.A(exu_n16591), .B(div_x[42]), .Y(div_adderin2[42]));
XNOR2X1 exu_div_U253(.A(exu_n16591), .B(div_x[43]), .Y(div_adderin2[43]));
XNOR2X1 exu_div_U252(.A(exu_n16591), .B(div_x[44]), .Y(div_adderin2[44]));
XNOR2X1 exu_div_U251(.A(exu_n15987), .B(div_x[45]), .Y(div_adderin2[45]));
XNOR2X1 exu_div_U250(.A(exu_n16591), .B(div_x[46]), .Y(div_adderin2[46]));
XNOR2X1 exu_div_U249(.A(exu_n15987), .B(div_x[47]), .Y(div_adderin2[47]));
XNOR2X1 exu_div_U248(.A(exu_n16591), .B(div_x[48]), .Y(div_adderin2[48]));
XNOR2X1 exu_div_U247(.A(exu_n16591), .B(div_x[49]), .Y(div_adderin2[49]));
XNOR2X1 exu_div_U246(.A(exu_n16591), .B(div_x[4]), .Y(div_adderin2[4]));
XNOR2X1 exu_div_U245(.A(exu_n15987), .B(div_x[50]), .Y(div_adderin2[50]));
XNOR2X1 exu_div_U244(.A(exu_n15987), .B(div_x[51]), .Y(div_adderin2[51]));
XNOR2X1 exu_div_U243(.A(exu_n16591), .B(div_x[52]), .Y(div_adderin2[52]));
XNOR2X1 exu_div_U242(.A(exu_n15987), .B(div_x[53]), .Y(div_adderin2[53]));
XNOR2X1 exu_div_U241(.A(exu_n15987), .B(div_x[54]), .Y(div_adderin2[54]));
XNOR2X1 exu_div_U240(.A(exu_n15987), .B(div_x[55]), .Y(div_adderin2[55]));
XNOR2X1 exu_div_U239(.A(exu_n16591), .B(div_x[56]), .Y(div_adderin2[56]));
XNOR2X1 exu_div_U238(.A(exu_n15987), .B(div_x[57]), .Y(div_adderin2[57]));
XNOR2X1 exu_div_U237(.A(exu_n15987), .B(div_x[58]), .Y(div_adderin2[58]));
XNOR2X1 exu_div_U236(.A(exu_n16591), .B(div_x[59]), .Y(div_adderin2[59]));
XNOR2X1 exu_div_U235(.A(exu_n16591), .B(div_x[5]), .Y(div_adderin2[5]));
XNOR2X1 exu_div_U234(.A(exu_n15987), .B(div_x[60]), .Y(div_adderin2[60]));
XNOR2X1 exu_div_U233(.A(exu_n16591), .B(div_x[61]), .Y(div_adderin2[61]));
XNOR2X1 exu_div_U232(.A(exu_n15987), .B(div_x[62]), .Y(div_adderin2[62]));
XNOR2X1 exu_div_U231(.A(exu_n15987), .B(div_ecl_x_msb), .Y(div_adderin2[63]));
XNOR2X1 exu_div_U230(.A(exu_n16591), .B(div_x[6]), .Y(div_adderin2[6]));
XNOR2X1 exu_div_U229(.A(exu_n16591), .B(div_x[7]), .Y(div_adderin2[7]));
XNOR2X1 exu_div_U228(.A(exu_n15987), .B(div_x[8]), .Y(div_adderin2[8]));
XNOR2X1 exu_div_U227(.A(exu_n16591), .B(div_x[9]), .Y(div_adderin2[9]));
XOR2X1 exu_rml_U174(.A(rml_rml_ecl_cleanwin_e[1]), .B(rml_rml_ecl_canrestore_e[1]), .Y(rml_n122));
XOR2X1 exu_rml_U173(.A(rml_rml_ecl_cleanwin_e[0]), .B(rml_rml_ecl_canrestore_e[0]), .Y(rml_n123));
XOR2X1 exu_rml_U171(.A(rml_rml_ecl_cleanwin_e[2]), .B(rml_rml_ecl_canrestore_e[2]), .Y(rml_n117));
XOR2X1 exu_rml_U106(.A(exu_n15548), .B(exu_n15553), .Y(rml_irf_new_e_cwp_e[0]));
XNOR2X1 exu_rml_U104(.A(exu_n15392), .B(exu_n15120), .Y(rml_irf_new_e_cwp_e[1]));
XOR2X1 exu_rml_U103(.A(exu_n15547), .B(exu_n15857), .Y(rml_irf_old_e_cwp_e[0]));
XNOR2X1 exu_rml_U101(.A(exu_n15391), .B(exu_n15119), .Y(rml_irf_old_e_cwp_e[1]));
NAND2X1 exu_rml_U97(.A(exu_n11854), .B(exu_n10686), .Y(rml_irf_swap_even_e));
NAND2X1 exu_rml_U93(.A(exu_n11853), .B(exu_n10685), .Y(rml_irf_swap_odd_e));
XOR2X1 exu_rml_U92(.A(rml_rml_ecl_cleanwin_e[1]), .B(rml_rml_ecl_cleanwin_e[0]), .Y(rml_rml_next_cleanwin_e[1]));
XOR2X1 exu_rml_U89(.A(exu_n16587), .B(rml_rml_ecl_otherwin_e[1]), .Y(rml_rml_next_otherwin_e[1]));
XOR2X1 exu_rml_U88(.A(rml_rml_ecl_cwp_e[0]), .B(rml_rml_ecl_cansave_e[0]), .Y(rml_spill_cwp_e[0]));
XOR2X1 exu_rml_U86(.A(rml_rml_ecl_cwp_e[1]), .B(rml_rml_ecl_cansave_e[1]), .Y(rml_n43));
XOR2X1 exu_rml_U85(.A(exu_n15683), .B(rml_n43), .Y(rml_spill_cwp_e[1]));
XNOR2X1 exu_rml_U79(.A(rml_rml_ecl_cansave_e[2]), .B(rml_rml_ecl_cwp_e[2]), .Y(rml_n37));
XOR2X1 exu_rml_U78(.A(exu_n15117), .B(rml_n37), .Y(rml_spill_cwp_e[2]));
AND2X2 exu_bypass_irf_write_clkbuf_U2(.A(bypass_irf_write_clkbuf_clken), .B(rclk), .Y(bypass_sehold_clk));
LATCH bypass_irf_write_clkbuf_clken_reg(.D(exu_n2), .CLK(bypass_irf_write_clkbuf_n1), .Q(bypass_irf_write_clkbuf_clken));
DFFPOSX1 bypass_dfill_data_dff_q_reg[0](.D(bypass_dfill_data_dff_n89), .CLK(rclk), .Q(bypass_dfill_data_g2[0]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[1](.D(bypass_dfill_data_dff_n67), .CLK(rclk), .Q(bypass_dfill_data_g2[1]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[2](.D(bypass_dfill_data_dff_n45), .CLK(rclk), .Q(bypass_dfill_data_g2[2]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[3](.D(bypass_dfill_data_dff_n23), .CLK(rclk), .Q(bypass_dfill_data_g2[3]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[4](.D(bypass_dfill_data_dff_n7), .CLK(rclk), .Q(bypass_dfill_data_g2[4]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[5](.D(bypass_dfill_data_dff_n5), .CLK(rclk), .Q(bypass_dfill_data_g2[5]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[6](.D(bypass_dfill_data_dff_n3), .CLK(rclk), .Q(bypass_dfill_data_g2[6]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[7](.D(bypass_dfill_data_dff_n129), .CLK(rclk), .Q(bypass_dfill_data_g2[7]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[8](.D(bypass_dfill_data_dff_n127), .CLK(rclk), .Q(bypass_dfill_data_g2[8]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[9](.D(bypass_dfill_data_dff_n125), .CLK(rclk), .Q(bypass_dfill_data_g2[9]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[10](.D(bypass_dfill_data_dff_n123), .CLK(rclk), .Q(bypass_dfill_data_g2[10]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[11](.D(bypass_dfill_data_dff_n121), .CLK(rclk), .Q(bypass_dfill_data_g2[11]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[12](.D(bypass_dfill_data_dff_n119), .CLK(rclk), .Q(bypass_dfill_data_g2[12]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[13](.D(bypass_dfill_data_dff_n117), .CLK(rclk), .Q(bypass_dfill_data_g2[13]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[14](.D(bypass_dfill_data_dff_n115), .CLK(rclk), .Q(bypass_dfill_data_g2[14]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[15](.D(bypass_dfill_data_dff_n113), .CLK(rclk), .Q(bypass_dfill_data_g2[15]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[16](.D(bypass_dfill_data_dff_n111), .CLK(rclk), .Q(bypass_dfill_data_g2[16]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[17](.D(bypass_dfill_data_dff_n109), .CLK(rclk), .Q(bypass_dfill_data_g2[17]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[18](.D(bypass_dfill_data_dff_n107), .CLK(rclk), .Q(bypass_dfill_data_g2[18]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[19](.D(bypass_dfill_data_dff_n105), .CLK(rclk), .Q(bypass_dfill_data_g2[19]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[20](.D(bypass_dfill_data_dff_n103), .CLK(rclk), .Q(bypass_dfill_data_g2[20]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[21](.D(bypass_dfill_data_dff_n101), .CLK(rclk), .Q(bypass_dfill_data_g2[21]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[22](.D(bypass_dfill_data_dff_n99), .CLK(rclk), .Q(bypass_dfill_data_g2[22]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[23](.D(bypass_dfill_data_dff_n97), .CLK(rclk), .Q(bypass_dfill_data_g2[23]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[24](.D(bypass_dfill_data_dff_n95), .CLK(rclk), .Q(bypass_dfill_data_g2[24]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[25](.D(bypass_dfill_data_dff_n93), .CLK(rclk), .Q(bypass_dfill_data_g2[25]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[26](.D(bypass_dfill_data_dff_n91), .CLK(rclk), .Q(bypass_dfill_data_g2[26]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[27](.D(bypass_dfill_data_dff_n87), .CLK(rclk), .Q(bypass_dfill_data_g2[27]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[28](.D(bypass_dfill_data_dff_n85), .CLK(rclk), .Q(bypass_dfill_data_g2[28]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[29](.D(bypass_dfill_data_dff_n83), .CLK(rclk), .Q(bypass_dfill_data_g2[29]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[30](.D(bypass_dfill_data_dff_n81), .CLK(rclk), .Q(bypass_dfill_data_g2[30]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[31](.D(bypass_dfill_data_dff_n79), .CLK(rclk), .Q(bypass_dfill_data_g2[31]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[32](.D(bypass_dfill_data_dff_n77), .CLK(rclk), .Q(bypass_dfill_data_g2[32]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[33](.D(bypass_dfill_data_dff_n75), .CLK(rclk), .Q(bypass_dfill_data_g2[33]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[34](.D(bypass_dfill_data_dff_n73), .CLK(rclk), .Q(bypass_dfill_data_g2[34]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[35](.D(bypass_dfill_data_dff_n71), .CLK(rclk), .Q(bypass_dfill_data_g2[35]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[36](.D(bypass_dfill_data_dff_n69), .CLK(rclk), .Q(bypass_dfill_data_g2[36]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[37](.D(bypass_dfill_data_dff_n65), .CLK(rclk), .Q(bypass_dfill_data_g2[37]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[38](.D(bypass_dfill_data_dff_n63), .CLK(rclk), .Q(bypass_dfill_data_g2[38]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[39](.D(bypass_dfill_data_dff_n61), .CLK(rclk), .Q(bypass_dfill_data_g2[39]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[40](.D(bypass_dfill_data_dff_n59), .CLK(rclk), .Q(bypass_dfill_data_g2[40]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[41](.D(bypass_dfill_data_dff_n57), .CLK(rclk), .Q(bypass_dfill_data_g2[41]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[42](.D(bypass_dfill_data_dff_n55), .CLK(rclk), .Q(bypass_dfill_data_g2[42]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[43](.D(bypass_dfill_data_dff_n53), .CLK(rclk), .Q(bypass_dfill_data_g2[43]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[44](.D(bypass_dfill_data_dff_n51), .CLK(rclk), .Q(bypass_dfill_data_g2[44]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[45](.D(bypass_dfill_data_dff_n49), .CLK(rclk), .Q(bypass_dfill_data_g2[45]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[46](.D(bypass_dfill_data_dff_n47), .CLK(rclk), .Q(bypass_dfill_data_g2[46]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[47](.D(bypass_dfill_data_dff_n43), .CLK(rclk), .Q(bypass_dfill_data_g2[47]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[48](.D(bypass_dfill_data_dff_n41), .CLK(rclk), .Q(bypass_dfill_data_g2[48]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[49](.D(bypass_dfill_data_dff_n39), .CLK(rclk), .Q(bypass_dfill_data_g2[49]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[50](.D(bypass_dfill_data_dff_n37), .CLK(rclk), .Q(bypass_dfill_data_g2[50]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[51](.D(bypass_dfill_data_dff_n35), .CLK(rclk), .Q(bypass_dfill_data_g2[51]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[52](.D(bypass_dfill_data_dff_n33), .CLK(rclk), .Q(bypass_dfill_data_g2[52]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[53](.D(bypass_dfill_data_dff_n31), .CLK(rclk), .Q(bypass_dfill_data_g2[53]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[54](.D(bypass_dfill_data_dff_n29), .CLK(rclk), .Q(bypass_dfill_data_g2[54]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[55](.D(bypass_dfill_data_dff_n27), .CLK(rclk), .Q(bypass_dfill_data_g2[55]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[56](.D(bypass_dfill_data_dff_n25), .CLK(rclk), .Q(bypass_dfill_data_g2[56]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[57](.D(bypass_dfill_data_dff_n21), .CLK(rclk), .Q(bypass_dfill_data_g2[57]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[58](.D(bypass_dfill_data_dff_n19), .CLK(rclk), .Q(bypass_dfill_data_g2[58]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[59](.D(bypass_dfill_data_dff_n17), .CLK(rclk), .Q(bypass_dfill_data_g2[59]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[60](.D(bypass_dfill_data_dff_n15), .CLK(rclk), .Q(bypass_dfill_data_g2[60]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[61](.D(bypass_dfill_data_dff_n13), .CLK(rclk), .Q(bypass_dfill_data_g2[61]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[62](.D(bypass_dfill_data_dff_n11), .CLK(rclk), .Q(bypass_dfill_data_g2[62]));
DFFPOSX1 bypass_dfill_data_dff_q_reg[63](.D(bypass_dfill_data_dff_n9), .CLK(rclk), .Q(bypass_dfill_data_g2[63]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[0](.D(bypass_rs3h_data_dff_n25), .CLK(rclk), .Q(bypass_rs3h_data_e[0]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[1](.D(bypass_rs3h_data_dff_n13), .CLK(rclk), .Q(bypass_rs3h_data_e[1]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[2](.D(bypass_rs3h_data_dff_n11), .CLK(rclk), .Q(bypass_rs3h_data_e[2]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[3](.D(bypass_rs3h_data_dff_n9), .CLK(rclk), .Q(bypass_rs3h_data_e[3]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[4](.D(bypass_rs3h_data_dff_n7), .CLK(rclk), .Q(bypass_rs3h_data_e[4]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[5](.D(bypass_rs3h_data_dff_n5), .CLK(rclk), .Q(bypass_rs3h_data_e[5]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[6](.D(bypass_rs3h_data_dff_n3), .CLK(rclk), .Q(bypass_rs3h_data_e[6]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[7](.D(bypass_rs3h_data_dff_n65), .CLK(rclk), .Q(bypass_rs3h_data_e[7]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[8](.D(bypass_rs3h_data_dff_n63), .CLK(rclk), .Q(bypass_rs3h_data_e[8]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[9](.D(bypass_rs3h_data_dff_n61), .CLK(rclk), .Q(bypass_rs3h_data_e[9]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[10](.D(bypass_rs3h_data_dff_n59), .CLK(rclk), .Q(bypass_rs3h_data_e[10]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[11](.D(bypass_rs3h_data_dff_n57), .CLK(rclk), .Q(bypass_rs3h_data_e[11]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[12](.D(bypass_rs3h_data_dff_n55), .CLK(rclk), .Q(bypass_rs3h_data_e[12]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[13](.D(bypass_rs3h_data_dff_n53), .CLK(rclk), .Q(bypass_rs3h_data_e[13]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[14](.D(bypass_rs3h_data_dff_n51), .CLK(rclk), .Q(bypass_rs3h_data_e[14]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[15](.D(bypass_rs3h_data_dff_n49), .CLK(rclk), .Q(bypass_rs3h_data_e[15]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[16](.D(bypass_rs3h_data_dff_n47), .CLK(rclk), .Q(bypass_rs3h_data_e[16]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[17](.D(bypass_rs3h_data_dff_n45), .CLK(rclk), .Q(bypass_rs3h_data_e[17]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[18](.D(bypass_rs3h_data_dff_n43), .CLK(rclk), .Q(bypass_rs3h_data_e[18]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[19](.D(bypass_rs3h_data_dff_n41), .CLK(rclk), .Q(bypass_rs3h_data_e[19]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[20](.D(bypass_rs3h_data_dff_n39), .CLK(rclk), .Q(bypass_rs3h_data_e[20]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[21](.D(bypass_rs3h_data_dff_n37), .CLK(rclk), .Q(bypass_rs3h_data_e[21]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[22](.D(bypass_rs3h_data_dff_n35), .CLK(rclk), .Q(bypass_rs3h_data_e[22]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[23](.D(bypass_rs3h_data_dff_n33), .CLK(rclk), .Q(bypass_rs3h_data_e[23]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[24](.D(bypass_rs3h_data_dff_n31), .CLK(rclk), .Q(bypass_rs3h_data_e[24]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[25](.D(bypass_rs3h_data_dff_n29), .CLK(rclk), .Q(bypass_rs3h_data_e[25]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[26](.D(bypass_rs3h_data_dff_n27), .CLK(rclk), .Q(bypass_rs3h_data_e[26]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[27](.D(bypass_rs3h_data_dff_n23), .CLK(rclk), .Q(bypass_rs3h_data_e[27]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[28](.D(bypass_rs3h_data_dff_n21), .CLK(rclk), .Q(bypass_rs3h_data_e[28]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[29](.D(bypass_rs3h_data_dff_n19), .CLK(rclk), .Q(bypass_rs3h_data_e[29]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[30](.D(bypass_rs3h_data_dff_n17), .CLK(rclk), .Q(bypass_rs3h_data_e[30]));
DFFPOSX1 bypass_rs3h_data_dff_q_reg[31](.D(bypass_rs3h_data_dff_n15), .CLK(rclk), .Q(bypass_rs3h_data_e[31]));
XOR2X1 exu_bypass_w1_eccgen_U183(.A(bypass_w1_eccgen_n2), .B(bypass_w1_eccgen_n1), .Y(bypass_rd_synd_w_l[0]));
XOR2X1 exu_bypass_w1_eccgen_U182(.A(bypass_w1_eccgen_n4), .B(bypass_w1_eccgen_n3), .Y(bypass_w1_eccgen_n1));
XOR2X1 exu_bypass_w1_eccgen_U181(.A(bypass_w1_eccgen_n6), .B(bypass_w1_eccgen_n5), .Y(bypass_w1_eccgen_n2));
XOR2X1 exu_bypass_w1_eccgen_U180(.A(bypass_w1_eccgen_p0_w[1]), .B(bypass_w1_eccgen_p0_w[0]), .Y(bypass_w1_eccgen_n3));
XOR2X1 exu_bypass_w1_eccgen_U179(.A(bypass_w1_eccgen_p0_w[3]), .B(bypass_w1_eccgen_p0_w[2]), .Y(bypass_w1_eccgen_n4));
XOR2X1 exu_bypass_w1_eccgen_U178(.A(bypass_w1_eccgen_p0_w[5]), .B(bypass_w1_eccgen_p0_w[4]), .Y(bypass_w1_eccgen_n5));
XOR2X1 exu_bypass_w1_eccgen_U177(.A(bypass_w1_eccgen_p0_w[7]), .B(bypass_w1_eccgen_p0_w[6]), .Y(bypass_w1_eccgen_n6));
XOR2X1 exu_bypass_w1_eccgen_U176(.A(bypass_w1_eccgen_n8), .B(bypass_w1_eccgen_n7), .Y(bypass_rd_synd_w_l[1]));
XOR2X1 exu_bypass_w1_eccgen_U175(.A(bypass_w1_eccgen_n10), .B(bypass_w1_eccgen_n9), .Y(bypass_w1_eccgen_n7));
XOR2X1 exu_bypass_w1_eccgen_U174(.A(bypass_w1_eccgen_n12), .B(bypass_w1_eccgen_n11), .Y(bypass_w1_eccgen_n8));
XOR2X1 exu_bypass_w1_eccgen_U173(.A(bypass_w1_eccgen_p1_w[1]), .B(bypass_w1_eccgen_p1_w[0]), .Y(bypass_w1_eccgen_n9));
XOR2X1 exu_bypass_w1_eccgen_U172(.A(bypass_w1_eccgen_p1_w[3]), .B(bypass_w1_eccgen_p1_w[2]), .Y(bypass_w1_eccgen_n10));
XOR2X1 exu_bypass_w1_eccgen_U171(.A(bypass_w1_eccgen_p1_w[5]), .B(bypass_w1_eccgen_p1_w[4]), .Y(bypass_w1_eccgen_n11));
XOR2X1 exu_bypass_w1_eccgen_U170(.A(bypass_w1_eccgen_p1_w[7]), .B(bypass_w1_eccgen_p1_w[6]), .Y(bypass_w1_eccgen_n12));
XOR2X1 exu_bypass_w1_eccgen_U169(.A(bypass_w1_eccgen_n14), .B(bypass_w1_eccgen_n13), .Y(bypass_rd_synd_w_l[2]));
XOR2X1 exu_bypass_w1_eccgen_U168(.A(bypass_w1_eccgen_n16), .B(bypass_w1_eccgen_n15), .Y(bypass_w1_eccgen_n13));
XOR2X1 exu_bypass_w1_eccgen_U167(.A(bypass_w1_eccgen_n18), .B(bypass_w1_eccgen_n17), .Y(bypass_w1_eccgen_n14));
XOR2X1 exu_bypass_w1_eccgen_U166(.A(bypass_w1_eccgen_p2_w[1]), .B(bypass_w1_eccgen_p2_w[0]), .Y(bypass_w1_eccgen_n15));
XOR2X1 exu_bypass_w1_eccgen_U165(.A(bypass_w1_eccgen_p2_w[3]), .B(bypass_w1_eccgen_p2_w[2]), .Y(bypass_w1_eccgen_n16));
XOR2X1 exu_bypass_w1_eccgen_U164(.A(bypass_w1_eccgen_p2_w[5]), .B(bypass_w1_eccgen_p2_w[4]), .Y(bypass_w1_eccgen_n17));
XOR2X1 exu_bypass_w1_eccgen_U163(.A(bypass_w1_eccgen_p2_w[7]), .B(bypass_w1_eccgen_p2_w[6]), .Y(bypass_w1_eccgen_n18));
XOR2X1 exu_bypass_w1_eccgen_U162(.A(bypass_w1_eccgen_n20), .B(bypass_w1_eccgen_n19), .Y(bypass_rd_synd_w_l[3]));
XOR2X1 exu_bypass_w1_eccgen_U161(.A(bypass_w1_eccgen_n22), .B(bypass_w1_eccgen_n21), .Y(bypass_w1_eccgen_n19));
XOR2X1 exu_bypass_w1_eccgen_U160(.A(bypass_w1_eccgen_n24), .B(bypass_w1_eccgen_n23), .Y(bypass_w1_eccgen_n20));
XOR2X1 exu_bypass_w1_eccgen_U159(.A(bypass_w1_eccgen_p3_w[1]), .B(bypass_w1_eccgen_p3_w[0]), .Y(bypass_w1_eccgen_n21));
XOR2X1 exu_bypass_w1_eccgen_U158(.A(bypass_w1_eccgen_p3_w[3]), .B(bypass_w1_eccgen_p3_w[2]), .Y(bypass_w1_eccgen_n22));
XOR2X1 exu_bypass_w1_eccgen_U157(.A(bypass_w1_eccgen_p3_w[5]), .B(bypass_w1_eccgen_p3_w[4]), .Y(bypass_w1_eccgen_n23));
XOR2X1 exu_bypass_w1_eccgen_U156(.A(bypass_w1_eccgen_p3_w[7]), .B(bypass_w1_eccgen_p3_w[6]), .Y(bypass_w1_eccgen_n24));
XOR2X1 exu_bypass_w1_eccgen_U155(.A(bypass_w1_eccgen_n26), .B(bypass_w1_eccgen_n25), .Y(bypass_rd_synd_w_l[4]));
XOR2X1 exu_bypass_w1_eccgen_U154(.A(bypass_w1_eccgen_p4_w[0]), .B(bypass_w1_eccgen_n27), .Y(bypass_w1_eccgen_n25));
XOR2X1 exu_bypass_w1_eccgen_U153(.A(bypass_w1_eccgen_p4_w[2]), .B(bypass_w1_eccgen_p4_w[1]), .Y(bypass_w1_eccgen_n26));
XOR2X1 exu_bypass_w1_eccgen_U152(.A(bypass_w1_eccgen_msk_w4), .B(bypass_w1_eccgen_p4_w[3]), .Y(bypass_w1_eccgen_n27));
XOR2X1 exu_bypass_w1_eccgen_U151(.A(bypass_w1_eccgen_n29), .B(bypass_w1_eccgen_n28), .Y(bypass_rd_synd_w_l[5]));
XOR2X1 exu_bypass_w1_eccgen_U150(.A(bypass_w1_eccgen_p5_w[0]), .B(bypass_w1_eccgen_n30), .Y(bypass_w1_eccgen_n28));
XOR2X1 exu_bypass_w1_eccgen_U149(.A(bypass_w1_eccgen_p4_w[2]), .B(bypass_w1_eccgen_p5_w[1]), .Y(bypass_w1_eccgen_n29));
XOR2X1 exu_bypass_w1_eccgen_U148(.A(bypass_w1_eccgen_msk_w5), .B(bypass_w1_eccgen_p4_w[3]), .Y(bypass_w1_eccgen_n30));
XOR2X1 exu_bypass_w1_eccgen_U147(.A(bypass_w1_eccgen_n32), .B(bypass_w1_eccgen_n31), .Y(bypass_rd_synd_w_l[7]));
XOR2X1 exu_bypass_w1_eccgen_U146(.A(bypass_w1_eccgen_n34), .B(bypass_w1_eccgen_n33), .Y(bypass_w1_eccgen_n31));
XOR2X1 exu_bypass_w1_eccgen_U145(.A(bypass_w1_eccgen_n36), .B(bypass_w1_eccgen_n35), .Y(bypass_w1_eccgen_n32));
XOR2X1 exu_bypass_w1_eccgen_U144(.A(bypass_w1_eccgen_p7_w[1]), .B(bypass_w1_eccgen_p7_w[0]), .Y(bypass_w1_eccgen_n33));
XOR2X1 exu_bypass_w1_eccgen_U143(.A(bypass_w1_eccgen_p7_w[3]), .B(bypass_w1_eccgen_p7_w[2]), .Y(bypass_w1_eccgen_n34));
XOR2X1 exu_bypass_w1_eccgen_U142(.A(bypass_w1_eccgen_p7_w[5]), .B(bypass_w1_eccgen_p7_w[4]), .Y(bypass_w1_eccgen_n35));
XOR2X1 exu_bypass_w1_eccgen_U141(.A(bypass_w1_eccgen_p7_w[7]), .B(bypass_w1_eccgen_p7_w[6]), .Y(bypass_w1_eccgen_n36));
XOR2X1 exu_bypass_w1_eccgen_U140(.A(bypass_byp_irf_rd_data_m[0]), .B(bypass_w1_eccgen_n37), .Y(bypass_w1_eccgen_n124));
XOR2X1 exu_bypass_w1_eccgen_U139(.A(bypass_byp_irf_rd_data_m[4]), .B(bypass_byp_irf_rd_data_m[1]), .Y(bypass_w1_eccgen_n37));
XOR2X1 exu_bypass_w1_eccgen_U138(.A(bypass_byp_irf_rd_data_m[2]), .B(bypass_w1_eccgen_n124), .Y(bypass_w1_eccgen_p7_g[0]));
XOR2X1 exu_bypass_w1_eccgen_U137(.A(bypass_w1_eccgen_n39), .B(bypass_w1_eccgen_n38), .Y(bypass_w1_eccgen_p7_g[1]));
XOR2X1 exu_bypass_w1_eccgen_U136(.A(bypass_byp_irf_rd_data_m[7]), .B(bypass_byp_irf_rd_data_m[5]), .Y(bypass_w1_eccgen_n38));
XOR2X1 exu_bypass_w1_eccgen_U135(.A(bypass_byp_irf_rd_data_m[11]), .B(bypass_byp_irf_rd_data_m[10]), .Y(bypass_w1_eccgen_n39));
XOR2X1 exu_bypass_w1_eccgen_U134(.A(bypass_w1_eccgen_n41), .B(bypass_w1_eccgen_n40), .Y(bypass_w1_eccgen_p7_g[2]));
XOR2X1 exu_bypass_w1_eccgen_U133(.A(bypass_byp_irf_rd_data_m[14]), .B(bypass_byp_irf_rd_data_m[12]), .Y(bypass_w1_eccgen_n40));
XOR2X1 exu_bypass_w1_eccgen_U132(.A(bypass_byp_irf_rd_data_m[18]), .B(bypass_byp_irf_rd_data_m[17]), .Y(bypass_w1_eccgen_n41));
XOR2X1 exu_bypass_w1_eccgen_U131(.A(bypass_byp_irf_rd_data_m[21]), .B(bypass_w1_eccgen_n42), .Y(bypass_w1_eccgen_n125));
XOR2X1 exu_bypass_w1_eccgen_U130(.A(bypass_byp_irf_rd_data_m[26]), .B(bypass_byp_irf_rd_data_m[23]), .Y(bypass_w1_eccgen_n42));
XOR2X1 exu_bypass_w1_eccgen_U129(.A(bypass_byp_irf_rd_data_m[24]), .B(bypass_w1_eccgen_n125), .Y(bypass_w1_eccgen_p7_g[3]));
XOR2X1 exu_bypass_w1_eccgen_U128(.A(bypass_w1_eccgen_n44), .B(bypass_w1_eccgen_n43), .Y(bypass_w1_eccgen_p7_g[4]));
XOR2X1 exu_bypass_w1_eccgen_U127(.A(bypass_byp_irf_rd_data_m[29]), .B(bypass_byp_irf_rd_data_m[27]), .Y(bypass_w1_eccgen_n43));
XOR2X1 exu_bypass_w1_eccgen_U126(.A(bypass_byp_irf_rd_data_m[33]), .B(bypass_byp_irf_rd_data_m[32]), .Y(bypass_w1_eccgen_n44));
XOR2X1 exu_bypass_w1_eccgen_U125(.A(bypass_w1_eccgen_n46), .B(bypass_w1_eccgen_n45), .Y(bypass_w1_eccgen_p7_g[5]));
XOR2X1 exu_bypass_w1_eccgen_U124(.A(bypass_byp_irf_rd_data_m[38]), .B(bypass_byp_irf_rd_data_m[36]), .Y(bypass_w1_eccgen_n45));
XOR2X1 exu_bypass_w1_eccgen_U123(.A(bypass_byp_irf_rd_data_m[41]), .B(bypass_byp_irf_rd_data_m[39]), .Y(bypass_w1_eccgen_n46));
XOR2X1 exu_bypass_w1_eccgen_U122(.A(bypass_byp_irf_rd_data_m[44]), .B(bypass_w1_eccgen_n47), .Y(bypass_w1_eccgen_n126));
XOR2X1 exu_bypass_w1_eccgen_U121(.A(bypass_byp_irf_rd_data_m[50]), .B(bypass_byp_irf_rd_data_m[46]), .Y(bypass_w1_eccgen_n47));
XOR2X1 exu_bypass_w1_eccgen_U120(.A(bypass_byp_irf_rd_data_m[47]), .B(bypass_w1_eccgen_n126), .Y(bypass_w1_eccgen_p7_g[6]));
XOR2X1 exu_bypass_w1_eccgen_U119(.A(bypass_byp_irf_rd_data_m[57]), .B(bypass_w1_eccgen_n48), .Y(bypass_w1_eccgen_n117));
XOR2X1 exu_bypass_w1_eccgen_U118(.A(bypass_byp_irf_rd_data_m[60]), .B(bypass_byp_irf_rd_data_m[58]), .Y(bypass_w1_eccgen_n48));
XOR2X1 exu_bypass_w1_eccgen_U117(.A(bypass_w1_eccgen_n50), .B(bypass_w1_eccgen_n49), .Y(bypass_w1_eccgen_p7_g[7]));
XOR2X1 exu_bypass_w1_eccgen_U116(.A(bypass_w1_eccgen_n52), .B(bypass_w1_eccgen_n51), .Y(bypass_w1_eccgen_n49));
XOR2X1 exu_bypass_w1_eccgen_U115(.A(exu_n15513), .B(bypass_w1_eccgen_n117), .Y(bypass_w1_eccgen_n50));
XOR2X1 exu_bypass_w1_eccgen_U114(.A(bypass_byp_irf_rd_data_m[53]), .B(bypass_byp_irf_rd_data_m[51]), .Y(bypass_w1_eccgen_n51));
XOR2X1 exu_bypass_w1_eccgen_U113(.A(bypass_byp_irf_rd_data_m[63]), .B(bypass_byp_irf_rd_data_m[56]), .Y(bypass_w1_eccgen_n52));
XOR2X1 exu_bypass_w1_eccgen_U112(.A(bypass_byp_irf_rd_data_m[59]), .B(bypass_w1_eccgen_n117), .Y(bypass_w1_eccgen_p6_g[0]));
XOR2X1 exu_bypass_w1_eccgen_U111(.A(bypass_byp_irf_rd_data_m[61]), .B(bypass_w1_eccgen_n53), .Y(bypass_w1_eccgen_n120));
XOR2X1 exu_bypass_w1_eccgen_U110(.A(bypass_byp_irf_rd_data_m[63]), .B(bypass_byp_irf_rd_data_m[62]), .Y(bypass_w1_eccgen_n53));
XOR2X1 exu_bypass_w1_eccgen_U109(.A(exu_n15514), .B(bypass_w1_eccgen_n120), .Y(bypass_w1_eccgen_p6_g[1]));
XOR2X1 exu_bypass_w1_eccgen_U108(.A(bypass_w1_eccgen_n55), .B(bypass_w1_eccgen_n54), .Y(bypass_w1_eccgen_p5_g[0]));
XOR2X1 exu_bypass_w1_eccgen_U107(.A(bypass_w1_eccgen_p7_g[4]), .B(bypass_w1_eccgen_n56), .Y(bypass_w1_eccgen_n54));
XOR2X1 exu_bypass_w1_eccgen_U106(.A(bypass_byp_irf_rd_data_m[28]), .B(bypass_byp_irf_rd_data_m[26]), .Y(bypass_w1_eccgen_n55));
XOR2X1 exu_bypass_w1_eccgen_U105(.A(bypass_byp_irf_rd_data_m[31]), .B(bypass_byp_irf_rd_data_m[30]), .Y(bypass_w1_eccgen_n56));
XOR2X1 exu_bypass_w1_eccgen_U104(.A(bypass_w1_eccgen_n58), .B(bypass_w1_eccgen_n57), .Y(bypass_w1_eccgen_p3_g[4]));
XOR2X1 exu_bypass_w1_eccgen_U103(.A(bypass_byp_irf_rd_data_m[35]), .B(bypass_byp_irf_rd_data_m[34]), .Y(bypass_w1_eccgen_n57));
XOR2X1 exu_bypass_w1_eccgen_U102(.A(bypass_byp_irf_rd_data_m[37]), .B(bypass_byp_irf_rd_data_m[36]), .Y(bypass_w1_eccgen_n58));
XOR2X1 exu_bypass_w1_eccgen_U101(.A(bypass_byp_irf_rd_data_m[38]), .B(bypass_w1_eccgen_n59), .Y(bypass_w1_eccgen_n119));
XOR2X1 exu_bypass_w1_eccgen_U100(.A(bypass_byp_irf_rd_data_m[40]), .B(bypass_byp_irf_rd_data_m[39]), .Y(bypass_w1_eccgen_n59));
XOR2X1 exu_bypass_w1_eccgen_U99(.A(bypass_w1_eccgen_n119), .B(bypass_w1_eccgen_n60), .Y(bypass_w1_eccgen_p5_g[1]));
XOR2X1 exu_bypass_w1_eccgen_U98(.A(bypass_byp_irf_rd_data_m[41]), .B(bypass_w1_eccgen_p3_g[4]), .Y(bypass_w1_eccgen_n60));
XOR2X1 exu_bypass_w1_eccgen_U97(.A(bypass_w1_eccgen_n62), .B(bypass_w1_eccgen_n61), .Y(bypass_w1_eccgen_p4_g[0]));
XOR2X1 exu_bypass_w1_eccgen_U96(.A(bypass_w1_eccgen_p7_g[2]), .B(bypass_w1_eccgen_n63), .Y(bypass_w1_eccgen_n61));
XOR2X1 exu_bypass_w1_eccgen_U95(.A(bypass_byp_irf_rd_data_m[13]), .B(bypass_byp_irf_rd_data_m[11]), .Y(bypass_w1_eccgen_n62));
XOR2X1 exu_bypass_w1_eccgen_U94(.A(bypass_byp_irf_rd_data_m[16]), .B(bypass_byp_irf_rd_data_m[15]), .Y(bypass_w1_eccgen_n63));
XOR2X1 exu_bypass_w1_eccgen_U93(.A(bypass_w1_eccgen_n65), .B(bypass_w1_eccgen_n64), .Y(bypass_w1_eccgen_p3_g[2]));
XOR2X1 exu_bypass_w1_eccgen_U92(.A(bypass_byp_irf_rd_data_m[20]), .B(bypass_byp_irf_rd_data_m[19]), .Y(bypass_w1_eccgen_n64));
XOR2X1 exu_bypass_w1_eccgen_U91(.A(bypass_byp_irf_rd_data_m[22]), .B(bypass_byp_irf_rd_data_m[21]), .Y(bypass_w1_eccgen_n65));
XOR2X1 exu_bypass_w1_eccgen_U90(.A(bypass_byp_irf_rd_data_m[23]), .B(bypass_w1_eccgen_n66), .Y(bypass_w1_eccgen_n118));
XOR2X1 exu_bypass_w1_eccgen_U89(.A(bypass_byp_irf_rd_data_m[25]), .B(bypass_byp_irf_rd_data_m[24]), .Y(bypass_w1_eccgen_n66));
XOR2X1 exu_bypass_w1_eccgen_U88(.A(bypass_w1_eccgen_n118), .B(bypass_w1_eccgen_n67), .Y(bypass_w1_eccgen_p4_g[1]));
XOR2X1 exu_bypass_w1_eccgen_U87(.A(bypass_byp_irf_rd_data_m[41]), .B(bypass_w1_eccgen_p3_g[2]), .Y(bypass_w1_eccgen_n67));
XOR2X1 exu_bypass_w1_eccgen_U86(.A(bypass_byp_irf_rd_data_m[48]), .B(bypass_byp_irf_rd_data_m[47]), .Y(bypass_w1_eccgen_n123));
XOR2X1 exu_bypass_w1_eccgen_U85(.A(bypass_w1_eccgen_n69), .B(bypass_w1_eccgen_n68), .Y(bypass_w1_eccgen_p4_g[2]));
XOR2X1 exu_bypass_w1_eccgen_U84(.A(bypass_w1_eccgen_n71), .B(bypass_w1_eccgen_n70), .Y(bypass_w1_eccgen_n68));
XOR2X1 exu_bypass_w1_eccgen_U83(.A(bypass_w1_eccgen_n123), .B(bypass_w1_eccgen_n72), .Y(bypass_w1_eccgen_n69));
XOR2X1 exu_bypass_w1_eccgen_U82(.A(bypass_byp_irf_rd_data_m[43]), .B(bypass_byp_irf_rd_data_m[42]), .Y(bypass_w1_eccgen_n70));
XOR2X1 exu_bypass_w1_eccgen_U81(.A(bypass_byp_irf_rd_data_m[45]), .B(bypass_byp_irf_rd_data_m[44]), .Y(bypass_w1_eccgen_n71));
XOR2X1 exu_bypass_w1_eccgen_U80(.A(bypass_byp_irf_rd_data_m[49]), .B(bypass_byp_irf_rd_data_m[46]), .Y(bypass_w1_eccgen_n72));
XOR2X1 exu_bypass_w1_eccgen_U79(.A(bypass_w1_eccgen_n74), .B(bypass_w1_eccgen_n73), .Y(bypass_w1_eccgen_p3_g[6]));
XOR2X1 exu_bypass_w1_eccgen_U78(.A(bypass_byp_irf_rd_data_m[51]), .B(bypass_byp_irf_rd_data_m[50]), .Y(bypass_w1_eccgen_n73));
XOR2X1 exu_bypass_w1_eccgen_U77(.A(bypass_byp_irf_rd_data_m[53]), .B(bypass_byp_irf_rd_data_m[52]), .Y(bypass_w1_eccgen_n74));
XOR2X1 exu_bypass_w1_eccgen_U76(.A(bypass_byp_irf_rd_data_m[54]), .B(bypass_w1_eccgen_n75), .Y(bypass_w1_eccgen_n121));
XOR2X1 exu_bypass_w1_eccgen_U75(.A(bypass_byp_irf_rd_data_m[56]), .B(bypass_byp_irf_rd_data_m[55]), .Y(bypass_w1_eccgen_n75));
XOR2X1 exu_bypass_w1_eccgen_U74(.A(bypass_w1_eccgen_p3_g[6]), .B(bypass_w1_eccgen_n121), .Y(bypass_w1_eccgen_p4_g[3]));
XOR2X1 exu_bypass_w1_eccgen_U73(.A(bypass_w1_eccgen_n77), .B(bypass_w1_eccgen_n76), .Y(bypass_w1_eccgen_p3_g[0]));
XOR2X1 exu_bypass_w1_eccgen_U72(.A(bypass_byp_irf_rd_data_m[5]), .B(bypass_byp_irf_rd_data_m[4]), .Y(bypass_w1_eccgen_n76));
XOR2X1 exu_bypass_w1_eccgen_U71(.A(bypass_byp_irf_rd_data_m[7]), .B(bypass_byp_irf_rd_data_m[6]), .Y(bypass_w1_eccgen_n77));
XOR2X1 exu_bypass_w1_eccgen_U70(.A(bypass_byp_irf_rd_data_m[10]), .B(bypass_byp_irf_rd_data_m[9]), .Y(bypass_w1_eccgen_n122));
XOR2X1 exu_bypass_w1_eccgen_U69(.A(bypass_w1_eccgen_n122), .B(bypass_w1_eccgen_n78), .Y(bypass_w1_eccgen_p3_g[1]));
XOR2X1 exu_bypass_w1_eccgen_U68(.A(bypass_byp_irf_rd_data_m[18]), .B(bypass_byp_irf_rd_data_m[8]), .Y(bypass_w1_eccgen_n78));
XOR2X1 exu_bypass_w1_eccgen_U67(.A(bypass_byp_irf_rd_data_m[33]), .B(bypass_w1_eccgen_n118), .Y(bypass_w1_eccgen_p3_g[3]));
XOR2X1 exu_bypass_w1_eccgen_U66(.A(bypass_byp_irf_rd_data_m[49]), .B(bypass_w1_eccgen_n119), .Y(bypass_w1_eccgen_p3_g[5]));
XOR2X1 exu_bypass_w1_eccgen_U65(.A(exu_n15515), .B(bypass_w1_eccgen_n121), .Y(bypass_w1_eccgen_p3_g[7]));
XOR2X1 exu_bypass_w1_eccgen_U64(.A(bypass_w1_eccgen_n80), .B(bypass_w1_eccgen_n79), .Y(bypass_w1_eccgen_p2_g[0]));
XOR2X1 exu_bypass_w1_eccgen_U63(.A(bypass_byp_irf_rd_data_m[2]), .B(bypass_byp_irf_rd_data_m[1]), .Y(bypass_w1_eccgen_n79));
XOR2X1 exu_bypass_w1_eccgen_U62(.A(bypass_byp_irf_rd_data_m[7]), .B(bypass_byp_irf_rd_data_m[3]), .Y(bypass_w1_eccgen_n80));
XOR2X1 exu_bypass_w1_eccgen_U61(.A(bypass_w1_eccgen_n122), .B(bypass_w1_eccgen_n81), .Y(bypass_w1_eccgen_p2_g[1]));
XOR2X1 exu_bypass_w1_eccgen_U60(.A(bypass_byp_irf_rd_data_m[14]), .B(bypass_byp_irf_rd_data_m[8]), .Y(bypass_w1_eccgen_n81));
XOR2X1 exu_bypass_w1_eccgen_U59(.A(bypass_w1_eccgen_n83), .B(bypass_w1_eccgen_n82), .Y(bypass_w1_eccgen_p2_g[2]));
XOR2X1 exu_bypass_w1_eccgen_U58(.A(bypass_byp_irf_rd_data_m[16]), .B(bypass_byp_irf_rd_data_m[15]), .Y(bypass_w1_eccgen_n82));
XOR2X1 exu_bypass_w1_eccgen_U57(.A(bypass_byp_irf_rd_data_m[22]), .B(bypass_byp_irf_rd_data_m[17]), .Y(bypass_w1_eccgen_n83));
XOR2X1 exu_bypass_w1_eccgen_U56(.A(bypass_byp_irf_rd_data_m[29]), .B(bypass_w1_eccgen_n118), .Y(bypass_w1_eccgen_p2_g[3]));
XOR2X1 exu_bypass_w1_eccgen_U55(.A(bypass_w1_eccgen_n85), .B(bypass_w1_eccgen_n84), .Y(bypass_w1_eccgen_p2_g[4]));
XOR2X1 exu_bypass_w1_eccgen_U54(.A(bypass_byp_irf_rd_data_m[31]), .B(bypass_byp_irf_rd_data_m[30]), .Y(bypass_w1_eccgen_n84));
XOR2X1 exu_bypass_w1_eccgen_U53(.A(bypass_byp_irf_rd_data_m[37]), .B(bypass_byp_irf_rd_data_m[32]), .Y(bypass_w1_eccgen_n85));
XOR2X1 exu_bypass_w1_eccgen_U52(.A(bypass_byp_irf_rd_data_m[45]), .B(bypass_w1_eccgen_n119), .Y(bypass_w1_eccgen_p2_g[5]));
XOR2X1 exu_bypass_w1_eccgen_U51(.A(bypass_w1_eccgen_n123), .B(bypass_w1_eccgen_n86), .Y(bypass_w1_eccgen_p2_g[6]));
XOR2X1 exu_bypass_w1_eccgen_U50(.A(bypass_byp_irf_rd_data_m[53]), .B(bypass_byp_irf_rd_data_m[46]), .Y(bypass_w1_eccgen_n86));
XOR2X1 exu_bypass_w1_eccgen_U49(.A(bypass_w1_eccgen_n88), .B(bypass_w1_eccgen_n87), .Y(bypass_w1_eccgen_p2_g[7]));
XOR2X1 exu_bypass_w1_eccgen_U48(.A(bypass_w1_eccgen_n121), .B(bypass_w1_eccgen_n120), .Y(bypass_w1_eccgen_n87));
XOR2X1 exu_bypass_w1_eccgen_U47(.A(bypass_byp_irf_rd_data_m[60]), .B(exu_n15550), .Y(bypass_w1_eccgen_n88));
XOR2X1 exu_bypass_w1_eccgen_U46(.A(bypass_w1_eccgen_n90), .B(bypass_w1_eccgen_n89), .Y(bypass_w1_eccgen_p1_g[0]));
XOR2X1 exu_bypass_w1_eccgen_U45(.A(bypass_byp_irf_rd_data_m[2]), .B(bypass_byp_irf_rd_data_m[0]), .Y(bypass_w1_eccgen_n89));
XOR2X1 exu_bypass_w1_eccgen_U44(.A(bypass_byp_irf_rd_data_m[5]), .B(bypass_byp_irf_rd_data_m[3]), .Y(bypass_w1_eccgen_n90));
XOR2X1 exu_bypass_w1_eccgen_U43(.A(bypass_w1_eccgen_n122), .B(bypass_w1_eccgen_n91), .Y(bypass_w1_eccgen_p1_g[1]));
XOR2X1 exu_bypass_w1_eccgen_U42(.A(bypass_byp_irf_rd_data_m[12]), .B(bypass_byp_irf_rd_data_m[6]), .Y(bypass_w1_eccgen_n91));
XOR2X1 exu_bypass_w1_eccgen_U41(.A(bypass_w1_eccgen_n93), .B(bypass_w1_eccgen_n92), .Y(bypass_w1_eccgen_p1_g[2]));
XOR2X1 exu_bypass_w1_eccgen_U40(.A(bypass_byp_irf_rd_data_m[16]), .B(bypass_byp_irf_rd_data_m[13]), .Y(bypass_w1_eccgen_n92));
XOR2X1 exu_bypass_w1_eccgen_U39(.A(bypass_byp_irf_rd_data_m[20]), .B(bypass_byp_irf_rd_data_m[17]), .Y(bypass_w1_eccgen_n93));
XOR2X1 exu_bypass_w1_eccgen_U38(.A(bypass_w1_eccgen_n95), .B(bypass_w1_eccgen_n94), .Y(bypass_w1_eccgen_p1_g[3]));
XOR2X1 exu_bypass_w1_eccgen_U37(.A(bypass_byp_irf_rd_data_m[24]), .B(bypass_byp_irf_rd_data_m[21]), .Y(bypass_w1_eccgen_n94));
XOR2X1 exu_bypass_w1_eccgen_U36(.A(bypass_byp_irf_rd_data_m[27]), .B(bypass_byp_irf_rd_data_m[25]), .Y(bypass_w1_eccgen_n95));
XOR2X1 exu_bypass_w1_eccgen_U35(.A(bypass_w1_eccgen_n97), .B(bypass_w1_eccgen_n96), .Y(bypass_w1_eccgen_p1_g[4]));
XOR2X1 exu_bypass_w1_eccgen_U34(.A(bypass_byp_irf_rd_data_m[31]), .B(bypass_byp_irf_rd_data_m[28]), .Y(bypass_w1_eccgen_n96));
XOR2X1 exu_bypass_w1_eccgen_U33(.A(bypass_byp_irf_rd_data_m[35]), .B(bypass_byp_irf_rd_data_m[32]), .Y(bypass_w1_eccgen_n97));
XOR2X1 exu_bypass_w1_eccgen_U32(.A(bypass_w1_eccgen_n99), .B(bypass_w1_eccgen_n98), .Y(bypass_w1_eccgen_p1_g[5]));
XOR2X1 exu_bypass_w1_eccgen_U31(.A(bypass_byp_irf_rd_data_m[39]), .B(bypass_byp_irf_rd_data_m[36]), .Y(bypass_w1_eccgen_n98));
XOR2X1 exu_bypass_w1_eccgen_U30(.A(bypass_byp_irf_rd_data_m[43]), .B(bypass_byp_irf_rd_data_m[40]), .Y(bypass_w1_eccgen_n99));
XOR2X1 exu_bypass_w1_eccgen_U29(.A(bypass_w1_eccgen_n123), .B(bypass_w1_eccgen_n100), .Y(bypass_w1_eccgen_p1_g[6]));
XOR2X1 exu_bypass_w1_eccgen_U28(.A(bypass_byp_irf_rd_data_m[51]), .B(bypass_byp_irf_rd_data_m[44]), .Y(bypass_w1_eccgen_n100));
XOR2X1 exu_bypass_w1_eccgen_U27(.A(bypass_w1_eccgen_n102), .B(bypass_w1_eccgen_n101), .Y(bypass_w1_eccgen_n127));
XOR2X1 exu_bypass_w1_eccgen_U26(.A(bypass_byp_irf_rd_data_m[56]), .B(bypass_byp_irf_rd_data_m[52]), .Y(bypass_w1_eccgen_n101));
XOR2X1 exu_bypass_w1_eccgen_U25(.A(bypass_byp_irf_rd_data_m[63]), .B(bypass_byp_irf_rd_data_m[59]), .Y(bypass_w1_eccgen_n102));
XOR2X1 exu_bypass_w1_eccgen_U24(.A(bypass_w1_eccgen_n104), .B(bypass_w1_eccgen_n103), .Y(bypass_w1_eccgen_p1_g[7]));
XOR2X1 exu_bypass_w1_eccgen_U23(.A(bypass_w1_eccgen_n127), .B(bypass_w1_eccgen_n105), .Y(bypass_w1_eccgen_n103));
XOR2X1 exu_bypass_w1_eccgen_U22(.A(bypass_byp_irf_rd_data_m[55]), .B(exu_n15551), .Y(bypass_w1_eccgen_n104));
XOR2X1 exu_bypass_w1_eccgen_U21(.A(bypass_byp_irf_rd_data_m[62]), .B(bypass_byp_irf_rd_data_m[58]), .Y(bypass_w1_eccgen_n105));
XOR2X1 exu_bypass_w1_eccgen_U20(.A(bypass_byp_irf_rd_data_m[3]), .B(bypass_w1_eccgen_n124), .Y(bypass_w1_eccgen_p0_g[0]));
XOR2X1 exu_bypass_w1_eccgen_U19(.A(bypass_w1_eccgen_n107), .B(bypass_w1_eccgen_n106), .Y(bypass_w1_eccgen_p0_g[1]));
XOR2X1 exu_bypass_w1_eccgen_U18(.A(bypass_byp_irf_rd_data_m[8]), .B(bypass_byp_irf_rd_data_m[6]), .Y(bypass_w1_eccgen_n106));
XOR2X1 exu_bypass_w1_eccgen_U17(.A(bypass_byp_irf_rd_data_m[11]), .B(bypass_byp_irf_rd_data_m[10]), .Y(bypass_w1_eccgen_n107));
XOR2X1 exu_bypass_w1_eccgen_U16(.A(bypass_w1_eccgen_n109), .B(bypass_w1_eccgen_n108), .Y(bypass_w1_eccgen_p0_g[2]));
XOR2X1 exu_bypass_w1_eccgen_U15(.A(bypass_byp_irf_rd_data_m[15]), .B(bypass_byp_irf_rd_data_m[13]), .Y(bypass_w1_eccgen_n108));
XOR2X1 exu_bypass_w1_eccgen_U14(.A(bypass_byp_irf_rd_data_m[19]), .B(bypass_byp_irf_rd_data_m[17]), .Y(bypass_w1_eccgen_n109));
XOR2X1 exu_bypass_w1_eccgen_U13(.A(bypass_byp_irf_rd_data_m[25]), .B(bypass_w1_eccgen_n125), .Y(bypass_w1_eccgen_p0_g[3]));
XOR2X1 exu_bypass_w1_eccgen_U12(.A(bypass_w1_eccgen_n111), .B(bypass_w1_eccgen_n110), .Y(bypass_w1_eccgen_p0_g[4]));
XOR2X1 exu_bypass_w1_eccgen_U11(.A(bypass_byp_irf_rd_data_m[30]), .B(bypass_byp_irf_rd_data_m[28]), .Y(bypass_w1_eccgen_n110));
XOR2X1 exu_bypass_w1_eccgen_U10(.A(bypass_byp_irf_rd_data_m[34]), .B(bypass_byp_irf_rd_data_m[32]), .Y(bypass_w1_eccgen_n111));
XOR2X1 exu_bypass_w1_eccgen_U9(.A(bypass_w1_eccgen_n113), .B(bypass_w1_eccgen_n112), .Y(bypass_w1_eccgen_p0_g[5]));
XOR2X1 exu_bypass_w1_eccgen_U8(.A(bypass_byp_irf_rd_data_m[38]), .B(bypass_byp_irf_rd_data_m[36]), .Y(bypass_w1_eccgen_n112));
XOR2X1 exu_bypass_w1_eccgen_U7(.A(bypass_byp_irf_rd_data_m[42]), .B(bypass_byp_irf_rd_data_m[40]), .Y(bypass_w1_eccgen_n113));
XOR2X1 exu_bypass_w1_eccgen_U6(.A(bypass_byp_irf_rd_data_m[48]), .B(bypass_w1_eccgen_n126), .Y(bypass_w1_eccgen_p0_g[6]));
XOR2X1 exu_bypass_w1_eccgen_U5(.A(bypass_w1_eccgen_n115), .B(bypass_w1_eccgen_n114), .Y(bypass_w1_eccgen_p0_g[7]));
XOR2X1 exu_bypass_w1_eccgen_U4(.A(bypass_w1_eccgen_n127), .B(bypass_w1_eccgen_n116), .Y(bypass_w1_eccgen_n114));
XOR2X1 exu_bypass_w1_eccgen_U3(.A(bypass_byp_irf_rd_data_m[54]), .B(exu_n15552), .Y(bypass_w1_eccgen_n115));
XOR2X1 exu_bypass_w1_eccgen_U2(.A(bypass_byp_irf_rd_data_m[61]), .B(bypass_byp_irf_rd_data_m[57]), .Y(bypass_w1_eccgen_n116));
XOR2X1 exu_bypass_w1_eccgen_U1(.A(bypass_w1_eccgen_p6_w[1]), .B(bypass_w1_eccgen_p6_w[0]), .Y(bypass_rd_synd_w_l[6]));
DFFPOSX1 ecc_rs1_ecc_d2e_q_reg[0](.D(ecc_rs1_ecc_d2e_n15), .CLK(rclk), .Q(ecc_rs1_ecc_e[0]));
DFFPOSX1 ecc_rs1_ecc_d2e_q_reg[1](.D(ecc_rs1_ecc_d2e_n13), .CLK(rclk), .Q(ecc_rs1_ecc_e[1]));
DFFPOSX1 ecc_rs1_ecc_d2e_q_reg[2](.D(ecc_rs1_ecc_d2e_n11), .CLK(rclk), .Q(ecc_rs1_ecc_e[2]));
DFFPOSX1 ecc_rs1_ecc_d2e_q_reg[3](.D(ecc_rs1_ecc_d2e_n9), .CLK(rclk), .Q(ecc_rs1_ecc_e[3]));
DFFPOSX1 ecc_rs1_ecc_d2e_q_reg[4](.D(ecc_rs1_ecc_d2e_n7), .CLK(rclk), .Q(ecc_rs1_ecc_e[4]));
DFFPOSX1 ecc_rs1_ecc_d2e_q_reg[5](.D(ecc_rs1_ecc_d2e_n5), .CLK(rclk), .Q(ecc_rs1_ecc_e[5]));
DFFPOSX1 ecc_rs1_ecc_d2e_q_reg[6](.D(ecc_rs1_ecc_d2e_n3), .CLK(rclk), .Q(ecc_rs1_ecc_e[6]));
DFFPOSX1 ecc_rs1_ecc_d2e_q_reg[7](.D(ecc_rs1_ecc_d2e_n17), .CLK(rclk), .Q(ecc_rs1_ecc_e[7]));
XOR2X1 exu_ecc_chk_rs1_U149(.A(ecc_chk_rs1_n11), .B(ecc_chk_rs1_n10), .Y(ecc_chk_rs1_n133));
XOR2X1 exu_ecc_chk_rs1_U148(.A(byp_alu_rcc_data_e[52]), .B(byp_alu_rcc_data_e[50]), .Y(ecc_chk_rs1_n10));
XOR2X1 exu_ecc_chk_rs1_U147(.A(byp_alu_rcc_data_e[56]), .B(byp_alu_rcc_data_e[54]), .Y(ecc_chk_rs1_n11));
XOR2X1 exu_ecc_chk_rs1_U146(.A(ecc_chk_rs1_n13), .B(ecc_chk_rs1_n12), .Y(ecc_chk_rs1_n137));
XOR2X1 exu_ecc_chk_rs1_U145(.A(byp_alu_rcc_data_e[36]), .B(byp_alu_rcc_data_e[34]), .Y(ecc_chk_rs1_n12));
XOR2X1 exu_ecc_chk_rs1_U144(.A(byp_alu_rcc_data_e[40]), .B(byp_alu_rcc_data_e[38]), .Y(ecc_chk_rs1_n13));
XOR2X1 exu_ecc_chk_rs1_U143(.A(ecc_chk_rs1_n15), .B(ecc_chk_rs1_n14), .Y(ecc_chk_rs1_n135));
XOR2X1 exu_ecc_chk_rs1_U142(.A(byp_alu_rcc_data_e[21]), .B(byp_alu_rcc_data_e[19]), .Y(ecc_chk_rs1_n14));
XOR2X1 exu_ecc_chk_rs1_U141(.A(byp_alu_rcc_data_e[25]), .B(byp_alu_rcc_data_e[23]), .Y(ecc_chk_rs1_n15));
XOR2X1 exu_ecc_chk_rs1_U140(.A(ecc_chk_rs1_n17), .B(ecc_chk_rs1_n16), .Y(ecc_chk_rs1_n131));
XOR2X1 exu_ecc_chk_rs1_U139(.A(ecc_chk_rs1_n19), .B(ecc_chk_rs1_n18), .Y(ecc_chk_rs1_n16));
XOR2X1 exu_ecc_chk_rs1_U138(.A(ecc_chk_rs1_n135), .B(ecc_chk_rs1_n20), .Y(ecc_chk_rs1_n17));
XOR2X1 exu_ecc_chk_rs1_U137(.A(ecc_chk_rs1_n133), .B(ecc_chk_rs1_n137), .Y(ecc_chk_rs1_n18));
XOR2X1 exu_ecc_chk_rs1_U136(.A(byp_alu_rcc_data_e[6]), .B(byp_alu_rcc_data_e[4]), .Y(ecc_chk_rs1_n19));
XOR2X1 exu_ecc_chk_rs1_U135(.A(byp_alu_rcc_data_e[10]), .B(byp_alu_rcc_data_e[8]), .Y(ecc_chk_rs1_n20));
XOR2X1 exu_ecc_chk_rs1_U134(.A(ecc_chk_rs1_n22), .B(ecc_chk_rs1_n21), .Y(ecc_chk_rs1_n124));
XOR2X1 exu_ecc_chk_rs1_U133(.A(byp_alu_rcc_data_e[3]), .B(ecc_chk_rs1_n23), .Y(ecc_chk_rs1_n21));
XOR2X1 exu_ecc_chk_rs1_U132(.A(byp_alu_rcc_data_e[32]), .B(byp_alu_rcc_data_e[17]), .Y(ecc_chk_rs1_n22));
XOR2X1 exu_ecc_chk_rs1_U131(.A(exu_ifu_regn_e), .B(byp_alu_rcc_data_e[48]), .Y(ecc_chk_rs1_n23));
XOR2X1 exu_ecc_chk_rs1_U130(.A(ecc_chk_rs1_n25), .B(ecc_chk_rs1_n24), .Y(ecc_chk_rs1_n128));
XOR2X1 exu_ecc_chk_rs1_U129(.A(byp_alu_rcc_data_e[1]), .B(ecc_chk_rs1_n26), .Y(ecc_chk_rs1_n24));
XOR2X1 exu_ecc_chk_rs1_U128(.A(byp_alu_rcc_data_e[30]), .B(byp_alu_rcc_data_e[15]), .Y(ecc_chk_rs1_n25));
XOR2X1 exu_ecc_chk_rs1_U127(.A(byp_alu_rcc_data_e[61]), .B(byp_alu_rcc_data_e[46]), .Y(ecc_chk_rs1_n26));
XOR2X1 exu_ecc_chk_rs1_U126(.A(ecc_chk_rs1_n28), .B(ecc_chk_rs1_n27), .Y(ecc_chk_rs1_n126));
XOR2X1 exu_ecc_chk_rs1_U125(.A(byp_alu_rcc_data_e[0]), .B(ecc_chk_rs1_n29), .Y(ecc_chk_rs1_n27));
XOR2X1 exu_ecc_chk_rs1_U124(.A(byp_alu_rcc_data_e[28]), .B(byp_alu_rcc_data_e[13]), .Y(ecc_chk_rs1_n28));
XOR2X1 exu_ecc_chk_rs1_U123(.A(byp_alu_rcc_data_e[59]), .B(byp_alu_rcc_data_e[44]), .Y(ecc_chk_rs1_n29));
XOR2X1 exu_ecc_chk_rs1_U122(.A(ecc_chk_rs1_n31), .B(ecc_chk_rs1_n30), .Y(ecc_rs1_err_e[0]));
XOR2X1 exu_ecc_chk_rs1_U121(.A(ecc_chk_rs1_n33), .B(ecc_chk_rs1_n32), .Y(ecc_chk_rs1_n30));
XOR2X1 exu_ecc_chk_rs1_U120(.A(ecc_chk_rs1_n35), .B(ecc_chk_rs1_n34), .Y(ecc_chk_rs1_n31));
XOR2X1 exu_ecc_chk_rs1_U119(.A(ecc_chk_rs1_n126), .B(ecc_chk_rs1_n36), .Y(ecc_chk_rs1_n32));
XOR2X1 exu_ecc_chk_rs1_U118(.A(ecc_chk_rs1_n124), .B(ecc_chk_rs1_n128), .Y(ecc_chk_rs1_n33));
XOR2X1 exu_ecc_chk_rs1_U117(.A(ecc_rs1_ecc_e[0]), .B(ecc_chk_rs1_n131), .Y(ecc_chk_rs1_n34));
XOR2X1 exu_ecc_chk_rs1_U116(.A(byp_alu_rcc_data_e[26]), .B(byp_alu_rcc_data_e[11]), .Y(ecc_chk_rs1_n35));
XOR2X1 exu_ecc_chk_rs1_U115(.A(byp_alu_rcc_data_e[57]), .B(byp_alu_rcc_data_e[42]), .Y(ecc_chk_rs1_n36));
XOR2X1 exu_ecc_chk_rs1_U114(.A(ecc_chk_rs1_n38), .B(ecc_chk_rs1_n37), .Y(ecc_chk_rs1_n132));
XOR2X1 exu_ecc_chk_rs1_U113(.A(byp_alu_rcc_data_e[51]), .B(byp_alu_rcc_data_e[49]), .Y(ecc_chk_rs1_n37));
XOR2X1 exu_ecc_chk_rs1_U112(.A(byp_alu_rcc_data_e[55]), .B(byp_alu_rcc_data_e[53]), .Y(ecc_chk_rs1_n38));
XOR2X1 exu_ecc_chk_rs1_U111(.A(ecc_chk_rs1_n40), .B(ecc_chk_rs1_n39), .Y(ecc_chk_rs1_n136));
XOR2X1 exu_ecc_chk_rs1_U110(.A(byp_alu_rcc_data_e[35]), .B(byp_alu_rcc_data_e[33]), .Y(ecc_chk_rs1_n39));
XOR2X1 exu_ecc_chk_rs1_U109(.A(byp_alu_rcc_data_e[39]), .B(byp_alu_rcc_data_e[37]), .Y(ecc_chk_rs1_n40));
XOR2X1 exu_ecc_chk_rs1_U108(.A(ecc_chk_rs1_n42), .B(ecc_chk_rs1_n41), .Y(ecc_chk_rs1_n134));
XOR2X1 exu_ecc_chk_rs1_U107(.A(byp_alu_rcc_data_e[20]), .B(byp_alu_rcc_data_e[18]), .Y(ecc_chk_rs1_n41));
XOR2X1 exu_ecc_chk_rs1_U106(.A(byp_alu_rcc_data_e[24]), .B(byp_alu_rcc_data_e[22]), .Y(ecc_chk_rs1_n42));
XOR2X1 exu_ecc_chk_rs1_U105(.A(ecc_chk_rs1_n44), .B(ecc_chk_rs1_n43), .Y(ecc_chk_rs1_n130));
XOR2X1 exu_ecc_chk_rs1_U104(.A(ecc_chk_rs1_n46), .B(ecc_chk_rs1_n45), .Y(ecc_chk_rs1_n43));
XOR2X1 exu_ecc_chk_rs1_U103(.A(ecc_chk_rs1_n134), .B(ecc_chk_rs1_n47), .Y(ecc_chk_rs1_n44));
XOR2X1 exu_ecc_chk_rs1_U102(.A(ecc_chk_rs1_n132), .B(ecc_chk_rs1_n136), .Y(ecc_chk_rs1_n45));
XOR2X1 exu_ecc_chk_rs1_U101(.A(byp_alu_rcc_data_e[5]), .B(ecc_rs1_ecc_e[3]), .Y(ecc_chk_rs1_n46));
XOR2X1 exu_ecc_chk_rs1_U100(.A(byp_alu_rcc_data_e[9]), .B(byp_alu_rcc_data_e[7]), .Y(ecc_chk_rs1_n47));
XOR2X1 exu_ecc_chk_rs1_U99(.A(ecc_chk_rs1_n49), .B(ecc_chk_rs1_n48), .Y(ecc_chk_rs1_n123));
XOR2X1 exu_ecc_chk_rs1_U98(.A(byp_alu_rcc_data_e[2]), .B(ecc_chk_rs1_n50), .Y(ecc_chk_rs1_n48));
XOR2X1 exu_ecc_chk_rs1_U97(.A(byp_alu_rcc_data_e[31]), .B(byp_alu_rcc_data_e[16]), .Y(ecc_chk_rs1_n49));
XOR2X1 exu_ecc_chk_rs1_U96(.A(byp_alu_rcc_data_e[62]), .B(byp_alu_rcc_data_e[47]), .Y(ecc_chk_rs1_n50));
XOR2X1 exu_ecc_chk_rs1_U95(.A(ecc_chk_rs1_n52), .B(ecc_chk_rs1_n51), .Y(ecc_chk_rs1_n127));
XOR2X1 exu_ecc_chk_rs1_U94(.A(ecc_rs1_ecc_e[2]), .B(ecc_chk_rs1_n53), .Y(ecc_chk_rs1_n51));
XOR2X1 exu_ecc_chk_rs1_U93(.A(byp_alu_rcc_data_e[29]), .B(byp_alu_rcc_data_e[14]), .Y(ecc_chk_rs1_n52));
XOR2X1 exu_ecc_chk_rs1_U92(.A(byp_alu_rcc_data_e[60]), .B(byp_alu_rcc_data_e[45]), .Y(ecc_chk_rs1_n53));
XOR2X1 exu_ecc_chk_rs1_U91(.A(ecc_chk_rs1_n55), .B(ecc_chk_rs1_n54), .Y(ecc_chk_rs1_n125));
XOR2X1 exu_ecc_chk_rs1_U90(.A(ecc_rs1_ecc_e[1]), .B(ecc_chk_rs1_n56), .Y(ecc_chk_rs1_n54));
XOR2X1 exu_ecc_chk_rs1_U89(.A(byp_alu_rcc_data_e[27]), .B(byp_alu_rcc_data_e[12]), .Y(ecc_chk_rs1_n55));
XOR2X1 exu_ecc_chk_rs1_U88(.A(byp_alu_rcc_data_e[58]), .B(byp_alu_rcc_data_e[43]), .Y(ecc_chk_rs1_n56));
XOR2X1 exu_ecc_chk_rs1_U87(.A(ecc_chk_rs1_n58), .B(ecc_chk_rs1_n57), .Y(ecc_chk_rs1_parity));
XOR2X1 exu_ecc_chk_rs1_U86(.A(ecc_chk_rs1_n60), .B(ecc_chk_rs1_n59), .Y(ecc_chk_rs1_n57));
XOR2X1 exu_ecc_chk_rs1_U85(.A(ecc_chk_rs1_n62), .B(ecc_chk_rs1_n61), .Y(ecc_chk_rs1_n58));
XOR2X1 exu_ecc_chk_rs1_U84(.A(ecc_chk_rs1_n64), .B(ecc_chk_rs1_n63), .Y(ecc_chk_rs1_n59));
XOR2X1 exu_ecc_chk_rs1_U83(.A(ecc_chk_rs1_n127), .B(ecc_chk_rs1_n125), .Y(ecc_chk_rs1_n60));
XOR2X1 exu_ecc_chk_rs1_U82(.A(ecc_chk_rs1_n130), .B(ecc_chk_rs1_n123), .Y(ecc_chk_rs1_n61));
XOR2X1 exu_ecc_chk_rs1_U81(.A(ecc_rs1_ecc_e[4]), .B(ecc_rs1_err_e[0]), .Y(ecc_chk_rs1_n62));
XOR2X1 exu_ecc_chk_rs1_U80(.A(ecc_rs1_ecc_e[6]), .B(ecc_rs1_ecc_e[5]), .Y(ecc_chk_rs1_n63));
XOR2X1 exu_ecc_chk_rs1_U79(.A(byp_alu_rcc_data_e[41]), .B(ecc_rs1_ecc_e[7]), .Y(ecc_chk_rs1_n64));
XOR2X1 exu_ecc_chk_rs1_U78(.A(ecc_chk_rs1_n66), .B(ecc_chk_rs1_n65), .Y(ecc_chk_rs1_n129));
XOR2X1 exu_ecc_chk_rs1_U77(.A(ecc_chk_rs1_n68), .B(ecc_chk_rs1_n67), .Y(ecc_chk_rs1_n65));
XOR2X1 exu_ecc_chk_rs1_U76(.A(ecc_chk_rs1_n70), .B(ecc_chk_rs1_n69), .Y(ecc_chk_rs1_n66));
XOR2X1 exu_ecc_chk_rs1_U75(.A(ecc_chk_rs1_n72), .B(ecc_chk_rs1_n71), .Y(ecc_chk_rs1_n67));
XOR2X1 exu_ecc_chk_rs1_U74(.A(ecc_chk_rs1_n124), .B(ecc_chk_rs1_n123), .Y(ecc_chk_rs1_n68));
XOR2X1 exu_ecc_chk_rs1_U73(.A(byp_alu_rcc_data_e[10]), .B(byp_alu_rcc_data_e[9]), .Y(ecc_chk_rs1_n69));
XOR2X1 exu_ecc_chk_rs1_U72(.A(byp_alu_rcc_data_e[25]), .B(byp_alu_rcc_data_e[24]), .Y(ecc_chk_rs1_n70));
XOR2X1 exu_ecc_chk_rs1_U71(.A(byp_alu_rcc_data_e[40]), .B(byp_alu_rcc_data_e[39]), .Y(ecc_chk_rs1_n71));
XOR2X1 exu_ecc_chk_rs1_U70(.A(byp_alu_rcc_data_e[56]), .B(byp_alu_rcc_data_e[55]), .Y(ecc_chk_rs1_n72));
XOR2X1 exu_ecc_chk_rs1_U69(.A(ecc_chk_rs1_n74), .B(ecc_chk_rs1_n73), .Y(ecc_rs1_err_e[1]));
XOR2X1 exu_ecc_chk_rs1_U68(.A(ecc_chk_rs1_n76), .B(ecc_chk_rs1_n75), .Y(ecc_chk_rs1_n73));
XOR2X1 exu_ecc_chk_rs1_U67(.A(ecc_chk_rs1_n78), .B(ecc_chk_rs1_n77), .Y(ecc_chk_rs1_n74));
XOR2X1 exu_ecc_chk_rs1_U66(.A(ecc_chk_rs1_n80), .B(ecc_chk_rs1_n79), .Y(ecc_chk_rs1_n75));
XOR2X1 exu_ecc_chk_rs1_U65(.A(ecc_chk_rs1_n125), .B(ecc_chk_rs1_n81), .Y(ecc_chk_rs1_n76));
XOR2X1 exu_ecc_chk_rs1_U64(.A(ecc_chk_rs1_n129), .B(ecc_chk_rs1_n126), .Y(ecc_chk_rs1_n77));
XOR2X1 exu_ecc_chk_rs1_U63(.A(byp_alu_rcc_data_e[6]), .B(byp_alu_rcc_data_e[5]), .Y(ecc_chk_rs1_n78));
XOR2X1 exu_ecc_chk_rs1_U62(.A(byp_alu_rcc_data_e[21]), .B(byp_alu_rcc_data_e[20]), .Y(ecc_chk_rs1_n79));
XOR2X1 exu_ecc_chk_rs1_U61(.A(byp_alu_rcc_data_e[36]), .B(byp_alu_rcc_data_e[35]), .Y(ecc_chk_rs1_n80));
XOR2X1 exu_ecc_chk_rs1_U60(.A(byp_alu_rcc_data_e[52]), .B(byp_alu_rcc_data_e[51]), .Y(ecc_chk_rs1_n81));
XOR2X1 exu_ecc_chk_rs1_U59(.A(ecc_chk_rs1_n83), .B(ecc_chk_rs1_n82), .Y(ecc_rs1_err_e[2]));
XOR2X1 exu_ecc_chk_rs1_U58(.A(ecc_chk_rs1_n85), .B(ecc_chk_rs1_n84), .Y(ecc_chk_rs1_n82));
XOR2X1 exu_ecc_chk_rs1_U57(.A(ecc_chk_rs1_n87), .B(ecc_chk_rs1_n86), .Y(ecc_chk_rs1_n83));
XOR2X1 exu_ecc_chk_rs1_U56(.A(ecc_chk_rs1_n89), .B(ecc_chk_rs1_n88), .Y(ecc_chk_rs1_n84));
XOR2X1 exu_ecc_chk_rs1_U55(.A(ecc_chk_rs1_n127), .B(ecc_chk_rs1_n90), .Y(ecc_chk_rs1_n85));
XOR2X1 exu_ecc_chk_rs1_U54(.A(ecc_chk_rs1_n129), .B(ecc_chk_rs1_n128), .Y(ecc_chk_rs1_n86));
XOR2X1 exu_ecc_chk_rs1_U53(.A(byp_alu_rcc_data_e[8]), .B(byp_alu_rcc_data_e[7]), .Y(ecc_chk_rs1_n87));
XOR2X1 exu_ecc_chk_rs1_U52(.A(byp_alu_rcc_data_e[23]), .B(byp_alu_rcc_data_e[22]), .Y(ecc_chk_rs1_n88));
XOR2X1 exu_ecc_chk_rs1_U51(.A(byp_alu_rcc_data_e[38]), .B(byp_alu_rcc_data_e[37]), .Y(ecc_chk_rs1_n89));
XOR2X1 exu_ecc_chk_rs1_U50(.A(byp_alu_rcc_data_e[54]), .B(byp_alu_rcc_data_e[53]), .Y(ecc_chk_rs1_n90));
XOR2X1 exu_ecc_chk_rs1_U49(.A(ecc_chk_rs1_n131), .B(ecc_chk_rs1_n130), .Y(ecc_rs1_err_e[3]));
XOR2X1 exu_ecc_chk_rs1_U48(.A(ecc_chk_rs1_n92), .B(ecc_chk_rs1_n91), .Y(ecc_chk_rs1_n138));
XOR2X1 exu_ecc_chk_rs1_U47(.A(ecc_chk_rs1_n94), .B(ecc_chk_rs1_n93), .Y(ecc_chk_rs1_n91));
XOR2X1 exu_ecc_chk_rs1_U46(.A(ecc_chk_rs1_n96), .B(ecc_chk_rs1_n95), .Y(ecc_chk_rs1_n92));
XOR2X1 exu_ecc_chk_rs1_U45(.A(ecc_chk_rs1_n98), .B(ecc_chk_rs1_n97), .Y(ecc_chk_rs1_n93));
XOR2X1 exu_ecc_chk_rs1_U44(.A(ecc_chk_rs1_n133), .B(ecc_chk_rs1_n132), .Y(ecc_chk_rs1_n94));
XOR2X1 exu_ecc_chk_rs1_U43(.A(byp_alu_rcc_data_e[42]), .B(byp_alu_rcc_data_e[41]), .Y(ecc_chk_rs1_n95));
XOR2X1 exu_ecc_chk_rs1_U42(.A(byp_alu_rcc_data_e[44]), .B(byp_alu_rcc_data_e[43]), .Y(ecc_chk_rs1_n96));
XOR2X1 exu_ecc_chk_rs1_U41(.A(byp_alu_rcc_data_e[46]), .B(byp_alu_rcc_data_e[45]), .Y(ecc_chk_rs1_n97));
XOR2X1 exu_ecc_chk_rs1_U40(.A(byp_alu_rcc_data_e[48]), .B(byp_alu_rcc_data_e[47]), .Y(ecc_chk_rs1_n98));
XOR2X1 exu_ecc_chk_rs1_U39(.A(ecc_chk_rs1_n100), .B(ecc_chk_rs1_n99), .Y(ecc_rs1_err_e[4]));
XOR2X1 exu_ecc_chk_rs1_U38(.A(ecc_chk_rs1_n102), .B(ecc_chk_rs1_n101), .Y(ecc_chk_rs1_n99));
XOR2X1 exu_ecc_chk_rs1_U37(.A(ecc_chk_rs1_n104), .B(ecc_chk_rs1_n103), .Y(ecc_chk_rs1_n100));
XOR2X1 exu_ecc_chk_rs1_U36(.A(ecc_chk_rs1_n106), .B(ecc_chk_rs1_n105), .Y(ecc_chk_rs1_n101));
XOR2X1 exu_ecc_chk_rs1_U35(.A(ecc_chk_rs1_n134), .B(ecc_chk_rs1_n107), .Y(ecc_chk_rs1_n102));
XOR2X1 exu_ecc_chk_rs1_U34(.A(ecc_chk_rs1_n138), .B(ecc_chk_rs1_n135), .Y(ecc_chk_rs1_n103));
XOR2X1 exu_ecc_chk_rs1_U33(.A(byp_alu_rcc_data_e[11]), .B(ecc_rs1_ecc_e[4]), .Y(ecc_chk_rs1_n104));
XOR2X1 exu_ecc_chk_rs1_U32(.A(byp_alu_rcc_data_e[13]), .B(byp_alu_rcc_data_e[12]), .Y(ecc_chk_rs1_n105));
XOR2X1 exu_ecc_chk_rs1_U31(.A(byp_alu_rcc_data_e[15]), .B(byp_alu_rcc_data_e[14]), .Y(ecc_chk_rs1_n106));
XOR2X1 exu_ecc_chk_rs1_U30(.A(byp_alu_rcc_data_e[17]), .B(byp_alu_rcc_data_e[16]), .Y(ecc_chk_rs1_n107));
XOR2X1 exu_ecc_chk_rs1_U29(.A(ecc_chk_rs1_n109), .B(ecc_chk_rs1_n108), .Y(ecc_rs1_err_e[5]));
XOR2X1 exu_ecc_chk_rs1_U28(.A(ecc_chk_rs1_n111), .B(ecc_chk_rs1_n110), .Y(ecc_chk_rs1_n108));
XOR2X1 exu_ecc_chk_rs1_U27(.A(ecc_chk_rs1_n113), .B(ecc_chk_rs1_n112), .Y(ecc_chk_rs1_n109));
XOR2X1 exu_ecc_chk_rs1_U26(.A(ecc_chk_rs1_n115), .B(ecc_chk_rs1_n114), .Y(ecc_chk_rs1_n110));
XOR2X1 exu_ecc_chk_rs1_U25(.A(ecc_chk_rs1_n136), .B(ecc_chk_rs1_n116), .Y(ecc_chk_rs1_n111));
XOR2X1 exu_ecc_chk_rs1_U24(.A(ecc_chk_rs1_n138), .B(ecc_chk_rs1_n137), .Y(ecc_chk_rs1_n112));
XOR2X1 exu_ecc_chk_rs1_U23(.A(byp_alu_rcc_data_e[26]), .B(ecc_rs1_ecc_e[5]), .Y(ecc_chk_rs1_n113));
XOR2X1 exu_ecc_chk_rs1_U22(.A(byp_alu_rcc_data_e[28]), .B(byp_alu_rcc_data_e[27]), .Y(ecc_chk_rs1_n114));
XOR2X1 exu_ecc_chk_rs1_U21(.A(byp_alu_rcc_data_e[30]), .B(byp_alu_rcc_data_e[29]), .Y(ecc_chk_rs1_n115));
XOR2X1 exu_ecc_chk_rs1_U20(.A(byp_alu_rcc_data_e[32]), .B(byp_alu_rcc_data_e[31]), .Y(ecc_chk_rs1_n116));
XOR2X1 exu_ecc_chk_rs1_U19(.A(ecc_chk_rs1_n118), .B(ecc_chk_rs1_n117), .Y(ecc_rs1_err_e[6]));
XOR2X1 exu_ecc_chk_rs1_U18(.A(ecc_chk_rs1_n120), .B(ecc_chk_rs1_n119), .Y(ecc_chk_rs1_n117));
XOR2X1 exu_ecc_chk_rs1_U17(.A(ecc_chk_rs1_n122), .B(ecc_chk_rs1_n121), .Y(ecc_chk_rs1_n118));
XOR2X1 exu_ecc_chk_rs1_U16(.A(byp_alu_rcc_data_e[57]), .B(ecc_rs1_ecc_e[6]), .Y(ecc_chk_rs1_n119));
XOR2X1 exu_ecc_chk_rs1_U15(.A(byp_alu_rcc_data_e[59]), .B(byp_alu_rcc_data_e[58]), .Y(ecc_chk_rs1_n120));
XOR2X1 exu_ecc_chk_rs1_U14(.A(byp_alu_rcc_data_e[61]), .B(byp_alu_rcc_data_e[60]), .Y(ecc_chk_rs1_n121));
XOR2X1 exu_ecc_chk_rs1_U13(.A(exu_ifu_regn_e), .B(byp_alu_rcc_data_e[62]), .Y(ecc_chk_rs1_n122));
DFFPOSX1 ecc_rs1_err_e2m_q_reg[0](.D(ecc_rs1_err_e2m_n15), .CLK(rclk), .Q(ecc_rs1_err_m[0]));
DFFPOSX1 ecc_rs1_err_e2m_q_reg[1](.D(ecc_rs1_err_e2m_n13), .CLK(rclk), .Q(ecc_rs1_err_m[1]));
DFFPOSX1 ecc_rs1_err_e2m_q_reg[2](.D(ecc_rs1_err_e2m_n11), .CLK(rclk), .Q(ecc_rs1_err_m[2]));
DFFPOSX1 ecc_rs1_err_e2m_q_reg[3](.D(ecc_rs1_err_e2m_n9), .CLK(rclk), .Q(ecc_rs1_err_m[3]));
DFFPOSX1 ecc_rs1_err_e2m_q_reg[4](.D(ecc_rs1_err_e2m_n7), .CLK(rclk), .Q(ecc_rs1_err_m[4]));
DFFPOSX1 ecc_rs1_err_e2m_q_reg[5](.D(ecc_rs1_err_e2m_n5), .CLK(rclk), .Q(ecc_rs1_err_m[5]));
DFFPOSX1 ecc_rs1_err_e2m_q_reg[6](.D(ecc_rs1_err_e2m_n3), .CLK(rclk), .Q(ecc_rs1_err_m[6]));
DFFSR ecl_rstff_q_reg[0](.D(exu_n19921), .CLK(rclk), .Q(ecl_ecl_reset_l));
DFFPOSX1 ecl_dff_rs1_s2d_q_reg[0](.D(ecl_dff_rs1_s2d_n11), .CLK(rclk), .Q(ecl_ifu_exu_rs1_d[0]));
DFFPOSX1 ecl_dff_rs1_s2d_q_reg[1](.D(ecl_dff_rs1_s2d_n9), .CLK(rclk), .Q(ecl_ifu_exu_rs1_d[1]));
DFFPOSX1 ecl_dff_rs1_s2d_q_reg[2](.D(ecl_dff_rs1_s2d_n7), .CLK(rclk), .Q(ecl_ifu_exu_rs1_d[2]));
DFFPOSX1 ecl_dff_rs1_s2d_q_reg[3](.D(ecl_dff_rs1_s2d_n5), .CLK(rclk), .Q(ecl_ifu_exu_rs1_d[3]));
DFFPOSX1 ecl_dff_rs1_s2d_q_reg[4](.D(ecl_dff_rs1_s2d_n3), .CLK(rclk), .Q(ecl_ifu_exu_rs1_d[4]));
DFFPOSX1 ecl_dff_ld_tid_m2g_q_reg[0](.D(ecl_dff_ld_tid_m2g_n5), .CLK(rclk), .Q(ecl_ld_tid_g[0]));
DFFPOSX1 ecl_dff_ld_tid_m2g_q_reg[1](.D(ecl_dff_ld_tid_m2g_n3), .CLK(rclk), .Q(ecl_ld_tid_g[1]));
DFFPOSX1 ecl_dff_aluop_d2e_q_reg[0](.D(ecl_dff_aluop_d2e_n7), .CLK(rclk), .Q(ecl_ifu_exu_aluop_e[0]));
DFFPOSX1 ecl_dff_aluop_d2e_q_reg[1](.D(ecl_dff_aluop_d2e_n5), .CLK(rclk), .Q(ecl_ifu_exu_aluop_e[1]));
DFFPOSX1 ecl_dff_aluop_d2e_q_reg[2](.D(ecl_dff_aluop_d2e_n3), .CLK(rclk), .Q(ecl_ifu_exu_aluop_e[2]));
DFFPOSX1 ecl_dff_enshift_d2e_q_reg[0](.D(ecl_dff_enshift_d2e_n3), .CLK(rclk), .Q(ecl_enshift_e));
DFFPOSX1 ecl_perr_dff_q_reg[0](.D(ecl_perr_dff_n9), .CLK(rclk), .Q(ecl_perr_store[0]));
DFFPOSX1 ecl_perr_dff_q_reg[1](.D(ecl_perr_dff_n7), .CLK(rclk), .Q(ecl_perr_store[1]));
DFFPOSX1 ecl_perr_dff_q_reg[2](.D(ecl_perr_dff_n5), .CLK(rclk), .Q(ecl_perr_store[2]));
DFFPOSX1 ecl_perr_dff_q_reg[3](.D(ecl_perr_dff_n2), .CLK(rclk), .Q(ecl_perr_store[3]));
DFFPOSX1 ecl_ttype_e2m_q_reg[0](.D(ecl_ttype_e2m_n15), .CLK(rclk), .Q(ecl_early_ttype_m[0]));
DFFPOSX1 ecl_ttype_e2m_q_reg[1](.D(ecl_ttype_e2m_n13), .CLK(rclk), .Q(ecl_early_ttype_m[1]));
DFFPOSX1 ecl_ttype_e2m_q_reg[2](.D(ecl_ttype_e2m_n11), .CLK(rclk), .Q(ecl_early_ttype_m[2]));
DFFPOSX1 ecl_ttype_e2m_q_reg[3](.D(ecl_ttype_e2m_n9), .CLK(rclk), .Q(ecl_early_ttype_m[3]));
DFFPOSX1 ecl_ttype_e2m_q_reg[4](.D(ecl_ttype_e2m_n7), .CLK(rclk), .Q(ecl_early_ttype_m[4]));
DFFPOSX1 ecl_ttype_e2m_q_reg[5](.D(ecl_ttype_e2m_n5), .CLK(rclk), .Q(ecl_early_ttype_m[5]));
DFFPOSX1 ecl_ttype_e2m_q_reg[6](.D(ecl_ttype_e2m_n3), .CLK(rclk), .Q(ecl_early_ttype_m[6]));
DFFPOSX1 ecl_ttype_e2m_q_reg[7](.D(ecl_ttype_e2m_n19), .CLK(rclk), .Q(ecl_early_ttype_m[7]));
DFFPOSX1 ecl_ttype_e2m_q_reg[8](.D(ecl_ttype_e2m_n17), .CLK(rclk), .Q(ecl_early_ttype_m[8]));
XOR2X1 exu_ecl_ccr_U33(.A(ecl_tid_w[1]), .B(ecl_tid_d[1]), .Y(ecl_ccr_n25));
XOR2X1 exu_ecl_ccr_U32(.A(ecl_tid_w[0]), .B(ecl_tid_d[0]), .Y(ecl_ccr_n26));
NAND2X1 exu_ecl_writeback_U207(.A(exu_n11689), .B(exu_n10553), .Y(ecl_irf_tid_m[0]));
NAND2X1 exu_ecl_writeback_U201(.A(exu_n11686), .B(exu_n10552), .Y(ecl_irf_tid_m[1]));
XOR2X1 exu_ecl_writeback_U191(.A(ecl_tid_w1[0]), .B(ecl_writeback_dfill_tid_g2[0]), .Y(ecl_writeback_n157));
XNOR2X1 exu_ecl_writeback_U190(.A(ecl_writeback_dfill_tid_g2[1]), .B(ecl_tid_w1[1]), .Y(ecl_writeback_n159));
NAND2X1 exu_ecl_writeback_U180(.A(exu_n11680), .B(exu_n10550), .Y(ecl_irf_wen_w));
NAND2X1 exu_ecl_writeback_U149(.A(ecl_writeback_n118), .B(exu_n10549), .Y(exu_ifu_longop_done_g[0]));
NAND2X1 exu_ecl_writeback_U142(.A(ecl_writeback_n111), .B(exu_n10548), .Y(exu_ifu_longop_done_g[1]));
NAND2X1 exu_ecl_writeback_U135(.A(ecl_writeback_n103), .B(exu_n10547), .Y(exu_ifu_longop_done_g[2]));
NAND2X1 exu_ecl_writeback_U129(.A(ecl_writeback_n92), .B(exu_n10546), .Y(exu_ifu_longop_done_g[3]));
NOR2X1 exu_ecl_eccctl_U58(.A(exu_n16273), .B(exu_ifu_ecc_ue_m), .Y(exu_ifu_ecc_ce_m));
NAND2X1 exu_ecl_eccctl_U54(.A(exu_n11672), .B(exu_n10542), .Y(exu_ifu_err_reg_m[5]));
NAND2X1 exu_ecl_eccctl_U51(.A(exu_n11671), .B(exu_n10541), .Y(exu_ifu_err_reg_m[6]));
XOR2X1 exu_ecl_divcntl_U90(.A(div_xin[63]), .B(exu_n15814), .Y(ecl_divcntl_n59));
XOR2X1 exu_ecl_divcntl_U83(.A(exu_n15077), .B(div_ecl_x_msb), .Y(ecl_divcntl_n50));
XOR2X1 exu_ecl_divcntl_U81(.A(ecl_divcntl_subtract), .B(div_ecl_d_msb), .Y(ecl_divcntl_subnext_mux_in1[0]));
XOR2X1 exu_ecl_mdqctl_U94(.A(ecl_tid_w1[0]), .B(ecl_mdqctl_wb_divthr_g[0]), .Y(ecl_mdqctl_n62));
XNOR2X1 exu_ecl_mdqctl_U92(.A(ecl_tid_w1[1]), .B(ecl_mdqctl_wb_divthr_g[1]), .Y(ecl_mdqctl_n61));
XOR2X1 exu_ecl_mdqctl_U81(.A(ecl_tid_w1[0]), .B(ecl_mdqctl_wb_multhr_g[0]), .Y(ecl_mdqctl_n50));
XNOR2X1 exu_ecl_mdqctl_U79(.A(ecl_mdqctl_wb_multhr_g[1]), .B(ecl_tid_w1[1]), .Y(ecl_mdqctl_n49));
XOR2X1 exu_alu_addsub_U65(.A(alu_addsub_subtract_e[31]), .B(div_input_data_e[95]), .Y(alu_ecl_adderin2_31_e));
XOR2X1 exu_alu_addsub_U64(.A(alu_addsub_subtract_e[63]), .B(div_input_data_e[127]), .Y(alu_ecl_adderin2_63_e));
XOR2X1 exu_alu_addsub_U63(.A(alu_addsub_subtract_e[32]), .B(div_input_data_e[96]), .Y(alu_addsub_rs2_data[32]));
XOR2X1 exu_alu_addsub_U62(.A(alu_addsub_subtract_e[33]), .B(div_input_data_e[97]), .Y(alu_addsub_rs2_data[33]));
XOR2X1 exu_alu_addsub_U61(.A(alu_addsub_subtract_e[34]), .B(div_input_data_e[98]), .Y(alu_addsub_rs2_data[34]));
XOR2X1 exu_alu_addsub_U60(.A(alu_addsub_subtract_e[35]), .B(div_input_data_e[99]), .Y(alu_addsub_rs2_data[35]));
XOR2X1 exu_alu_addsub_U59(.A(alu_addsub_subtract_e[36]), .B(div_input_data_e[100]), .Y(alu_addsub_rs2_data[36]));
XOR2X1 exu_alu_addsub_U58(.A(alu_addsub_subtract_e[37]), .B(div_input_data_e[101]), .Y(alu_addsub_rs2_data[37]));
XOR2X1 exu_alu_addsub_U57(.A(alu_addsub_subtract_e[38]), .B(div_input_data_e[102]), .Y(alu_addsub_rs2_data[38]));
XOR2X1 exu_alu_addsub_U56(.A(alu_addsub_subtract_e[39]), .B(div_input_data_e[103]), .Y(alu_addsub_rs2_data[39]));
XOR2X1 exu_alu_addsub_U55(.A(alu_addsub_subtract_e[40]), .B(div_input_data_e[104]), .Y(alu_addsub_rs2_data[40]));
XOR2X1 exu_alu_addsub_U54(.A(alu_addsub_subtract_e[41]), .B(div_input_data_e[105]), .Y(alu_addsub_rs2_data[41]));
XOR2X1 exu_alu_addsub_U53(.A(alu_addsub_subtract_e[42]), .B(div_input_data_e[106]), .Y(alu_addsub_rs2_data[42]));
XOR2X1 exu_alu_addsub_U52(.A(alu_addsub_subtract_e[43]), .B(div_input_data_e[107]), .Y(alu_addsub_rs2_data[43]));
XOR2X1 exu_alu_addsub_U51(.A(alu_addsub_subtract_e[44]), .B(div_input_data_e[108]), .Y(alu_addsub_rs2_data[44]));
XOR2X1 exu_alu_addsub_U50(.A(alu_addsub_subtract_e[45]), .B(div_input_data_e[109]), .Y(alu_addsub_rs2_data[45]));
XOR2X1 exu_alu_addsub_U49(.A(alu_addsub_subtract_e[46]), .B(div_input_data_e[110]), .Y(alu_addsub_rs2_data[46]));
XOR2X1 exu_alu_addsub_U48(.A(alu_addsub_subtract_e[47]), .B(div_input_data_e[111]), .Y(alu_addsub_rs2_data[47]));
XOR2X1 exu_alu_addsub_U47(.A(alu_addsub_subtract_e[48]), .B(div_input_data_e[112]), .Y(alu_addsub_rs2_data[48]));
XOR2X1 exu_alu_addsub_U46(.A(alu_addsub_subtract_e[49]), .B(div_input_data_e[113]), .Y(alu_addsub_rs2_data[49]));
XOR2X1 exu_alu_addsub_U45(.A(alu_addsub_subtract_e[50]), .B(div_input_data_e[114]), .Y(alu_addsub_rs2_data[50]));
XOR2X1 exu_alu_addsub_U44(.A(alu_addsub_subtract_e[51]), .B(div_input_data_e[115]), .Y(alu_addsub_rs2_data[51]));
XOR2X1 exu_alu_addsub_U43(.A(alu_addsub_subtract_e[52]), .B(div_input_data_e[116]), .Y(alu_addsub_rs2_data[52]));
XOR2X1 exu_alu_addsub_U42(.A(alu_addsub_subtract_e[53]), .B(div_input_data_e[117]), .Y(alu_addsub_rs2_data[53]));
XOR2X1 exu_alu_addsub_U41(.A(alu_addsub_subtract_e[54]), .B(div_input_data_e[118]), .Y(alu_addsub_rs2_data[54]));
XOR2X1 exu_alu_addsub_U40(.A(alu_addsub_subtract_e[55]), .B(div_input_data_e[119]), .Y(alu_addsub_rs2_data[55]));
XOR2X1 exu_alu_addsub_U39(.A(alu_addsub_subtract_e[56]), .B(div_input_data_e[120]), .Y(alu_addsub_rs2_data[56]));
XOR2X1 exu_alu_addsub_U38(.A(alu_addsub_subtract_e[57]), .B(div_input_data_e[121]), .Y(alu_addsub_rs2_data[57]));
XOR2X1 exu_alu_addsub_U37(.A(alu_addsub_subtract_e[58]), .B(div_input_data_e[122]), .Y(alu_addsub_rs2_data[58]));
XOR2X1 exu_alu_addsub_U36(.A(alu_addsub_subtract_e[59]), .B(div_input_data_e[123]), .Y(alu_addsub_rs2_data[59]));
XOR2X1 exu_alu_addsub_U35(.A(alu_addsub_subtract_e[60]), .B(div_input_data_e[124]), .Y(alu_addsub_rs2_data[60]));
XOR2X1 exu_alu_addsub_U34(.A(alu_addsub_subtract_e[61]), .B(div_input_data_e[125]), .Y(alu_addsub_rs2_data[61]));
XOR2X1 exu_alu_addsub_U33(.A(alu_addsub_subtract_e[62]), .B(div_input_data_e[126]), .Y(alu_addsub_rs2_data[62]));
XOR2X1 exu_alu_addsub_U32(.A(alu_addsub_subtract_e[0]), .B(div_input_data_e[64]), .Y(alu_addsub_rs2_data_0));
XOR2X1 exu_alu_addsub_U31(.A(alu_addsub_subtract_e[1]), .B(div_input_data_e[65]), .Y(alu_addsub_rs2_data_1));
XOR2X1 exu_alu_addsub_U30(.A(alu_addsub_subtract_e[10]), .B(div_input_data_e[74]), .Y(alu_addsub_rs2_data_10));
XOR2X1 exu_alu_addsub_U29(.A(alu_addsub_subtract_e[11]), .B(div_input_data_e[75]), .Y(alu_addsub_rs2_data_11));
XOR2X1 exu_alu_addsub_U28(.A(alu_addsub_subtract_e[12]), .B(div_input_data_e[76]), .Y(alu_addsub_rs2_data_12));
XOR2X1 exu_alu_addsub_U27(.A(alu_addsub_subtract_e[13]), .B(div_input_data_e[77]), .Y(alu_addsub_rs2_data_13));
XOR2X1 exu_alu_addsub_U26(.A(alu_addsub_subtract_e[14]), .B(div_input_data_e[78]), .Y(alu_addsub_rs2_data_14));
XOR2X1 exu_alu_addsub_U25(.A(alu_addsub_subtract_e[15]), .B(div_input_data_e[79]), .Y(alu_addsub_rs2_data_15));
XOR2X1 exu_alu_addsub_U24(.A(alu_addsub_subtract_e[16]), .B(div_input_data_e[80]), .Y(alu_addsub_rs2_data_16));
XOR2X1 exu_alu_addsub_U23(.A(alu_addsub_subtract_e[17]), .B(div_input_data_e[81]), .Y(alu_addsub_rs2_data_17));
XOR2X1 exu_alu_addsub_U22(.A(alu_addsub_subtract_e[18]), .B(div_input_data_e[82]), .Y(alu_addsub_rs2_data_18));
XOR2X1 exu_alu_addsub_U21(.A(alu_addsub_subtract_e[19]), .B(div_input_data_e[83]), .Y(alu_addsub_rs2_data_19));
XOR2X1 exu_alu_addsub_U20(.A(alu_addsub_subtract_e[2]), .B(div_input_data_e[66]), .Y(alu_addsub_rs2_data_2));
XOR2X1 exu_alu_addsub_U19(.A(alu_addsub_subtract_e[20]), .B(div_input_data_e[84]), .Y(alu_addsub_rs2_data_20));
XOR2X1 exu_alu_addsub_U18(.A(alu_addsub_subtract_e[21]), .B(div_input_data_e[85]), .Y(alu_addsub_rs2_data_21));
XOR2X1 exu_alu_addsub_U17(.A(alu_addsub_subtract_e[22]), .B(div_input_data_e[86]), .Y(alu_addsub_rs2_data_22));
XOR2X1 exu_alu_addsub_U16(.A(alu_addsub_subtract_e[23]), .B(div_input_data_e[87]), .Y(alu_addsub_rs2_data_23));
XOR2X1 exu_alu_addsub_U15(.A(alu_addsub_subtract_e[24]), .B(div_input_data_e[88]), .Y(alu_addsub_rs2_data_24));
XOR2X1 exu_alu_addsub_U14(.A(alu_addsub_subtract_e[25]), .B(div_input_data_e[89]), .Y(alu_addsub_rs2_data_25));
XOR2X1 exu_alu_addsub_U13(.A(alu_addsub_subtract_e[26]), .B(div_input_data_e[90]), .Y(alu_addsub_rs2_data_26));
XOR2X1 exu_alu_addsub_U12(.A(alu_addsub_subtract_e[27]), .B(div_input_data_e[91]), .Y(alu_addsub_rs2_data_27));
XOR2X1 exu_alu_addsub_U11(.A(alu_addsub_subtract_e[28]), .B(div_input_data_e[92]), .Y(alu_addsub_rs2_data_28));
XOR2X1 exu_alu_addsub_U10(.A(alu_addsub_subtract_e[29]), .B(div_input_data_e[93]), .Y(alu_addsub_rs2_data_29));
XOR2X1 exu_alu_addsub_U9(.A(alu_addsub_subtract_e[3]), .B(div_input_data_e[67]), .Y(alu_addsub_rs2_data_3));
XOR2X1 exu_alu_addsub_U8(.A(alu_addsub_subtract_e[30]), .B(div_input_data_e[94]), .Y(alu_addsub_rs2_data_30));
XOR2X1 exu_alu_addsub_U7(.A(alu_addsub_subtract_e[4]), .B(div_input_data_e[68]), .Y(alu_addsub_rs2_data_4));
XOR2X1 exu_alu_addsub_U6(.A(alu_addsub_subtract_e[5]), .B(div_input_data_e[69]), .Y(alu_addsub_rs2_data_5));
XOR2X1 exu_alu_addsub_U5(.A(alu_addsub_subtract_e[6]), .B(div_input_data_e[70]), .Y(alu_addsub_rs2_data_6));
XOR2X1 exu_alu_addsub_U4(.A(alu_addsub_subtract_e[7]), .B(div_input_data_e[71]), .Y(alu_addsub_rs2_data_7));
XOR2X1 exu_alu_addsub_U3(.A(alu_addsub_subtract_e[8]), .B(div_input_data_e[72]), .Y(alu_addsub_rs2_data_8));
XOR2X1 exu_alu_addsub_U2(.A(alu_addsub_subtract_e[9]), .B(div_input_data_e[73]), .Y(alu_addsub_rs2_data_9));
XOR2X1 exu_alu_logic_U352(.A(div_input_data_e[64]), .B(alu_invert_e), .Y(alu_logic_n160));
XOR2X1 exu_alu_logic_U351(.A(div_input_data_e[74]), .B(alu_invert_e), .Y(alu_logic_n159));
XOR2X1 exu_alu_logic_U350(.A(div_input_data_e[75]), .B(exu_n16150), .Y(alu_logic_n158));
XOR2X1 exu_alu_logic_U349(.A(div_input_data_e[76]), .B(alu_invert_e), .Y(alu_logic_n157));
XOR2X1 exu_alu_logic_U348(.A(div_input_data_e[77]), .B(alu_invert_e), .Y(alu_logic_n156));
XOR2X1 exu_alu_logic_U347(.A(div_input_data_e[78]), .B(alu_invert_e), .Y(alu_logic_n155));
XOR2X1 exu_alu_logic_U346(.A(div_input_data_e[79]), .B(exu_n16150), .Y(alu_logic_n154));
XOR2X1 exu_alu_logic_U345(.A(div_input_data_e[80]), .B(alu_invert_e), .Y(alu_logic_n153));
XOR2X1 exu_alu_logic_U344(.A(div_input_data_e[81]), .B(exu_n16150), .Y(alu_logic_n152));
XOR2X1 exu_alu_logic_U343(.A(div_input_data_e[82]), .B(alu_invert_e), .Y(alu_logic_n151));
XOR2X1 exu_alu_logic_U342(.A(div_input_data_e[83]), .B(exu_n16150), .Y(alu_logic_n150));
XOR2X1 exu_alu_logic_U341(.A(div_input_data_e[65]), .B(alu_invert_e), .Y(alu_logic_n149));
XOR2X1 exu_alu_logic_U340(.A(div_input_data_e[84]), .B(alu_invert_e), .Y(alu_logic_n148));
XOR2X1 exu_alu_logic_U339(.A(div_input_data_e[85]), .B(alu_invert_e), .Y(alu_logic_n147));
XOR2X1 exu_alu_logic_U338(.A(div_input_data_e[86]), .B(alu_invert_e), .Y(alu_logic_n146));
XOR2X1 exu_alu_logic_U337(.A(div_input_data_e[87]), .B(alu_invert_e), .Y(alu_logic_n145));
XOR2X1 exu_alu_logic_U336(.A(div_input_data_e[88]), .B(alu_invert_e), .Y(alu_logic_n144));
XOR2X1 exu_alu_logic_U335(.A(div_input_data_e[89]), .B(alu_invert_e), .Y(alu_logic_n143));
XOR2X1 exu_alu_logic_U334(.A(div_input_data_e[90]), .B(alu_invert_e), .Y(alu_logic_n142));
XOR2X1 exu_alu_logic_U333(.A(div_input_data_e[91]), .B(alu_invert_e), .Y(alu_logic_n141));
XOR2X1 exu_alu_logic_U332(.A(div_input_data_e[92]), .B(alu_invert_e), .Y(alu_logic_n140));
XOR2X1 exu_alu_logic_U331(.A(div_input_data_e[93]), .B(alu_invert_e), .Y(alu_logic_n139));
XOR2X1 exu_alu_logic_U330(.A(div_input_data_e[66]), .B(alu_invert_e), .Y(alu_logic_n138));
XOR2X1 exu_alu_logic_U329(.A(div_input_data_e[94]), .B(alu_invert_e), .Y(alu_logic_n137));
XOR2X1 exu_alu_logic_U328(.A(div_input_data_e[95]), .B(alu_invert_e), .Y(alu_logic_n136));
XNOR2X1 exu_alu_logic_U327(.A(exu_n16520), .B(alu_invert_e), .Y(alu_logic_n135));
XNOR2X1 exu_alu_logic_U326(.A(exu_n16521), .B(exu_n16150), .Y(alu_logic_n134));
XNOR2X1 exu_alu_logic_U325(.A(exu_n16522), .B(alu_invert_e), .Y(alu_logic_n133));
XNOR2X1 exu_alu_logic_U324(.A(exu_n16523), .B(exu_n16150), .Y(alu_logic_n132));
XNOR2X1 exu_alu_logic_U323(.A(exu_n16524), .B(exu_n16150), .Y(alu_logic_n131));
XNOR2X1 exu_alu_logic_U322(.A(exu_n16525), .B(exu_n16150), .Y(alu_logic_n130));
XNOR2X1 exu_alu_logic_U321(.A(exu_n16526), .B(exu_n16150), .Y(alu_logic_n129));
XNOR2X1 exu_alu_logic_U320(.A(exu_n16527), .B(exu_n16150), .Y(alu_logic_n128));
XOR2X1 exu_alu_logic_U319(.A(div_input_data_e[67]), .B(alu_invert_e), .Y(alu_logic_n127));
XNOR2X1 exu_alu_logic_U318(.A(exu_n16528), .B(exu_n16150), .Y(alu_logic_n126));
XNOR2X1 exu_alu_logic_U317(.A(exu_n16529), .B(exu_n16150), .Y(alu_logic_n125));
XNOR2X1 exu_alu_logic_U316(.A(exu_n16530), .B(exu_n16150), .Y(alu_logic_n124));
XNOR2X1 exu_alu_logic_U315(.A(exu_n16531), .B(exu_n16150), .Y(alu_logic_n123));
XNOR2X1 exu_alu_logic_U314(.A(exu_n16532), .B(exu_n16150), .Y(alu_logic_n122));
XNOR2X1 exu_alu_logic_U313(.A(exu_n16533), .B(exu_n16150), .Y(alu_logic_n121));
XNOR2X1 exu_alu_logic_U312(.A(exu_n16534), .B(exu_n16150), .Y(alu_logic_n120));
XNOR2X1 exu_alu_logic_U311(.A(exu_n16535), .B(alu_invert_e), .Y(alu_logic_n119));
XNOR2X1 exu_alu_logic_U310(.A(exu_n16536), .B(alu_invert_e), .Y(alu_logic_n118));
XNOR2X1 exu_alu_logic_U309(.A(exu_n16537), .B(alu_invert_e), .Y(alu_logic_n117));
XOR2X1 exu_alu_logic_U308(.A(div_input_data_e[68]), .B(alu_invert_e), .Y(alu_logic_n116));
XNOR2X1 exu_alu_logic_U307(.A(exu_n16538), .B(alu_invert_e), .Y(alu_logic_n115));
XNOR2X1 exu_alu_logic_U306(.A(exu_n16539), .B(alu_invert_e), .Y(alu_logic_n114));
XNOR2X1 exu_alu_logic_U305(.A(exu_n16540), .B(exu_n16150), .Y(alu_logic_n113));
XNOR2X1 exu_alu_logic_U304(.A(exu_n16541), .B(alu_invert_e), .Y(alu_logic_n112));
XNOR2X1 exu_alu_logic_U303(.A(exu_n16542), .B(alu_invert_e), .Y(alu_logic_n111));
XNOR2X1 exu_alu_logic_U302(.A(exu_n16543), .B(alu_invert_e), .Y(alu_logic_n110));
XNOR2X1 exu_alu_logic_U301(.A(exu_n16544), .B(exu_n16150), .Y(alu_logic_n109));
XNOR2X1 exu_alu_logic_U300(.A(exu_n16545), .B(alu_invert_e), .Y(alu_logic_n108));
XNOR2X1 exu_alu_logic_U299(.A(exu_n16546), .B(alu_invert_e), .Y(alu_logic_n107));
XNOR2X1 exu_alu_logic_U298(.A(exu_n16547), .B(alu_invert_e), .Y(alu_logic_n106));
XOR2X1 exu_alu_logic_U297(.A(div_input_data_e[69]), .B(exu_n16150), .Y(alu_logic_n105));
XNOR2X1 exu_alu_logic_U296(.A(exu_n16548), .B(exu_n16150), .Y(alu_logic_n104));
XNOR2X1 exu_alu_logic_U295(.A(exu_n16549), .B(exu_n16150), .Y(alu_logic_n103));
XNOR2X1 exu_alu_logic_U294(.A(exu_n16550), .B(alu_invert_e), .Y(alu_logic_n102));
XNOR2X1 exu_alu_logic_U293(.A(exu_n16551), .B(exu_n16150), .Y(alu_logic_n101));
XOR2X1 exu_alu_logic_U292(.A(div_input_data_e[70]), .B(exu_n16150), .Y(alu_logic_n100));
XOR2X1 exu_alu_logic_U291(.A(div_input_data_e[71]), .B(alu_invert_e), .Y(alu_logic_n99));
XOR2X1 exu_alu_logic_U290(.A(div_input_data_e[72]), .B(exu_n16150), .Y(alu_logic_n98));
XOR2X1 exu_alu_logic_U289(.A(div_input_data_e[73]), .B(alu_invert_e), .Y(alu_logic_n97));
XOR2X1 exu_alu_logic_U288(.A(div_input_data_e[64]), .B(alu_logic_rs1_data_bf1[0]), .Y(alu_logic_n96));
XOR2X1 exu_alu_logic_U287(.A(exu_n16150), .B(alu_logic_n96), .Y(alu_logic_result_xor[0]));
XOR2X1 exu_alu_logic_U286(.A(div_input_data_e[74]), .B(alu_logic_rs1_data_bf1[10]), .Y(alu_logic_n95));
XOR2X1 exu_alu_logic_U285(.A(alu_invert_e), .B(alu_logic_n95), .Y(alu_logic_result_xor[10]));
XOR2X1 exu_alu_logic_U284(.A(div_input_data_e[75]), .B(alu_logic_rs1_data_bf1[11]), .Y(alu_logic_n94));
XOR2X1 exu_alu_logic_U283(.A(alu_invert_e), .B(alu_logic_n94), .Y(alu_logic_result_xor[11]));
XOR2X1 exu_alu_logic_U282(.A(div_input_data_e[76]), .B(alu_logic_rs1_data_bf1[12]), .Y(alu_logic_n93));
XOR2X1 exu_alu_logic_U281(.A(exu_n16150), .B(alu_logic_n93), .Y(alu_logic_result_xor[12]));
XOR2X1 exu_alu_logic_U280(.A(div_input_data_e[77]), .B(alu_logic_rs1_data_bf1[13]), .Y(alu_logic_n92));
XOR2X1 exu_alu_logic_U279(.A(alu_invert_e), .B(alu_logic_n92), .Y(alu_logic_result_xor[13]));
XOR2X1 exu_alu_logic_U278(.A(div_input_data_e[78]), .B(alu_logic_rs1_data_bf1[14]), .Y(alu_logic_n91));
XOR2X1 exu_alu_logic_U277(.A(alu_invert_e), .B(alu_logic_n91), .Y(alu_logic_result_xor[14]));
XOR2X1 exu_alu_logic_U276(.A(div_input_data_e[79]), .B(alu_logic_rs1_data_bf1[15]), .Y(alu_logic_n90));
XOR2X1 exu_alu_logic_U275(.A(exu_n16150), .B(alu_logic_n90), .Y(alu_logic_result_xor[15]));
XOR2X1 exu_alu_logic_U274(.A(div_input_data_e[80]), .B(alu_logic_rs1_data_bf1[16]), .Y(alu_logic_n89));
XOR2X1 exu_alu_logic_U273(.A(alu_invert_e), .B(alu_logic_n89), .Y(alu_logic_result_xor[16]));
XOR2X1 exu_alu_logic_U272(.A(div_input_data_e[81]), .B(alu_logic_rs1_data_bf1[17]), .Y(alu_logic_n88));
XOR2X1 exu_alu_logic_U271(.A(alu_invert_e), .B(alu_logic_n88), .Y(alu_logic_result_xor[17]));
XOR2X1 exu_alu_logic_U270(.A(div_input_data_e[82]), .B(alu_logic_rs1_data_bf1[18]), .Y(alu_logic_n87));
XOR2X1 exu_alu_logic_U269(.A(exu_n16150), .B(alu_logic_n87), .Y(alu_logic_result_xor[18]));
XOR2X1 exu_alu_logic_U268(.A(div_input_data_e[83]), .B(alu_logic_rs1_data_bf1[19]), .Y(alu_logic_n86));
XOR2X1 exu_alu_logic_U267(.A(alu_invert_e), .B(alu_logic_n86), .Y(alu_logic_result_xor[19]));
XOR2X1 exu_alu_logic_U266(.A(div_input_data_e[65]), .B(alu_logic_rs1_data_bf1[1]), .Y(alu_logic_n85));
XOR2X1 exu_alu_logic_U265(.A(alu_invert_e), .B(alu_logic_n85), .Y(alu_logic_result_xor[1]));
XOR2X1 exu_alu_logic_U264(.A(div_input_data_e[84]), .B(alu_logic_rs1_data_bf1[20]), .Y(alu_logic_n84));
XOR2X1 exu_alu_logic_U263(.A(exu_n16150), .B(alu_logic_n84), .Y(alu_logic_result_xor[20]));
XOR2X1 exu_alu_logic_U262(.A(div_input_data_e[85]), .B(alu_logic_rs1_data_bf1[21]), .Y(alu_logic_n83));
XOR2X1 exu_alu_logic_U261(.A(alu_invert_e), .B(alu_logic_n83), .Y(alu_logic_result_xor[21]));
XOR2X1 exu_alu_logic_U260(.A(div_input_data_e[86]), .B(alu_logic_rs1_data_bf1[22]), .Y(alu_logic_n82));
XOR2X1 exu_alu_logic_U259(.A(alu_invert_e), .B(alu_logic_n82), .Y(alu_logic_result_xor[22]));
XOR2X1 exu_alu_logic_U258(.A(div_input_data_e[87]), .B(alu_logic_rs1_data_bf1[23]), .Y(alu_logic_n81));
XOR2X1 exu_alu_logic_U257(.A(alu_invert_e), .B(alu_logic_n81), .Y(alu_logic_result_xor[23]));
XOR2X1 exu_alu_logic_U256(.A(div_input_data_e[88]), .B(alu_logic_rs1_data_bf1[24]), .Y(alu_logic_n80));
XOR2X1 exu_alu_logic_U255(.A(alu_invert_e), .B(alu_logic_n80), .Y(alu_logic_result_xor[24]));
XOR2X1 exu_alu_logic_U254(.A(div_input_data_e[89]), .B(alu_logic_rs1_data_bf1[25]), .Y(alu_logic_n79));
XOR2X1 exu_alu_logic_U253(.A(alu_invert_e), .B(alu_logic_n79), .Y(alu_logic_result_xor[25]));
XOR2X1 exu_alu_logic_U252(.A(div_input_data_e[90]), .B(alu_logic_rs1_data_bf1[26]), .Y(alu_logic_n78));
XOR2X1 exu_alu_logic_U251(.A(exu_n16150), .B(alu_logic_n78), .Y(alu_logic_result_xor[26]));
XOR2X1 exu_alu_logic_U250(.A(div_input_data_e[91]), .B(alu_logic_rs1_data_bf1[27]), .Y(alu_logic_n77));
XOR2X1 exu_alu_logic_U249(.A(exu_n16150), .B(alu_logic_n77), .Y(alu_logic_result_xor[27]));
XOR2X1 exu_alu_logic_U248(.A(div_input_data_e[92]), .B(alu_logic_rs1_data_bf1[28]), .Y(alu_logic_n76));
XOR2X1 exu_alu_logic_U247(.A(exu_n16150), .B(alu_logic_n76), .Y(alu_logic_result_xor[28]));
XOR2X1 exu_alu_logic_U246(.A(div_input_data_e[93]), .B(alu_logic_rs1_data_bf1[29]), .Y(alu_logic_n75));
XOR2X1 exu_alu_logic_U245(.A(alu_invert_e), .B(alu_logic_n75), .Y(alu_logic_result_xor[29]));
XOR2X1 exu_alu_logic_U244(.A(div_input_data_e[66]), .B(alu_logic_rs1_data_bf1[2]), .Y(alu_logic_n74));
XOR2X1 exu_alu_logic_U243(.A(alu_invert_e), .B(alu_logic_n74), .Y(alu_logic_result_xor[2]));
XOR2X1 exu_alu_logic_U242(.A(div_input_data_e[94]), .B(alu_logic_rs1_data_bf1[30]), .Y(alu_logic_n73));
XOR2X1 exu_alu_logic_U241(.A(alu_invert_e), .B(alu_logic_n73), .Y(alu_logic_result_xor[30]));
XOR2X1 exu_alu_logic_U240(.A(div_input_data_e[95]), .B(alu_logic_rs1_data_bf1[31]), .Y(alu_logic_n72));
XOR2X1 exu_alu_logic_U239(.A(alu_invert_e), .B(alu_logic_n72), .Y(alu_logic_result_xor[31]));
XOR2X1 exu_alu_logic_U238(.A(div_input_data_e[96]), .B(alu_logic_rs1_data_bf1[32]), .Y(alu_logic_n71));
XOR2X1 exu_alu_logic_U237(.A(alu_invert_e), .B(alu_logic_n71), .Y(alu_logic_result_xor[32]));
XOR2X1 exu_alu_logic_U236(.A(div_input_data_e[97]), .B(alu_logic_rs1_data_bf1[33]), .Y(alu_logic_n70));
XOR2X1 exu_alu_logic_U235(.A(alu_invert_e), .B(alu_logic_n70), .Y(alu_logic_result_xor[33]));
XOR2X1 exu_alu_logic_U234(.A(div_input_data_e[98]), .B(alu_logic_rs1_data_bf1[34]), .Y(alu_logic_n69));
XOR2X1 exu_alu_logic_U233(.A(alu_invert_e), .B(alu_logic_n69), .Y(alu_logic_result_xor[34]));
XOR2X1 exu_alu_logic_U232(.A(div_input_data_e[99]), .B(alu_logic_rs1_data_bf1[35]), .Y(alu_logic_n68));
XOR2X1 exu_alu_logic_U231(.A(exu_n16150), .B(alu_logic_n68), .Y(alu_logic_result_xor[35]));
XOR2X1 exu_alu_logic_U230(.A(div_input_data_e[100]), .B(alu_logic_rs1_data_bf1[36]), .Y(alu_logic_n67));
XOR2X1 exu_alu_logic_U229(.A(alu_invert_e), .B(alu_logic_n67), .Y(alu_logic_result_xor[36]));
XOR2X1 exu_alu_logic_U228(.A(div_input_data_e[101]), .B(alu_logic_rs1_data_bf1[37]), .Y(alu_logic_n66));
XOR2X1 exu_alu_logic_U227(.A(exu_n16150), .B(alu_logic_n66), .Y(alu_logic_result_xor[37]));
XOR2X1 exu_alu_logic_U226(.A(div_input_data_e[102]), .B(alu_logic_rs1_data_bf1[38]), .Y(alu_logic_n65));
XOR2X1 exu_alu_logic_U225(.A(alu_invert_e), .B(alu_logic_n65), .Y(alu_logic_result_xor[38]));
XOR2X1 exu_alu_logic_U224(.A(div_input_data_e[103]), .B(alu_logic_rs1_data_bf1[39]), .Y(alu_logic_n64));
XOR2X1 exu_alu_logic_U223(.A(alu_invert_e), .B(alu_logic_n64), .Y(alu_logic_result_xor[39]));
XOR2X1 exu_alu_logic_U222(.A(div_input_data_e[67]), .B(alu_logic_rs1_data_bf1[3]), .Y(alu_logic_n63));
XOR2X1 exu_alu_logic_U221(.A(alu_invert_e), .B(alu_logic_n63), .Y(alu_logic_result_xor[3]));
XOR2X1 exu_alu_logic_U220(.A(div_input_data_e[104]), .B(alu_logic_rs1_data_bf1[40]), .Y(alu_logic_n62));
XOR2X1 exu_alu_logic_U219(.A(alu_invert_e), .B(alu_logic_n62), .Y(alu_logic_result_xor[40]));
XOR2X1 exu_alu_logic_U218(.A(div_input_data_e[105]), .B(alu_logic_rs1_data_bf1[41]), .Y(alu_logic_n61));
XOR2X1 exu_alu_logic_U217(.A(alu_invert_e), .B(alu_logic_n61), .Y(alu_logic_result_xor[41]));
XOR2X1 exu_alu_logic_U216(.A(div_input_data_e[106]), .B(alu_logic_rs1_data_bf1[42]), .Y(alu_logic_n60));
XOR2X1 exu_alu_logic_U215(.A(exu_n16150), .B(alu_logic_n60), .Y(alu_logic_result_xor[42]));
XOR2X1 exu_alu_logic_U214(.A(div_input_data_e[107]), .B(alu_logic_rs1_data_bf1[43]), .Y(alu_logic_n59));
XOR2X1 exu_alu_logic_U213(.A(alu_invert_e), .B(alu_logic_n59), .Y(alu_logic_result_xor[43]));
XOR2X1 exu_alu_logic_U212(.A(div_input_data_e[108]), .B(alu_logic_rs1_data_bf1[44]), .Y(alu_logic_n58));
XOR2X1 exu_alu_logic_U211(.A(alu_invert_e), .B(alu_logic_n58), .Y(alu_logic_result_xor[44]));
XOR2X1 exu_alu_logic_U210(.A(div_input_data_e[109]), .B(alu_logic_rs1_data_bf1[45]), .Y(alu_logic_n57));
XOR2X1 exu_alu_logic_U209(.A(alu_invert_e), .B(alu_logic_n57), .Y(alu_logic_result_xor[45]));
XOR2X1 exu_alu_logic_U208(.A(div_input_data_e[110]), .B(alu_logic_rs1_data_bf1[46]), .Y(alu_logic_n56));
XOR2X1 exu_alu_logic_U207(.A(alu_invert_e), .B(alu_logic_n56), .Y(alu_logic_result_xor[46]));
XOR2X1 exu_alu_logic_U206(.A(div_input_data_e[111]), .B(alu_logic_rs1_data_bf1[47]), .Y(alu_logic_n55));
XOR2X1 exu_alu_logic_U205(.A(alu_invert_e), .B(alu_logic_n55), .Y(alu_logic_result_xor[47]));
XOR2X1 exu_alu_logic_U204(.A(div_input_data_e[112]), .B(alu_logic_rs1_data_bf1[48]), .Y(alu_logic_n54));
XOR2X1 exu_alu_logic_U203(.A(alu_invert_e), .B(alu_logic_n54), .Y(alu_logic_result_xor[48]));
XOR2X1 exu_alu_logic_U202(.A(div_input_data_e[113]), .B(alu_logic_rs1_data_bf1[49]), .Y(alu_logic_n53));
XOR2X1 exu_alu_logic_U201(.A(exu_n16150), .B(alu_logic_n53), .Y(alu_logic_result_xor[49]));
XOR2X1 exu_alu_logic_U200(.A(div_input_data_e[68]), .B(alu_logic_rs1_data_bf1[4]), .Y(alu_logic_n52));
XOR2X1 exu_alu_logic_U199(.A(alu_invert_e), .B(alu_logic_n52), .Y(alu_logic_result_xor[4]));
XOR2X1 exu_alu_logic_U198(.A(div_input_data_e[114]), .B(alu_logic_rs1_data_bf1[50]), .Y(alu_logic_n51));
XOR2X1 exu_alu_logic_U197(.A(exu_n16150), .B(alu_logic_n51), .Y(alu_logic_result_xor[50]));
XOR2X1 exu_alu_logic_U196(.A(div_input_data_e[115]), .B(alu_logic_rs1_data_bf1[51]), .Y(alu_logic_n50));
XOR2X1 exu_alu_logic_U195(.A(exu_n16150), .B(alu_logic_n50), .Y(alu_logic_result_xor[51]));
XOR2X1 exu_alu_logic_U194(.A(div_input_data_e[116]), .B(alu_logic_rs1_data_bf1[52]), .Y(alu_logic_n49));
XOR2X1 exu_alu_logic_U193(.A(alu_invert_e), .B(alu_logic_n49), .Y(alu_logic_result_xor[52]));
XOR2X1 exu_alu_logic_U192(.A(div_input_data_e[117]), .B(alu_logic_rs1_data_bf1[53]), .Y(alu_logic_n48));
XOR2X1 exu_alu_logic_U191(.A(alu_invert_e), .B(alu_logic_n48), .Y(alu_logic_result_xor[53]));
XOR2X1 exu_alu_logic_U190(.A(div_input_data_e[118]), .B(alu_logic_rs1_data_bf1[54]), .Y(alu_logic_n47));
XOR2X1 exu_alu_logic_U189(.A(alu_invert_e), .B(alu_logic_n47), .Y(alu_logic_result_xor[54]));
XOR2X1 exu_alu_logic_U188(.A(div_input_data_e[119]), .B(alu_logic_rs1_data_bf1[55]), .Y(alu_logic_n46));
XOR2X1 exu_alu_logic_U187(.A(alu_invert_e), .B(alu_logic_n46), .Y(alu_logic_result_xor[55]));
XOR2X1 exu_alu_logic_U186(.A(div_input_data_e[120]), .B(alu_logic_rs1_data_bf1[56]), .Y(alu_logic_n45));
XOR2X1 exu_alu_logic_U185(.A(alu_invert_e), .B(alu_logic_n45), .Y(alu_logic_result_xor[56]));
XOR2X1 exu_alu_logic_U184(.A(div_input_data_e[121]), .B(alu_logic_rs1_data_bf1[57]), .Y(alu_logic_n44));
XOR2X1 exu_alu_logic_U183(.A(exu_n16150), .B(alu_logic_n44), .Y(alu_logic_result_xor[57]));
XOR2X1 exu_alu_logic_U182(.A(div_input_data_e[122]), .B(alu_logic_rs1_data_bf1[58]), .Y(alu_logic_n43));
XOR2X1 exu_alu_logic_U181(.A(exu_n16150), .B(alu_logic_n43), .Y(alu_logic_result_xor[58]));
XOR2X1 exu_alu_logic_U180(.A(div_input_data_e[123]), .B(alu_logic_rs1_data_bf1[59]), .Y(alu_logic_n42));
XOR2X1 exu_alu_logic_U179(.A(exu_n16150), .B(alu_logic_n42), .Y(alu_logic_result_xor[59]));
XOR2X1 exu_alu_logic_U178(.A(div_input_data_e[69]), .B(alu_logic_rs1_data_bf1[5]), .Y(alu_logic_n41));
XOR2X1 exu_alu_logic_U177(.A(alu_invert_e), .B(alu_logic_n41), .Y(alu_logic_result_xor[5]));
XOR2X1 exu_alu_logic_U176(.A(div_input_data_e[124]), .B(alu_logic_rs1_data_bf1[60]), .Y(alu_logic_n40));
XOR2X1 exu_alu_logic_U175(.A(alu_invert_e), .B(alu_logic_n40), .Y(alu_logic_result_xor[60]));
XOR2X1 exu_alu_logic_U174(.A(div_input_data_e[125]), .B(alu_logic_rs1_data_bf1[61]), .Y(alu_logic_n39));
XOR2X1 exu_alu_logic_U173(.A(alu_invert_e), .B(alu_logic_n39), .Y(alu_logic_result_xor[61]));
XOR2X1 exu_alu_logic_U172(.A(div_input_data_e[126]), .B(alu_logic_rs1_data_bf1[62]), .Y(alu_logic_n38));
XOR2X1 exu_alu_logic_U171(.A(alu_invert_e), .B(alu_logic_n38), .Y(alu_logic_result_xor[62]));
XOR2X1 exu_alu_logic_U170(.A(div_input_data_e[127]), .B(alu_logic_rs1_data_bf1[63]), .Y(alu_logic_n37));
XOR2X1 exu_alu_logic_U169(.A(alu_invert_e), .B(alu_logic_n37), .Y(alu_logic_result_xor[63]));
XOR2X1 exu_alu_logic_U168(.A(div_input_data_e[70]), .B(alu_logic_rs1_data_bf1[6]), .Y(alu_logic_n36));
XOR2X1 exu_alu_logic_U167(.A(alu_invert_e), .B(alu_logic_n36), .Y(alu_logic_result_xor[6]));
XOR2X1 exu_alu_logic_U166(.A(div_input_data_e[71]), .B(alu_logic_rs1_data_bf1[7]), .Y(alu_logic_n35));
XOR2X1 exu_alu_logic_U165(.A(alu_invert_e), .B(alu_logic_n35), .Y(alu_logic_result_xor[7]));
XOR2X1 exu_alu_logic_U164(.A(div_input_data_e[72]), .B(alu_logic_rs1_data_bf1[8]), .Y(alu_logic_n34));
XOR2X1 exu_alu_logic_U163(.A(alu_invert_e), .B(alu_logic_n34), .Y(alu_logic_result_xor[8]));
XOR2X1 exu_alu_logic_U162(.A(div_input_data_e[73]), .B(alu_logic_rs1_data_bf1[9]), .Y(alu_logic_n33));
XOR2X1 exu_alu_logic_U161(.A(exu_n16150), .B(alu_logic_n33), .Y(alu_logic_result_xor[9]));
XNOR2X1 exu_alu_chk_mem_addr_U31(.A(exu_n15505), .B(exu_n15504), .Y(alu_chk_mem_addr_n29));
XNOR2X1 exu_alu_chk_mem_addr_U30(.A(exu_n15479), .B(exu_n15505), .Y(alu_chk_mem_addr_n30));
XNOR2X1 exu_alu_chk_mem_addr_U28(.A(exu_n15479), .B(exu_lsu_ldst_va_e[47]), .Y(alu_chk_mem_addr_n27));
XNOR2X1 exu_alu_chk_mem_addr_U27(.A(exu_n15494), .B(exu_n15118), .Y(alu_chk_mem_addr_n28));
XNOR2X1 exu_alu_chk_mem_addr_U24(.A(exu_n15501), .B(exu_n15500), .Y(alu_chk_mem_addr_n23));
XNOR2X1 exu_alu_chk_mem_addr_U23(.A(exu_n15502), .B(exu_n15501), .Y(alu_chk_mem_addr_n24));
XNOR2X1 exu_alu_chk_mem_addr_U21(.A(exu_n15503), .B(exu_n15502), .Y(alu_chk_mem_addr_n21));
XNOR2X1 exu_alu_chk_mem_addr_U20(.A(exu_n15504), .B(exu_n15503), .Y(alu_chk_mem_addr_n22));
XNOR2X1 exu_alu_chk_mem_addr_U16(.A(exu_n15478), .B(exu_n15498), .Y(alu_chk_mem_addr_n15));
XNOR2X1 exu_alu_chk_mem_addr_U15(.A(exu_n15478), .B(exu_n15546), .Y(alu_chk_mem_addr_n16));
XNOR2X1 exu_alu_chk_mem_addr_U13(.A(exu_n15499), .B(exu_n15546), .Y(alu_chk_mem_addr_n13));
XNOR2X1 exu_alu_chk_mem_addr_U12(.A(exu_n15500), .B(exu_n15499), .Y(alu_chk_mem_addr_n14));
XNOR2X1 exu_alu_chk_mem_addr_U9(.A(exu_n15495), .B(exu_n15494), .Y(alu_chk_mem_addr_n9));
XNOR2X1 exu_alu_chk_mem_addr_U8(.A(exu_n15496), .B(exu_n15495), .Y(alu_chk_mem_addr_n10));
XNOR2X1 exu_alu_chk_mem_addr_U6(.A(exu_n15497), .B(exu_n15496), .Y(alu_chk_mem_addr_n7));
XNOR2X1 exu_alu_chk_mem_addr_U5(.A(exu_n15498), .B(exu_n15497), .Y(alu_chk_mem_addr_n8));
XOR2X1 exu_div_u32eql_U32(.A(exu_n15526), .B(exu_n15527), .Y(div_u32eql_inxor[11]));
XOR2X1 exu_div_u32eql_U31(.A(exu_n15527), .B(exu_n15528), .Y(div_u32eql_inxor[12]));
XOR2X1 exu_div_u32eql_U30(.A(exu_n15528), .B(exu_n15529), .Y(div_u32eql_inxor[13]));
XOR2X1 exu_div_u32eql_U29(.A(exu_n15529), .B(exu_n15530), .Y(div_u32eql_inxor[14]));
XOR2X1 exu_div_u32eql_U28(.A(exu_n15530), .B(exu_n15531), .Y(div_u32eql_inxor[15]));
XOR2X1 exu_div_u32eql_U27(.A(exu_n15531), .B(exu_n15532), .Y(div_u32eql_inxor[16]));
XOR2X1 exu_div_u32eql_U26(.A(exu_n15532), .B(exu_n15533), .Y(div_u32eql_inxor[17]));
XOR2X1 exu_div_u32eql_U25(.A(exu_n15533), .B(exu_n15534), .Y(div_u32eql_inxor[18]));
XOR2X1 exu_div_u32eql_U24(.A(exu_n15534), .B(exu_n15535), .Y(div_u32eql_inxor[19]));
XOR2X1 exu_div_u32eql_U23(.A(exu_n15419), .B(exu_n15517), .Y(div_u32eql_inxor[1]));
XOR2X1 exu_div_u32eql_U22(.A(exu_n15535), .B(exu_n15536), .Y(div_u32eql_inxor[20]));
XOR2X1 exu_div_u32eql_U21(.A(exu_n15536), .B(exu_n15549), .Y(div_u32eql_inxor[21]));
XOR2X1 exu_div_u32eql_U20(.A(exu_n15512), .B(exu_n15549), .Y(div_u32eql_inxor[22]));
XOR2X1 exu_div_u32eql_U19(.A(exu_n15512), .B(exu_n15537), .Y(div_u32eql_inxor[23]));
XOR2X1 exu_div_u32eql_U18(.A(exu_n15537), .B(exu_n15538), .Y(div_u32eql_inxor[24]));
XOR2X1 exu_div_u32eql_U17(.A(exu_n15538), .B(exu_n15539), .Y(div_u32eql_inxor[25]));
XOR2X1 exu_div_u32eql_U16(.A(exu_n15539), .B(exu_n15540), .Y(div_u32eql_inxor[26]));
XOR2X1 exu_div_u32eql_U15(.A(exu_n15540), .B(exu_n15541), .Y(div_u32eql_inxor[27]));
XOR2X1 exu_div_u32eql_U14(.A(exu_n15541), .B(exu_n15542), .Y(div_u32eql_inxor[28]));
XOR2X1 exu_div_u32eql_U13(.A(exu_n15542), .B(exu_n15543), .Y(div_u32eql_inxor[29]));
XOR2X1 exu_div_u32eql_U12(.A(exu_n15517), .B(exu_n15518), .Y(div_u32eql_inxor[2]));
XOR2X1 exu_div_u32eql_U11(.A(exu_n15543), .B(exu_n15544), .Y(div_u32eql_inxor[30]));
XOR2X1 exu_div_u32eql_U10(.A(exu_n15544), .B(exu_n15187), .Y(div_u32eql_inxor[31]));
XOR2X1 exu_div_u32eql_U9(.A(exu_n15518), .B(exu_n15519), .Y(div_u32eql_inxor[3]));
XOR2X1 exu_div_u32eql_U8(.A(exu_n15519), .B(exu_n15520), .Y(div_u32eql_inxor[4]));
XOR2X1 exu_div_u32eql_U7(.A(exu_n15520), .B(exu_n15521), .Y(div_u32eql_inxor[5]));
XOR2X1 exu_div_u32eql_U6(.A(exu_n15521), .B(exu_n15522), .Y(div_u32eql_inxor[6]));
XOR2X1 exu_div_u32eql_U5(.A(exu_n15522), .B(exu_n15523), .Y(div_u32eql_inxor[7]));
XOR2X1 exu_div_u32eql_U4(.A(exu_n15523), .B(exu_n15524), .Y(div_u32eql_inxor[8]));
XOR2X1 exu_div_u32eql_U3(.A(exu_n15524), .B(exu_n15525), .Y(div_u32eql_inxor[9]));
DFFPOSX1 div_d_dff_q_reg[0](.D(div_d_dff_n155), .CLK(rclk), .Q(div_d[0]));
DFFPOSX1 div_d_dff_q_reg[1](.D(div_d_dff_n133), .CLK(rclk), .Q(div_d[1]));
DFFPOSX1 div_d_dff_q_reg[2](.D(div_d_dff_n111), .CLK(rclk), .Q(div_d[2]));
DFFPOSX1 div_d_dff_q_reg[3](.D(div_d_dff_n89), .CLK(rclk), .Q(div_d[3]));
DFFPOSX1 div_d_dff_q_reg[4](.D(div_d_dff_n67), .CLK(rclk), .Q(div_d[4]));
DFFPOSX1 div_d_dff_q_reg[5](.D(div_d_dff_n45), .CLK(rclk), .Q(div_d[5]));
DFFPOSX1 div_d_dff_q_reg[6](.D(div_d_dff_n23), .CLK(rclk), .Q(div_d[6]));
DFFPOSX1 div_d_dff_q_reg[7](.D(div_d_dff_n257), .CLK(rclk), .Q(div_d[7]));
DFFPOSX1 div_d_dff_q_reg[8](.D(div_d_dff_n235), .CLK(rclk), .Q(div_d[8]));
DFFPOSX1 div_d_dff_q_reg[9](.D(div_d_dff_n213), .CLK(rclk), .Q(div_d[9]));
DFFPOSX1 div_d_dff_q_reg[10](.D(div_d_dff_n191), .CLK(rclk), .Q(div_d[10]));
DFFPOSX1 div_d_dff_q_reg[11](.D(div_d_dff_n187), .CLK(rclk), .Q(div_d[11]));
DFFPOSX1 div_d_dff_q_reg[12](.D(div_d_dff_n185), .CLK(rclk), .Q(div_d[12]));
DFFPOSX1 div_d_dff_q_reg[13](.D(div_d_dff_n183), .CLK(rclk), .Q(div_d[13]));
DFFPOSX1 div_d_dff_q_reg[14](.D(div_d_dff_n181), .CLK(rclk), .Q(div_d[14]));
DFFPOSX1 div_d_dff_q_reg[15](.D(div_d_dff_n179), .CLK(rclk), .Q(div_d[15]));
DFFPOSX1 div_d_dff_q_reg[16](.D(div_d_dff_n177), .CLK(rclk), .Q(div_d[16]));
DFFPOSX1 div_d_dff_q_reg[17](.D(div_d_dff_n175), .CLK(rclk), .Q(div_d[17]));
DFFPOSX1 div_d_dff_q_reg[18](.D(div_d_dff_n173), .CLK(rclk), .Q(div_d[18]));
DFFPOSX1 div_d_dff_q_reg[19](.D(div_d_dff_n171), .CLK(rclk), .Q(div_d[19]));
DFFPOSX1 div_d_dff_q_reg[20](.D(div_d_dff_n169), .CLK(rclk), .Q(div_d[20]));
DFFPOSX1 div_d_dff_q_reg[21](.D(div_d_dff_n167), .CLK(rclk), .Q(div_d[21]));
DFFPOSX1 div_d_dff_q_reg[22](.D(div_d_dff_n165), .CLK(rclk), .Q(div_d[22]));
DFFPOSX1 div_d_dff_q_reg[23](.D(div_d_dff_n163), .CLK(rclk), .Q(div_d[23]));
DFFPOSX1 div_d_dff_q_reg[24](.D(div_d_dff_n161), .CLK(rclk), .Q(div_d[24]));
DFFPOSX1 div_d_dff_q_reg[25](.D(div_d_dff_n159), .CLK(rclk), .Q(div_d[25]));
DFFPOSX1 div_d_dff_q_reg[26](.D(div_d_dff_n157), .CLK(rclk), .Q(div_d[26]));
DFFPOSX1 div_d_dff_q_reg[27](.D(div_d_dff_n153), .CLK(rclk), .Q(div_d[27]));
DFFPOSX1 div_d_dff_q_reg[28](.D(div_d_dff_n151), .CLK(rclk), .Q(div_d[28]));
DFFPOSX1 div_d_dff_q_reg[29](.D(div_d_dff_n149), .CLK(rclk), .Q(div_d[29]));
DFFPOSX1 div_d_dff_q_reg[30](.D(div_d_dff_n147), .CLK(rclk), .Q(div_d[30]));
DFFPOSX1 div_d_dff_q_reg[31](.D(div_d_dff_n145), .CLK(rclk), .Q(div_d[31]));
DFFPOSX1 div_d_dff_q_reg[32](.D(div_d_dff_n143), .CLK(rclk), .Q(div_d[32]));
DFFPOSX1 div_d_dff_q_reg[33](.D(div_d_dff_n141), .CLK(rclk), .Q(div_d[33]));
DFFPOSX1 div_d_dff_q_reg[34](.D(div_d_dff_n139), .CLK(rclk), .Q(div_d[34]));
DFFPOSX1 div_d_dff_q_reg[35](.D(div_d_dff_n137), .CLK(rclk), .Q(div_d[35]));
DFFPOSX1 div_d_dff_q_reg[36](.D(div_d_dff_n135), .CLK(rclk), .Q(div_d[36]));
DFFPOSX1 div_d_dff_q_reg[37](.D(div_d_dff_n131), .CLK(rclk), .Q(div_d[37]));
DFFPOSX1 div_d_dff_q_reg[38](.D(div_d_dff_n129), .CLK(rclk), .Q(div_d[38]));
DFFPOSX1 div_d_dff_q_reg[39](.D(div_d_dff_n127), .CLK(rclk), .Q(div_d[39]));
DFFPOSX1 div_d_dff_q_reg[40](.D(div_d_dff_n125), .CLK(rclk), .Q(div_d[40]));
DFFPOSX1 div_d_dff_q_reg[41](.D(div_d_dff_n123), .CLK(rclk), .Q(div_d[41]));
DFFPOSX1 div_d_dff_q_reg[42](.D(div_d_dff_n121), .CLK(rclk), .Q(div_d[42]));
DFFPOSX1 div_d_dff_q_reg[43](.D(div_d_dff_n119), .CLK(rclk), .Q(div_d[43]));
DFFPOSX1 div_d_dff_q_reg[44](.D(div_d_dff_n117), .CLK(rclk), .Q(div_d[44]));
DFFPOSX1 div_d_dff_q_reg[45](.D(div_d_dff_n115), .CLK(rclk), .Q(div_d[45]));
DFFPOSX1 div_d_dff_q_reg[46](.D(div_d_dff_n113), .CLK(rclk), .Q(div_d[46]));
DFFPOSX1 div_d_dff_q_reg[47](.D(div_d_dff_n109), .CLK(rclk), .Q(div_d[47]));
DFFPOSX1 div_d_dff_q_reg[48](.D(div_d_dff_n107), .CLK(rclk), .Q(div_d[48]));
DFFPOSX1 div_d_dff_q_reg[49](.D(div_d_dff_n105), .CLK(rclk), .Q(div_d[49]));
DFFPOSX1 div_d_dff_q_reg[50](.D(div_d_dff_n103), .CLK(rclk), .Q(div_d[50]));
DFFPOSX1 div_d_dff_q_reg[51](.D(div_d_dff_n101), .CLK(rclk), .Q(div_d[51]));
DFFPOSX1 div_d_dff_q_reg[52](.D(div_d_dff_n99), .CLK(rclk), .Q(div_d[52]));
DFFPOSX1 div_d_dff_q_reg[53](.D(div_d_dff_n97), .CLK(rclk), .Q(div_d[53]));
DFFPOSX1 div_d_dff_q_reg[54](.D(div_d_dff_n95), .CLK(rclk), .Q(div_d[54]));
DFFPOSX1 div_d_dff_q_reg[55](.D(div_d_dff_n93), .CLK(rclk), .Q(div_d[55]));
DFFPOSX1 div_d_dff_q_reg[56](.D(div_d_dff_n91), .CLK(rclk), .Q(div_d[56]));
DFFPOSX1 div_d_dff_q_reg[57](.D(div_d_dff_n87), .CLK(rclk), .Q(div_d[57]));
DFFPOSX1 div_d_dff_q_reg[58](.D(div_d_dff_n85), .CLK(rclk), .Q(div_d[58]));
DFFPOSX1 div_d_dff_q_reg[59](.D(div_d_dff_n83), .CLK(rclk), .Q(div_d[59]));
DFFPOSX1 div_d_dff_q_reg[60](.D(div_d_dff_n81), .CLK(rclk), .Q(div_d[60]));
DFFPOSX1 div_d_dff_q_reg[61](.D(div_d_dff_n79), .CLK(rclk), .Q(div_d[61]));
DFFPOSX1 div_d_dff_q_reg[62](.D(div_d_dff_n77), .CLK(rclk), .Q(div_ecl_d_62));
DFFPOSX1 div_d_dff_q_reg[63](.D(div_d_dff_n75), .CLK(rclk), .Q(div_d_63));
DFFPOSX1 div_d_dff_q_reg[64](.D(div_d_dff_n73), .CLK(rclk), .Q(div_curr_q[0]));
DFFPOSX1 div_d_dff_q_reg[65](.D(div_d_dff_n71), .CLK(rclk), .Q(div_curr_q[1]));
DFFPOSX1 div_d_dff_q_reg[66](.D(div_d_dff_n69), .CLK(rclk), .Q(div_curr_q[2]));
DFFPOSX1 div_d_dff_q_reg[67](.D(div_d_dff_n65), .CLK(rclk), .Q(div_curr_q[3]));
DFFPOSX1 div_d_dff_q_reg[68](.D(div_d_dff_n63), .CLK(rclk), .Q(div_curr_q[4]));
DFFPOSX1 div_d_dff_q_reg[69](.D(div_d_dff_n61), .CLK(rclk), .Q(div_curr_q[5]));
DFFPOSX1 div_d_dff_q_reg[70](.D(div_d_dff_n59), .CLK(rclk), .Q(div_curr_q[6]));
DFFPOSX1 div_d_dff_q_reg[71](.D(div_d_dff_n57), .CLK(rclk), .Q(div_curr_q[7]));
DFFPOSX1 div_d_dff_q_reg[72](.D(div_d_dff_n55), .CLK(rclk), .Q(div_curr_q[8]));
DFFPOSX1 div_d_dff_q_reg[73](.D(div_d_dff_n53), .CLK(rclk), .Q(div_curr_q[9]));
DFFPOSX1 div_d_dff_q_reg[74](.D(div_d_dff_n51), .CLK(rclk), .Q(div_curr_q[10]));
DFFPOSX1 div_d_dff_q_reg[75](.D(div_d_dff_n49), .CLK(rclk), .Q(div_curr_q[11]));
DFFPOSX1 div_d_dff_q_reg[76](.D(div_d_dff_n47), .CLK(rclk), .Q(div_curr_q[12]));
DFFPOSX1 div_d_dff_q_reg[77](.D(div_d_dff_n43), .CLK(rclk), .Q(div_curr_q[13]));
DFFPOSX1 div_d_dff_q_reg[78](.D(div_d_dff_n41), .CLK(rclk), .Q(div_curr_q[14]));
DFFPOSX1 div_d_dff_q_reg[79](.D(div_d_dff_n39), .CLK(rclk), .Q(div_curr_q[15]));
DFFPOSX1 div_d_dff_q_reg[80](.D(div_d_dff_n37), .CLK(rclk), .Q(div_curr_q[16]));
DFFPOSX1 div_d_dff_q_reg[81](.D(div_d_dff_n35), .CLK(rclk), .Q(div_curr_q[17]));
DFFPOSX1 div_d_dff_q_reg[82](.D(div_d_dff_n33), .CLK(rclk), .Q(div_curr_q[18]));
DFFPOSX1 div_d_dff_q_reg[83](.D(div_d_dff_n31), .CLK(rclk), .Q(div_curr_q[19]));
DFFPOSX1 div_d_dff_q_reg[84](.D(div_d_dff_n29), .CLK(rclk), .Q(div_curr_q[20]));
DFFPOSX1 div_d_dff_q_reg[85](.D(div_d_dff_n27), .CLK(rclk), .Q(div_curr_q[21]));
DFFPOSX1 div_d_dff_q_reg[86](.D(div_d_dff_n25), .CLK(rclk), .Q(div_curr_q[22]));
DFFPOSX1 div_d_dff_q_reg[87](.D(div_d_dff_n21), .CLK(rclk), .Q(div_curr_q[23]));
DFFPOSX1 div_d_dff_q_reg[88](.D(div_d_dff_n19), .CLK(rclk), .Q(div_curr_q[24]));
DFFPOSX1 div_d_dff_q_reg[89](.D(div_d_dff_n17), .CLK(rclk), .Q(div_curr_q[25]));
DFFPOSX1 div_d_dff_q_reg[90](.D(div_d_dff_n15), .CLK(rclk), .Q(div_curr_q[26]));
DFFPOSX1 div_d_dff_q_reg[91](.D(div_d_dff_n13), .CLK(rclk), .Q(div_curr_q[27]));
DFFPOSX1 div_d_dff_q_reg[92](.D(div_d_dff_n11), .CLK(rclk), .Q(div_curr_q[28]));
DFFPOSX1 div_d_dff_q_reg[93](.D(div_d_dff_n9), .CLK(rclk), .Q(div_curr_q[29]));
DFFPOSX1 div_d_dff_q_reg[94](.D(div_d_dff_n7), .CLK(rclk), .Q(div_curr_q[30]));
DFFPOSX1 div_d_dff_q_reg[95](.D(div_d_dff_n5), .CLK(rclk), .Q(div_curr_q[31]));
DFFPOSX1 div_d_dff_q_reg[96](.D(div_d_dff_n3), .CLK(rclk), .Q(div_curr_q[32]));
DFFPOSX1 div_d_dff_q_reg[97](.D(div_d_dff_n255), .CLK(rclk), .Q(div_curr_q[33]));
DFFPOSX1 div_d_dff_q_reg[98](.D(div_d_dff_n253), .CLK(rclk), .Q(div_curr_q[34]));
DFFPOSX1 div_d_dff_q_reg[99](.D(div_d_dff_n251), .CLK(rclk), .Q(div_curr_q[35]));
DFFPOSX1 div_d_dff_q_reg[100](.D(div_d_dff_n249), .CLK(rclk), .Q(div_curr_q[36]));
DFFPOSX1 div_d_dff_q_reg[101](.D(div_d_dff_n247), .CLK(rclk), .Q(div_curr_q[37]));
DFFPOSX1 div_d_dff_q_reg[102](.D(div_d_dff_n245), .CLK(rclk), .Q(div_curr_q[38]));
DFFPOSX1 div_d_dff_q_reg[103](.D(div_d_dff_n243), .CLK(rclk), .Q(div_curr_q[39]));
DFFPOSX1 div_d_dff_q_reg[104](.D(div_d_dff_n241), .CLK(rclk), .Q(div_curr_q[40]));
DFFPOSX1 div_d_dff_q_reg[105](.D(div_d_dff_n239), .CLK(rclk), .Q(div_curr_q[41]));
DFFPOSX1 div_d_dff_q_reg[106](.D(div_d_dff_n237), .CLK(rclk), .Q(div_curr_q[42]));
DFFPOSX1 div_d_dff_q_reg[107](.D(div_d_dff_n233), .CLK(rclk), .Q(div_curr_q[43]));
DFFPOSX1 div_d_dff_q_reg[108](.D(div_d_dff_n231), .CLK(rclk), .Q(div_curr_q[44]));
DFFPOSX1 div_d_dff_q_reg[109](.D(div_d_dff_n229), .CLK(rclk), .Q(div_curr_q[45]));
DFFPOSX1 div_d_dff_q_reg[110](.D(div_d_dff_n227), .CLK(rclk), .Q(div_curr_q[46]));
DFFPOSX1 div_d_dff_q_reg[111](.D(div_d_dff_n225), .CLK(rclk), .Q(div_curr_q[47]));
DFFPOSX1 div_d_dff_q_reg[112](.D(div_d_dff_n223), .CLK(rclk), .Q(div_curr_q[48]));
DFFPOSX1 div_d_dff_q_reg[113](.D(div_d_dff_n221), .CLK(rclk), .Q(div_curr_q[49]));
DFFPOSX1 div_d_dff_q_reg[114](.D(div_d_dff_n219), .CLK(rclk), .Q(div_curr_q[50]));
DFFPOSX1 div_d_dff_q_reg[115](.D(div_d_dff_n217), .CLK(rclk), .Q(div_curr_q[51]));
DFFPOSX1 div_d_dff_q_reg[116](.D(div_d_dff_n215), .CLK(rclk), .Q(div_curr_q[52]));
DFFPOSX1 div_d_dff_q_reg[117](.D(div_d_dff_n211), .CLK(rclk), .Q(div_curr_q[53]));
DFFPOSX1 div_d_dff_q_reg[118](.D(div_d_dff_n209), .CLK(rclk), .Q(div_curr_q[54]));
DFFPOSX1 div_d_dff_q_reg[119](.D(div_d_dff_n207), .CLK(rclk), .Q(div_curr_q[55]));
DFFPOSX1 div_d_dff_q_reg[120](.D(div_d_dff_n205), .CLK(rclk), .Q(div_curr_q[56]));
DFFPOSX1 div_d_dff_q_reg[121](.D(div_d_dff_n203), .CLK(rclk), .Q(div_curr_q[57]));
DFFPOSX1 div_d_dff_q_reg[122](.D(div_d_dff_n201), .CLK(rclk), .Q(div_curr_q[58]));
DFFPOSX1 div_d_dff_q_reg[123](.D(div_d_dff_n199), .CLK(rclk), .Q(div_curr_q[59]));
DFFPOSX1 div_d_dff_q_reg[124](.D(div_d_dff_n197), .CLK(rclk), .Q(div_curr_q[60]));
DFFPOSX1 div_d_dff_q_reg[125](.D(div_d_dff_n195), .CLK(rclk), .Q(div_curr_q[61]));
DFFPOSX1 div_d_dff_q_reg[126](.D(div_d_dff_n193), .CLK(rclk), .Q(div_curr_q[62]));
DFFPOSX1 div_d_dff_q_reg[127](.D(div_d_dff_n189), .CLK(rclk), .Q(div_ecl_d_msb));
XOR2X1 exu_div_spr_U191(.A(div_adderin2[0]), .B(exu_n15859), .Y(div_spr_n127));
XOR2X1 exu_div_spr_U190(.A(exu_n15794), .B(div_spr_n127), .Y(div_spr_out[0]));
XOR2X1 exu_div_spr_U189(.A(div_adderin2[10]), .B(exu_n15920), .Y(div_spr_n126));
XOR2X1 exu_div_spr_U188(.A(div_spr_n125), .B(div_spr_n126), .Y(div_spr_out[10]));
XOR2X1 exu_div_spr_U187(.A(div_adderin2[11]), .B(exu_n15919), .Y(div_spr_n124));
XOR2X1 exu_div_spr_U186(.A(div_spr_n123), .B(div_spr_n124), .Y(div_spr_out[11]));
XOR2X1 exu_div_spr_U185(.A(div_adderin2[12]), .B(exu_n15918), .Y(div_spr_n122));
XOR2X1 exu_div_spr_U184(.A(div_spr_n121), .B(div_spr_n122), .Y(div_spr_out[12]));
XOR2X1 exu_div_spr_U183(.A(div_adderin2[13]), .B(exu_n15917), .Y(div_spr_n120));
XOR2X1 exu_div_spr_U182(.A(div_spr_n119), .B(div_spr_n120), .Y(div_spr_out[13]));
XOR2X1 exu_div_spr_U181(.A(div_adderin2[14]), .B(exu_n15916), .Y(div_spr_n118));
XOR2X1 exu_div_spr_U180(.A(div_spr_n117), .B(div_spr_n118), .Y(div_spr_out[14]));
XOR2X1 exu_div_spr_U179(.A(div_adderin2[15]), .B(exu_n15915), .Y(div_spr_n116));
XOR2X1 exu_div_spr_U178(.A(div_spr_n115), .B(div_spr_n116), .Y(div_spr_out[15]));
XOR2X1 exu_div_spr_U177(.A(div_adderin2[16]), .B(exu_n15914), .Y(div_spr_n114));
XOR2X1 exu_div_spr_U176(.A(div_spr_n113), .B(div_spr_n114), .Y(div_spr_out[16]));
XOR2X1 exu_div_spr_U175(.A(div_adderin2[17]), .B(exu_n15913), .Y(div_spr_n112));
XOR2X1 exu_div_spr_U174(.A(div_spr_n111), .B(div_spr_n112), .Y(div_spr_out[17]));
XOR2X1 exu_div_spr_U173(.A(div_adderin2[18]), .B(exu_n15912), .Y(div_spr_n110));
XOR2X1 exu_div_spr_U172(.A(div_spr_n109), .B(div_spr_n110), .Y(div_spr_out[18]));
XOR2X1 exu_div_spr_U171(.A(div_adderin2[19]), .B(exu_n15911), .Y(div_spr_n108));
XOR2X1 exu_div_spr_U170(.A(div_spr_n107), .B(div_spr_n108), .Y(div_spr_out[19]));
XOR2X1 exu_div_spr_U169(.A(div_adderin2[1]), .B(exu_n15910), .Y(div_spr_n106));
XOR2X1 exu_div_spr_U168(.A(div_spr_n105), .B(div_spr_n106), .Y(div_spr_out[1]));
XOR2X1 exu_div_spr_U167(.A(div_adderin2[20]), .B(exu_n15909), .Y(div_spr_n104));
XOR2X1 exu_div_spr_U166(.A(div_spr_n103), .B(div_spr_n104), .Y(div_spr_out[20]));
XOR2X1 exu_div_spr_U165(.A(div_adderin2[21]), .B(exu_n15908), .Y(div_spr_n102));
XOR2X1 exu_div_spr_U164(.A(div_spr_n101), .B(div_spr_n102), .Y(div_spr_out[21]));
XOR2X1 exu_div_spr_U163(.A(div_adderin2[22]), .B(exu_n15907), .Y(div_spr_n100));
XOR2X1 exu_div_spr_U162(.A(div_spr_n99), .B(div_spr_n100), .Y(div_spr_out[22]));
XOR2X1 exu_div_spr_U161(.A(div_adderin2[23]), .B(exu_n15906), .Y(div_spr_n98));
XOR2X1 exu_div_spr_U160(.A(div_spr_n97), .B(div_spr_n98), .Y(div_spr_out[23]));
XOR2X1 exu_div_spr_U159(.A(div_adderin2[24]), .B(exu_n15905), .Y(div_spr_n96));
XOR2X1 exu_div_spr_U158(.A(div_spr_n95), .B(div_spr_n96), .Y(div_spr_out[24]));
XOR2X1 exu_div_spr_U157(.A(div_adderin2[25]), .B(exu_n15904), .Y(div_spr_n94));
XOR2X1 exu_div_spr_U156(.A(div_spr_n93), .B(div_spr_n94), .Y(div_spr_out[25]));
XOR2X1 exu_div_spr_U155(.A(div_adderin2[26]), .B(exu_n15903), .Y(div_spr_n92));
XOR2X1 exu_div_spr_U154(.A(div_spr_n91), .B(div_spr_n92), .Y(div_spr_out[26]));
XOR2X1 exu_div_spr_U153(.A(div_adderin2[27]), .B(exu_n15902), .Y(div_spr_n90));
XOR2X1 exu_div_spr_U152(.A(div_spr_n89), .B(div_spr_n90), .Y(div_spr_out[27]));
XOR2X1 exu_div_spr_U151(.A(div_adderin2[28]), .B(exu_n15901), .Y(div_spr_n88));
XOR2X1 exu_div_spr_U150(.A(div_spr_n87), .B(div_spr_n88), .Y(div_spr_out[28]));
XOR2X1 exu_div_spr_U149(.A(div_adderin2[29]), .B(exu_n15900), .Y(div_spr_n86));
XOR2X1 exu_div_spr_U148(.A(div_spr_n85), .B(div_spr_n86), .Y(div_spr_out[29]));
XOR2X1 exu_div_spr_U147(.A(div_adderin2[2]), .B(exu_n15899), .Y(div_spr_n84));
XOR2X1 exu_div_spr_U146(.A(div_spr_n83), .B(div_spr_n84), .Y(div_spr_out[2]));
XOR2X1 exu_div_spr_U145(.A(div_adderin2[30]), .B(exu_n15898), .Y(div_spr_n82));
XOR2X1 exu_div_spr_U144(.A(div_spr_n81), .B(div_spr_n82), .Y(div_spr_out[30]));
XOR2X1 exu_div_spr_U143(.A(div_adderin2[31]), .B(exu_n15897), .Y(div_spr_n80));
XOR2X1 exu_div_spr_U142(.A(div_spr_n79), .B(div_spr_n80), .Y(div_spr_out[31]));
XOR2X1 exu_div_spr_U141(.A(div_adderin2[32]), .B(exu_n15858), .Y(div_spr_n78));
XOR2X1 exu_div_spr_U140(.A(div_spr_n77), .B(div_spr_n78), .Y(div_spr_out[32]));
XOR2X1 exu_div_spr_U139(.A(div_adderin2[33]), .B(exu_n15896), .Y(div_spr_n76));
XOR2X1 exu_div_spr_U138(.A(div_spr_n75), .B(div_spr_n76), .Y(div_spr_out[33]));
XOR2X1 exu_div_spr_U137(.A(div_adderin2[34]), .B(exu_n15895), .Y(div_spr_n74));
XOR2X1 exu_div_spr_U136(.A(div_spr_n73), .B(div_spr_n74), .Y(div_spr_out[34]));
XOR2X1 exu_div_spr_U135(.A(div_adderin2[35]), .B(exu_n15894), .Y(div_spr_n72));
XOR2X1 exu_div_spr_U134(.A(div_spr_n71), .B(div_spr_n72), .Y(div_spr_out[35]));
XOR2X1 exu_div_spr_U133(.A(div_adderin2[36]), .B(exu_n15893), .Y(div_spr_n70));
XOR2X1 exu_div_spr_U132(.A(div_spr_n69), .B(div_spr_n70), .Y(div_spr_out[36]));
XOR2X1 exu_div_spr_U131(.A(div_adderin2[37]), .B(exu_n15892), .Y(div_spr_n68));
XOR2X1 exu_div_spr_U130(.A(div_spr_n67), .B(div_spr_n68), .Y(div_spr_out[37]));
XOR2X1 exu_div_spr_U129(.A(div_adderin2[38]), .B(exu_n15891), .Y(div_spr_n66));
XOR2X1 exu_div_spr_U128(.A(div_spr_n65), .B(div_spr_n66), .Y(div_spr_out[38]));
XOR2X1 exu_div_spr_U127(.A(div_adderin2[39]), .B(exu_n15890), .Y(div_spr_n64));
XOR2X1 exu_div_spr_U126(.A(div_spr_n63), .B(div_spr_n64), .Y(div_spr_out[39]));
XOR2X1 exu_div_spr_U125(.A(div_adderin2[3]), .B(exu_n15889), .Y(div_spr_n62));
XOR2X1 exu_div_spr_U124(.A(div_spr_n61), .B(div_spr_n62), .Y(div_spr_out[3]));
XOR2X1 exu_div_spr_U123(.A(div_adderin2[40]), .B(exu_n15888), .Y(div_spr_n60));
XOR2X1 exu_div_spr_U122(.A(div_spr_n59), .B(div_spr_n60), .Y(div_spr_out[40]));
XOR2X1 exu_div_spr_U121(.A(div_adderin2[41]), .B(exu_n15887), .Y(div_spr_n58));
XOR2X1 exu_div_spr_U120(.A(div_spr_n57), .B(div_spr_n58), .Y(div_spr_out[41]));
XOR2X1 exu_div_spr_U119(.A(div_adderin2[42]), .B(exu_n15886), .Y(div_spr_n56));
XOR2X1 exu_div_spr_U118(.A(div_spr_n55), .B(div_spr_n56), .Y(div_spr_out[42]));
XOR2X1 exu_div_spr_U117(.A(div_adderin2[43]), .B(exu_n15885), .Y(div_spr_n54));
XOR2X1 exu_div_spr_U116(.A(div_spr_n53), .B(div_spr_n54), .Y(div_spr_out[43]));
XOR2X1 exu_div_spr_U115(.A(div_adderin2[44]), .B(exu_n15884), .Y(div_spr_n52));
XOR2X1 exu_div_spr_U114(.A(div_spr_n51), .B(div_spr_n52), .Y(div_spr_out[44]));
XOR2X1 exu_div_spr_U113(.A(div_adderin2[45]), .B(exu_n15883), .Y(div_spr_n50));
XOR2X1 exu_div_spr_U112(.A(div_spr_n49), .B(div_spr_n50), .Y(div_spr_out[45]));
XOR2X1 exu_div_spr_U111(.A(div_adderin2[46]), .B(exu_n15882), .Y(div_spr_n48));
XOR2X1 exu_div_spr_U110(.A(div_spr_n47), .B(div_spr_n48), .Y(div_spr_out[46]));
XOR2X1 exu_div_spr_U109(.A(div_adderin2[47]), .B(exu_n15881), .Y(div_spr_n46));
XOR2X1 exu_div_spr_U108(.A(div_spr_n45), .B(div_spr_n46), .Y(div_spr_out[47]));
XOR2X1 exu_div_spr_U107(.A(div_adderin2[48]), .B(exu_n15880), .Y(div_spr_n44));
XOR2X1 exu_div_spr_U106(.A(div_spr_n43), .B(div_spr_n44), .Y(div_spr_out[48]));
XOR2X1 exu_div_spr_U105(.A(div_adderin2[49]), .B(exu_n15879), .Y(div_spr_n42));
XOR2X1 exu_div_spr_U104(.A(div_spr_n41), .B(div_spr_n42), .Y(div_spr_out[49]));
XOR2X1 exu_div_spr_U103(.A(div_adderin2[4]), .B(exu_n15878), .Y(div_spr_n40));
XOR2X1 exu_div_spr_U102(.A(div_spr_n39), .B(div_spr_n40), .Y(div_spr_out[4]));
XOR2X1 exu_div_spr_U101(.A(div_adderin2[50]), .B(exu_n15877), .Y(div_spr_n38));
XOR2X1 exu_div_spr_U100(.A(div_spr_n37), .B(div_spr_n38), .Y(div_spr_out[50]));
XOR2X1 exu_div_spr_U99(.A(div_adderin2[51]), .B(exu_n15876), .Y(div_spr_n36));
XOR2X1 exu_div_spr_U98(.A(div_spr_n35), .B(div_spr_n36), .Y(div_spr_out[51]));
XOR2X1 exu_div_spr_U97(.A(div_adderin2[52]), .B(exu_n15875), .Y(div_spr_n34));
XOR2X1 exu_div_spr_U96(.A(div_spr_n33), .B(div_spr_n34), .Y(div_spr_out[52]));
XOR2X1 exu_div_spr_U95(.A(div_adderin2[53]), .B(exu_n15874), .Y(div_spr_n32));
XOR2X1 exu_div_spr_U94(.A(div_spr_n31), .B(div_spr_n32), .Y(div_spr_out[53]));
XOR2X1 exu_div_spr_U93(.A(div_adderin2[54]), .B(exu_n15873), .Y(div_spr_n30));
XOR2X1 exu_div_spr_U92(.A(div_spr_n29), .B(div_spr_n30), .Y(div_spr_out[54]));
XOR2X1 exu_div_spr_U91(.A(div_adderin2[55]), .B(exu_n15872), .Y(div_spr_n28));
XOR2X1 exu_div_spr_U90(.A(div_spr_n27), .B(div_spr_n28), .Y(div_spr_out[55]));
XOR2X1 exu_div_spr_U89(.A(div_adderin2[56]), .B(exu_n15871), .Y(div_spr_n26));
XOR2X1 exu_div_spr_U88(.A(div_spr_n25), .B(div_spr_n26), .Y(div_spr_out[56]));
XOR2X1 exu_div_spr_U87(.A(div_adderin2[57]), .B(exu_n15870), .Y(div_spr_n24));
XOR2X1 exu_div_spr_U86(.A(div_spr_n23), .B(div_spr_n24), .Y(div_spr_out[57]));
XOR2X1 exu_div_spr_U85(.A(div_adderin2[58]), .B(exu_n15869), .Y(div_spr_n22));
XOR2X1 exu_div_spr_U84(.A(div_spr_n21), .B(div_spr_n22), .Y(div_spr_out[58]));
XOR2X1 exu_div_spr_U83(.A(div_adderin2[59]), .B(exu_n15868), .Y(div_spr_n20));
XOR2X1 exu_div_spr_U82(.A(div_spr_n19), .B(div_spr_n20), .Y(div_spr_out[59]));
XOR2X1 exu_div_spr_U81(.A(div_adderin2[5]), .B(exu_n15867), .Y(div_spr_n18));
XOR2X1 exu_div_spr_U80(.A(div_spr_n17), .B(div_spr_n18), .Y(div_spr_out[5]));
XOR2X1 exu_div_spr_U79(.A(div_adderin2[60]), .B(exu_n15866), .Y(div_spr_n16));
XOR2X1 exu_div_spr_U78(.A(div_spr_n15), .B(div_spr_n16), .Y(div_spr_out[60]));
XOR2X1 exu_div_spr_U77(.A(div_adderin2[61]), .B(exu_n15865), .Y(div_spr_n14));
XOR2X1 exu_div_spr_U76(.A(div_spr_n13), .B(div_spr_n14), .Y(div_spr_out[61]));
XOR2X1 exu_div_spr_U75(.A(div_adderin2[62]), .B(exu_n15864), .Y(div_spr_n12));
XOR2X1 exu_div_spr_U74(.A(div_spr_n11), .B(div_spr_n12), .Y(div_spr_out[62]));
XOR2X1 exu_div_spr_U73(.A(div_adderin2[63]), .B(exu_n15823), .Y(div_spr_n10));
XOR2X1 exu_div_spr_U72(.A(div_spr_n9), .B(div_spr_n10), .Y(div_spr_out[63]));
XOR2X1 exu_div_spr_U71(.A(div_adderin2[6]), .B(exu_n15863), .Y(div_spr_n8));
XOR2X1 exu_div_spr_U70(.A(div_spr_n7), .B(div_spr_n8), .Y(div_spr_out[6]));
XOR2X1 exu_div_spr_U69(.A(div_adderin2[7]), .B(exu_n15862), .Y(div_spr_n6));
XOR2X1 exu_div_spr_U68(.A(div_spr_n5), .B(div_spr_n6), .Y(div_spr_out[7]));
XOR2X1 exu_div_spr_U67(.A(div_adderin2[8]), .B(exu_n15861), .Y(div_spr_n4));
XOR2X1 exu_div_spr_U66(.A(div_spr_n3), .B(div_spr_n4), .Y(div_spr_out[8]));
XOR2X1 exu_div_spr_U65(.A(div_adderin2[9]), .B(exu_n15860), .Y(div_spr_n2));
XOR2X1 exu_div_spr_U64(.A(div_spr_n1), .B(div_spr_n2), .Y(div_spr_out[9]));
XNOR2X1 exu_rml_cwp_inc_U8(.A(exu_n16569), .B(rml_rml_ecl_cwp_e[1]), .Y(rml_cwp_inc_n6));
XNOR2X1 exu_rml_cwp_inc_U7(.A(rml_save_e), .B(rml_cwp_inc_n6), .Y(rml_rml_next_cwp_e[1]));
XOR2X1 exu_rml_cwp_inc_U3(.A(exu_n15076), .B(rml_rml_ecl_cwp_e[2]), .Y(rml_cwp_inc_n2));
XOR2X1 exu_rml_cwp_inc_U2(.A(rml_rml_next_cwp_e[1]), .B(rml_cwp_inc_n2), .Y(rml_rml_next_cwp_e[2]));
DFFPOSX1 rml_oddwin_dff_q_reg[0](.D(rml_oddwin_dff_n9), .CLK(rclk), .Q(exu_ifu_oddwin_s[0]));
DFFPOSX1 rml_oddwin_dff_q_reg[1](.D(rml_oddwin_dff_n7), .CLK(rclk), .Q(exu_ifu_oddwin_s[1]));
DFFPOSX1 rml_oddwin_dff_q_reg[2](.D(rml_oddwin_dff_n5), .CLK(rclk), .Q(exu_ifu_oddwin_s[2]));
DFFPOSX1 rml_oddwin_dff_q_reg[3](.D(rml_oddwin_dff_n3), .CLK(rclk), .Q(exu_ifu_oddwin_s[3]));
XNOR2X1 exu_rml_cwp_U155(.A(rml_cwp_trap_old_cwp_m[2]), .B(tlu_exu_cwp_m[2]), .Y(rml_cwp_n101));
XNOR2X1 exu_rml_cwp_U153(.A(rml_cwp_trap_old_cwp_m[0]), .B(tlu_exu_cwp_m[0]), .Y(rml_cwp_n99));
XNOR2X1 exu_rml_cwp_U152(.A(rml_cwp_trap_old_cwp_m[1]), .B(tlu_exu_cwp_m[1]), .Y(rml_cwp_n100));
NAND2X1 exu_rml_cwp_U108(.A(exu_n11617), .B(exu_n10384), .Y(rml_irf_new_lo_cwp_e[0]));
NAND2X1 exu_rml_cwp_U105(.A(exu_n11616), .B(exu_n10383), .Y(rml_irf_new_lo_cwp_e[1]));
NAND2X1 exu_rml_cwp_U102(.A(exu_n11615), .B(exu_n10382), .Y(rml_irf_new_lo_cwp_e[2]));
NAND2X1 exu_rml_cwp_U99(.A(exu_n11614), .B(exu_n10381), .Y(rml_irf_old_lo_cwp_e[0]));
NAND2X1 exu_rml_cwp_U96(.A(exu_n11613), .B(exu_n10380), .Y(rml_irf_old_lo_cwp_e[1]));
NAND2X1 exu_rml_cwp_U93(.A(exu_n11612), .B(exu_n10379), .Y(rml_irf_old_lo_cwp_e[2]));
DFFPOSX1 ecl_writeback_dff_wb_m2w_q_reg[0](.D(ecl_writeback_dff_wb_m2w_n2), .CLK(rclk), .Q(ecl_writeback_wb_w));
DFFPOSX1 ecl_writeback_restore_tid_dff_q_reg[0](.D(exu_n4977), .CLK(rclk), .Q(ecl_writeback_restore_tid[0]));
DFFPOSX1 ecl_writeback_restore_tid_dff_q_reg[1](.D(exu_n4978), .CLK(rclk), .Q(ecl_writeback_restore_tid[1]));
DFFPOSX1 ecl_writeback_restore_rd_dff_q_reg[0](.D(exu_n4972), .CLK(rclk), .Q(ecl_writeback_restore_rd[0]));
DFFPOSX1 ecl_writeback_restore_rd_dff_q_reg[1](.D(exu_n4973), .CLK(rclk), .Q(ecl_writeback_restore_rd[1]));
DFFPOSX1 ecl_writeback_restore_rd_dff_q_reg[2](.D(exu_n4974), .CLK(rclk), .Q(ecl_writeback_restore_rd[2]));
DFFPOSX1 ecl_writeback_restore_rd_dff_q_reg[3](.D(exu_n4975), .CLK(rclk), .Q(ecl_writeback_restore_rd[3]));
DFFPOSX1 ecl_writeback_restore_rd_dff_q_reg[4](.D(exu_n4976), .CLK(rclk), .Q(ecl_writeback_restore_rd[4]));
NAND2X1 exu_ecl_eccctl_ecc_synd7_mux_U2(.A(ecl_eccctl_ecc_synd7_mux_n1), .B(exu_n10346), .Y(exu_ifu_err_synd_m[7]));
XOR2X1 exu_ecl_byplog_rs1_w_comp7_U13(.A(ecl_ecl_irf_rd_w[4]), .B(ecl_ifu_exu_rs1_d[4]), .Y(ecl_byplog_rs1_w_comp7_n9));
XNOR2X1 exu_ecl_byplog_rs1_w_comp7_U12(.A(ecl_ecl_irf_rd_w[3]), .B(ecl_ifu_exu_rs1_d[3]), .Y(ecl_byplog_rs1_w_comp7_n11));
XNOR2X1 exu_ecl_byplog_rs1_w_comp7_U11(.A(ecl_ecl_irf_tid_w[0]), .B(ecl_tid_d[0]), .Y(ecl_byplog_rs1_w_comp7_n12));
XNOR2X1 exu_ecl_byplog_rs1_w_comp7_U8(.A(ecl_ecl_irf_rd_w[0]), .B(ecl_ifu_exu_rs1_d[0]), .Y(ecl_byplog_rs1_w_comp7_n7));
XNOR2X1 exu_ecl_byplog_rs1_w_comp7_U7(.A(ecl_ecl_irf_tid_w[1]), .B(ecl_tid_d[1]), .Y(ecl_byplog_rs1_w_comp7_n8));
XNOR2X1 exu_ecl_byplog_rs1_w_comp7_U5(.A(ecl_ecl_irf_rd_w[2]), .B(ecl_ifu_exu_rs1_d[2]), .Y(ecl_byplog_rs1_w_comp7_n5));
XNOR2X1 exu_ecl_byplog_rs1_w_comp7_U4(.A(ecl_ecl_irf_rd_w[1]), .B(ecl_ifu_exu_rs1_d[1]), .Y(ecl_byplog_rs1_w_comp7_n6));
DFFPOSX1 ecl_divcntl_divstate_dff_q_reg[0](.D(ecl_divcntl_divstate_dff_n13), .CLK(rclk), .Q(ecl_divcntl_div_state_0));
DFFPOSX1 ecl_divcntl_divstate_dff_q_reg[1](.D(ecl_divcntl_divstate_dff_n11), .CLK(rclk), .Q(ecl_divcntl_div_state_1));
DFFPOSX1 ecl_divcntl_divstate_dff_q_reg[2](.D(ecl_divcntl_divstate_dff_n9), .CLK(rclk), .Q(ecl_div_last_cycle));
DFFPOSX1 ecl_divcntl_divstate_dff_q_reg[3](.D(ecl_divcntl_divstate_dff_n7), .CLK(rclk), .Q(ecl_divcntl_div_state[3]));
DFFPOSX1 ecl_divcntl_divstate_dff_q_reg[4](.D(ecl_divcntl_divstate_dff_n5), .CLK(rclk), .Q(ecl_divcntl_div_state[4]));
DFFPOSX1 ecl_divcntl_divstate_dff_q_reg[5](.D(ecl_divcntl_divstate_dff_n3), .CLK(rclk), .Q(ecl_divcntl_div_state[5]));
XOR2X1 exu_ecl_divcntl_cnt6_U36(.A(ecl_divcntl_cntr[1]), .B(ecl_divcntl_cntr[0]), .Y(ecl_divcntl_cnt6_n32));
XOR2X1 exu_ecl_divcntl_cnt6_U16(.A(exu_n15075), .B(ecl_divcntl_cntr[5]), .Y(ecl_divcntl_cnt6_n9));
DFFPOSX1 ecl_divcntl_inputs_neg_dff_q_reg[0](.D(exu_n4971), .CLK(rclk), .Q(ecl_divcntl_inputs_neg_q));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[0](.D(ecl_mdqctl_div_data_dff_n25), .CLK(rclk), .Q(ecl_mdqctl_wb_divthr_g[0]));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[1](.D(ecl_mdqctl_div_data_dff_n23), .CLK(rclk), .Q(ecl_mdqctl_wb_divthr_g[1]));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[2](.D(ecl_mdqctl_div_data_dff_n21), .CLK(rclk), .Q(ecl_mdqctl_wb_divrd_g[0]));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[3](.D(ecl_mdqctl_div_data_dff_n19), .CLK(rclk), .Q(ecl_mdqctl_wb_divrd_g[1]));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[4](.D(ecl_mdqctl_div_data_dff_n17), .CLK(rclk), .Q(ecl_mdqctl_wb_divrd_g[2]));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[5](.D(ecl_mdqctl_div_data_dff_n15), .CLK(rclk), .Q(ecl_mdqctl_wb_divrd_g[3]));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[6](.D(ecl_mdqctl_div_data_dff_n13), .CLK(rclk), .Q(ecl_mdqctl_wb_divrd_g[4]));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[7](.D(ecl_mdqctl_div_data_dff_n11), .CLK(rclk), .Q(ecl_mdqctl_div_data_7));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[8](.D(ecl_mdqctl_div_data_dff_n9), .CLK(rclk), .Q(ecl_ecl_div_signed_div));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[9](.D(ecl_mdqctl_div_data_dff_n7), .CLK(rclk), .Q(ecl_div_div64));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[10](.D(ecl_mdqctl_div_data_dff_n5), .CLK(rclk), .Q(ecl_div_muls));
DFFPOSX1 ecl_mdqctl_div_data_dff_q_reg[11](.D(ecl_mdqctl_div_data_dff_n2), .CLK(rclk), .Q(ecl_mdqctl_div_data[11]));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[0](.D(ecl_mdqctl_mul_data_dff_n15), .CLK(rclk), .Q(ecl_mdqctl_wb_multhr_g[0]));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[1](.D(ecl_mdqctl_mul_data_dff_n13), .CLK(rclk), .Q(ecl_mdqctl_wb_multhr_g[1]));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[2](.D(ecl_mdqctl_mul_data_dff_n11), .CLK(rclk), .Q(ecl_mdqctl_wb_mulrd_g[0]));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[3](.D(ecl_mdqctl_mul_data_dff_n9), .CLK(rclk), .Q(ecl_mdqctl_wb_mulrd_g[1]));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[4](.D(ecl_mdqctl_mul_data_dff_n7), .CLK(rclk), .Q(ecl_mdqctl_wb_mulrd_g[2]));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[5](.D(ecl_mdqctl_mul_data_dff_n5), .CLK(rclk), .Q(ecl_mdqctl_wb_mulrd_g[3]));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[6](.D(ecl_mdqctl_mul_data_dff_n3), .CLK(rclk), .Q(ecl_mdqctl_wb_mulrd_g[4]));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[7](.D(ecl_mdqctl_mul_data_dff_n21), .CLK(rclk), .Q(ecl_mdqctl_wb_mulsetcc_g));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[8](.D(ecl_mdqctl_mul_data_dff_n19), .CLK(rclk), .Q(ecl_mdqctl_mul_data[8]));
DFFPOSX1 ecl_mdqctl_mul_data_dff_q_reg[9](.D(ecl_mdqctl_mul_data_dff_n17), .CLK(rclk), .Q(ecl_mdqctl_mul_data[9]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[0](.D(rml_cwp_slot0_data_dff_n31), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[0]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[1](.D(rml_cwp_slot0_data_dff_n29), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[1]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[2](.D(rml_cwp_slot0_data_dff_n27), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[2]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[3](.D(rml_cwp_slot0_data_dff_n25), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[3]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[4](.D(rml_cwp_slot0_data_dff_n23), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[4]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[5](.D(rml_cwp_slot0_data_dff_n21), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[5]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[6](.D(rml_cwp_slot0_data_dff_n19), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[6]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[7](.D(rml_cwp_slot0_data_dff_n17), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[7]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[8](.D(rml_cwp_slot0_data_dff_n15), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[8]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[9](.D(rml_cwp_slot0_data_dff_n13), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[9]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[10](.D(rml_cwp_slot0_data_dff_n11), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[10]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[11](.D(rml_cwp_slot0_data_dff_n9), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[11]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[12](.D(rml_cwp_slot0_data_dff_n7), .CLK(rclk), .Q(rml_cwp_swap_slot0_data[12]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[13](.D(rml_cwp_slot0_data_dff_n5), .CLK(rclk), .Q(rml_cwp_swap_slot0_state_valid[0]));
DFFPOSX1 rml_cwp_slot0_data_dff_q_reg[14](.D(rml_cwp_slot0_data_dff_n2), .CLK(rclk), .Q(rml_cwp_swap_slot0_state[1]));
XOR2X1 exu_alu_addsub_spr_U191(.A(alu_addsub_rs2_data_0), .B(alu_logic_rs1_data_bf1[0]), .Y(exu_n31615));
XOR2X1 exu_alu_addsub_spr_U190(.A(ecl_alu_cin_e), .B(exu_n31615), .Y(alu_spr_out[0]));
XOR2X1 exu_alu_addsub_spr_U189(.A(alu_addsub_rs2_data_10), .B(alu_logic_rs1_data_bf1[10]), .Y(exu_n31614));
XOR2X1 exu_alu_addsub_spr_U188(.A(exu_n31613), .B(exu_n31614), .Y(alu_spr_out[10]));
XOR2X1 exu_alu_addsub_spr_U187(.A(alu_addsub_rs2_data_11), .B(alu_logic_rs1_data_bf1[11]), .Y(exu_n31612));
XOR2X1 exu_alu_addsub_spr_U186(.A(exu_n31611), .B(exu_n31612), .Y(alu_spr_out[11]));
XOR2X1 exu_alu_addsub_spr_U185(.A(alu_addsub_rs2_data_12), .B(alu_logic_rs1_data_bf1[12]), .Y(exu_n31610));
XOR2X1 exu_alu_addsub_spr_U184(.A(exu_n31609), .B(exu_n31610), .Y(alu_spr_out[12]));
XOR2X1 exu_alu_addsub_spr_U183(.A(alu_addsub_rs2_data_13), .B(alu_logic_rs1_data_bf1[13]), .Y(exu_n31608));
XOR2X1 exu_alu_addsub_spr_U182(.A(exu_n31607), .B(exu_n31608), .Y(alu_spr_out[13]));
XOR2X1 exu_alu_addsub_spr_U181(.A(alu_addsub_rs2_data_14), .B(alu_logic_rs1_data_bf1[14]), .Y(exu_n31606));
XOR2X1 exu_alu_addsub_spr_U180(.A(exu_n31605), .B(exu_n31606), .Y(alu_spr_out[14]));
XOR2X1 exu_alu_addsub_spr_U179(.A(alu_addsub_rs2_data_15), .B(alu_logic_rs1_data_bf1[15]), .Y(exu_n31604));
XOR2X1 exu_alu_addsub_spr_U178(.A(exu_n31603), .B(exu_n31604), .Y(alu_spr_out[15]));
XOR2X1 exu_alu_addsub_spr_U177(.A(alu_addsub_rs2_data_16), .B(alu_logic_rs1_data_bf1[16]), .Y(exu_n31602));
XOR2X1 exu_alu_addsub_spr_U176(.A(exu_n31601), .B(exu_n31602), .Y(alu_spr_out[16]));
XOR2X1 exu_alu_addsub_spr_U175(.A(alu_addsub_rs2_data_17), .B(alu_logic_rs1_data_bf1[17]), .Y(exu_n31600));
XOR2X1 exu_alu_addsub_spr_U174(.A(exu_n31599), .B(exu_n31600), .Y(alu_spr_out[17]));
XOR2X1 exu_alu_addsub_spr_U173(.A(alu_addsub_rs2_data_18), .B(alu_logic_rs1_data_bf1[18]), .Y(exu_n31598));
XOR2X1 exu_alu_addsub_spr_U172(.A(exu_n31597), .B(exu_n31598), .Y(alu_spr_out[18]));
XOR2X1 exu_alu_addsub_spr_U171(.A(alu_addsub_rs2_data_19), .B(alu_logic_rs1_data_bf1[19]), .Y(exu_n31596));
XOR2X1 exu_alu_addsub_spr_U170(.A(exu_n31595), .B(exu_n31596), .Y(alu_spr_out[19]));
XOR2X1 exu_alu_addsub_spr_U169(.A(alu_addsub_rs2_data_1), .B(alu_logic_rs1_data_bf1[1]), .Y(exu_n31594));
XOR2X1 exu_alu_addsub_spr_U168(.A(exu_n31593), .B(exu_n31594), .Y(alu_spr_out[1]));
XOR2X1 exu_alu_addsub_spr_U167(.A(alu_addsub_rs2_data_20), .B(alu_logic_rs1_data_bf1[20]), .Y(exu_n31592));
XOR2X1 exu_alu_addsub_spr_U166(.A(exu_n31591), .B(exu_n31592), .Y(alu_spr_out[20]));
XOR2X1 exu_alu_addsub_spr_U165(.A(alu_addsub_rs2_data_21), .B(alu_logic_rs1_data_bf1[21]), .Y(exu_n31590));
XOR2X1 exu_alu_addsub_spr_U164(.A(exu_n31589), .B(exu_n31590), .Y(alu_spr_out[21]));
XOR2X1 exu_alu_addsub_spr_U163(.A(alu_addsub_rs2_data_22), .B(alu_logic_rs1_data_bf1[22]), .Y(exu_n31588));
XOR2X1 exu_alu_addsub_spr_U162(.A(exu_n31587), .B(exu_n31588), .Y(alu_spr_out[22]));
XOR2X1 exu_alu_addsub_spr_U161(.A(alu_addsub_rs2_data_23), .B(alu_logic_rs1_data_bf1[23]), .Y(exu_n31586));
XOR2X1 exu_alu_addsub_spr_U160(.A(exu_n31585), .B(exu_n31586), .Y(alu_spr_out[23]));
XOR2X1 exu_alu_addsub_spr_U159(.A(alu_addsub_rs2_data_24), .B(alu_logic_rs1_data_bf1[24]), .Y(exu_n31584));
XOR2X1 exu_alu_addsub_spr_U158(.A(exu_n31583), .B(exu_n31584), .Y(alu_spr_out[24]));
XOR2X1 exu_alu_addsub_spr_U157(.A(alu_addsub_rs2_data_25), .B(alu_logic_rs1_data_bf1[25]), .Y(exu_n31582));
XOR2X1 exu_alu_addsub_spr_U156(.A(exu_n31581), .B(exu_n31582), .Y(alu_spr_out[25]));
XOR2X1 exu_alu_addsub_spr_U155(.A(alu_addsub_rs2_data_26), .B(alu_logic_rs1_data_bf1[26]), .Y(exu_n31580));
XOR2X1 exu_alu_addsub_spr_U154(.A(exu_n31579), .B(exu_n31580), .Y(alu_spr_out[26]));
XOR2X1 exu_alu_addsub_spr_U153(.A(alu_addsub_rs2_data_27), .B(alu_logic_rs1_data_bf1[27]), .Y(exu_n31578));
XOR2X1 exu_alu_addsub_spr_U152(.A(exu_n31577), .B(exu_n31578), .Y(alu_spr_out[27]));
XOR2X1 exu_alu_addsub_spr_U151(.A(alu_addsub_rs2_data_28), .B(alu_logic_rs1_data_bf1[28]), .Y(exu_n31576));
XOR2X1 exu_alu_addsub_spr_U150(.A(exu_n31575), .B(exu_n31576), .Y(alu_spr_out[28]));
XOR2X1 exu_alu_addsub_spr_U149(.A(alu_addsub_rs2_data_29), .B(alu_logic_rs1_data_bf1[29]), .Y(exu_n31574));
XOR2X1 exu_alu_addsub_spr_U148(.A(exu_n31573), .B(exu_n31574), .Y(alu_spr_out[29]));
XOR2X1 exu_alu_addsub_spr_U147(.A(alu_addsub_rs2_data_2), .B(alu_logic_rs1_data_bf1[2]), .Y(exu_n31572));
XOR2X1 exu_alu_addsub_spr_U146(.A(exu_n31571), .B(exu_n31572), .Y(alu_spr_out[2]));
XOR2X1 exu_alu_addsub_spr_U145(.A(alu_addsub_rs2_data_30), .B(alu_logic_rs1_data_bf1[30]), .Y(exu_n31570));
XOR2X1 exu_alu_addsub_spr_U144(.A(exu_n31569), .B(exu_n31570), .Y(alu_spr_out[30]));
XOR2X1 exu_alu_addsub_spr_U143(.A(alu_ecl_adderin2_31_e), .B(alu_logic_rs1_data_bf1[31]), .Y(exu_n31568));
XOR2X1 exu_alu_addsub_spr_U142(.A(exu_n31567), .B(exu_n31568), .Y(alu_spr_out[31]));
XOR2X1 exu_alu_addsub_spr_U141(.A(alu_addsub_rs2_data[32]), .B(alu_logic_rs1_data_bf1[32]), .Y(exu_n31566));
XOR2X1 exu_alu_addsub_spr_U140(.A(exu_n31565), .B(exu_n31566), .Y(alu_spr_out[32]));
XOR2X1 exu_alu_addsub_spr_U139(.A(alu_addsub_rs2_data[33]), .B(alu_logic_rs1_data_bf1[33]), .Y(exu_n31564));
XOR2X1 exu_alu_addsub_spr_U138(.A(exu_n31563), .B(exu_n31564), .Y(alu_spr_out[33]));
XOR2X1 exu_alu_addsub_spr_U137(.A(alu_addsub_rs2_data[34]), .B(alu_logic_rs1_data_bf1[34]), .Y(exu_n31562));
XOR2X1 exu_alu_addsub_spr_U136(.A(exu_n31561), .B(exu_n31562), .Y(alu_spr_out[34]));
XOR2X1 exu_alu_addsub_spr_U135(.A(alu_addsub_rs2_data[35]), .B(alu_logic_rs1_data_bf1[35]), .Y(exu_n31560));
XOR2X1 exu_alu_addsub_spr_U134(.A(exu_n31559), .B(exu_n31560), .Y(alu_spr_out[35]));
XOR2X1 exu_alu_addsub_spr_U133(.A(alu_addsub_rs2_data[36]), .B(alu_logic_rs1_data_bf1[36]), .Y(exu_n31558));
XOR2X1 exu_alu_addsub_spr_U132(.A(exu_n31557), .B(exu_n31558), .Y(alu_spr_out[36]));
XOR2X1 exu_alu_addsub_spr_U131(.A(alu_addsub_rs2_data[37]), .B(alu_logic_rs1_data_bf1[37]), .Y(exu_n31556));
XOR2X1 exu_alu_addsub_spr_U130(.A(exu_n31555), .B(exu_n31556), .Y(alu_spr_out[37]));
XOR2X1 exu_alu_addsub_spr_U129(.A(alu_addsub_rs2_data[38]), .B(alu_logic_rs1_data_bf1[38]), .Y(exu_n31554));
XOR2X1 exu_alu_addsub_spr_U128(.A(exu_n31553), .B(exu_n31554), .Y(alu_spr_out[38]));
XOR2X1 exu_alu_addsub_spr_U127(.A(alu_addsub_rs2_data[39]), .B(alu_logic_rs1_data_bf1[39]), .Y(exu_n31552));
XOR2X1 exu_alu_addsub_spr_U126(.A(exu_n31551), .B(exu_n31552), .Y(alu_spr_out[39]));
XOR2X1 exu_alu_addsub_spr_U125(.A(alu_addsub_rs2_data_3), .B(alu_logic_rs1_data_bf1[3]), .Y(exu_n31550));
XOR2X1 exu_alu_addsub_spr_U124(.A(exu_n31549), .B(exu_n31550), .Y(alu_spr_out[3]));
XOR2X1 exu_alu_addsub_spr_U123(.A(alu_addsub_rs2_data[40]), .B(alu_logic_rs1_data_bf1[40]), .Y(exu_n31548));
XOR2X1 exu_alu_addsub_spr_U122(.A(exu_n31547), .B(exu_n31548), .Y(alu_spr_out[40]));
XOR2X1 exu_alu_addsub_spr_U121(.A(alu_addsub_rs2_data[41]), .B(alu_logic_rs1_data_bf1[41]), .Y(exu_n31546));
XOR2X1 exu_alu_addsub_spr_U120(.A(exu_n31545), .B(exu_n31546), .Y(alu_spr_out[41]));
XOR2X1 exu_alu_addsub_spr_U119(.A(alu_addsub_rs2_data[42]), .B(alu_logic_rs1_data_bf1[42]), .Y(exu_n31544));
XOR2X1 exu_alu_addsub_spr_U118(.A(exu_n31543), .B(exu_n31544), .Y(alu_spr_out[42]));
XOR2X1 exu_alu_addsub_spr_U117(.A(alu_addsub_rs2_data[43]), .B(alu_logic_rs1_data_bf1[43]), .Y(exu_n31542));
XOR2X1 exu_alu_addsub_spr_U116(.A(exu_n31541), .B(exu_n31542), .Y(alu_spr_out[43]));
XOR2X1 exu_alu_addsub_spr_U115(.A(alu_addsub_rs2_data[44]), .B(alu_logic_rs1_data_bf1[44]), .Y(exu_n31540));
XOR2X1 exu_alu_addsub_spr_U114(.A(exu_n31539), .B(exu_n31540), .Y(alu_spr_out[44]));
XOR2X1 exu_alu_addsub_spr_U113(.A(alu_addsub_rs2_data[45]), .B(alu_logic_rs1_data_bf1[45]), .Y(exu_n31538));
XOR2X1 exu_alu_addsub_spr_U112(.A(exu_n31537), .B(exu_n31538), .Y(alu_spr_out[45]));
XOR2X1 exu_alu_addsub_spr_U111(.A(alu_addsub_rs2_data[46]), .B(alu_logic_rs1_data_bf1[46]), .Y(exu_n31536));
XOR2X1 exu_alu_addsub_spr_U110(.A(exu_n31535), .B(exu_n31536), .Y(alu_spr_out[46]));
XOR2X1 exu_alu_addsub_spr_U109(.A(alu_addsub_rs2_data[47]), .B(alu_logic_rs1_data_bf1[47]), .Y(exu_n31534));
XOR2X1 exu_alu_addsub_spr_U108(.A(exu_n31533), .B(exu_n31534), .Y(alu_spr_out[47]));
XOR2X1 exu_alu_addsub_spr_U107(.A(alu_addsub_rs2_data[48]), .B(alu_logic_rs1_data_bf1[48]), .Y(exu_n31532));
XOR2X1 exu_alu_addsub_spr_U106(.A(exu_n31531), .B(exu_n31532), .Y(alu_spr_out[48]));
XOR2X1 exu_alu_addsub_spr_U105(.A(alu_addsub_rs2_data[49]), .B(alu_logic_rs1_data_bf1[49]), .Y(exu_n31530));
XOR2X1 exu_alu_addsub_spr_U104(.A(exu_n31529), .B(exu_n31530), .Y(alu_spr_out[49]));
XOR2X1 exu_alu_addsub_spr_U103(.A(alu_addsub_rs2_data_4), .B(alu_logic_rs1_data_bf1[4]), .Y(exu_n31528));
XOR2X1 exu_alu_addsub_spr_U102(.A(exu_n31527), .B(exu_n31528), .Y(alu_spr_out[4]));
XOR2X1 exu_alu_addsub_spr_U101(.A(alu_addsub_rs2_data[50]), .B(alu_logic_rs1_data_bf1[50]), .Y(exu_n31526));
XOR2X1 exu_alu_addsub_spr_U100(.A(exu_n31525), .B(exu_n31526), .Y(alu_spr_out[50]));
XOR2X1 exu_alu_addsub_spr_U99(.A(alu_addsub_rs2_data[51]), .B(alu_logic_rs1_data_bf1[51]), .Y(exu_n31524));
XOR2X1 exu_alu_addsub_spr_U98(.A(exu_n31523), .B(exu_n31524), .Y(alu_spr_out[51]));
XOR2X1 exu_alu_addsub_spr_U97(.A(alu_addsub_rs2_data[52]), .B(alu_logic_rs1_data_bf1[52]), .Y(exu_n31522));
XOR2X1 exu_alu_addsub_spr_U96(.A(exu_n31521), .B(exu_n31522), .Y(alu_spr_out[52]));
XOR2X1 exu_alu_addsub_spr_U95(.A(alu_addsub_rs2_data[53]), .B(alu_logic_rs1_data_bf1[53]), .Y(exu_n31520));
XOR2X1 exu_alu_addsub_spr_U94(.A(exu_n31519), .B(exu_n31520), .Y(alu_spr_out[53]));
XOR2X1 exu_alu_addsub_spr_U93(.A(alu_addsub_rs2_data[54]), .B(alu_logic_rs1_data_bf1[54]), .Y(exu_n31518));
XOR2X1 exu_alu_addsub_spr_U92(.A(exu_n31517), .B(exu_n31518), .Y(alu_spr_out[54]));
XOR2X1 exu_alu_addsub_spr_U91(.A(alu_addsub_rs2_data[55]), .B(alu_logic_rs1_data_bf1[55]), .Y(exu_n31516));
XOR2X1 exu_alu_addsub_spr_U90(.A(exu_n31515), .B(exu_n31516), .Y(alu_spr_out[55]));
XOR2X1 exu_alu_addsub_spr_U89(.A(alu_addsub_rs2_data[56]), .B(alu_logic_rs1_data_bf1[56]), .Y(exu_n31514));
XOR2X1 exu_alu_addsub_spr_U88(.A(exu_n31513), .B(exu_n31514), .Y(alu_spr_out[56]));
XOR2X1 exu_alu_addsub_spr_U87(.A(alu_addsub_rs2_data[57]), .B(alu_logic_rs1_data_bf1[57]), .Y(exu_n31512));
XOR2X1 exu_alu_addsub_spr_U86(.A(exu_n31511), .B(exu_n31512), .Y(alu_spr_out[57]));
XOR2X1 exu_alu_addsub_spr_U85(.A(alu_addsub_rs2_data[58]), .B(alu_logic_rs1_data_bf1[58]), .Y(exu_n31510));
XOR2X1 exu_alu_addsub_spr_U84(.A(exu_n31509), .B(exu_n31510), .Y(alu_spr_out[58]));
XOR2X1 exu_alu_addsub_spr_U83(.A(alu_addsub_rs2_data[59]), .B(alu_logic_rs1_data_bf1[59]), .Y(exu_n31508));
XOR2X1 exu_alu_addsub_spr_U82(.A(exu_n31507), .B(exu_n31508), .Y(alu_spr_out[59]));
XOR2X1 exu_alu_addsub_spr_U81(.A(alu_addsub_rs2_data_5), .B(alu_logic_rs1_data_bf1[5]), .Y(exu_n31506));
XOR2X1 exu_alu_addsub_spr_U80(.A(exu_n31505), .B(exu_n31506), .Y(alu_spr_out[5]));
XOR2X1 exu_alu_addsub_spr_U79(.A(alu_addsub_rs2_data[60]), .B(alu_logic_rs1_data_bf1[60]), .Y(exu_n31504));
XOR2X1 exu_alu_addsub_spr_U78(.A(exu_n31503), .B(exu_n31504), .Y(alu_spr_out[60]));
XOR2X1 exu_alu_addsub_spr_U77(.A(alu_addsub_rs2_data[61]), .B(alu_logic_rs1_data_bf1[61]), .Y(exu_n31502));
XOR2X1 exu_alu_addsub_spr_U76(.A(exu_n31501), .B(exu_n31502), .Y(alu_spr_out[61]));
XOR2X1 exu_alu_addsub_spr_U75(.A(alu_addsub_rs2_data[62]), .B(alu_logic_rs1_data_bf1[62]), .Y(exu_n31500));
XOR2X1 exu_alu_addsub_spr_U74(.A(exu_n31499), .B(exu_n31500), .Y(alu_spr_out[62]));
XOR2X1 exu_alu_addsub_spr_U73(.A(alu_ecl_adderin2_63_e), .B(alu_logic_rs1_data_bf1[63]), .Y(exu_n31498));
XOR2X1 exu_alu_addsub_spr_U72(.A(exu_n31497), .B(exu_n31498), .Y(alu_spr_out[63]));
XOR2X1 exu_alu_addsub_spr_U71(.A(alu_addsub_rs2_data_6), .B(alu_logic_rs1_data_bf1[6]), .Y(exu_n31496));
XOR2X1 exu_alu_addsub_spr_U70(.A(exu_n31495), .B(exu_n31496), .Y(alu_spr_out[6]));
XOR2X1 exu_alu_addsub_spr_U69(.A(alu_addsub_rs2_data_7), .B(alu_logic_rs1_data_bf1[7]), .Y(exu_n31494));
XOR2X1 exu_alu_addsub_spr_U68(.A(exu_n31493), .B(exu_n31494), .Y(alu_spr_out[7]));
XOR2X1 exu_alu_addsub_spr_U67(.A(alu_addsub_rs2_data_8), .B(alu_logic_rs1_data_bf1[8]), .Y(exu_n31492));
XOR2X1 exu_alu_addsub_spr_U66(.A(exu_n31491), .B(exu_n31492), .Y(alu_spr_out[8]));
XOR2X1 exu_alu_addsub_spr_U65(.A(alu_addsub_rs2_data_9), .B(alu_logic_rs1_data_bf1[9]), .Y(exu_n31490));
XOR2X1 exu_alu_addsub_spr_U64(.A(exu_n31489), .B(exu_n31490), .Y(alu_spr_out[9]));
NAND2X1 exu_alu_lsu_va_mux_U191(.A(exu_n11233), .B(exu_n10239), .Y(exu_lsu_ldst_va_e[0]));
NAND2X1 exu_alu_lsu_va_mux_U188(.A(exu_n11232), .B(exu_n10238), .Y(exu_lsu_ldst_va_e[10]));
NAND2X1 exu_alu_lsu_va_mux_U185(.A(exu_n11231), .B(exu_n10237), .Y(exu_lsu_ldst_va_e[11]));
NAND2X1 exu_alu_lsu_va_mux_U182(.A(exu_n11230), .B(exu_n10236), .Y(exu_lsu_ldst_va_e[12]));
NAND2X1 exu_alu_lsu_va_mux_U179(.A(exu_n11229), .B(exu_n10235), .Y(exu_lsu_ldst_va_e[13]));
NAND2X1 exu_alu_lsu_va_mux_U176(.A(exu_n11228), .B(exu_n10234), .Y(exu_lsu_ldst_va_e[14]));
NAND2X1 exu_alu_lsu_va_mux_U173(.A(exu_n11227), .B(exu_n10233), .Y(exu_lsu_ldst_va_e[15]));
NAND2X1 exu_alu_lsu_va_mux_U170(.A(exu_n11226), .B(exu_n10232), .Y(exu_lsu_ldst_va_e[16]));
NAND2X1 exu_alu_lsu_va_mux_U167(.A(exu_n11225), .B(exu_n10231), .Y(exu_lsu_ldst_va_e[17]));
NAND2X1 exu_alu_lsu_va_mux_U164(.A(exu_n11224), .B(exu_n10230), .Y(exu_lsu_ldst_va_e[18]));
NAND2X1 exu_alu_lsu_va_mux_U161(.A(exu_n11223), .B(exu_n10229), .Y(exu_lsu_ldst_va_e[19]));
NAND2X1 exu_alu_lsu_va_mux_U158(.A(exu_n11222), .B(exu_n10228), .Y(exu_lsu_ldst_va_e[1]));
NAND2X1 exu_alu_lsu_va_mux_U155(.A(exu_n11221), .B(exu_n10227), .Y(exu_lsu_ldst_va_e[20]));
NAND2X1 exu_alu_lsu_va_mux_U152(.A(exu_n11220), .B(exu_n10226), .Y(exu_lsu_ldst_va_e[21]));
NAND2X1 exu_alu_lsu_va_mux_U149(.A(exu_n11219), .B(exu_n10225), .Y(exu_lsu_ldst_va_e[22]));
NAND2X1 exu_alu_lsu_va_mux_U146(.A(exu_n11218), .B(exu_n10224), .Y(exu_lsu_ldst_va_e[23]));
NAND2X1 exu_alu_lsu_va_mux_U143(.A(exu_n11217), .B(exu_n10223), .Y(exu_lsu_ldst_va_e[24]));
NAND2X1 exu_alu_lsu_va_mux_U140(.A(exu_n11216), .B(exu_n10222), .Y(exu_lsu_ldst_va_e[25]));
NAND2X1 exu_alu_lsu_va_mux_U137(.A(exu_n11215), .B(exu_n10221), .Y(exu_lsu_ldst_va_e[26]));
NAND2X1 exu_alu_lsu_va_mux_U134(.A(exu_n11214), .B(exu_n10220), .Y(exu_lsu_ldst_va_e[27]));
NAND2X1 exu_alu_lsu_va_mux_U131(.A(exu_n11213), .B(exu_n10219), .Y(exu_lsu_ldst_va_e[28]));
NAND2X1 exu_alu_lsu_va_mux_U128(.A(exu_n11212), .B(exu_n10218), .Y(exu_lsu_ldst_va_e[29]));
NAND2X1 exu_alu_lsu_va_mux_U125(.A(exu_n11211), .B(exu_n10217), .Y(exu_lsu_ldst_va_e[2]));
NAND2X1 exu_alu_lsu_va_mux_U122(.A(exu_n11210), .B(exu_n10216), .Y(exu_lsu_ldst_va_e[30]));
NAND2X1 exu_alu_lsu_va_mux_U119(.A(exu_n11209), .B(exu_n10215), .Y(exu_lsu_ldst_va_e[31]));
NAND2X1 exu_alu_lsu_va_mux_U116(.A(exu_n11208), .B(exu_n10214), .Y(exu_lsu_ldst_va_e[32]));
NAND2X1 exu_alu_lsu_va_mux_U113(.A(exu_n11207), .B(exu_n10213), .Y(exu_lsu_ldst_va_e[33]));
NAND2X1 exu_alu_lsu_va_mux_U110(.A(exu_n11206), .B(exu_n10212), .Y(exu_lsu_ldst_va_e[34]));
NAND2X1 exu_alu_lsu_va_mux_U107(.A(exu_n11205), .B(exu_n10211), .Y(exu_lsu_ldst_va_e[35]));
NAND2X1 exu_alu_lsu_va_mux_U104(.A(exu_n11204), .B(exu_n10210), .Y(exu_lsu_ldst_va_e[36]));
NAND2X1 exu_alu_lsu_va_mux_U101(.A(exu_n11203), .B(exu_n10209), .Y(exu_lsu_ldst_va_e[37]));
NAND2X1 exu_alu_lsu_va_mux_U98(.A(exu_n11202), .B(exu_n10208), .Y(exu_lsu_ldst_va_e[38]));
NAND2X1 exu_alu_lsu_va_mux_U95(.A(exu_n11201), .B(exu_n10207), .Y(exu_lsu_ldst_va_e[39]));
NAND2X1 exu_alu_lsu_va_mux_U92(.A(exu_n11200), .B(exu_n10206), .Y(exu_lsu_ldst_va_e[3]));
NAND2X1 exu_alu_lsu_va_mux_U89(.A(exu_n11199), .B(exu_n10205), .Y(exu_lsu_ldst_va_e[40]));
NAND2X1 exu_alu_lsu_va_mux_U86(.A(exu_n11198), .B(exu_n10204), .Y(exu_lsu_ldst_va_e[41]));
NAND2X1 exu_alu_lsu_va_mux_U83(.A(exu_n11197), .B(exu_n10203), .Y(exu_lsu_ldst_va_e[42]));
NAND2X1 exu_alu_lsu_va_mux_U80(.A(exu_n11196), .B(exu_n10202), .Y(exu_lsu_ldst_va_e[43]));
NAND2X1 exu_alu_lsu_va_mux_U77(.A(exu_n11195), .B(exu_n10201), .Y(exu_lsu_ldst_va_e[44]));
NAND2X1 exu_alu_lsu_va_mux_U74(.A(exu_n11194), .B(exu_n10200), .Y(exu_lsu_ldst_va_e[45]));
NAND2X1 exu_alu_lsu_va_mux_U71(.A(exu_n11193), .B(exu_n10199), .Y(exu_lsu_ldst_va_e[46]));
NAND2X1 exu_alu_lsu_va_mux_U59(.A(exu_n11192), .B(exu_n10198), .Y(exu_lsu_ldst_va_e[4]));
NAND2X1 exu_alu_lsu_va_mux_U26(.A(exu_n11191), .B(exu_n10197), .Y(exu_lsu_ldst_va_e[5]));
NAND2X1 exu_alu_lsu_va_mux_U11(.A(exu_n11190), .B(exu_n10196), .Y(exu_lsu_ldst_va_e[6]));
NAND2X1 exu_alu_lsu_va_mux_U8(.A(exu_n11189), .B(exu_n10195), .Y(exu_lsu_ldst_va_e[7]));
NAND2X1 exu_alu_lsu_va_mux_U5(.A(exu_n11188), .B(exu_n10194), .Y(exu_lsu_ldst_va_e[8]));
NAND2X1 exu_alu_lsu_va_mux_U2(.A(exu_n11187), .B(exu_n10193), .Y(exu_lsu_ldst_va_e[9]));
NAND2X1 exu_bypass_rs2_data_out_mux_U191(.A(exu_n11186), .B(exu_n10192), .Y(exu_lsu_rs2_data_e[0]));
NAND2X1 exu_bypass_rs2_data_out_mux_U188(.A(exu_n11185), .B(exu_n10191), .Y(exu_lsu_rs2_data_e[10]));
NAND2X1 exu_bypass_rs2_data_out_mux_U185(.A(exu_n11184), .B(exu_n10190), .Y(exu_lsu_rs2_data_e[11]));
NAND2X1 exu_bypass_rs2_data_out_mux_U182(.A(exu_n11183), .B(exu_n10189), .Y(exu_lsu_rs2_data_e[12]));
NAND2X1 exu_bypass_rs2_data_out_mux_U179(.A(exu_n11182), .B(exu_n10188), .Y(exu_lsu_rs2_data_e[13]));
NAND2X1 exu_bypass_rs2_data_out_mux_U176(.A(exu_n11181), .B(exu_n10187), .Y(exu_lsu_rs2_data_e[14]));
NAND2X1 exu_bypass_rs2_data_out_mux_U173(.A(exu_n11180), .B(exu_n10186), .Y(exu_lsu_rs2_data_e[15]));
NAND2X1 exu_bypass_rs2_data_out_mux_U170(.A(exu_n11179), .B(exu_n10185), .Y(exu_lsu_rs2_data_e[16]));
NAND2X1 exu_bypass_rs2_data_out_mux_U167(.A(exu_n11178), .B(exu_n10184), .Y(exu_lsu_rs2_data_e[17]));
NAND2X1 exu_bypass_rs2_data_out_mux_U164(.A(exu_n11177), .B(exu_n10183), .Y(exu_lsu_rs2_data_e[18]));
NAND2X1 exu_bypass_rs2_data_out_mux_U161(.A(exu_n11176), .B(exu_n10182), .Y(exu_lsu_rs2_data_e[19]));
NAND2X1 exu_bypass_rs2_data_out_mux_U158(.A(exu_n11175), .B(exu_n10181), .Y(exu_lsu_rs2_data_e[1]));
NAND2X1 exu_bypass_rs2_data_out_mux_U155(.A(exu_n11174), .B(exu_n10180), .Y(exu_lsu_rs2_data_e[20]));
NAND2X1 exu_bypass_rs2_data_out_mux_U152(.A(exu_n11173), .B(exu_n10179), .Y(exu_lsu_rs2_data_e[21]));
NAND2X1 exu_bypass_rs2_data_out_mux_U149(.A(exu_n11172), .B(exu_n10178), .Y(exu_lsu_rs2_data_e[22]));
NAND2X1 exu_bypass_rs2_data_out_mux_U146(.A(exu_n11171), .B(exu_n10177), .Y(exu_lsu_rs2_data_e[23]));
NAND2X1 exu_bypass_rs2_data_out_mux_U143(.A(exu_n11170), .B(exu_n10176), .Y(exu_lsu_rs2_data_e[24]));
NAND2X1 exu_bypass_rs2_data_out_mux_U140(.A(exu_n11169), .B(exu_n10175), .Y(exu_lsu_rs2_data_e[25]));
NAND2X1 exu_bypass_rs2_data_out_mux_U137(.A(exu_n11168), .B(exu_n10174), .Y(exu_lsu_rs2_data_e[26]));
NAND2X1 exu_bypass_rs2_data_out_mux_U134(.A(exu_n11167), .B(exu_n10173), .Y(exu_lsu_rs2_data_e[27]));
NAND2X1 exu_bypass_rs2_data_out_mux_U131(.A(exu_n11166), .B(exu_n10172), .Y(exu_lsu_rs2_data_e[28]));
NAND2X1 exu_bypass_rs2_data_out_mux_U128(.A(exu_n11165), .B(exu_n10171), .Y(exu_lsu_rs2_data_e[29]));
NAND2X1 exu_bypass_rs2_data_out_mux_U125(.A(exu_n11164), .B(exu_n10170), .Y(exu_lsu_rs2_data_e[2]));
NAND2X1 exu_bypass_rs2_data_out_mux_U122(.A(exu_n11163), .B(exu_n10169), .Y(exu_lsu_rs2_data_e[30]));
NAND2X1 exu_bypass_rs2_data_out_mux_U119(.A(exu_n11162), .B(exu_n10168), .Y(exu_lsu_rs2_data_e[31]));
NAND2X1 exu_bypass_rs2_data_out_mux_U116(.A(exu_n11161), .B(exu_n10167), .Y(exu_lsu_rs2_data_e[32]));
NAND2X1 exu_bypass_rs2_data_out_mux_U113(.A(exu_n11160), .B(exu_n10166), .Y(exu_lsu_rs2_data_e[33]));
NAND2X1 exu_bypass_rs2_data_out_mux_U110(.A(exu_n11159), .B(exu_n10165), .Y(exu_lsu_rs2_data_e[34]));
NAND2X1 exu_bypass_rs2_data_out_mux_U107(.A(exu_n11158), .B(exu_n10164), .Y(exu_lsu_rs2_data_e[35]));
NAND2X1 exu_bypass_rs2_data_out_mux_U104(.A(exu_n11157), .B(exu_n10163), .Y(exu_lsu_rs2_data_e[36]));
NAND2X1 exu_bypass_rs2_data_out_mux_U101(.A(exu_n11156), .B(exu_n10162), .Y(exu_lsu_rs2_data_e[37]));
NAND2X1 exu_bypass_rs2_data_out_mux_U98(.A(exu_n11155), .B(exu_n10161), .Y(exu_lsu_rs2_data_e[38]));
NAND2X1 exu_bypass_rs2_data_out_mux_U95(.A(exu_n11154), .B(exu_n10160), .Y(exu_lsu_rs2_data_e[39]));
NAND2X1 exu_bypass_rs2_data_out_mux_U92(.A(exu_n11153), .B(exu_n10159), .Y(exu_lsu_rs2_data_e[3]));
NAND2X1 exu_bypass_rs2_data_out_mux_U89(.A(exu_n11152), .B(exu_n10158), .Y(exu_lsu_rs2_data_e[40]));
NAND2X1 exu_bypass_rs2_data_out_mux_U86(.A(exu_n11151), .B(exu_n10157), .Y(exu_lsu_rs2_data_e[41]));
NAND2X1 exu_bypass_rs2_data_out_mux_U83(.A(exu_n11150), .B(exu_n10156), .Y(exu_lsu_rs2_data_e[42]));
NAND2X1 exu_bypass_rs2_data_out_mux_U80(.A(exu_n11149), .B(exu_n10155), .Y(exu_lsu_rs2_data_e[43]));
NAND2X1 exu_bypass_rs2_data_out_mux_U77(.A(exu_n11148), .B(exu_n10154), .Y(exu_lsu_rs2_data_e[44]));
NAND2X1 exu_bypass_rs2_data_out_mux_U74(.A(exu_n11147), .B(exu_n10153), .Y(exu_lsu_rs2_data_e[45]));
NAND2X1 exu_bypass_rs2_data_out_mux_U71(.A(exu_n11146), .B(exu_n10152), .Y(exu_lsu_rs2_data_e[46]));
NAND2X1 exu_bypass_rs2_data_out_mux_U68(.A(exu_n11145), .B(exu_n10151), .Y(exu_lsu_rs2_data_e[47]));
NAND2X1 exu_bypass_rs2_data_out_mux_U65(.A(exu_n11144), .B(exu_n10150), .Y(exu_lsu_rs2_data_e[48]));
NAND2X1 exu_bypass_rs2_data_out_mux_U62(.A(exu_n11143), .B(exu_n10149), .Y(exu_lsu_rs2_data_e[49]));
NAND2X1 exu_bypass_rs2_data_out_mux_U59(.A(exu_n11142), .B(exu_n10148), .Y(exu_lsu_rs2_data_e[4]));
NAND2X1 exu_bypass_rs2_data_out_mux_U56(.A(exu_n11141), .B(exu_n10147), .Y(exu_lsu_rs2_data_e[50]));
NAND2X1 exu_bypass_rs2_data_out_mux_U53(.A(exu_n11140), .B(exu_n10146), .Y(exu_lsu_rs2_data_e[51]));
NAND2X1 exu_bypass_rs2_data_out_mux_U50(.A(exu_n11139), .B(exu_n10145), .Y(exu_lsu_rs2_data_e[52]));
NAND2X1 exu_bypass_rs2_data_out_mux_U47(.A(exu_n11138), .B(exu_n10144), .Y(exu_lsu_rs2_data_e[53]));
NAND2X1 exu_bypass_rs2_data_out_mux_U44(.A(exu_n11137), .B(exu_n10143), .Y(exu_lsu_rs2_data_e[54]));
NAND2X1 exu_bypass_rs2_data_out_mux_U41(.A(exu_n11136), .B(exu_n10142), .Y(exu_lsu_rs2_data_e[55]));
NAND2X1 exu_bypass_rs2_data_out_mux_U38(.A(exu_n11135), .B(exu_n10141), .Y(exu_lsu_rs2_data_e[56]));
NAND2X1 exu_bypass_rs2_data_out_mux_U35(.A(exu_n11134), .B(exu_n10140), .Y(exu_lsu_rs2_data_e[57]));
NAND2X1 exu_bypass_rs2_data_out_mux_U32(.A(exu_n11133), .B(exu_n10139), .Y(exu_lsu_rs2_data_e[58]));
NAND2X1 exu_bypass_rs2_data_out_mux_U29(.A(exu_n11132), .B(exu_n10138), .Y(exu_lsu_rs2_data_e[59]));
NAND2X1 exu_bypass_rs2_data_out_mux_U26(.A(exu_n11131), .B(exu_n10137), .Y(exu_lsu_rs2_data_e[5]));
NAND2X1 exu_bypass_rs2_data_out_mux_U23(.A(exu_n11130), .B(exu_n10136), .Y(exu_lsu_rs2_data_e[60]));
NAND2X1 exu_bypass_rs2_data_out_mux_U20(.A(exu_n11129), .B(exu_n10135), .Y(exu_lsu_rs2_data_e[61]));
NAND2X1 exu_bypass_rs2_data_out_mux_U17(.A(exu_n11128), .B(exu_n10134), .Y(exu_lsu_rs2_data_e[62]));
NAND2X1 exu_bypass_rs2_data_out_mux_U14(.A(exu_n11127), .B(exu_n10133), .Y(exu_lsu_rs2_data_e[63]));
NAND2X1 exu_bypass_rs2_data_out_mux_U11(.A(exu_n11126), .B(exu_n10132), .Y(exu_lsu_rs2_data_e[6]));
NAND2X1 exu_bypass_rs2_data_out_mux_U8(.A(exu_n11125), .B(exu_n10131), .Y(exu_lsu_rs2_data_e[7]));
NAND2X1 exu_bypass_rs2_data_out_mux_U5(.A(exu_n11124), .B(exu_n10130), .Y(exu_lsu_rs2_data_e[8]));
NAND2X1 exu_bypass_rs2_data_out_mux_U2(.A(exu_n11123), .B(exu_n10129), .Y(exu_lsu_rs2_data_e[9]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[0](.D(exu_n16357), .CLK(rclk), .Q(alu_addsub_subtract_e[0]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[1](.D(exu_n16350), .CLK(rclk), .Q(alu_addsub_subtract_e[1]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[2](.D(exu_n16341), .CLK(rclk), .Q(alu_addsub_subtract_e[2]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[3](.D(exu_n16332), .CLK(rclk), .Q(alu_addsub_subtract_e[3]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[4](.D(exu_n16324), .CLK(rclk), .Q(alu_addsub_subtract_e[4]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[5](.D(exu_n16323), .CLK(rclk), .Q(alu_addsub_subtract_e[5]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[6](.D(exu_n16322), .CLK(rclk), .Q(alu_addsub_subtract_e[6]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[7](.D(exu_n19280), .CLK(rclk), .Q(alu_addsub_subtract_e[7]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[8](.D(exu_n16340), .CLK(rclk), .Q(alu_addsub_subtract_e[8]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[9](.D(exu_n16369), .CLK(rclk), .Q(alu_addsub_subtract_e[9]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[10](.D(exu_n16368), .CLK(rclk), .Q(alu_addsub_subtract_e[10]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[11](.D(exu_n19338), .CLK(rclk), .Q(alu_addsub_subtract_e[11]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[12](.D(exu_n16367), .CLK(rclk), .Q(alu_addsub_subtract_e[12]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[13](.D(exu_n16339), .CLK(rclk), .Q(alu_addsub_subtract_e[13]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[14](.D(exu_n16366), .CLK(rclk), .Q(alu_addsub_subtract_e[14]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[15](.D(exu_n16365), .CLK(rclk), .Q(alu_addsub_subtract_e[15]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[16](.D(exu_n16364), .CLK(rclk), .Q(alu_addsub_subtract_e[16]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[17](.D(exu_n16363), .CLK(rclk), .Q(alu_addsub_subtract_e[17]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[18](.D(exu_n16362), .CLK(rclk), .Q(alu_addsub_subtract_e[18]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[19](.D(exu_n16361), .CLK(rclk), .Q(alu_addsub_subtract_e[19]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[20](.D(exu_n16328), .CLK(rclk), .Q(alu_addsub_subtract_e[20]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[21](.D(exu_n16322), .CLK(rclk), .Q(alu_addsub_subtract_e[21]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[22](.D(exu_n16360), .CLK(rclk), .Q(alu_addsub_subtract_e[22]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[23](.D(exu_n16325), .CLK(rclk), .Q(alu_addsub_subtract_e[23]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[24](.D(exu_n16332), .CLK(rclk), .Q(alu_addsub_subtract_e[24]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[25](.D(exu_n16359), .CLK(rclk), .Q(alu_addsub_subtract_e[25]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[26](.D(exu_n16358), .CLK(rclk), .Q(alu_addsub_subtract_e[26]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[27](.D(exu_n16356), .CLK(rclk), .Q(alu_addsub_subtract_e[27]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[28](.D(exu_n16355), .CLK(rclk), .Q(alu_addsub_subtract_e[28]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[29](.D(exu_n16354), .CLK(rclk), .Q(alu_addsub_subtract_e[29]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[30](.D(exu_n16353), .CLK(rclk), .Q(alu_addsub_subtract_e[30]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[31](.D(exu_n16352), .CLK(rclk), .Q(alu_addsub_subtract_e[31]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[32](.D(exu_n16337), .CLK(rclk), .Q(alu_addsub_subtract_e[32]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[33](.D(exu_n16333), .CLK(rclk), .Q(alu_addsub_subtract_e[33]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[34](.D(exu_n16351), .CLK(rclk), .Q(alu_addsub_subtract_e[34]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[35](.D(exu_n16336), .CLK(rclk), .Q(alu_addsub_subtract_e[35]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[36](.D(exu_n16334), .CLK(rclk), .Q(alu_addsub_subtract_e[36]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[37](.D(exu_n16349), .CLK(rclk), .Q(alu_addsub_subtract_e[37]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[38](.D(exu_n16348), .CLK(rclk), .Q(alu_addsub_subtract_e[38]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[39](.D(exu_n16347), .CLK(rclk), .Q(alu_addsub_subtract_e[39]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[40](.D(exu_n16346), .CLK(rclk), .Q(alu_addsub_subtract_e[40]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[41](.D(exu_n16345), .CLK(rclk), .Q(alu_addsub_subtract_e[41]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[42](.D(exu_n16344), .CLK(rclk), .Q(alu_addsub_subtract_e[42]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[43](.D(exu_n16343), .CLK(rclk), .Q(alu_addsub_subtract_e[43]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[44](.D(exu_n16330), .CLK(rclk), .Q(alu_addsub_subtract_e[44]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[45](.D(exu_n16326), .CLK(rclk), .Q(alu_addsub_subtract_e[45]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[46](.D(exu_n16342), .CLK(rclk), .Q(alu_addsub_subtract_e[46]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[47](.D(exu_n16340), .CLK(rclk), .Q(alu_addsub_subtract_e[47]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[48](.D(exu_n16327), .CLK(rclk), .Q(alu_addsub_subtract_e[48]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[49](.D(exu_n16339), .CLK(rclk), .Q(alu_addsub_subtract_e[49]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[50](.D(exu_n16338), .CLK(rclk), .Q(alu_addsub_subtract_e[50]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[51](.D(exu_n16337), .CLK(rclk), .Q(alu_addsub_subtract_e[51]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[52](.D(exu_n16336), .CLK(rclk), .Q(alu_addsub_subtract_e[52]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[53](.D(exu_n16335), .CLK(rclk), .Q(alu_addsub_subtract_e[53]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[54](.D(exu_n16334), .CLK(rclk), .Q(alu_addsub_subtract_e[54]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[55](.D(exu_n16333), .CLK(rclk), .Q(alu_addsub_subtract_e[55]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[56](.D(exu_n16335), .CLK(rclk), .Q(alu_addsub_subtract_e[56]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[57](.D(exu_n16331), .CLK(rclk), .Q(alu_addsub_subtract_e[57]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[58](.D(exu_n16330), .CLK(rclk), .Q(alu_addsub_subtract_e[58]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[59](.D(exu_n16329), .CLK(rclk), .Q(alu_addsub_subtract_e[59]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[60](.D(exu_n16328), .CLK(rclk), .Q(alu_addsub_subtract_e[60]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[61](.D(exu_n16327), .CLK(rclk), .Q(alu_addsub_subtract_e[61]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[62](.D(exu_n16326), .CLK(rclk), .Q(alu_addsub_subtract_e[62]));
DFFPOSX1 alu_addsub_sub_dff_q_reg[63](.D(exu_n16325), .CLK(rclk), .Q(alu_addsub_subtract_e[63]));
DFFPOSX1 div_mul_result_dff_q_reg[0](.D(exu_n30124), .CLK(rclk), .Q(div_mul_result[0]));
DFFPOSX1 div_mul_result_dff_q_reg[1](.D(exu_n30113), .CLK(rclk), .Q(div_mul_result[1]));
DFFPOSX1 div_mul_result_dff_q_reg[2](.D(exu_n30102), .CLK(rclk), .Q(div_mul_result[2]));
DFFPOSX1 div_mul_result_dff_q_reg[3](.D(exu_n30091), .CLK(rclk), .Q(div_mul_result[3]));
DFFPOSX1 div_mul_result_dff_q_reg[4](.D(exu_n30083), .CLK(rclk), .Q(div_mul_result[4]));
DFFPOSX1 div_mul_result_dff_q_reg[5](.D(exu_n30082), .CLK(rclk), .Q(div_mul_result[5]));
DFFPOSX1 div_mul_result_dff_q_reg[6](.D(exu_n30081), .CLK(rclk), .Q(div_mul_result[6]));
DFFPOSX1 div_mul_result_dff_q_reg[7](.D(exu_n30144), .CLK(rclk), .Q(div_mul_result[7]));
DFFPOSX1 div_mul_result_dff_q_reg[8](.D(exu_n30143), .CLK(rclk), .Q(div_mul_result[8]));
DFFPOSX1 div_mul_result_dff_q_reg[9](.D(exu_n30142), .CLK(rclk), .Q(div_mul_result[9]));
DFFPOSX1 div_mul_result_dff_q_reg[10](.D(exu_n30141), .CLK(rclk), .Q(div_mul_result[10]));
DFFPOSX1 div_mul_result_dff_q_reg[11](.D(exu_n30140), .CLK(rclk), .Q(div_mul_result[11]));
DFFPOSX1 div_mul_result_dff_q_reg[12](.D(exu_n30139), .CLK(rclk), .Q(div_mul_result[12]));
DFFPOSX1 div_mul_result_dff_q_reg[13](.D(exu_n30138), .CLK(rclk), .Q(div_mul_result[13]));
DFFPOSX1 div_mul_result_dff_q_reg[14](.D(exu_n30137), .CLK(rclk), .Q(div_mul_result[14]));
DFFPOSX1 div_mul_result_dff_q_reg[15](.D(exu_n30136), .CLK(rclk), .Q(div_mul_result[15]));
DFFPOSX1 div_mul_result_dff_q_reg[16](.D(exu_n30135), .CLK(rclk), .Q(div_mul_result[16]));
DFFPOSX1 div_mul_result_dff_q_reg[17](.D(exu_n30134), .CLK(rclk), .Q(div_mul_result[17]));
DFFPOSX1 div_mul_result_dff_q_reg[18](.D(exu_n30133), .CLK(rclk), .Q(div_mul_result[18]));
DFFPOSX1 div_mul_result_dff_q_reg[19](.D(exu_n30132), .CLK(rclk), .Q(div_mul_result[19]));
DFFPOSX1 div_mul_result_dff_q_reg[20](.D(exu_n30131), .CLK(rclk), .Q(div_mul_result[20]));
DFFPOSX1 div_mul_result_dff_q_reg[21](.D(exu_n30130), .CLK(rclk), .Q(div_mul_result[21]));
DFFPOSX1 div_mul_result_dff_q_reg[22](.D(exu_n30129), .CLK(rclk), .Q(div_mul_result[22]));
DFFPOSX1 div_mul_result_dff_q_reg[23](.D(exu_n30128), .CLK(rclk), .Q(div_mul_result[23]));
DFFPOSX1 div_mul_result_dff_q_reg[24](.D(exu_n30127), .CLK(rclk), .Q(div_mul_result[24]));
DFFPOSX1 div_mul_result_dff_q_reg[25](.D(exu_n30126), .CLK(rclk), .Q(div_mul_result[25]));
DFFPOSX1 div_mul_result_dff_q_reg[26](.D(exu_n30125), .CLK(rclk), .Q(div_mul_result[26]));
DFFPOSX1 div_mul_result_dff_q_reg[27](.D(exu_n30123), .CLK(rclk), .Q(div_mul_result[27]));
DFFPOSX1 div_mul_result_dff_q_reg[28](.D(exu_n30122), .CLK(rclk), .Q(div_mul_result[28]));
DFFPOSX1 div_mul_result_dff_q_reg[29](.D(exu_n30121), .CLK(rclk), .Q(div_mul_result[29]));
DFFPOSX1 div_mul_result_dff_q_reg[30](.D(exu_n30120), .CLK(rclk), .Q(div_mul_result[30]));
DFFPOSX1 div_mul_result_dff_q_reg[31](.D(exu_n30119), .CLK(rclk), .Q(div_mul_result[31]));
DFFPOSX1 div_mul_result_dff_q_reg[32](.D(exu_n30118), .CLK(rclk), .Q(div_mul_result[32]));
DFFPOSX1 div_mul_result_dff_q_reg[33](.D(exu_n30117), .CLK(rclk), .Q(div_mul_result[33]));
DFFPOSX1 div_mul_result_dff_q_reg[34](.D(exu_n30116), .CLK(rclk), .Q(div_mul_result[34]));
DFFPOSX1 div_mul_result_dff_q_reg[35](.D(exu_n30115), .CLK(rclk), .Q(div_mul_result[35]));
DFFPOSX1 div_mul_result_dff_q_reg[36](.D(exu_n30114), .CLK(rclk), .Q(div_mul_result[36]));
DFFPOSX1 div_mul_result_dff_q_reg[37](.D(exu_n30112), .CLK(rclk), .Q(div_mul_result[37]));
DFFPOSX1 div_mul_result_dff_q_reg[38](.D(exu_n30111), .CLK(rclk), .Q(div_mul_result[38]));
DFFPOSX1 div_mul_result_dff_q_reg[39](.D(exu_n30110), .CLK(rclk), .Q(div_mul_result[39]));
DFFPOSX1 div_mul_result_dff_q_reg[40](.D(exu_n30109), .CLK(rclk), .Q(div_mul_result[40]));
DFFPOSX1 div_mul_result_dff_q_reg[41](.D(exu_n30108), .CLK(rclk), .Q(div_mul_result[41]));
DFFPOSX1 div_mul_result_dff_q_reg[42](.D(exu_n30107), .CLK(rclk), .Q(div_mul_result[42]));
DFFPOSX1 div_mul_result_dff_q_reg[43](.D(exu_n30106), .CLK(rclk), .Q(div_mul_result[43]));
DFFPOSX1 div_mul_result_dff_q_reg[44](.D(exu_n30105), .CLK(rclk), .Q(div_mul_result[44]));
DFFPOSX1 div_mul_result_dff_q_reg[45](.D(exu_n30104), .CLK(rclk), .Q(div_mul_result[45]));
DFFPOSX1 div_mul_result_dff_q_reg[46](.D(exu_n30103), .CLK(rclk), .Q(div_mul_result[46]));
DFFPOSX1 div_mul_result_dff_q_reg[47](.D(exu_n30101), .CLK(rclk), .Q(div_mul_result[47]));
DFFPOSX1 div_mul_result_dff_q_reg[48](.D(exu_n30100), .CLK(rclk), .Q(div_mul_result[48]));
DFFPOSX1 div_mul_result_dff_q_reg[49](.D(exu_n30099), .CLK(rclk), .Q(div_mul_result[49]));
DFFPOSX1 div_mul_result_dff_q_reg[50](.D(exu_n30098), .CLK(rclk), .Q(div_mul_result[50]));
DFFPOSX1 div_mul_result_dff_q_reg[51](.D(exu_n30097), .CLK(rclk), .Q(div_mul_result[51]));
DFFPOSX1 div_mul_result_dff_q_reg[52](.D(exu_n30096), .CLK(rclk), .Q(div_mul_result[52]));
DFFPOSX1 div_mul_result_dff_q_reg[53](.D(exu_n30095), .CLK(rclk), .Q(div_mul_result[53]));
DFFPOSX1 div_mul_result_dff_q_reg[54](.D(exu_n30094), .CLK(rclk), .Q(div_mul_result[54]));
DFFPOSX1 div_mul_result_dff_q_reg[55](.D(exu_n30093), .CLK(rclk), .Q(div_mul_result[55]));
DFFPOSX1 div_mul_result_dff_q_reg[56](.D(exu_n30092), .CLK(rclk), .Q(div_mul_result[56]));
DFFPOSX1 div_mul_result_dff_q_reg[57](.D(exu_n30090), .CLK(rclk), .Q(div_mul_result[57]));
DFFPOSX1 div_mul_result_dff_q_reg[58](.D(exu_n30089), .CLK(rclk), .Q(div_mul_result[58]));
DFFPOSX1 div_mul_result_dff_q_reg[59](.D(exu_n30088), .CLK(rclk), .Q(div_mul_result[59]));
DFFPOSX1 div_mul_result_dff_q_reg[60](.D(exu_n30087), .CLK(rclk), .Q(div_mul_result[60]));
DFFPOSX1 div_mul_result_dff_q_reg[61](.D(exu_n30086), .CLK(rclk), .Q(div_mul_result[61]));
DFFPOSX1 div_mul_result_dff_q_reg[62](.D(exu_n30085), .CLK(rclk), .Q(div_mul_result[62]));
DFFPOSX1 div_mul_result_dff_q_reg[63](.D(exu_n30084), .CLK(rclk), .Q(div_mul_result[63]));
DFFPOSX1 div_x_dff_q_reg[0](.D(exu_n30059), .CLK(rclk), .Q(div_x[0]));
DFFPOSX1 div_x_dff_q_reg[1](.D(exu_n30048), .CLK(rclk), .Q(div_x[1]));
DFFPOSX1 div_x_dff_q_reg[2](.D(exu_n30037), .CLK(rclk), .Q(div_x[2]));
DFFPOSX1 div_x_dff_q_reg[3](.D(exu_n30026), .CLK(rclk), .Q(div_x[3]));
DFFPOSX1 div_x_dff_q_reg[4](.D(exu_n30018), .CLK(rclk), .Q(div_x[4]));
DFFPOSX1 div_x_dff_q_reg[5](.D(exu_n30017), .CLK(rclk), .Q(div_x[5]));
DFFPOSX1 div_x_dff_q_reg[6](.D(exu_n30016), .CLK(rclk), .Q(div_x[6]));
DFFPOSX1 div_x_dff_q_reg[7](.D(exu_n30079), .CLK(rclk), .Q(div_x[7]));
DFFPOSX1 div_x_dff_q_reg[8](.D(exu_n30078), .CLK(rclk), .Q(div_x[8]));
DFFPOSX1 div_x_dff_q_reg[9](.D(exu_n30077), .CLK(rclk), .Q(div_x[9]));
DFFPOSX1 div_x_dff_q_reg[10](.D(exu_n30076), .CLK(rclk), .Q(div_x[10]));
DFFPOSX1 div_x_dff_q_reg[11](.D(exu_n30075), .CLK(rclk), .Q(div_x[11]));
DFFPOSX1 div_x_dff_q_reg[12](.D(exu_n30074), .CLK(rclk), .Q(div_x[12]));
DFFPOSX1 div_x_dff_q_reg[13](.D(exu_n30073), .CLK(rclk), .Q(div_x[13]));
DFFPOSX1 div_x_dff_q_reg[14](.D(exu_n30072), .CLK(rclk), .Q(div_x[14]));
DFFPOSX1 div_x_dff_q_reg[15](.D(exu_n30071), .CLK(rclk), .Q(div_x[15]));
DFFPOSX1 div_x_dff_q_reg[16](.D(exu_n30070), .CLK(rclk), .Q(div_x[16]));
DFFPOSX1 div_x_dff_q_reg[17](.D(exu_n30069), .CLK(rclk), .Q(div_x[17]));
DFFPOSX1 div_x_dff_q_reg[18](.D(exu_n30068), .CLK(rclk), .Q(div_x[18]));
DFFPOSX1 div_x_dff_q_reg[19](.D(exu_n30067), .CLK(rclk), .Q(div_x[19]));
DFFPOSX1 div_x_dff_q_reg[20](.D(exu_n30066), .CLK(rclk), .Q(div_x[20]));
DFFPOSX1 div_x_dff_q_reg[21](.D(exu_n30065), .CLK(rclk), .Q(div_x[21]));
DFFPOSX1 div_x_dff_q_reg[22](.D(exu_n30064), .CLK(rclk), .Q(div_x[22]));
DFFPOSX1 div_x_dff_q_reg[23](.D(exu_n30063), .CLK(rclk), .Q(div_x[23]));
DFFPOSX1 div_x_dff_q_reg[24](.D(exu_n30062), .CLK(rclk), .Q(div_x[24]));
DFFPOSX1 div_x_dff_q_reg[25](.D(exu_n30061), .CLK(rclk), .Q(div_x[25]));
DFFPOSX1 div_x_dff_q_reg[26](.D(exu_n30060), .CLK(rclk), .Q(div_x[26]));
DFFPOSX1 div_x_dff_q_reg[27](.D(exu_n30058), .CLK(rclk), .Q(div_x[27]));
DFFPOSX1 div_x_dff_q_reg[28](.D(exu_n30057), .CLK(rclk), .Q(div_x[28]));
DFFPOSX1 div_x_dff_q_reg[29](.D(exu_n30056), .CLK(rclk), .Q(div_x[29]));
DFFPOSX1 div_x_dff_q_reg[30](.D(exu_n30055), .CLK(rclk), .Q(div_x[30]));
DFFPOSX1 div_x_dff_q_reg[31](.D(exu_n30054), .CLK(rclk), .Q(div_x[31]));
DFFPOSX1 div_x_dff_q_reg[32](.D(exu_n30053), .CLK(rclk), .Q(div_x[32]));
DFFPOSX1 div_x_dff_q_reg[33](.D(exu_n30052), .CLK(rclk), .Q(div_x[33]));
DFFPOSX1 div_x_dff_q_reg[34](.D(exu_n30051), .CLK(rclk), .Q(div_x[34]));
DFFPOSX1 div_x_dff_q_reg[35](.D(exu_n30050), .CLK(rclk), .Q(div_x[35]));
DFFPOSX1 div_x_dff_q_reg[36](.D(exu_n30049), .CLK(rclk), .Q(div_x[36]));
DFFPOSX1 div_x_dff_q_reg[37](.D(exu_n30047), .CLK(rclk), .Q(div_x[37]));
DFFPOSX1 div_x_dff_q_reg[38](.D(exu_n30046), .CLK(rclk), .Q(div_x[38]));
DFFPOSX1 div_x_dff_q_reg[39](.D(exu_n30045), .CLK(rclk), .Q(div_x[39]));
DFFPOSX1 div_x_dff_q_reg[40](.D(exu_n30044), .CLK(rclk), .Q(div_x[40]));
DFFPOSX1 div_x_dff_q_reg[41](.D(exu_n30043), .CLK(rclk), .Q(div_x[41]));
DFFPOSX1 div_x_dff_q_reg[42](.D(exu_n30042), .CLK(rclk), .Q(div_x[42]));
DFFPOSX1 div_x_dff_q_reg[43](.D(exu_n30041), .CLK(rclk), .Q(div_x[43]));
DFFPOSX1 div_x_dff_q_reg[44](.D(exu_n30040), .CLK(rclk), .Q(div_x[44]));
DFFPOSX1 div_x_dff_q_reg[45](.D(exu_n30039), .CLK(rclk), .Q(div_x[45]));
DFFPOSX1 div_x_dff_q_reg[46](.D(exu_n30038), .CLK(rclk), .Q(div_x[46]));
DFFPOSX1 div_x_dff_q_reg[47](.D(exu_n30036), .CLK(rclk), .Q(div_x[47]));
DFFPOSX1 div_x_dff_q_reg[48](.D(exu_n30035), .CLK(rclk), .Q(div_x[48]));
DFFPOSX1 div_x_dff_q_reg[49](.D(exu_n30034), .CLK(rclk), .Q(div_x[49]));
DFFPOSX1 div_x_dff_q_reg[50](.D(exu_n30033), .CLK(rclk), .Q(div_x[50]));
DFFPOSX1 div_x_dff_q_reg[51](.D(exu_n30032), .CLK(rclk), .Q(div_x[51]));
DFFPOSX1 div_x_dff_q_reg[52](.D(exu_n30031), .CLK(rclk), .Q(div_x[52]));
DFFPOSX1 div_x_dff_q_reg[53](.D(exu_n30030), .CLK(rclk), .Q(div_x[53]));
DFFPOSX1 div_x_dff_q_reg[54](.D(exu_n30029), .CLK(rclk), .Q(div_x[54]));
DFFPOSX1 div_x_dff_q_reg[55](.D(exu_n30028), .CLK(rclk), .Q(div_x[55]));
DFFPOSX1 div_x_dff_q_reg[56](.D(exu_n30027), .CLK(rclk), .Q(div_x[56]));
DFFPOSX1 div_x_dff_q_reg[57](.D(exu_n30025), .CLK(rclk), .Q(div_x[57]));
DFFPOSX1 div_x_dff_q_reg[58](.D(exu_n30024), .CLK(rclk), .Q(div_x[58]));
DFFPOSX1 div_x_dff_q_reg[59](.D(exu_n30023), .CLK(rclk), .Q(div_x[59]));
DFFPOSX1 div_x_dff_q_reg[60](.D(exu_n30022), .CLK(rclk), .Q(div_x[60]));
DFFPOSX1 div_x_dff_q_reg[61](.D(exu_n30021), .CLK(rclk), .Q(div_x[61]));
DFFPOSX1 div_x_dff_q_reg[62](.D(exu_n30020), .CLK(rclk), .Q(div_x[62]));
DFFPOSX1 div_x_dff_q_reg[63](.D(exu_n30019), .CLK(rclk), .Q(div_ecl_x_msb));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[0](.D(exu_n29994), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[0]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[1](.D(exu_n29983), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[1]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[2](.D(exu_n29972), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[2]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[3](.D(exu_n29961), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[3]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[4](.D(exu_n29953), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[4]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[5](.D(exu_n29952), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[5]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[6](.D(exu_n29951), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[6]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[7](.D(exu_n30014), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[7]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[8](.D(exu_n30013), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[8]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[9](.D(exu_n30012), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[9]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[10](.D(exu_n30011), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[10]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[11](.D(exu_n30010), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[11]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[12](.D(exu_n30009), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[12]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[13](.D(exu_n30008), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[13]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[14](.D(exu_n30007), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[14]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[15](.D(exu_n30006), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[15]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[16](.D(exu_n30005), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[16]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[17](.D(exu_n30004), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[17]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[18](.D(exu_n30003), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[18]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[19](.D(exu_n30002), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[19]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[20](.D(exu_n30001), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[20]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[21](.D(exu_n30000), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[21]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[22](.D(exu_n29999), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[22]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[23](.D(exu_n29998), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[23]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[24](.D(exu_n29997), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[24]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[25](.D(exu_n29996), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[25]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[26](.D(exu_n29995), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[26]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[27](.D(exu_n29993), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[27]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[28](.D(exu_n29992), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[28]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[29](.D(exu_n29991), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[29]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[30](.D(exu_n29990), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[30]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[31](.D(exu_n29989), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[31]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[32](.D(exu_n29988), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[32]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[33](.D(exu_n29987), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[33]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[34](.D(exu_n29986), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[34]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[35](.D(exu_n29985), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[35]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[36](.D(exu_n29984), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[36]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[37](.D(exu_n29982), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[37]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[38](.D(exu_n29981), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[38]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[39](.D(exu_n29980), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[39]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[40](.D(exu_n29979), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[40]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[41](.D(exu_n29978), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[41]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[42](.D(exu_n29977), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[42]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[43](.D(exu_n29976), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[43]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[44](.D(exu_n29975), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[44]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[45](.D(exu_n29974), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[45]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[46](.D(exu_n29973), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[46]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[47](.D(exu_n29971), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[47]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[48](.D(exu_n29970), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[48]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[49](.D(exu_n29969), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[49]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[50](.D(exu_n29968), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[50]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[51](.D(exu_n29967), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[51]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[52](.D(exu_n29966), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[52]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[53](.D(exu_n29965), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[53]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[54](.D(exu_n29964), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[54]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[55](.D(exu_n29963), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[55]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[56](.D(exu_n29962), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[56]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[57](.D(exu_n29960), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[57]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[58](.D(exu_n29959), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[58]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[59](.D(exu_n29958), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[59]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[60](.D(exu_n29957), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[60]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[61](.D(exu_n29956), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[61]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[62](.D(exu_n29955), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[62]));
DFFPOSX1 ecc_rs3_data_e2m_q_reg[63](.D(exu_n29954), .CLK(rclk), .Q(ecc_exu_lsu_rs3_data_m[63]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[0](.D(exu_n29929), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[0]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[1](.D(exu_n29919), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[1]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[2](.D(exu_n29908), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[2]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[3](.D(exu_n29897), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[3]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[4](.D(exu_n29889), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[4]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[5](.D(exu_n29888), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[5]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[6](.D(exu_n29887), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[6]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[7](.D(exu_n29949), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[7]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[8](.D(exu_n29948), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[8]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[9](.D(exu_n29947), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[9]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[10](.D(exu_n29946), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[10]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[11](.D(exu_n29945), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[11]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[12](.D(exu_n29944), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[12]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[13](.D(exu_n29943), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[13]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[14](.D(exu_n29942), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[14]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[15](.D(exu_n29941), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[15]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[16](.D(exu_n29940), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[16]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[17](.D(exu_n29939), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[17]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[18](.D(exu_n29938), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[18]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[19](.D(exu_n29937), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[19]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[20](.D(exu_n29936), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[20]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[21](.D(exu_n29935), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[21]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[22](.D(exu_n29934), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[22]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[23](.D(exu_n29933), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[23]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[24](.D(exu_n29932), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[24]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[25](.D(exu_n29931), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[25]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[26](.D(exu_n29930), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[26]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[27](.D(exu_n29928), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[27]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[28](.D(exu_n29927), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[28]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[29](.D(exu_n29926), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[29]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[30](.D(exu_n29925), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[30]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[31](.D(exu_n19290), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[31]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[32](.D(exu_n29924), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[32]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[33](.D(exu_n29923), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[33]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[34](.D(exu_n29922), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[34]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[35](.D(exu_n29921), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[35]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[36](.D(exu_n29920), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[36]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[37](.D(exu_n29918), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[37]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[38](.D(exu_n29917), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[38]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[39](.D(exu_n29916), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[39]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[40](.D(exu_n29915), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[40]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[41](.D(exu_n29914), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[41]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[42](.D(exu_n29913), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[42]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[43](.D(exu_n29912), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[43]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[44](.D(exu_n29911), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[44]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[45](.D(exu_n29910), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[45]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[46](.D(exu_n29909), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[46]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[47](.D(exu_n29907), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[47]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[48](.D(exu_n29906), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[48]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[49](.D(exu_n29905), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[49]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[50](.D(exu_n29904), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[50]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[51](.D(exu_n29903), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[51]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[52](.D(exu_n29902), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[52]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[53](.D(exu_n29901), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[53]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[54](.D(exu_n29900), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[54]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[55](.D(exu_n29899), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[55]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[56](.D(exu_n29898), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[56]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[57](.D(exu_n29896), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[57]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[58](.D(exu_n29895), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[58]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[59](.D(exu_n29894), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[59]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[60](.D(exu_n29893), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[60]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[61](.D(exu_n29892), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[61]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[62](.D(exu_n29891), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[62]));
DFFPOSX1 ecc_rs2_data_e2m_q_reg[63](.D(exu_n29890), .CLK(rclk), .Q(ecc_byp_alu_rs2_data_m[63]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[0](.D(exu_n29865), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[0]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[1](.D(exu_n29854), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[1]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[2](.D(exu_n29843), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[2]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[3](.D(exu_n29832), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[3]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[4](.D(exu_n29824), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[4]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[5](.D(exu_n29823), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[5]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[6](.D(exu_n29822), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[6]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[7](.D(exu_n29885), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[7]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[8](.D(exu_n29884), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[8]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[9](.D(exu_n29883), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[9]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[10](.D(exu_n29882), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[10]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[11](.D(exu_n29881), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[11]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[12](.D(exu_n29880), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[12]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[13](.D(exu_n29879), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[13]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[14](.D(exu_n29878), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[14]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[15](.D(exu_n29877), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[15]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[16](.D(exu_n29876), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[16]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[17](.D(exu_n29875), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[17]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[18](.D(exu_n29874), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[18]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[19](.D(exu_n29873), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[19]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[20](.D(exu_n29872), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[20]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[21](.D(exu_n29871), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[21]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[22](.D(exu_n29870), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[22]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[23](.D(exu_n29869), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[23]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[24](.D(exu_n29868), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[24]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[25](.D(exu_n29867), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[25]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[26](.D(exu_n29866), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[26]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[27](.D(exu_n29864), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[27]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[28](.D(exu_n29863), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[28]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[29](.D(exu_n29862), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[29]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[30](.D(exu_n29861), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[30]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[31](.D(exu_n29860), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[31]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[32](.D(exu_n29859), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[32]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[33](.D(exu_n29858), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[33]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[34](.D(exu_n29857), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[34]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[35](.D(exu_n29856), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[35]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[36](.D(exu_n29855), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[36]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[37](.D(exu_n29853), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[37]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[38](.D(exu_n29852), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[38]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[39](.D(exu_n29851), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[39]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[40](.D(exu_n29850), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[40]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[41](.D(exu_n29849), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[41]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[42](.D(exu_n29848), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[42]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[43](.D(exu_n29847), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[43]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[44](.D(exu_n29846), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[44]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[45](.D(exu_n29845), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[45]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[46](.D(exu_n29844), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[46]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[47](.D(exu_n29842), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[47]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[48](.D(exu_n29841), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[48]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[49](.D(exu_n29840), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[49]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[50](.D(exu_n29839), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[50]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[51](.D(exu_n29838), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[51]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[52](.D(exu_n29837), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[52]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[53](.D(exu_n29836), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[53]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[54](.D(exu_n29835), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[54]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[55](.D(exu_n29834), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[55]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[56](.D(exu_n29833), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[56]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[57](.D(exu_n29831), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[57]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[58](.D(exu_n29830), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[58]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[59](.D(exu_n29829), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[59]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[60](.D(exu_n29828), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[60]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[61](.D(exu_n29827), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[61]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[62](.D(exu_n29826), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[62]));
DFFPOSX1 ecc_rs1_data_e2m_q_reg[63](.D(exu_n29825), .CLK(rclk), .Q(ecc_byp_ecc_rcc_data_m[63]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[0](.D(exu_n29800), .CLK(rclk), .Q(byp_alu_rcc_data_e[0]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[1](.D(exu_n29789), .CLK(rclk), .Q(byp_alu_rcc_data_e[1]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[2](.D(exu_n29778), .CLK(rclk), .Q(byp_alu_rcc_data_e[2]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[3](.D(exu_n29767), .CLK(rclk), .Q(byp_alu_rcc_data_e[3]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[4](.D(exu_n29759), .CLK(rclk), .Q(byp_alu_rcc_data_e[4]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[5](.D(exu_n29758), .CLK(rclk), .Q(byp_alu_rcc_data_e[5]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[6](.D(exu_n29757), .CLK(rclk), .Q(byp_alu_rcc_data_e[6]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[7](.D(exu_n29820), .CLK(rclk), .Q(byp_alu_rcc_data_e[7]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[8](.D(exu_n29819), .CLK(rclk), .Q(byp_alu_rcc_data_e[8]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[9](.D(exu_n29818), .CLK(rclk), .Q(byp_alu_rcc_data_e[9]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[10](.D(exu_n29817), .CLK(rclk), .Q(byp_alu_rcc_data_e[10]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[11](.D(exu_n29816), .CLK(rclk), .Q(byp_alu_rcc_data_e[11]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[12](.D(exu_n29815), .CLK(rclk), .Q(byp_alu_rcc_data_e[12]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[13](.D(exu_n29814), .CLK(rclk), .Q(byp_alu_rcc_data_e[13]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[14](.D(exu_n29813), .CLK(rclk), .Q(byp_alu_rcc_data_e[14]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[15](.D(exu_n29812), .CLK(rclk), .Q(byp_alu_rcc_data_e[15]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[16](.D(exu_n29811), .CLK(rclk), .Q(byp_alu_rcc_data_e[16]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[17](.D(exu_n29810), .CLK(rclk), .Q(byp_alu_rcc_data_e[17]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[18](.D(exu_n29809), .CLK(rclk), .Q(byp_alu_rcc_data_e[18]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[19](.D(exu_n29808), .CLK(rclk), .Q(byp_alu_rcc_data_e[19]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[20](.D(exu_n29807), .CLK(rclk), .Q(byp_alu_rcc_data_e[20]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[21](.D(exu_n29806), .CLK(rclk), .Q(byp_alu_rcc_data_e[21]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[22](.D(exu_n29805), .CLK(rclk), .Q(byp_alu_rcc_data_e[22]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[23](.D(exu_n29804), .CLK(rclk), .Q(byp_alu_rcc_data_e[23]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[24](.D(exu_n29803), .CLK(rclk), .Q(byp_alu_rcc_data_e[24]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[25](.D(exu_n29802), .CLK(rclk), .Q(byp_alu_rcc_data_e[25]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[26](.D(exu_n29801), .CLK(rclk), .Q(byp_alu_rcc_data_e[26]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[27](.D(exu_n29799), .CLK(rclk), .Q(byp_alu_rcc_data_e[27]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[28](.D(exu_n29798), .CLK(rclk), .Q(byp_alu_rcc_data_e[28]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[29](.D(exu_n29797), .CLK(rclk), .Q(byp_alu_rcc_data_e[29]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[30](.D(exu_n29796), .CLK(rclk), .Q(byp_alu_rcc_data_e[30]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[31](.D(exu_n29795), .CLK(rclk), .Q(byp_alu_rcc_data_e[31]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[32](.D(exu_n29794), .CLK(rclk), .Q(byp_alu_rcc_data_e[32]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[33](.D(exu_n29793), .CLK(rclk), .Q(byp_alu_rcc_data_e[33]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[34](.D(exu_n29792), .CLK(rclk), .Q(byp_alu_rcc_data_e[34]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[35](.D(exu_n29791), .CLK(rclk), .Q(byp_alu_rcc_data_e[35]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[36](.D(exu_n29790), .CLK(rclk), .Q(byp_alu_rcc_data_e[36]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[37](.D(exu_n29788), .CLK(rclk), .Q(byp_alu_rcc_data_e[37]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[38](.D(exu_n29787), .CLK(rclk), .Q(byp_alu_rcc_data_e[38]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[39](.D(exu_n29786), .CLK(rclk), .Q(byp_alu_rcc_data_e[39]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[40](.D(exu_n29785), .CLK(rclk), .Q(byp_alu_rcc_data_e[40]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[41](.D(exu_n29784), .CLK(rclk), .Q(byp_alu_rcc_data_e[41]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[42](.D(exu_n29783), .CLK(rclk), .Q(byp_alu_rcc_data_e[42]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[43](.D(exu_n29782), .CLK(rclk), .Q(byp_alu_rcc_data_e[43]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[44](.D(exu_n29781), .CLK(rclk), .Q(byp_alu_rcc_data_e[44]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[45](.D(exu_n29780), .CLK(rclk), .Q(byp_alu_rcc_data_e[45]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[46](.D(exu_n29779), .CLK(rclk), .Q(byp_alu_rcc_data_e[46]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[47](.D(exu_n29777), .CLK(rclk), .Q(byp_alu_rcc_data_e[47]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[48](.D(exu_n29776), .CLK(rclk), .Q(byp_alu_rcc_data_e[48]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[49](.D(exu_n29775), .CLK(rclk), .Q(byp_alu_rcc_data_e[49]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[50](.D(exu_n29774), .CLK(rclk), .Q(byp_alu_rcc_data_e[50]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[51](.D(exu_n29773), .CLK(rclk), .Q(byp_alu_rcc_data_e[51]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[52](.D(exu_n29772), .CLK(rclk), .Q(byp_alu_rcc_data_e[52]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[53](.D(exu_n29771), .CLK(rclk), .Q(byp_alu_rcc_data_e[53]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[54](.D(exu_n29770), .CLK(rclk), .Q(byp_alu_rcc_data_e[54]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[55](.D(exu_n29769), .CLK(rclk), .Q(byp_alu_rcc_data_e[55]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[56](.D(exu_n29768), .CLK(rclk), .Q(byp_alu_rcc_data_e[56]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[57](.D(exu_n29766), .CLK(rclk), .Q(byp_alu_rcc_data_e[57]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[58](.D(exu_n29765), .CLK(rclk), .Q(byp_alu_rcc_data_e[58]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[59](.D(exu_n29764), .CLK(rclk), .Q(byp_alu_rcc_data_e[59]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[60](.D(exu_n29763), .CLK(rclk), .Q(byp_alu_rcc_data_e[60]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[61](.D(exu_n29762), .CLK(rclk), .Q(byp_alu_rcc_data_e[61]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[62](.D(exu_n29761), .CLK(rclk), .Q(byp_alu_rcc_data_e[62]));
DFFPOSX1 bypass_rcc_data_dff_q_reg[63](.D(exu_n29760), .CLK(rclk), .Q(exu_ifu_regn_e));
DFFPOSX1 bypass_rs3_data_dff_q_reg[0](.D(exu_n29735), .CLK(rclk), .Q(exu_spu_rs3_data_e[0]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[1](.D(exu_n29724), .CLK(rclk), .Q(exu_spu_rs3_data_e[1]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[2](.D(exu_n29713), .CLK(rclk), .Q(exu_spu_rs3_data_e[2]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[3](.D(exu_n29702), .CLK(rclk), .Q(exu_spu_rs3_data_e[3]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[4](.D(exu_n29694), .CLK(rclk), .Q(exu_spu_rs3_data_e[4]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[5](.D(exu_n29693), .CLK(rclk), .Q(exu_spu_rs3_data_e[5]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[6](.D(exu_n29692), .CLK(rclk), .Q(exu_spu_rs3_data_e[6]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[7](.D(exu_n29755), .CLK(rclk), .Q(exu_spu_rs3_data_e[7]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[8](.D(exu_n29754), .CLK(rclk), .Q(exu_spu_rs3_data_e[8]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[9](.D(exu_n29753), .CLK(rclk), .Q(exu_spu_rs3_data_e[9]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[10](.D(exu_n29752), .CLK(rclk), .Q(exu_spu_rs3_data_e[10]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[11](.D(exu_n29751), .CLK(rclk), .Q(exu_spu_rs3_data_e[11]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[12](.D(exu_n29750), .CLK(rclk), .Q(exu_spu_rs3_data_e[12]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[13](.D(exu_n29749), .CLK(rclk), .Q(exu_spu_rs3_data_e[13]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[14](.D(exu_n29748), .CLK(rclk), .Q(exu_spu_rs3_data_e[14]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[15](.D(exu_n29747), .CLK(rclk), .Q(exu_spu_rs3_data_e[15]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[16](.D(exu_n29746), .CLK(rclk), .Q(exu_spu_rs3_data_e[16]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[17](.D(exu_n29745), .CLK(rclk), .Q(exu_spu_rs3_data_e[17]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[18](.D(exu_n29744), .CLK(rclk), .Q(exu_spu_rs3_data_e[18]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[19](.D(exu_n29743), .CLK(rclk), .Q(exu_spu_rs3_data_e[19]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[20](.D(exu_n29742), .CLK(rclk), .Q(exu_spu_rs3_data_e[20]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[21](.D(exu_n29741), .CLK(rclk), .Q(exu_spu_rs3_data_e[21]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[22](.D(exu_n29740), .CLK(rclk), .Q(exu_spu_rs3_data_e[22]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[23](.D(exu_n29739), .CLK(rclk), .Q(exu_spu_rs3_data_e[23]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[24](.D(exu_n29738), .CLK(rclk), .Q(exu_spu_rs3_data_e[24]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[25](.D(exu_n29737), .CLK(rclk), .Q(exu_spu_rs3_data_e[25]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[26](.D(exu_n29736), .CLK(rclk), .Q(exu_spu_rs3_data_e[26]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[27](.D(exu_n29734), .CLK(rclk), .Q(exu_spu_rs3_data_e[27]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[28](.D(exu_n29733), .CLK(rclk), .Q(exu_spu_rs3_data_e[28]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[29](.D(exu_n29732), .CLK(rclk), .Q(exu_spu_rs3_data_e[29]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[30](.D(exu_n29731), .CLK(rclk), .Q(exu_spu_rs3_data_e[30]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[31](.D(exu_n29730), .CLK(rclk), .Q(exu_spu_rs3_data_e[31]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[32](.D(exu_n29729), .CLK(rclk), .Q(exu_spu_rs3_data_e[32]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[33](.D(exu_n29728), .CLK(rclk), .Q(exu_spu_rs3_data_e[33]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[34](.D(exu_n29727), .CLK(rclk), .Q(exu_spu_rs3_data_e[34]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[35](.D(exu_n29726), .CLK(rclk), .Q(exu_spu_rs3_data_e[35]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[36](.D(exu_n29725), .CLK(rclk), .Q(exu_spu_rs3_data_e[36]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[37](.D(exu_n29723), .CLK(rclk), .Q(exu_spu_rs3_data_e[37]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[38](.D(exu_n29722), .CLK(rclk), .Q(exu_spu_rs3_data_e[38]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[39](.D(exu_n29721), .CLK(rclk), .Q(exu_spu_rs3_data_e[39]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[40](.D(exu_n29720), .CLK(rclk), .Q(exu_spu_rs3_data_e[40]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[41](.D(exu_n29719), .CLK(rclk), .Q(exu_spu_rs3_data_e[41]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[42](.D(exu_n29718), .CLK(rclk), .Q(exu_spu_rs3_data_e[42]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[43](.D(exu_n29717), .CLK(rclk), .Q(exu_spu_rs3_data_e[43]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[44](.D(exu_n29716), .CLK(rclk), .Q(exu_spu_rs3_data_e[44]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[45](.D(exu_n29715), .CLK(rclk), .Q(exu_spu_rs3_data_e[45]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[46](.D(exu_n29714), .CLK(rclk), .Q(exu_spu_rs3_data_e[46]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[47](.D(exu_n29712), .CLK(rclk), .Q(exu_spu_rs3_data_e[47]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[48](.D(exu_n29711), .CLK(rclk), .Q(exu_spu_rs3_data_e[48]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[49](.D(exu_n29710), .CLK(rclk), .Q(exu_spu_rs3_data_e[49]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[50](.D(exu_n29709), .CLK(rclk), .Q(exu_spu_rs3_data_e[50]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[51](.D(exu_n29708), .CLK(rclk), .Q(exu_spu_rs3_data_e[51]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[52](.D(exu_n29707), .CLK(rclk), .Q(exu_spu_rs3_data_e[52]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[53](.D(exu_n29706), .CLK(rclk), .Q(exu_spu_rs3_data_e[53]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[54](.D(exu_n29705), .CLK(rclk), .Q(exu_spu_rs3_data_e[54]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[55](.D(exu_n29704), .CLK(rclk), .Q(exu_spu_rs3_data_e[55]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[56](.D(exu_n29703), .CLK(rclk), .Q(exu_spu_rs3_data_e[56]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[57](.D(exu_n29701), .CLK(rclk), .Q(exu_spu_rs3_data_e[57]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[58](.D(exu_n29700), .CLK(rclk), .Q(exu_spu_rs3_data_e[58]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[59](.D(exu_n29699), .CLK(rclk), .Q(exu_spu_rs3_data_e[59]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[60](.D(exu_n29698), .CLK(rclk), .Q(exu_spu_rs3_data_e[60]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[61](.D(exu_n29697), .CLK(rclk), .Q(exu_spu_rs3_data_e[61]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[62](.D(exu_n29696), .CLK(rclk), .Q(exu_spu_rs3_data_e[62]));
DFFPOSX1 bypass_rs3_data_dff_q_reg[63](.D(exu_n29695), .CLK(rclk), .Q(exu_spu_rs3_data_e[63]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[0](.D(exu_n29670), .CLK(rclk), .Q(div_input_data_e[64]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[1](.D(exu_n29659), .CLK(rclk), .Q(div_input_data_e[65]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[2](.D(exu_n29648), .CLK(rclk), .Q(div_input_data_e[66]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[3](.D(exu_n29637), .CLK(rclk), .Q(div_input_data_e[67]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[4](.D(exu_n29629), .CLK(rclk), .Q(div_input_data_e[68]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[5](.D(exu_n29628), .CLK(rclk), .Q(div_input_data_e[69]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[6](.D(exu_n29627), .CLK(rclk), .Q(div_input_data_e[70]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[7](.D(exu_n29690), .CLK(rclk), .Q(div_input_data_e[71]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[8](.D(exu_n29689), .CLK(rclk), .Q(div_input_data_e[72]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[9](.D(exu_n29688), .CLK(rclk), .Q(div_input_data_e[73]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[10](.D(exu_n29687), .CLK(rclk), .Q(div_input_data_e[74]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[11](.D(exu_n29686), .CLK(rclk), .Q(div_input_data_e[75]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[12](.D(exu_n29685), .CLK(rclk), .Q(div_input_data_e[76]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[13](.D(exu_n29684), .CLK(rclk), .Q(div_input_data_e[77]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[14](.D(exu_n29683), .CLK(rclk), .Q(div_input_data_e[78]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[15](.D(exu_n29682), .CLK(rclk), .Q(div_input_data_e[79]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[16](.D(exu_n29681), .CLK(rclk), .Q(div_input_data_e[80]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[17](.D(exu_n29680), .CLK(rclk), .Q(div_input_data_e[81]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[18](.D(exu_n29679), .CLK(rclk), .Q(div_input_data_e[82]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[19](.D(exu_n29678), .CLK(rclk), .Q(div_input_data_e[83]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[20](.D(exu_n29677), .CLK(rclk), .Q(div_input_data_e[84]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[21](.D(exu_n29676), .CLK(rclk), .Q(div_input_data_e[85]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[22](.D(exu_n29675), .CLK(rclk), .Q(div_input_data_e[86]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[23](.D(exu_n29674), .CLK(rclk), .Q(div_input_data_e[87]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[24](.D(exu_n29673), .CLK(rclk), .Q(div_input_data_e[88]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[25](.D(exu_n29672), .CLK(rclk), .Q(div_input_data_e[89]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[26](.D(exu_n29671), .CLK(rclk), .Q(div_input_data_e[90]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[27](.D(exu_n29669), .CLK(rclk), .Q(div_input_data_e[91]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[28](.D(exu_n29668), .CLK(rclk), .Q(div_input_data_e[92]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[29](.D(exu_n29667), .CLK(rclk), .Q(div_input_data_e[93]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[30](.D(exu_n29666), .CLK(rclk), .Q(div_input_data_e[94]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[31](.D(exu_n29665), .CLK(rclk), .Q(div_input_data_e[95]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[32](.D(exu_n29664), .CLK(rclk), .Q(div_input_data_e[96]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[33](.D(exu_n29663), .CLK(rclk), .Q(div_input_data_e[97]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[34](.D(exu_n29662), .CLK(rclk), .Q(div_input_data_e[98]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[35](.D(exu_n29661), .CLK(rclk), .Q(div_input_data_e[99]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[36](.D(exu_n29660), .CLK(rclk), .Q(div_input_data_e[100]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[37](.D(exu_n29658), .CLK(rclk), .Q(div_input_data_e[101]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[38](.D(exu_n29657), .CLK(rclk), .Q(div_input_data_e[102]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[39](.D(exu_n29656), .CLK(rclk), .Q(div_input_data_e[103]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[40](.D(exu_n29655), .CLK(rclk), .Q(div_input_data_e[104]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[41](.D(exu_n29654), .CLK(rclk), .Q(div_input_data_e[105]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[42](.D(exu_n29653), .CLK(rclk), .Q(div_input_data_e[106]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[43](.D(exu_n29652), .CLK(rclk), .Q(div_input_data_e[107]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[44](.D(exu_n29651), .CLK(rclk), .Q(div_input_data_e[108]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[45](.D(exu_n29650), .CLK(rclk), .Q(div_input_data_e[109]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[46](.D(exu_n29649), .CLK(rclk), .Q(div_input_data_e[110]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[47](.D(exu_n29647), .CLK(rclk), .Q(div_input_data_e[111]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[48](.D(exu_n29646), .CLK(rclk), .Q(div_input_data_e[112]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[49](.D(exu_n29645), .CLK(rclk), .Q(div_input_data_e[113]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[50](.D(exu_n29644), .CLK(rclk), .Q(div_input_data_e[114]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[51](.D(exu_n29643), .CLK(rclk), .Q(div_input_data_e[115]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[52](.D(exu_n29642), .CLK(rclk), .Q(div_input_data_e[116]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[53](.D(exu_n29641), .CLK(rclk), .Q(div_input_data_e[117]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[54](.D(exu_n29640), .CLK(rclk), .Q(div_input_data_e[118]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[55](.D(exu_n29639), .CLK(rclk), .Q(div_input_data_e[119]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[56](.D(exu_n29638), .CLK(rclk), .Q(div_input_data_e[120]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[57](.D(exu_n29636), .CLK(rclk), .Q(div_input_data_e[121]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[58](.D(exu_n29635), .CLK(rclk), .Q(div_input_data_e[122]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[59](.D(exu_n29634), .CLK(rclk), .Q(div_input_data_e[123]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[60](.D(exu_n29633), .CLK(rclk), .Q(div_input_data_e[124]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[61](.D(exu_n29632), .CLK(rclk), .Q(div_input_data_e[125]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[62](.D(exu_n29631), .CLK(rclk), .Q(div_input_data_e[126]));
DFFPOSX1 bypass_rs2_data_dff_q_reg[63](.D(exu_n29630), .CLK(rclk), .Q(div_input_data_e[127]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[0](.D(exu_n29605), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[0]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[1](.D(exu_n29594), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[1]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[2](.D(exu_n29583), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[2]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[3](.D(exu_n29572), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[3]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[4](.D(exu_n29564), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[4]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[5](.D(exu_n29563), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[5]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[6](.D(exu_n29562), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[6]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[7](.D(exu_n29625), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[7]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[8](.D(exu_n29624), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[8]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[9](.D(exu_n29623), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[9]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[10](.D(exu_n29622), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[10]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[11](.D(exu_n29621), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[11]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[12](.D(exu_n29620), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[12]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[13](.D(exu_n29619), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[13]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[14](.D(exu_n29618), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[14]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[15](.D(exu_n29617), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[15]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[16](.D(exu_n29616), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[16]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[17](.D(exu_n29615), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[17]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[18](.D(exu_n29614), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[18]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[19](.D(exu_n29613), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[19]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[20](.D(exu_n29612), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[20]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[21](.D(exu_n29611), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[21]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[22](.D(exu_n29610), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[22]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[23](.D(exu_n29609), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[23]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[24](.D(exu_n29608), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[24]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[25](.D(exu_n29607), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[25]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[26](.D(exu_n29606), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[26]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[27](.D(exu_n29604), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[27]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[28](.D(exu_n29603), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[28]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[29](.D(exu_n29602), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[29]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[30](.D(exu_n29601), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[30]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[31](.D(exu_n29600), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[31]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[32](.D(exu_n29599), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[32]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[33](.D(exu_n29598), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[33]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[34](.D(exu_n29597), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[34]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[35](.D(exu_n29596), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[35]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[36](.D(exu_n29595), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[36]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[37](.D(exu_n29593), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[37]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[38](.D(exu_n29592), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[38]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[39](.D(exu_n29591), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[39]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[40](.D(exu_n29590), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[40]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[41](.D(exu_n29589), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[41]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[42](.D(exu_n29588), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[42]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[43](.D(exu_n29587), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[43]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[44](.D(exu_n29586), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[44]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[45](.D(exu_n29585), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[45]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[46](.D(exu_n29584), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[46]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[47](.D(exu_n29582), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[47]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[48](.D(exu_n29581), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[48]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[49](.D(exu_n29580), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[49]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[50](.D(exu_n29579), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[50]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[51](.D(exu_n29578), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[51]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[52](.D(exu_n29577), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[52]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[53](.D(exu_n29576), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[53]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[54](.D(exu_n29575), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[54]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[55](.D(exu_n29574), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[55]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[56](.D(exu_n29573), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[56]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[57](.D(exu_n29571), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[57]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[58](.D(exu_n29570), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[58]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[59](.D(exu_n29569), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[59]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[60](.D(exu_n29568), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[60]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[61](.D(exu_n29567), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[61]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[62](.D(exu_n29566), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[62]));
DFFPOSX1 bypass_rs1_data_dff_q_reg[63](.D(exu_n29565), .CLK(rclk), .Q(alu_logic_rs1_data_bf1[63]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[0](.D(exu_n29540), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[0]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[1](.D(exu_n29529), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[1]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[2](.D(exu_n29518), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[2]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[3](.D(exu_n29507), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[3]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[4](.D(exu_n29499), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[4]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[5](.D(exu_n29498), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[5]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[6](.D(exu_n29497), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[6]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[7](.D(exu_n29560), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[7]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[8](.D(exu_n29559), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[8]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[9](.D(exu_n29558), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[9]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[10](.D(exu_n29557), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[10]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[11](.D(exu_n29556), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[11]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[12](.D(exu_n29555), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[12]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[13](.D(exu_n29554), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[13]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[14](.D(exu_n29553), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[14]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[15](.D(exu_n29552), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[15]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[16](.D(exu_n29551), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[16]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[17](.D(exu_n29550), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[17]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[18](.D(exu_n29549), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[18]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[19](.D(exu_n29548), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[19]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[20](.D(exu_n29547), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[20]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[21](.D(exu_n29546), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[21]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[22](.D(exu_n29545), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[22]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[23](.D(exu_n29544), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[23]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[24](.D(exu_n29543), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[24]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[25](.D(exu_n29542), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[25]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[26](.D(exu_n29541), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[26]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[27](.D(exu_n29539), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[27]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[28](.D(exu_n29538), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[28]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[29](.D(exu_n29537), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[29]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[30](.D(exu_n29536), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[30]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[31](.D(exu_n29535), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[31]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[32](.D(exu_n29534), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[32]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[33](.D(exu_n29533), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[33]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[34](.D(exu_n29532), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[34]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[35](.D(exu_n29531), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[35]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[36](.D(exu_n29530), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[36]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[37](.D(exu_n29528), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[37]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[38](.D(exu_n29527), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[38]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[39](.D(exu_n29526), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[39]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[40](.D(exu_n29525), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[40]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[41](.D(exu_n29524), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[41]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[42](.D(exu_n29523), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[42]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[43](.D(exu_n29522), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[43]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[44](.D(exu_n29521), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[44]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[45](.D(exu_n29520), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[45]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[46](.D(exu_n29519), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[46]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[47](.D(exu_n29517), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[47]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[48](.D(exu_n29516), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[48]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[49](.D(exu_n29515), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[49]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[50](.D(exu_n29514), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[50]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[51](.D(exu_n29513), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[51]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[52](.D(exu_n29512), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[52]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[53](.D(exu_n29511), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[53]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[54](.D(exu_n29510), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[54]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[55](.D(exu_n29509), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[55]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[56](.D(exu_n29508), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[56]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[57](.D(exu_n29506), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[57]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[58](.D(exu_n29505), .CLK(bypass_sehold_clk), .Q(byp_irf_rd_data_w2[58]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[59](.D(exu_n29504), .CLK(exu_n16184), .Q(byp_irf_rd_data_w2[59]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[60](.D(exu_n29503), .CLK(exu_n16184), .Q(byp_irf_rd_data_w2[60]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[61](.D(exu_n29502), .CLK(exu_n16184), .Q(byp_irf_rd_data_w2[61]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[62](.D(exu_n29501), .CLK(exu_n16184), .Q(byp_irf_rd_data_w2[62]));
DFFPOSX1 bypass_dff_rd_data_g2w_q_reg[63](.D(exu_n29500), .CLK(exu_n16184), .Q(byp_irf_rd_data_w2[63]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[0](.D(exu_n29475), .CLK(exu_n16184), .Q(byp_irf_rd_data_w[0]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[1](.D(exu_n29464), .CLK(exu_n16184), .Q(byp_irf_rd_data_w[1]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[2](.D(exu_n29453), .CLK(exu_n16184), .Q(byp_irf_rd_data_w[2]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[3](.D(exu_n29442), .CLK(exu_n16184), .Q(byp_irf_rd_data_w[3]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[4](.D(exu_n29434), .CLK(exu_n16184), .Q(byp_irf_rd_data_w[4]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[5](.D(exu_n29433), .CLK(exu_n16184), .Q(byp_irf_rd_data_w[5]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[6](.D(exu_n29432), .CLK(exu_n16184), .Q(byp_irf_rd_data_w[6]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[7](.D(exu_n29495), .CLK(exu_n16184), .Q(byp_irf_rd_data_w[7]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[8](.D(exu_n29494), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[8]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[9](.D(exu_n29493), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[9]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[10](.D(exu_n29492), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[10]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[11](.D(exu_n29491), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[11]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[12](.D(exu_n29490), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[12]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[13](.D(exu_n29489), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[13]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[14](.D(exu_n29488), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[14]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[15](.D(exu_n29487), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[15]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[16](.D(exu_n29486), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[16]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[17](.D(exu_n29485), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[17]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[18](.D(exu_n29484), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[18]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[19](.D(exu_n29483), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[19]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[20](.D(exu_n29482), .CLK(exu_n16183), .Q(byp_irf_rd_data_w[20]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[21](.D(exu_n29481), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[21]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[22](.D(exu_n29480), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[22]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[23](.D(exu_n29479), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[23]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[24](.D(exu_n29478), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[24]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[25](.D(exu_n29477), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[25]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[26](.D(exu_n29476), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[26]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[27](.D(exu_n29474), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[27]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[28](.D(exu_n29473), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[28]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[29](.D(exu_n29472), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[29]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[30](.D(exu_n29471), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[30]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[31](.D(exu_n29470), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[31]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[32](.D(exu_n29469), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[32]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[33](.D(exu_n29468), .CLK(exu_n16182), .Q(byp_irf_rd_data_w[33]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[34](.D(exu_n29467), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[34]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[35](.D(exu_n29466), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[35]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[36](.D(exu_n29465), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[36]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[37](.D(exu_n29463), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[37]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[38](.D(exu_n29462), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[38]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[39](.D(exu_n29461), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[39]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[40](.D(exu_n29460), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[40]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[41](.D(exu_n29459), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[41]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[42](.D(exu_n29458), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[42]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[43](.D(exu_n29457), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[43]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[44](.D(exu_n29456), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[44]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[45](.D(exu_n29455), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[45]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[46](.D(exu_n29454), .CLK(exu_n16181), .Q(byp_irf_rd_data_w[46]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[47](.D(exu_n29452), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[47]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[48](.D(exu_n29451), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[48]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[49](.D(exu_n29450), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[49]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[50](.D(exu_n29449), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[50]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[51](.D(exu_n29448), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[51]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[52](.D(exu_n29447), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[52]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[53](.D(exu_n29446), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[53]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[54](.D(exu_n29445), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[54]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[55](.D(exu_n29444), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[55]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[56](.D(exu_n29443), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[56]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[57](.D(exu_n29441), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[57]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[58](.D(exu_n29440), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[58]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[59](.D(exu_n29439), .CLK(exu_n16180), .Q(byp_irf_rd_data_w[59]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[60](.D(exu_n29438), .CLK(exu_n16179), .Q(byp_irf_rd_data_w[60]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[61](.D(exu_n29437), .CLK(exu_n16179), .Q(byp_irf_rd_data_w[61]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[62](.D(exu_n29436), .CLK(exu_n16179), .Q(byp_irf_rd_data_w[62]));
DFFPOSX1 bypass_dff_rd_data_m2w_q_reg[63](.D(exu_n29435), .CLK(exu_n16179), .Q(byp_irf_rd_data_w[63]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[0](.D(exu_n29410), .CLK(rclk), .Q(bypass_restore_rd_data[0]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[1](.D(exu_n29399), .CLK(rclk), .Q(bypass_restore_rd_data[1]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[2](.D(exu_n29388), .CLK(rclk), .Q(bypass_restore_rd_data[2]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[3](.D(exu_n29377), .CLK(rclk), .Q(bypass_restore_rd_data[3]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[4](.D(exu_n29369), .CLK(rclk), .Q(bypass_restore_rd_data[4]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[5](.D(exu_n29368), .CLK(rclk), .Q(bypass_restore_rd_data[5]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[6](.D(exu_n29367), .CLK(rclk), .Q(bypass_restore_rd_data[6]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[7](.D(exu_n29430), .CLK(rclk), .Q(bypass_restore_rd_data[7]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[8](.D(exu_n29429), .CLK(rclk), .Q(bypass_restore_rd_data[8]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[9](.D(exu_n29428), .CLK(rclk), .Q(bypass_restore_rd_data[9]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[10](.D(exu_n29427), .CLK(rclk), .Q(bypass_restore_rd_data[10]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[11](.D(exu_n29426), .CLK(rclk), .Q(bypass_restore_rd_data[11]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[12](.D(exu_n29425), .CLK(rclk), .Q(bypass_restore_rd_data[12]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[13](.D(exu_n29424), .CLK(rclk), .Q(bypass_restore_rd_data[13]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[14](.D(exu_n29423), .CLK(rclk), .Q(bypass_restore_rd_data[14]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[15](.D(exu_n29422), .CLK(rclk), .Q(bypass_restore_rd_data[15]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[16](.D(exu_n29421), .CLK(rclk), .Q(bypass_restore_rd_data[16]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[17](.D(exu_n29420), .CLK(rclk), .Q(bypass_restore_rd_data[17]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[18](.D(exu_n29419), .CLK(rclk), .Q(bypass_restore_rd_data[18]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[19](.D(exu_n29418), .CLK(rclk), .Q(bypass_restore_rd_data[19]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[20](.D(exu_n29417), .CLK(rclk), .Q(bypass_restore_rd_data[20]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[21](.D(exu_n29416), .CLK(rclk), .Q(bypass_restore_rd_data[21]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[22](.D(exu_n29415), .CLK(rclk), .Q(bypass_restore_rd_data[22]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[23](.D(exu_n29414), .CLK(rclk), .Q(bypass_restore_rd_data[23]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[24](.D(exu_n29413), .CLK(rclk), .Q(bypass_restore_rd_data[24]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[25](.D(exu_n29412), .CLK(rclk), .Q(bypass_restore_rd_data[25]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[26](.D(exu_n29411), .CLK(rclk), .Q(bypass_restore_rd_data[26]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[27](.D(exu_n29409), .CLK(rclk), .Q(bypass_restore_rd_data[27]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[28](.D(exu_n29408), .CLK(rclk), .Q(bypass_restore_rd_data[28]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[29](.D(exu_n29407), .CLK(rclk), .Q(bypass_restore_rd_data[29]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[30](.D(exu_n29406), .CLK(rclk), .Q(bypass_restore_rd_data[30]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[31](.D(exu_n29405), .CLK(rclk), .Q(bypass_restore_rd_data[31]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[32](.D(exu_n29404), .CLK(rclk), .Q(bypass_restore_rd_data[32]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[33](.D(exu_n29403), .CLK(rclk), .Q(bypass_restore_rd_data[33]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[34](.D(exu_n29402), .CLK(rclk), .Q(bypass_restore_rd_data[34]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[35](.D(exu_n29401), .CLK(rclk), .Q(bypass_restore_rd_data[35]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[36](.D(exu_n29400), .CLK(rclk), .Q(bypass_restore_rd_data[36]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[37](.D(exu_n29398), .CLK(rclk), .Q(bypass_restore_rd_data[37]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[38](.D(exu_n29397), .CLK(rclk), .Q(bypass_restore_rd_data[38]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[39](.D(exu_n29396), .CLK(rclk), .Q(bypass_restore_rd_data[39]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[40](.D(exu_n29395), .CLK(rclk), .Q(bypass_restore_rd_data[40]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[41](.D(exu_n29394), .CLK(rclk), .Q(bypass_restore_rd_data[41]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[42](.D(exu_n29393), .CLK(rclk), .Q(bypass_restore_rd_data[42]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[43](.D(exu_n29392), .CLK(rclk), .Q(bypass_restore_rd_data[43]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[44](.D(exu_n29391), .CLK(rclk), .Q(bypass_restore_rd_data[44]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[45](.D(exu_n29390), .CLK(rclk), .Q(bypass_restore_rd_data[45]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[46](.D(exu_n29389), .CLK(rclk), .Q(bypass_restore_rd_data[46]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[47](.D(exu_n29387), .CLK(rclk), .Q(bypass_restore_rd_data[47]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[48](.D(exu_n29386), .CLK(rclk), .Q(bypass_restore_rd_data[48]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[49](.D(exu_n29385), .CLK(rclk), .Q(bypass_restore_rd_data[49]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[50](.D(exu_n29384), .CLK(rclk), .Q(bypass_restore_rd_data[50]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[51](.D(exu_n29383), .CLK(rclk), .Q(bypass_restore_rd_data[51]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[52](.D(exu_n29382), .CLK(rclk), .Q(bypass_restore_rd_data[52]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[53](.D(exu_n29381), .CLK(rclk), .Q(bypass_restore_rd_data[53]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[54](.D(exu_n29380), .CLK(rclk), .Q(bypass_restore_rd_data[54]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[55](.D(exu_n29379), .CLK(rclk), .Q(bypass_restore_rd_data[55]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[56](.D(exu_n29378), .CLK(rclk), .Q(bypass_restore_rd_data[56]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[57](.D(exu_n29376), .CLK(rclk), .Q(bypass_restore_rd_data[57]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[58](.D(exu_n29375), .CLK(rclk), .Q(bypass_restore_rd_data[58]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[59](.D(exu_n29374), .CLK(rclk), .Q(bypass_restore_rd_data[59]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[60](.D(exu_n29373), .CLK(rclk), .Q(bypass_restore_rd_data[60]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[61](.D(exu_n29372), .CLK(rclk), .Q(bypass_restore_rd_data[61]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[62](.D(exu_n29371), .CLK(rclk), .Q(bypass_restore_rd_data[62]));
DFFPOSX1 bypass_dff_restore_buf_q_reg[63](.D(exu_n29370), .CLK(rclk), .Q(bypass_restore_rd_data[63]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[0](.D(exu_n29345), .CLK(rclk), .Q(exu_tlu_wsr_data_m[0]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[1](.D(exu_n29334), .CLK(rclk), .Q(exu_tlu_wsr_data_m[1]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[2](.D(exu_n29323), .CLK(rclk), .Q(exu_tlu_wsr_data_m[2]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[3](.D(exu_n29312), .CLK(rclk), .Q(exu_tlu_wsr_data_m[3]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[4](.D(exu_n29304), .CLK(rclk), .Q(exu_tlu_wsr_data_m[4]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[5](.D(exu_n29303), .CLK(rclk), .Q(exu_tlu_wsr_data_m[5]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[6](.D(exu_n29302), .CLK(rclk), .Q(exu_tlu_wsr_data_m[6]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[7](.D(exu_n29365), .CLK(rclk), .Q(exu_tlu_wsr_data_m[7]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[8](.D(exu_n29364), .CLK(rclk), .Q(exu_tlu_wsr_data_m[8]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[9](.D(exu_n29363), .CLK(rclk), .Q(exu_tlu_wsr_data_m[9]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[10](.D(exu_n29362), .CLK(rclk), .Q(exu_tlu_wsr_data_m[10]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[11](.D(exu_n29361), .CLK(rclk), .Q(exu_tlu_wsr_data_m[11]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[12](.D(exu_n29360), .CLK(rclk), .Q(exu_tlu_wsr_data_m[12]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[13](.D(exu_n29359), .CLK(rclk), .Q(exu_tlu_wsr_data_m[13]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[14](.D(exu_n29358), .CLK(rclk), .Q(exu_tlu_wsr_data_m[14]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[15](.D(exu_n29357), .CLK(rclk), .Q(exu_tlu_wsr_data_m[15]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[16](.D(exu_n29356), .CLK(rclk), .Q(exu_tlu_wsr_data_m[16]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[17](.D(exu_n29355), .CLK(rclk), .Q(exu_tlu_wsr_data_m[17]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[18](.D(exu_n29354), .CLK(rclk), .Q(exu_tlu_wsr_data_m[18]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[19](.D(exu_n29353), .CLK(rclk), .Q(exu_tlu_wsr_data_m[19]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[20](.D(exu_n29352), .CLK(rclk), .Q(exu_tlu_wsr_data_m[20]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[21](.D(exu_n29351), .CLK(rclk), .Q(exu_tlu_wsr_data_m[21]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[22](.D(exu_n29350), .CLK(rclk), .Q(exu_tlu_wsr_data_m[22]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[23](.D(exu_n29349), .CLK(rclk), .Q(exu_tlu_wsr_data_m[23]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[24](.D(exu_n29348), .CLK(rclk), .Q(exu_tlu_wsr_data_m[24]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[25](.D(exu_n29347), .CLK(rclk), .Q(exu_tlu_wsr_data_m[25]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[26](.D(exu_n29346), .CLK(rclk), .Q(exu_tlu_wsr_data_m[26]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[27](.D(exu_n29344), .CLK(rclk), .Q(exu_tlu_wsr_data_m[27]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[28](.D(exu_n29343), .CLK(rclk), .Q(exu_tlu_wsr_data_m[28]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[29](.D(exu_n29342), .CLK(rclk), .Q(exu_tlu_wsr_data_m[29]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[30](.D(exu_n29341), .CLK(rclk), .Q(exu_tlu_wsr_data_m[30]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[31](.D(exu_n29340), .CLK(rclk), .Q(exu_tlu_wsr_data_m[31]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[32](.D(exu_n29339), .CLK(rclk), .Q(exu_tlu_wsr_data_m[32]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[33](.D(exu_n29338), .CLK(rclk), .Q(exu_tlu_wsr_data_m[33]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[34](.D(exu_n29337), .CLK(rclk), .Q(exu_tlu_wsr_data_m[34]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[35](.D(exu_n29336), .CLK(rclk), .Q(exu_tlu_wsr_data_m[35]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[36](.D(exu_n29335), .CLK(rclk), .Q(exu_tlu_wsr_data_m[36]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[37](.D(exu_n29333), .CLK(rclk), .Q(exu_tlu_wsr_data_m[37]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[38](.D(exu_n29332), .CLK(rclk), .Q(exu_tlu_wsr_data_m[38]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[39](.D(exu_n29331), .CLK(rclk), .Q(exu_tlu_wsr_data_m[39]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[40](.D(exu_n29330), .CLK(rclk), .Q(exu_tlu_wsr_data_m[40]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[41](.D(exu_n29329), .CLK(rclk), .Q(exu_tlu_wsr_data_m[41]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[42](.D(exu_n29328), .CLK(rclk), .Q(exu_tlu_wsr_data_m[42]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[43](.D(exu_n29327), .CLK(rclk), .Q(exu_tlu_wsr_data_m[43]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[44](.D(exu_n29326), .CLK(rclk), .Q(exu_tlu_wsr_data_m[44]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[45](.D(exu_n29325), .CLK(rclk), .Q(exu_tlu_wsr_data_m[45]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[46](.D(exu_n29324), .CLK(rclk), .Q(exu_tlu_wsr_data_m[46]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[47](.D(exu_n29322), .CLK(rclk), .Q(exu_tlu_wsr_data_m[47]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[48](.D(exu_n29321), .CLK(rclk), .Q(exu_tlu_wsr_data_m[48]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[49](.D(exu_n29320), .CLK(rclk), .Q(exu_tlu_wsr_data_m[49]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[50](.D(exu_n29319), .CLK(rclk), .Q(exu_tlu_wsr_data_m[50]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[51](.D(exu_n29318), .CLK(rclk), .Q(exu_tlu_wsr_data_m[51]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[52](.D(exu_n29317), .CLK(rclk), .Q(exu_tlu_wsr_data_m[52]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[53](.D(exu_n29316), .CLK(rclk), .Q(exu_tlu_wsr_data_m[53]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[54](.D(exu_n29315), .CLK(rclk), .Q(exu_tlu_wsr_data_m[54]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[55](.D(exu_n29314), .CLK(rclk), .Q(exu_tlu_wsr_data_m[55]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[56](.D(exu_n29313), .CLK(rclk), .Q(exu_tlu_wsr_data_m[56]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[57](.D(exu_n29311), .CLK(rclk), .Q(exu_tlu_wsr_data_m[57]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[58](.D(exu_n29310), .CLK(rclk), .Q(exu_tlu_wsr_data_m[58]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[59](.D(exu_n29309), .CLK(rclk), .Q(exu_tlu_wsr_data_m[59]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[60](.D(exu_n29308), .CLK(rclk), .Q(exu_tlu_wsr_data_m[60]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[61](.D(exu_n29307), .CLK(rclk), .Q(exu_tlu_wsr_data_m[61]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[62](.D(exu_n29306), .CLK(rclk), .Q(exu_tlu_wsr_data_m[62]));
DFFPOSX1 bypass_dff_rd_data_e2m_q_reg[63](.D(exu_n29305), .CLK(rclk), .Q(exu_tlu_wsr_data_m[63]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[0](.D(exu_n21772), .CLK(rclk), .Q(div_yreg_div_ecl_yreg_0[3]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[1](.D(exu_n21766), .CLK(rclk), .Q(div_yreg_yreg_thr3[1]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[2](.D(exu_n21765), .CLK(rclk), .Q(div_yreg_yreg_thr3[2]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[3](.D(exu_n21764), .CLK(rclk), .Q(div_yreg_yreg_thr3[3]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[4](.D(exu_n21763), .CLK(rclk), .Q(div_yreg_yreg_thr3[4]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[5](.D(exu_n21762), .CLK(rclk), .Q(div_yreg_yreg_thr3[5]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[6](.D(exu_n21761), .CLK(rclk), .Q(div_yreg_yreg_thr3[6]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[7](.D(exu_n21792), .CLK(rclk), .Q(div_yreg_yreg_thr3[7]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[8](.D(exu_n21791), .CLK(rclk), .Q(div_yreg_yreg_thr3[8]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[9](.D(exu_n21790), .CLK(rclk), .Q(div_yreg_yreg_thr3[9]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[10](.D(exu_n21789), .CLK(rclk), .Q(div_yreg_yreg_thr3[10]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[11](.D(exu_n21788), .CLK(rclk), .Q(div_yreg_yreg_thr3[11]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[12](.D(exu_n21787), .CLK(rclk), .Q(div_yreg_yreg_thr3[12]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[13](.D(exu_n21786), .CLK(rclk), .Q(div_yreg_yreg_thr3[13]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[14](.D(exu_n21785), .CLK(rclk), .Q(div_yreg_yreg_thr3[14]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[15](.D(exu_n21784), .CLK(rclk), .Q(div_yreg_yreg_thr3[15]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[16](.D(exu_n21783), .CLK(rclk), .Q(div_yreg_yreg_thr3[16]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[17](.D(exu_n21782), .CLK(rclk), .Q(div_yreg_yreg_thr3[17]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[18](.D(exu_n21781), .CLK(rclk), .Q(div_yreg_yreg_thr3[18]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[19](.D(exu_n21780), .CLK(rclk), .Q(div_yreg_yreg_thr3[19]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[20](.D(exu_n21779), .CLK(rclk), .Q(div_yreg_yreg_thr3[20]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[21](.D(exu_n21778), .CLK(rclk), .Q(div_yreg_yreg_thr3[21]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[22](.D(exu_n21777), .CLK(rclk), .Q(div_yreg_yreg_thr3[22]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[23](.D(exu_n21776), .CLK(rclk), .Q(div_yreg_yreg_thr3[23]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[24](.D(exu_n21775), .CLK(rclk), .Q(div_yreg_yreg_thr3[24]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[25](.D(exu_n21774), .CLK(rclk), .Q(div_yreg_yreg_thr3[25]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[26](.D(exu_n21773), .CLK(rclk), .Q(div_yreg_yreg_thr3[26]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[27](.D(exu_n21771), .CLK(rclk), .Q(div_yreg_yreg_thr3[27]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[28](.D(exu_n21770), .CLK(rclk), .Q(div_yreg_yreg_thr3[28]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[29](.D(exu_n21769), .CLK(rclk), .Q(div_yreg_yreg_thr3[29]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[30](.D(exu_n21768), .CLK(rclk), .Q(div_yreg_yreg_thr3[30]));
DFFPOSX1 div_yreg_dff_yreg_thr3_q_reg[31](.D(exu_n21767), .CLK(rclk), .Q(div_yreg_yreg_thr3[31]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[0](.D(exu_n21739), .CLK(rclk), .Q(div_yreg_div_ecl_yreg_0[2]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[1](.D(exu_n21733), .CLK(rclk), .Q(div_yreg_yreg_thr2[1]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[2](.D(exu_n21732), .CLK(rclk), .Q(div_yreg_yreg_thr2[2]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[3](.D(exu_n21731), .CLK(rclk), .Q(div_yreg_yreg_thr2[3]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[4](.D(exu_n21730), .CLK(rclk), .Q(div_yreg_yreg_thr2[4]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[5](.D(exu_n21729), .CLK(rclk), .Q(div_yreg_yreg_thr2[5]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[6](.D(exu_n21728), .CLK(rclk), .Q(div_yreg_yreg_thr2[6]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[7](.D(exu_n21759), .CLK(rclk), .Q(div_yreg_yreg_thr2[7]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[8](.D(exu_n21758), .CLK(rclk), .Q(div_yreg_yreg_thr2[8]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[9](.D(exu_n21757), .CLK(rclk), .Q(div_yreg_yreg_thr2[9]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[10](.D(exu_n21756), .CLK(rclk), .Q(div_yreg_yreg_thr2[10]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[11](.D(exu_n21755), .CLK(rclk), .Q(div_yreg_yreg_thr2[11]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[12](.D(exu_n21754), .CLK(rclk), .Q(div_yreg_yreg_thr2[12]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[13](.D(exu_n21753), .CLK(rclk), .Q(div_yreg_yreg_thr2[13]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[14](.D(exu_n21752), .CLK(rclk), .Q(div_yreg_yreg_thr2[14]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[15](.D(exu_n21751), .CLK(rclk), .Q(div_yreg_yreg_thr2[15]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[16](.D(exu_n21750), .CLK(rclk), .Q(div_yreg_yreg_thr2[16]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[17](.D(exu_n21749), .CLK(rclk), .Q(div_yreg_yreg_thr2[17]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[18](.D(exu_n21748), .CLK(rclk), .Q(div_yreg_yreg_thr2[18]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[19](.D(exu_n21747), .CLK(rclk), .Q(div_yreg_yreg_thr2[19]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[20](.D(exu_n21746), .CLK(rclk), .Q(div_yreg_yreg_thr2[20]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[21](.D(exu_n21745), .CLK(rclk), .Q(div_yreg_yreg_thr2[21]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[22](.D(exu_n21744), .CLK(rclk), .Q(div_yreg_yreg_thr2[22]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[23](.D(exu_n21743), .CLK(rclk), .Q(div_yreg_yreg_thr2[23]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[24](.D(exu_n21742), .CLK(rclk), .Q(div_yreg_yreg_thr2[24]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[25](.D(exu_n21741), .CLK(rclk), .Q(div_yreg_yreg_thr2[25]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[26](.D(exu_n21740), .CLK(rclk), .Q(div_yreg_yreg_thr2[26]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[27](.D(exu_n21738), .CLK(rclk), .Q(div_yreg_yreg_thr2[27]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[28](.D(exu_n21737), .CLK(rclk), .Q(div_yreg_yreg_thr2[28]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[29](.D(exu_n21736), .CLK(rclk), .Q(div_yreg_yreg_thr2[29]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[30](.D(exu_n21735), .CLK(rclk), .Q(div_yreg_yreg_thr2[30]));
DFFPOSX1 div_yreg_dff_yreg_thr2_q_reg[31](.D(exu_n21734), .CLK(rclk), .Q(div_yreg_yreg_thr2[31]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[0](.D(exu_n21706), .CLK(rclk), .Q(div_yreg_div_ecl_yreg_0[1]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[1](.D(exu_n21700), .CLK(rclk), .Q(div_yreg_yreg_thr1[1]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[2](.D(exu_n21699), .CLK(rclk), .Q(div_yreg_yreg_thr1[2]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[3](.D(exu_n21698), .CLK(rclk), .Q(div_yreg_yreg_thr1[3]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[4](.D(exu_n21697), .CLK(rclk), .Q(div_yreg_yreg_thr1[4]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[5](.D(exu_n21696), .CLK(rclk), .Q(div_yreg_yreg_thr1[5]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[6](.D(exu_n21695), .CLK(rclk), .Q(div_yreg_yreg_thr1[6]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[7](.D(exu_n21726), .CLK(rclk), .Q(div_yreg_yreg_thr1[7]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[8](.D(exu_n21725), .CLK(rclk), .Q(div_yreg_yreg_thr1[8]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[9](.D(exu_n21724), .CLK(rclk), .Q(div_yreg_yreg_thr1[9]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[10](.D(exu_n21723), .CLK(rclk), .Q(div_yreg_yreg_thr1[10]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[11](.D(exu_n21722), .CLK(rclk), .Q(div_yreg_yreg_thr1[11]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[12](.D(exu_n21721), .CLK(rclk), .Q(div_yreg_yreg_thr1[12]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[13](.D(exu_n21720), .CLK(rclk), .Q(div_yreg_yreg_thr1[13]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[14](.D(exu_n21719), .CLK(rclk), .Q(div_yreg_yreg_thr1[14]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[15](.D(exu_n21718), .CLK(rclk), .Q(div_yreg_yreg_thr1[15]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[16](.D(exu_n21717), .CLK(rclk), .Q(div_yreg_yreg_thr1[16]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[17](.D(exu_n21716), .CLK(rclk), .Q(div_yreg_yreg_thr1[17]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[18](.D(exu_n21715), .CLK(rclk), .Q(div_yreg_yreg_thr1[18]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[19](.D(exu_n21714), .CLK(rclk), .Q(div_yreg_yreg_thr1[19]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[20](.D(exu_n21713), .CLK(rclk), .Q(div_yreg_yreg_thr1[20]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[21](.D(exu_n21712), .CLK(rclk), .Q(div_yreg_yreg_thr1[21]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[22](.D(exu_n21711), .CLK(rclk), .Q(div_yreg_yreg_thr1[22]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[23](.D(exu_n21710), .CLK(rclk), .Q(div_yreg_yreg_thr1[23]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[24](.D(exu_n21709), .CLK(rclk), .Q(div_yreg_yreg_thr1[24]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[25](.D(exu_n21708), .CLK(rclk), .Q(div_yreg_yreg_thr1[25]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[26](.D(exu_n21707), .CLK(rclk), .Q(div_yreg_yreg_thr1[26]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[27](.D(exu_n21705), .CLK(rclk), .Q(div_yreg_yreg_thr1[27]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[28](.D(exu_n21704), .CLK(rclk), .Q(div_yreg_yreg_thr1[28]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[29](.D(exu_n21703), .CLK(rclk), .Q(div_yreg_yreg_thr1[29]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[30](.D(exu_n21702), .CLK(rclk), .Q(div_yreg_yreg_thr1[30]));
DFFPOSX1 div_yreg_dff_yreg_thr1_q_reg[31](.D(exu_n21701), .CLK(rclk), .Q(div_yreg_yreg_thr1[31]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[0](.D(exu_n21673), .CLK(rclk), .Q(div_yreg_div_ecl_yreg_0[0]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[1](.D(exu_n21667), .CLK(rclk), .Q(div_yreg_yreg_thr0[1]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[2](.D(exu_n21666), .CLK(rclk), .Q(div_yreg_yreg_thr0[2]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[3](.D(exu_n21665), .CLK(rclk), .Q(div_yreg_yreg_thr0[3]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[4](.D(exu_n21664), .CLK(rclk), .Q(div_yreg_yreg_thr0[4]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[5](.D(exu_n21663), .CLK(rclk), .Q(div_yreg_yreg_thr0[5]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[6](.D(exu_n21662), .CLK(rclk), .Q(div_yreg_yreg_thr0[6]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[7](.D(exu_n21693), .CLK(rclk), .Q(div_yreg_yreg_thr0[7]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[8](.D(exu_n21692), .CLK(rclk), .Q(div_yreg_yreg_thr0[8]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[9](.D(exu_n21691), .CLK(rclk), .Q(div_yreg_yreg_thr0[9]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[10](.D(exu_n21690), .CLK(rclk), .Q(div_yreg_yreg_thr0[10]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[11](.D(exu_n21689), .CLK(rclk), .Q(div_yreg_yreg_thr0[11]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[12](.D(exu_n21688), .CLK(rclk), .Q(div_yreg_yreg_thr0[12]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[13](.D(exu_n21687), .CLK(rclk), .Q(div_yreg_yreg_thr0[13]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[14](.D(exu_n21686), .CLK(rclk), .Q(div_yreg_yreg_thr0[14]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[15](.D(exu_n21685), .CLK(rclk), .Q(div_yreg_yreg_thr0[15]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[16](.D(exu_n21684), .CLK(rclk), .Q(div_yreg_yreg_thr0[16]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[17](.D(exu_n21683), .CLK(rclk), .Q(div_yreg_yreg_thr0[17]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[18](.D(exu_n21682), .CLK(rclk), .Q(div_yreg_yreg_thr0[18]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[19](.D(exu_n21681), .CLK(rclk), .Q(div_yreg_yreg_thr0[19]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[20](.D(exu_n21680), .CLK(rclk), .Q(div_yreg_yreg_thr0[20]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[21](.D(exu_n21679), .CLK(rclk), .Q(div_yreg_yreg_thr0[21]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[22](.D(exu_n21678), .CLK(rclk), .Q(div_yreg_yreg_thr0[22]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[23](.D(exu_n21677), .CLK(rclk), .Q(div_yreg_yreg_thr0[23]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[24](.D(exu_n21676), .CLK(rclk), .Q(div_yreg_yreg_thr0[24]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[25](.D(exu_n21675), .CLK(rclk), .Q(div_yreg_yreg_thr0[25]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[26](.D(exu_n21674), .CLK(rclk), .Q(div_yreg_yreg_thr0[26]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[27](.D(exu_n21672), .CLK(rclk), .Q(div_yreg_yreg_thr0[27]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[28](.D(exu_n21671), .CLK(rclk), .Q(div_yreg_yreg_thr0[28]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[29](.D(exu_n21670), .CLK(rclk), .Q(div_yreg_yreg_thr0[29]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[30](.D(exu_n21669), .CLK(rclk), .Q(div_yreg_yreg_thr0[30]));
DFFPOSX1 div_yreg_dff_yreg_thr0_q_reg[31](.D(exu_n21668), .CLK(rclk), .Q(div_yreg_yreg_thr0[31]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[0](.D(exu_n21640), .CLK(rclk), .Q(div_yreg_yreg_data_w1[0]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[1](.D(exu_n21634), .CLK(rclk), .Q(div_yreg_yreg_data_w1[1]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[2](.D(exu_n21633), .CLK(rclk), .Q(div_yreg_yreg_data_w1[2]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[3](.D(exu_n21632), .CLK(rclk), .Q(div_yreg_yreg_data_w1[3]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[4](.D(exu_n21631), .CLK(rclk), .Q(div_yreg_yreg_data_w1[4]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[5](.D(exu_n21630), .CLK(rclk), .Q(div_yreg_yreg_data_w1[5]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[6](.D(exu_n21629), .CLK(rclk), .Q(div_yreg_yreg_data_w1[6]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[7](.D(exu_n21660), .CLK(rclk), .Q(div_yreg_yreg_data_w1[7]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[8](.D(exu_n21659), .CLK(rclk), .Q(div_yreg_yreg_data_w1[8]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[9](.D(exu_n21658), .CLK(rclk), .Q(div_yreg_yreg_data_w1[9]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[10](.D(exu_n21657), .CLK(rclk), .Q(div_yreg_yreg_data_w1[10]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[11](.D(exu_n21656), .CLK(rclk), .Q(div_yreg_yreg_data_w1[11]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[12](.D(exu_n21655), .CLK(rclk), .Q(div_yreg_yreg_data_w1[12]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[13](.D(exu_n21654), .CLK(rclk), .Q(div_yreg_yreg_data_w1[13]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[14](.D(exu_n21653), .CLK(rclk), .Q(div_yreg_yreg_data_w1[14]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[15](.D(exu_n21652), .CLK(rclk), .Q(div_yreg_yreg_data_w1[15]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[16](.D(exu_n21651), .CLK(rclk), .Q(div_yreg_yreg_data_w1[16]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[17](.D(exu_n21650), .CLK(rclk), .Q(div_yreg_yreg_data_w1[17]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[18](.D(exu_n21649), .CLK(rclk), .Q(div_yreg_yreg_data_w1[18]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[19](.D(exu_n21648), .CLK(rclk), .Q(div_yreg_yreg_data_w1[19]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[20](.D(exu_n21647), .CLK(rclk), .Q(div_yreg_yreg_data_w1[20]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[21](.D(exu_n21646), .CLK(rclk), .Q(div_yreg_yreg_data_w1[21]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[22](.D(exu_n21645), .CLK(rclk), .Q(div_yreg_yreg_data_w1[22]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[23](.D(exu_n21644), .CLK(rclk), .Q(div_yreg_yreg_data_w1[23]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[24](.D(exu_n21643), .CLK(rclk), .Q(div_yreg_yreg_data_w1[24]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[25](.D(exu_n21642), .CLK(rclk), .Q(div_yreg_yreg_data_w1[25]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[26](.D(exu_n21641), .CLK(rclk), .Q(div_yreg_yreg_data_w1[26]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[27](.D(exu_n21639), .CLK(rclk), .Q(div_yreg_yreg_data_w1[27]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[28](.D(exu_n21638), .CLK(rclk), .Q(div_yreg_yreg_data_w1[28]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[29](.D(exu_n21637), .CLK(rclk), .Q(div_yreg_yreg_data_w1[29]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[30](.D(exu_n21636), .CLK(rclk), .Q(div_yreg_yreg_data_w1[30]));
DFFPOSX1 div_yreg_yreg_dff_w2w2_q_reg[31](.D(exu_n21635), .CLK(rclk), .Q(div_yreg_yreg_data_w1[31]));
XOR2X1 exu_bypass_w2_eccgen_U183(.A(exu_n20350), .B(exu_n20349), .Y(bypass_rd_synd_w2_l[0]));
XOR2X1 exu_bypass_w2_eccgen_U182(.A(exu_n20352), .B(exu_n20351), .Y(exu_n20349));
XOR2X1 exu_bypass_w2_eccgen_U181(.A(exu_n20354), .B(exu_n20353), .Y(exu_n20350));
XOR2X1 exu_bypass_w2_eccgen_U180(.A(bypass_w2_eccgen_p0_w[1]), .B(bypass_w2_eccgen_p0_w[0]), .Y(exu_n20351));
XOR2X1 exu_bypass_w2_eccgen_U179(.A(bypass_w2_eccgen_p0_w[3]), .B(bypass_w2_eccgen_p0_w[2]), .Y(exu_n20352));
XOR2X1 exu_bypass_w2_eccgen_U178(.A(bypass_w2_eccgen_p0_w[5]), .B(bypass_w2_eccgen_p0_w[4]), .Y(exu_n20353));
XOR2X1 exu_bypass_w2_eccgen_U177(.A(bypass_w2_eccgen_p0_w[7]), .B(bypass_w2_eccgen_p0_w[6]), .Y(exu_n20354));
XOR2X1 exu_bypass_w2_eccgen_U176(.A(exu_n20356), .B(exu_n20355), .Y(bypass_rd_synd_w2_l[1]));
XOR2X1 exu_bypass_w2_eccgen_U175(.A(exu_n20358), .B(exu_n20357), .Y(exu_n20355));
XOR2X1 exu_bypass_w2_eccgen_U174(.A(exu_n20360), .B(exu_n20359), .Y(exu_n20356));
XOR2X1 exu_bypass_w2_eccgen_U173(.A(bypass_w2_eccgen_p1_w[1]), .B(bypass_w2_eccgen_p1_w[0]), .Y(exu_n20357));
XOR2X1 exu_bypass_w2_eccgen_U172(.A(bypass_w2_eccgen_p1_w[3]), .B(bypass_w2_eccgen_p1_w[2]), .Y(exu_n20358));
XOR2X1 exu_bypass_w2_eccgen_U171(.A(bypass_w2_eccgen_p1_w[5]), .B(bypass_w2_eccgen_p1_w[4]), .Y(exu_n20359));
XOR2X1 exu_bypass_w2_eccgen_U170(.A(bypass_w2_eccgen_p1_w[7]), .B(bypass_w2_eccgen_p1_w[6]), .Y(exu_n20360));
XOR2X1 exu_bypass_w2_eccgen_U169(.A(exu_n20362), .B(exu_n20361), .Y(bypass_rd_synd_w2_l[2]));
XOR2X1 exu_bypass_w2_eccgen_U168(.A(exu_n20364), .B(exu_n20363), .Y(exu_n20361));
XOR2X1 exu_bypass_w2_eccgen_U167(.A(exu_n20366), .B(exu_n20365), .Y(exu_n20362));
XOR2X1 exu_bypass_w2_eccgen_U166(.A(bypass_w2_eccgen_p2_w[1]), .B(bypass_w2_eccgen_p2_w[0]), .Y(exu_n20363));
XOR2X1 exu_bypass_w2_eccgen_U165(.A(bypass_w2_eccgen_p2_w[3]), .B(bypass_w2_eccgen_p2_w[2]), .Y(exu_n20364));
XOR2X1 exu_bypass_w2_eccgen_U164(.A(bypass_w2_eccgen_p2_w[5]), .B(bypass_w2_eccgen_p2_w[4]), .Y(exu_n20365));
XOR2X1 exu_bypass_w2_eccgen_U163(.A(bypass_w2_eccgen_p2_w[7]), .B(bypass_w2_eccgen_p2_w[6]), .Y(exu_n20366));
XOR2X1 exu_bypass_w2_eccgen_U162(.A(exu_n20368), .B(exu_n20367), .Y(bypass_rd_synd_w2_l[3]));
XOR2X1 exu_bypass_w2_eccgen_U161(.A(exu_n20370), .B(exu_n20369), .Y(exu_n20367));
XOR2X1 exu_bypass_w2_eccgen_U160(.A(exu_n20372), .B(exu_n20371), .Y(exu_n20368));
XOR2X1 exu_bypass_w2_eccgen_U159(.A(bypass_w2_eccgen_p3_w[1]), .B(bypass_w2_eccgen_p3_w[0]), .Y(exu_n20369));
XOR2X1 exu_bypass_w2_eccgen_U158(.A(bypass_w2_eccgen_p3_w[3]), .B(bypass_w2_eccgen_p3_w[2]), .Y(exu_n20370));
XOR2X1 exu_bypass_w2_eccgen_U157(.A(bypass_w2_eccgen_p3_w[5]), .B(bypass_w2_eccgen_p3_w[4]), .Y(exu_n20371));
XOR2X1 exu_bypass_w2_eccgen_U156(.A(bypass_w2_eccgen_p3_w[7]), .B(bypass_w2_eccgen_p3_w[6]), .Y(exu_n20372));
XOR2X1 exu_bypass_w2_eccgen_U155(.A(exu_n20374), .B(exu_n20373), .Y(bypass_rd_synd_w2_l[4]));
XOR2X1 exu_bypass_w2_eccgen_U154(.A(bypass_w2_eccgen_p4_w[0]), .B(exu_n20375), .Y(exu_n20373));
XOR2X1 exu_bypass_w2_eccgen_U153(.A(bypass_w2_eccgen_p4_w[2]), .B(bypass_w2_eccgen_p4_w[1]), .Y(exu_n20374));
XOR2X1 exu_bypass_w2_eccgen_U152(.A(bypass_w2_eccgen_msk_w4), .B(bypass_w2_eccgen_p4_w[3]), .Y(exu_n20375));
XOR2X1 exu_bypass_w2_eccgen_U151(.A(exu_n20377), .B(exu_n20376), .Y(bypass_rd_synd_w2_l[5]));
XOR2X1 exu_bypass_w2_eccgen_U150(.A(bypass_w2_eccgen_p5_w[0]), .B(exu_n20378), .Y(exu_n20376));
XOR2X1 exu_bypass_w2_eccgen_U149(.A(bypass_w2_eccgen_p4_w[2]), .B(bypass_w2_eccgen_p5_w[1]), .Y(exu_n20377));
XOR2X1 exu_bypass_w2_eccgen_U148(.A(bypass_w2_eccgen_msk_w5), .B(bypass_w2_eccgen_p4_w[3]), .Y(exu_n20378));
XOR2X1 exu_bypass_w2_eccgen_U147(.A(exu_n20380), .B(exu_n20379), .Y(bypass_rd_synd_w2_l[7]));
XOR2X1 exu_bypass_w2_eccgen_U146(.A(exu_n20382), .B(exu_n20381), .Y(exu_n20379));
XOR2X1 exu_bypass_w2_eccgen_U145(.A(exu_n20384), .B(exu_n20383), .Y(exu_n20380));
XOR2X1 exu_bypass_w2_eccgen_U144(.A(bypass_w2_eccgen_p7_w[1]), .B(bypass_w2_eccgen_p7_w[0]), .Y(exu_n20381));
XOR2X1 exu_bypass_w2_eccgen_U143(.A(bypass_w2_eccgen_p7_w[3]), .B(bypass_w2_eccgen_p7_w[2]), .Y(exu_n20382));
XOR2X1 exu_bypass_w2_eccgen_U142(.A(bypass_w2_eccgen_p7_w[5]), .B(bypass_w2_eccgen_p7_w[4]), .Y(exu_n20383));
XOR2X1 exu_bypass_w2_eccgen_U141(.A(bypass_w2_eccgen_p7_w[7]), .B(bypass_w2_eccgen_p7_w[6]), .Y(exu_n20384));
XOR2X1 exu_bypass_w2_eccgen_U140(.A(exu_n15810), .B(exu_n20385), .Y(exu_n20472));
XOR2X1 exu_bypass_w2_eccgen_U139(.A(exu_n15801), .B(exu_n15813), .Y(exu_n20385));
XOR2X1 exu_bypass_w2_eccgen_U138(.A(exu_n15831), .B(exu_n20472), .Y(bypass_w2_eccgen_p7_g[0]));
XOR2X1 exu_bypass_w2_eccgen_U137(.A(exu_n20387), .B(exu_n20386), .Y(bypass_w2_eccgen_p7_g[1]));
XOR2X1 exu_bypass_w2_eccgen_U136(.A(exu_n15825), .B(exu_n15833), .Y(exu_n20386));
XOR2X1 exu_bypass_w2_eccgen_U135(.A(exu_n15838), .B(exu_n15850), .Y(exu_n20387));
XOR2X1 exu_bypass_w2_eccgen_U134(.A(exu_n20389), .B(exu_n20388), .Y(bypass_w2_eccgen_p7_g[2]));
XOR2X1 exu_bypass_w2_eccgen_U133(.A(exu_n15793), .B(exu_n15809), .Y(exu_n20388));
XOR2X1 exu_bypass_w2_eccgen_U132(.A(exu_n15792), .B(exu_n15929), .Y(exu_n20389));
XOR2X1 exu_bypass_w2_eccgen_U131(.A(exu_n15847), .B(exu_n20390), .Y(exu_n20473));
XOR2X1 exu_bypass_w2_eccgen_U130(.A(exu_n15806), .B(exu_n15807), .Y(exu_n20390));
XOR2X1 exu_bypass_w2_eccgen_U129(.A(exu_n15837), .B(exu_n20473), .Y(bypass_w2_eccgen_p7_g[3]));
XOR2X1 exu_bypass_w2_eccgen_U128(.A(exu_n20392), .B(exu_n20391), .Y(bypass_w2_eccgen_p7_g[4]));
XOR2X1 exu_bypass_w2_eccgen_U127(.A(exu_n15789), .B(exu_n15805), .Y(exu_n20391));
XOR2X1 exu_bypass_w2_eccgen_U126(.A(exu_n15788), .B(exu_n15928), .Y(exu_n20392));
XOR2X1 exu_bypass_w2_eccgen_U125(.A(exu_n20394), .B(exu_n20393), .Y(bypass_w2_eccgen_p7_g[5]));
XOR2X1 exu_bypass_w2_eccgen_U124(.A(exu_n15829), .B(exu_n15927), .Y(exu_n20393));
XOR2X1 exu_bypass_w2_eccgen_U123(.A(exu_n15828), .B(exu_n15844), .Y(exu_n20394));
XOR2X1 exu_bypass_w2_eccgen_U122(.A(exu_n15841), .B(exu_n20395), .Y(exu_n20474));
XOR2X1 exu_bypass_w2_eccgen_U121(.A(exu_n15800), .B(exu_n15855), .Y(exu_n20395));
XOR2X1 exu_bypass_w2_eccgen_U120(.A(exu_n15802), .B(exu_n20474), .Y(bypass_w2_eccgen_p7_g[6]));
XOR2X1 exu_bypass_w2_eccgen_U119(.A(exu_n15798), .B(exu_n20396), .Y(exu_n20465));
XOR2X1 exu_bypass_w2_eccgen_U118(.A(exu_n15780), .B(exu_n15811), .Y(exu_n20396));
XOR2X1 exu_bypass_w2_eccgen_U117(.A(exu_n20398), .B(exu_n20397), .Y(bypass_w2_eccgen_p7_g[7]));
XOR2X1 exu_bypass_w2_eccgen_U116(.A(exu_n20400), .B(exu_n20399), .Y(exu_n20397));
XOR2X1 exu_bypass_w2_eccgen_U115(.A(exu_n15513), .B(exu_n20465), .Y(exu_n20398));
XOR2X1 exu_bypass_w2_eccgen_U114(.A(exu_n15827), .B(exu_n15835), .Y(exu_n20399));
XOR2X1 exu_bypass_w2_eccgen_U113(.A(exu_n15826), .B(exu_n15834), .Y(exu_n20400));
XOR2X1 exu_bypass_w2_eccgen_U112(.A(exu_n15797), .B(exu_n20465), .Y(bypass_w2_eccgen_p6_g[0]));
XOR2X1 exu_bypass_w2_eccgen_U111(.A(exu_n15779), .B(exu_n20401), .Y(exu_n20468));
XOR2X1 exu_bypass_w2_eccgen_U110(.A(exu_n15826), .B(exu_n15796), .Y(exu_n20401));
XOR2X1 exu_bypass_w2_eccgen_U109(.A(exu_n15514), .B(exu_n20468), .Y(bypass_w2_eccgen_p6_g[1]));
XOR2X1 exu_bypass_w2_eccgen_U108(.A(exu_n20403), .B(exu_n20402), .Y(bypass_w2_eccgen_p5_g[0]));
XOR2X1 exu_bypass_w2_eccgen_U107(.A(bypass_w2_eccgen_p7_g[4]), .B(exu_n20404), .Y(exu_n20402));
XOR2X1 exu_bypass_w2_eccgen_U106(.A(exu_n15846), .B(exu_n15806), .Y(exu_n20403));
XOR2X1 exu_bypass_w2_eccgen_U105(.A(exu_n15830), .B(exu_n15845), .Y(exu_n20404));
XOR2X1 exu_bypass_w2_eccgen_U104(.A(exu_n20406), .B(exu_n20405), .Y(bypass_w2_eccgen_p3_g[4]));
XOR2X1 exu_bypass_w2_eccgen_U103(.A(exu_n15787), .B(exu_n15804), .Y(exu_n20405));
XOR2X1 exu_bypass_w2_eccgen_U102(.A(exu_n15786), .B(exu_n15927), .Y(exu_n20406));
XOR2X1 exu_bypass_w2_eccgen_U101(.A(exu_n15829), .B(exu_n20407), .Y(exu_n20467));
XOR2X1 exu_bypass_w2_eccgen_U100(.A(exu_n15842), .B(exu_n15844), .Y(exu_n20407));
XOR2X1 exu_bypass_w2_eccgen_U99(.A(exu_n20467), .B(exu_n20408), .Y(bypass_w2_eccgen_p5_g[1]));
XOR2X1 exu_bypass_w2_eccgen_U98(.A(exu_n15828), .B(bypass_w2_eccgen_p3_g[4]), .Y(exu_n20408));
XOR2X1 exu_bypass_w2_eccgen_U97(.A(exu_n20410), .B(exu_n20409), .Y(bypass_w2_eccgen_p4_g[0]));
XOR2X1 exu_bypass_w2_eccgen_U96(.A(bypass_w2_eccgen_p7_g[2]), .B(exu_n20411), .Y(exu_n20409));
XOR2X1 exu_bypass_w2_eccgen_U95(.A(exu_n15849), .B(exu_n15838), .Y(exu_n20410));
XOR2X1 exu_bypass_w2_eccgen_U94(.A(exu_n15832), .B(exu_n15848), .Y(exu_n20411));
XOR2X1 exu_bypass_w2_eccgen_U93(.A(exu_n20413), .B(exu_n20412), .Y(bypass_w2_eccgen_p3_g[2]));
XOR2X1 exu_bypass_w2_eccgen_U92(.A(exu_n15791), .B(exu_n15808), .Y(exu_n20412));
XOR2X1 exu_bypass_w2_eccgen_U91(.A(exu_n15790), .B(exu_n15847), .Y(exu_n20413));
XOR2X1 exu_bypass_w2_eccgen_U90(.A(exu_n15807), .B(exu_n20414), .Y(exu_n20466));
XOR2X1 exu_bypass_w2_eccgen_U89(.A(exu_n15836), .B(exu_n15837), .Y(exu_n20414));
XOR2X1 exu_bypass_w2_eccgen_U88(.A(exu_n20466), .B(exu_n20415), .Y(bypass_w2_eccgen_p4_g[1]));
XOR2X1 exu_bypass_w2_eccgen_U87(.A(exu_n15828), .B(bypass_w2_eccgen_p3_g[2]), .Y(exu_n20415));
XOR2X1 exu_bypass_w2_eccgen_U86(.A(exu_n15783), .B(exu_n15802), .Y(exu_n20471));
XOR2X1 exu_bypass_w2_eccgen_U85(.A(exu_n20417), .B(exu_n20416), .Y(bypass_w2_eccgen_p4_g[2]));
XOR2X1 exu_bypass_w2_eccgen_U84(.A(exu_n20419), .B(exu_n20418), .Y(exu_n20416));
XOR2X1 exu_bypass_w2_eccgen_U83(.A(exu_n20471), .B(exu_n20420), .Y(exu_n20417));
XOR2X1 exu_bypass_w2_eccgen_U82(.A(exu_n15785), .B(exu_n15803), .Y(exu_n20418));
XOR2X1 exu_bypass_w2_eccgen_U81(.A(exu_n15784), .B(exu_n15841), .Y(exu_n20419));
XOR2X1 exu_bypass_w2_eccgen_U80(.A(exu_n15782), .B(exu_n15855), .Y(exu_n20420));
XOR2X1 exu_bypass_w2_eccgen_U79(.A(exu_n20422), .B(exu_n20421), .Y(bypass_w2_eccgen_p3_g[6]));
XOR2X1 exu_bypass_w2_eccgen_U78(.A(exu_n15835), .B(exu_n15800), .Y(exu_n20421));
XOR2X1 exu_bypass_w2_eccgen_U77(.A(exu_n15827), .B(exu_n15812), .Y(exu_n20422));
XOR2X1 exu_bypass_w2_eccgen_U76(.A(exu_n15781), .B(exu_n20423), .Y(exu_n20469));
XOR2X1 exu_bypass_w2_eccgen_U75(.A(exu_n15834), .B(exu_n15799), .Y(exu_n20423));
XOR2X1 exu_bypass_w2_eccgen_U74(.A(bypass_w2_eccgen_p3_g[6]), .B(exu_n20469), .Y(bypass_w2_eccgen_p4_g[3]));
XOR2X1 exu_bypass_w2_eccgen_U73(.A(exu_n20425), .B(exu_n20424), .Y(bypass_w2_eccgen_p3_g[0]));
XOR2X1 exu_bypass_w2_eccgen_U72(.A(exu_n15833), .B(exu_n15801), .Y(exu_n20424));
XOR2X1 exu_bypass_w2_eccgen_U71(.A(exu_n15825), .B(exu_n15854), .Y(exu_n20425));
XOR2X1 exu_bypass_w2_eccgen_U70(.A(exu_n15850), .B(exu_n15418), .Y(exu_n20470));
XOR2X1 exu_bypass_w2_eccgen_U69(.A(exu_n20470), .B(exu_n20426), .Y(bypass_w2_eccgen_p3_g[1]));
XOR2X1 exu_bypass_w2_eccgen_U68(.A(exu_n15792), .B(exu_n15840), .Y(exu_n20426));
XOR2X1 exu_bypass_w2_eccgen_U67(.A(exu_n15788), .B(exu_n20466), .Y(bypass_w2_eccgen_p3_g[3]));
XOR2X1 exu_bypass_w2_eccgen_U66(.A(exu_n15782), .B(exu_n20467), .Y(bypass_w2_eccgen_p3_g[5]));
XOR2X1 exu_bypass_w2_eccgen_U65(.A(exu_n15515), .B(exu_n20469), .Y(bypass_w2_eccgen_p3_g[7]));
XOR2X1 exu_bypass_w2_eccgen_U64(.A(exu_n20428), .B(exu_n20427), .Y(bypass_w2_eccgen_p2_g[0]));
XOR2X1 exu_bypass_w2_eccgen_U63(.A(exu_n15831), .B(exu_n15813), .Y(exu_n20427));
XOR2X1 exu_bypass_w2_eccgen_U62(.A(exu_n15825), .B(exu_n15843), .Y(exu_n20428));
XOR2X1 exu_bypass_w2_eccgen_U61(.A(exu_n20470), .B(exu_n20429), .Y(bypass_w2_eccgen_p2_g[1]));
XOR2X1 exu_bypass_w2_eccgen_U60(.A(exu_n15793), .B(exu_n15840), .Y(exu_n20429));
XOR2X1 exu_bypass_w2_eccgen_U59(.A(exu_n20431), .B(exu_n20430), .Y(bypass_w2_eccgen_p2_g[2]));
XOR2X1 exu_bypass_w2_eccgen_U58(.A(exu_n15832), .B(exu_n15848), .Y(exu_n20430));
XOR2X1 exu_bypass_w2_eccgen_U57(.A(exu_n15790), .B(exu_n15929), .Y(exu_n20431));
XOR2X1 exu_bypass_w2_eccgen_U56(.A(exu_n15789), .B(exu_n20466), .Y(bypass_w2_eccgen_p2_g[3]));
XOR2X1 exu_bypass_w2_eccgen_U55(.A(exu_n20433), .B(exu_n20432), .Y(bypass_w2_eccgen_p2_g[4]));
XOR2X1 exu_bypass_w2_eccgen_U54(.A(exu_n15830), .B(exu_n15845), .Y(exu_n20432));
XOR2X1 exu_bypass_w2_eccgen_U53(.A(exu_n15786), .B(exu_n15928), .Y(exu_n20433));
XOR2X1 exu_bypass_w2_eccgen_U52(.A(exu_n15784), .B(exu_n20467), .Y(bypass_w2_eccgen_p2_g[5]));
XOR2X1 exu_bypass_w2_eccgen_U51(.A(exu_n20471), .B(exu_n20434), .Y(bypass_w2_eccgen_p2_g[6]));
XOR2X1 exu_bypass_w2_eccgen_U50(.A(exu_n15827), .B(exu_n15855), .Y(exu_n20434));
XOR2X1 exu_bypass_w2_eccgen_U49(.A(exu_n20436), .B(exu_n20435), .Y(bypass_w2_eccgen_p2_g[7]));
XOR2X1 exu_bypass_w2_eccgen_U48(.A(exu_n20469), .B(exu_n20468), .Y(exu_n20435));
XOR2X1 exu_bypass_w2_eccgen_U47(.A(exu_n15780), .B(exu_n15550), .Y(exu_n20436));
XOR2X1 exu_bypass_w2_eccgen_U46(.A(exu_n20438), .B(exu_n20437), .Y(bypass_w2_eccgen_p1_g[0]));
XOR2X1 exu_bypass_w2_eccgen_U45(.A(exu_n15831), .B(exu_n15810), .Y(exu_n20437));
XOR2X1 exu_bypass_w2_eccgen_U44(.A(exu_n15833), .B(exu_n15843), .Y(exu_n20438));
XOR2X1 exu_bypass_w2_eccgen_U43(.A(exu_n20470), .B(exu_n20439), .Y(bypass_w2_eccgen_p1_g[1]));
XOR2X1 exu_bypass_w2_eccgen_U42(.A(exu_n15809), .B(exu_n15854), .Y(exu_n20439));
XOR2X1 exu_bypass_w2_eccgen_U41(.A(exu_n20441), .B(exu_n20440), .Y(bypass_w2_eccgen_p1_g[2]));
XOR2X1 exu_bypass_w2_eccgen_U40(.A(exu_n15832), .B(exu_n15849), .Y(exu_n20440));
XOR2X1 exu_bypass_w2_eccgen_U39(.A(exu_n15791), .B(exu_n15929), .Y(exu_n20441));
XOR2X1 exu_bypass_w2_eccgen_U38(.A(exu_n20443), .B(exu_n20442), .Y(bypass_w2_eccgen_p1_g[3]));
XOR2X1 exu_bypass_w2_eccgen_U37(.A(exu_n15837), .B(exu_n15847), .Y(exu_n20442));
XOR2X1 exu_bypass_w2_eccgen_U36(.A(exu_n15805), .B(exu_n15836), .Y(exu_n20443));
XOR2X1 exu_bypass_w2_eccgen_U35(.A(exu_n20445), .B(exu_n20444), .Y(bypass_w2_eccgen_p1_g[4]));
XOR2X1 exu_bypass_w2_eccgen_U34(.A(exu_n15830), .B(exu_n15846), .Y(exu_n20444));
XOR2X1 exu_bypass_w2_eccgen_U33(.A(exu_n15787), .B(exu_n15928), .Y(exu_n20445));
XOR2X1 exu_bypass_w2_eccgen_U32(.A(exu_n20447), .B(exu_n20446), .Y(bypass_w2_eccgen_p1_g[5]));
XOR2X1 exu_bypass_w2_eccgen_U31(.A(exu_n15844), .B(exu_n15927), .Y(exu_n20446));
XOR2X1 exu_bypass_w2_eccgen_U30(.A(exu_n15785), .B(exu_n15842), .Y(exu_n20447));
XOR2X1 exu_bypass_w2_eccgen_U29(.A(exu_n20471), .B(exu_n20448), .Y(bypass_w2_eccgen_p1_g[6]));
XOR2X1 exu_bypass_w2_eccgen_U28(.A(exu_n15835), .B(exu_n15841), .Y(exu_n20448));
XOR2X1 exu_bypass_w2_eccgen_U27(.A(exu_n20450), .B(exu_n20449), .Y(exu_n20475));
XOR2X1 exu_bypass_w2_eccgen_U26(.A(exu_n15834), .B(exu_n15812), .Y(exu_n20449));
XOR2X1 exu_bypass_w2_eccgen_U25(.A(exu_n15826), .B(exu_n15797), .Y(exu_n20450));
XOR2X1 exu_bypass_w2_eccgen_U24(.A(exu_n20452), .B(exu_n20451), .Y(bypass_w2_eccgen_p1_g[7]));
XOR2X1 exu_bypass_w2_eccgen_U23(.A(exu_n20475), .B(exu_n20453), .Y(exu_n20451));
XOR2X1 exu_bypass_w2_eccgen_U22(.A(exu_n15799), .B(exu_n15551), .Y(exu_n20452));
XOR2X1 exu_bypass_w2_eccgen_U21(.A(exu_n15796), .B(exu_n15811), .Y(exu_n20453));
XOR2X1 exu_bypass_w2_eccgen_U20(.A(exu_n15843), .B(exu_n20472), .Y(bypass_w2_eccgen_p0_g[0]));
XOR2X1 exu_bypass_w2_eccgen_U19(.A(exu_n20455), .B(exu_n20454), .Y(bypass_w2_eccgen_p0_g[1]));
XOR2X1 exu_bypass_w2_eccgen_U18(.A(exu_n15840), .B(exu_n15854), .Y(exu_n20454));
XOR2X1 exu_bypass_w2_eccgen_U17(.A(exu_n15838), .B(exu_n15850), .Y(exu_n20455));
XOR2X1 exu_bypass_w2_eccgen_U16(.A(exu_n20457), .B(exu_n20456), .Y(bypass_w2_eccgen_p0_g[2]));
XOR2X1 exu_bypass_w2_eccgen_U15(.A(exu_n15848), .B(exu_n15849), .Y(exu_n20456));
XOR2X1 exu_bypass_w2_eccgen_U14(.A(exu_n15808), .B(exu_n15929), .Y(exu_n20457));
XOR2X1 exu_bypass_w2_eccgen_U13(.A(exu_n15836), .B(exu_n20473), .Y(bypass_w2_eccgen_p0_g[3]));
XOR2X1 exu_bypass_w2_eccgen_U12(.A(exu_n20459), .B(exu_n20458), .Y(bypass_w2_eccgen_p0_g[4]));
XOR2X1 exu_bypass_w2_eccgen_U11(.A(exu_n15845), .B(exu_n15846), .Y(exu_n20458));
XOR2X1 exu_bypass_w2_eccgen_U10(.A(exu_n15804), .B(exu_n15928), .Y(exu_n20459));
XOR2X1 exu_bypass_w2_eccgen_U9(.A(exu_n20461), .B(exu_n20460), .Y(bypass_w2_eccgen_p0_g[5]));
XOR2X1 exu_bypass_w2_eccgen_U8(.A(exu_n15829), .B(exu_n15927), .Y(exu_n20460));
XOR2X1 exu_bypass_w2_eccgen_U7(.A(exu_n15803), .B(exu_n15842), .Y(exu_n20461));
XOR2X1 exu_bypass_w2_eccgen_U6(.A(exu_n15783), .B(exu_n20474), .Y(bypass_w2_eccgen_p0_g[6]));
XOR2X1 exu_bypass_w2_eccgen_U5(.A(exu_n20463), .B(exu_n20462), .Y(bypass_w2_eccgen_p0_g[7]));
XOR2X1 exu_bypass_w2_eccgen_U4(.A(exu_n20475), .B(exu_n20464), .Y(exu_n20462));
XOR2X1 exu_bypass_w2_eccgen_U3(.A(exu_n15781), .B(exu_n15552), .Y(exu_n20463));
XOR2X1 exu_bypass_w2_eccgen_U2(.A(exu_n15779), .B(exu_n15798), .Y(exu_n20464));
XOR2X1 exu_bypass_w2_eccgen_U1(.A(bypass_w2_eccgen_p6_w[1]), .B(bypass_w2_eccgen_p6_w[0]), .Y(bypass_rd_synd_w2_l[6]));
DFFPOSX1 ecl_writeback_rdpr_dff_q_reg[0](.D(exu_n20347), .CLK(rclk), .Q(ecl_byp_eclpr_e[0]));
DFFPOSX1 ecl_writeback_rdpr_dff_q_reg[1](.D(exu_n20346), .CLK(rclk), .Q(ecl_byp_eclpr_e[1]));
DFFPOSX1 ecl_writeback_rdpr_dff_q_reg[2](.D(exu_n20345), .CLK(rclk), .Q(ecl_byp_eclpr_e[2]));
DFFPOSX1 ecl_writeback_rdpr_dff_q_reg[3](.D(exu_n20344), .CLK(rclk), .Q(ecl_byp_eclpr_e[3]));
DFFPOSX1 ecl_writeback_rdpr_dff_q_reg[4](.D(exu_n20343), .CLK(rclk), .Q(ecl_byp_eclpr_e[4]));
DFFPOSX1 ecl_writeback_rdpr_dff_q_reg[5](.D(exu_n20342), .CLK(rclk), .Q(ecl_byp_eclpr_e[5]));
DFFPOSX1 ecl_writeback_rdpr_dff_q_reg[6](.D(exu_n20341), .CLK(rclk), .Q(ecl_byp_eclpr_e[6]));
DFFPOSX1 ecl_writeback_rdpr_dff_q_reg[7](.D(exu_n20348), .CLK(rclk), .Q(ecl_byp_eclpr_e[7]));
DFFPOSX1 ecl_ccr_dff_ccr_thr3_q_reg[0](.D(exu_n20338), .CLK(rclk), .Q(exu_tlu_ccr3_w[0]));
DFFPOSX1 ecl_ccr_dff_ccr_thr3_q_reg[1](.D(exu_n20337), .CLK(rclk), .Q(exu_tlu_ccr3_w[1]));
DFFPOSX1 ecl_ccr_dff_ccr_thr3_q_reg[2](.D(exu_n20336), .CLK(rclk), .Q(exu_tlu_ccr3_w[2]));
DFFPOSX1 ecl_ccr_dff_ccr_thr3_q_reg[3](.D(exu_n20335), .CLK(rclk), .Q(exu_tlu_ccr3_w[3]));
DFFPOSX1 ecl_ccr_dff_ccr_thr3_q_reg[4](.D(exu_n20334), .CLK(rclk), .Q(exu_tlu_ccr3_w[4]));
DFFPOSX1 ecl_ccr_dff_ccr_thr3_q_reg[5](.D(exu_n20333), .CLK(rclk), .Q(exu_tlu_ccr3_w[5]));
DFFPOSX1 ecl_ccr_dff_ccr_thr3_q_reg[6](.D(exu_n20332), .CLK(rclk), .Q(exu_tlu_ccr3_w[6]));
DFFPOSX1 ecl_ccr_dff_ccr_thr3_q_reg[7](.D(exu_n20339), .CLK(rclk), .Q(exu_tlu_ccr3_w[7]));
DFFPOSX1 ecl_ccr_dff_ccr_thr2_q_reg[0](.D(exu_n20329), .CLK(rclk), .Q(exu_tlu_ccr2_w[0]));
DFFPOSX1 ecl_ccr_dff_ccr_thr2_q_reg[1](.D(exu_n20328), .CLK(rclk), .Q(exu_tlu_ccr2_w[1]));
DFFPOSX1 ecl_ccr_dff_ccr_thr2_q_reg[2](.D(exu_n20327), .CLK(rclk), .Q(exu_tlu_ccr2_w[2]));
DFFPOSX1 ecl_ccr_dff_ccr_thr2_q_reg[3](.D(exu_n20326), .CLK(rclk), .Q(exu_tlu_ccr2_w[3]));
DFFPOSX1 ecl_ccr_dff_ccr_thr2_q_reg[4](.D(exu_n20325), .CLK(rclk), .Q(exu_tlu_ccr2_w[4]));
DFFPOSX1 ecl_ccr_dff_ccr_thr2_q_reg[5](.D(exu_n20324), .CLK(rclk), .Q(exu_tlu_ccr2_w[5]));
DFFPOSX1 ecl_ccr_dff_ccr_thr2_q_reg[6](.D(exu_n20323), .CLK(rclk), .Q(exu_tlu_ccr2_w[6]));
DFFPOSX1 ecl_ccr_dff_ccr_thr2_q_reg[7](.D(exu_n20330), .CLK(rclk), .Q(exu_tlu_ccr2_w[7]));
DFFPOSX1 ecl_ccr_dff_ccr_thr1_q_reg[0](.D(exu_n20320), .CLK(rclk), .Q(exu_tlu_ccr1_w[0]));
DFFPOSX1 ecl_ccr_dff_ccr_thr1_q_reg[1](.D(exu_n20319), .CLK(rclk), .Q(exu_tlu_ccr1_w[1]));
DFFPOSX1 ecl_ccr_dff_ccr_thr1_q_reg[2](.D(exu_n20318), .CLK(rclk), .Q(exu_tlu_ccr1_w[2]));
DFFPOSX1 ecl_ccr_dff_ccr_thr1_q_reg[3](.D(exu_n20317), .CLK(rclk), .Q(exu_tlu_ccr1_w[3]));
DFFPOSX1 ecl_ccr_dff_ccr_thr1_q_reg[4](.D(exu_n20316), .CLK(rclk), .Q(exu_tlu_ccr1_w[4]));
DFFPOSX1 ecl_ccr_dff_ccr_thr1_q_reg[5](.D(exu_n20315), .CLK(rclk), .Q(exu_tlu_ccr1_w[5]));
DFFPOSX1 ecl_ccr_dff_ccr_thr1_q_reg[6](.D(exu_n20314), .CLK(rclk), .Q(exu_tlu_ccr1_w[6]));
DFFPOSX1 ecl_ccr_dff_ccr_thr1_q_reg[7](.D(exu_n20321), .CLK(rclk), .Q(exu_tlu_ccr1_w[7]));
DFFPOSX1 ecl_ccr_dff_ccr_thr0_q_reg[0](.D(exu_n20311), .CLK(rclk), .Q(exu_tlu_ccr0_w[0]));
DFFPOSX1 ecl_ccr_dff_ccr_thr0_q_reg[1](.D(exu_n20310), .CLK(rclk), .Q(exu_tlu_ccr0_w[1]));
DFFPOSX1 ecl_ccr_dff_ccr_thr0_q_reg[2](.D(exu_n20309), .CLK(rclk), .Q(exu_tlu_ccr0_w[2]));
DFFPOSX1 ecl_ccr_dff_ccr_thr0_q_reg[3](.D(exu_n20308), .CLK(rclk), .Q(exu_tlu_ccr0_w[3]));
DFFPOSX1 ecl_ccr_dff_ccr_thr0_q_reg[4](.D(exu_n20307), .CLK(rclk), .Q(exu_tlu_ccr0_w[4]));
DFFPOSX1 ecl_ccr_dff_ccr_thr0_q_reg[5](.D(exu_n20306), .CLK(rclk), .Q(exu_tlu_ccr0_w[5]));
DFFPOSX1 ecl_ccr_dff_ccr_thr0_q_reg[6](.D(exu_n20305), .CLK(rclk), .Q(exu_tlu_ccr0_w[6]));
DFFPOSX1 ecl_ccr_dff_ccr_thr0_q_reg[7](.D(exu_n20312), .CLK(rclk), .Q(exu_tlu_ccr0_w[7]));
DFFPOSX1 ecl_ccr_dff_cc_m2w_q_reg[0](.D(exu_n20302), .CLK(rclk), .Q(ecl_ccr_alu_cc_w[0]));
DFFPOSX1 ecl_ccr_dff_cc_m2w_q_reg[1](.D(exu_n20301), .CLK(rclk), .Q(ecl_ccr_alu_cc_w[1]));
DFFPOSX1 ecl_ccr_dff_cc_m2w_q_reg[2](.D(exu_n20300), .CLK(rclk), .Q(ecl_ccr_alu_cc_w[2]));
DFFPOSX1 ecl_ccr_dff_cc_m2w_q_reg[3](.D(exu_n20299), .CLK(rclk), .Q(ecl_ccr_alu_cc_w[3]));
DFFPOSX1 ecl_ccr_dff_cc_m2w_q_reg[4](.D(exu_n20298), .CLK(rclk), .Q(ecl_ccr_alu_cc_w[4]));
DFFPOSX1 ecl_ccr_dff_cc_m2w_q_reg[5](.D(exu_n20297), .CLK(rclk), .Q(ecl_ccr_alu_cc_w[5]));
DFFPOSX1 ecl_ccr_dff_cc_m2w_q_reg[6](.D(exu_n20296), .CLK(rclk), .Q(ecl_ccr_alu_cc_w[6]));
DFFPOSX1 ecl_ccr_dff_cc_m2w_q_reg[7](.D(exu_n20303), .CLK(rclk), .Q(ecl_ccr_alu_cc_w[7]));
DFFPOSX1 ecl_ccr_dff_cc_e2m_q_reg[0](.D(exu_n20293), .CLK(rclk), .Q(ecl_ccr_alu_cc_m[0]));
DFFPOSX1 ecl_ccr_dff_cc_e2m_q_reg[1](.D(exu_n20292), .CLK(rclk), .Q(ecl_ccr_alu_cc_m[1]));
DFFPOSX1 ecl_ccr_dff_cc_e2m_q_reg[2](.D(exu_n20291), .CLK(rclk), .Q(ecl_ccr_alu_cc_m[2]));
DFFPOSX1 ecl_ccr_dff_cc_e2m_q_reg[3](.D(exu_n20290), .CLK(rclk), .Q(ecl_ccr_alu_cc_m[3]));
DFFPOSX1 ecl_ccr_dff_cc_e2m_q_reg[4](.D(exu_n20289), .CLK(rclk), .Q(ecl_ccr_alu_cc_m[4]));
DFFPOSX1 ecl_ccr_dff_cc_e2m_q_reg[5](.D(exu_n20288), .CLK(rclk), .Q(ecl_ccr_alu_cc_m[5]));
DFFPOSX1 ecl_ccr_dff_cc_e2m_q_reg[6](.D(exu_n20287), .CLK(rclk), .Q(ecl_ccr_alu_cc_m[6]));
DFFPOSX1 ecl_ccr_dff_cc_e2m_q_reg[7](.D(exu_n20294), .CLK(rclk), .Q(ecl_ccr_alu_cc_m[7]));
DFFPOSX1 ecc_rs3_ecc_d2e_q_reg[0](.D(exu_n20284), .CLK(rclk), .Q(ecc_rs3_ecc_e[0]));
DFFPOSX1 ecc_rs3_ecc_d2e_q_reg[1](.D(exu_n20283), .CLK(rclk), .Q(ecc_rs3_ecc_e[1]));
DFFPOSX1 ecc_rs3_ecc_d2e_q_reg[2](.D(exu_n20282), .CLK(rclk), .Q(ecc_rs3_ecc_e[2]));
DFFPOSX1 ecc_rs3_ecc_d2e_q_reg[3](.D(exu_n20281), .CLK(rclk), .Q(ecc_rs3_ecc_e[3]));
DFFPOSX1 ecc_rs3_ecc_d2e_q_reg[4](.D(exu_n20280), .CLK(rclk), .Q(ecc_rs3_ecc_e[4]));
DFFPOSX1 ecc_rs3_ecc_d2e_q_reg[5](.D(exu_n20279), .CLK(rclk), .Q(ecc_rs3_ecc_e[5]));
DFFPOSX1 ecc_rs3_ecc_d2e_q_reg[6](.D(exu_n20278), .CLK(rclk), .Q(ecc_rs3_ecc_e[6]));
DFFPOSX1 ecc_rs3_ecc_d2e_q_reg[7](.D(exu_n20285), .CLK(rclk), .Q(ecc_rs3_ecc_e[7]));
DFFPOSX1 ecc_rs2_ecc_d2e_q_reg[0](.D(exu_n20275), .CLK(rclk), .Q(ecc_rs2_ecc_e[0]));
DFFPOSX1 ecc_rs2_ecc_d2e_q_reg[1](.D(exu_n20274), .CLK(rclk), .Q(ecc_rs2_ecc_e[1]));
DFFPOSX1 ecc_rs2_ecc_d2e_q_reg[2](.D(exu_n20273), .CLK(rclk), .Q(ecc_rs2_ecc_e[2]));
DFFPOSX1 ecc_rs2_ecc_d2e_q_reg[3](.D(exu_n20272), .CLK(rclk), .Q(ecc_rs2_ecc_e[3]));
DFFPOSX1 ecc_rs2_ecc_d2e_q_reg[4](.D(exu_n20271), .CLK(rclk), .Q(ecc_rs2_ecc_e[4]));
DFFPOSX1 ecc_rs2_ecc_d2e_q_reg[5](.D(exu_n20270), .CLK(rclk), .Q(ecc_rs2_ecc_e[5]));
DFFPOSX1 ecc_rs2_ecc_d2e_q_reg[6](.D(exu_n20269), .CLK(rclk), .Q(ecc_rs2_ecc_e[6]));
DFFPOSX1 ecc_rs2_ecc_d2e_q_reg[7](.D(exu_n20276), .CLK(rclk), .Q(ecc_rs2_ecc_e[7]));
XOR2X1 exu_ecc_chk_rs3_U149(.A(exu_n20140), .B(exu_n20139), .Y(exu_n20262));
XOR2X1 exu_ecc_chk_rs3_U148(.A(exu_spu_rs3_data_e[52]), .B(exu_spu_rs3_data_e[50]), .Y(exu_n20139));
XOR2X1 exu_ecc_chk_rs3_U147(.A(exu_spu_rs3_data_e[56]), .B(exu_spu_rs3_data_e[54]), .Y(exu_n20140));
XOR2X1 exu_ecc_chk_rs3_U146(.A(exu_n20142), .B(exu_n20141), .Y(exu_n20266));
XOR2X1 exu_ecc_chk_rs3_U145(.A(exu_spu_rs3_data_e[36]), .B(exu_spu_rs3_data_e[34]), .Y(exu_n20141));
XOR2X1 exu_ecc_chk_rs3_U144(.A(exu_spu_rs3_data_e[40]), .B(exu_spu_rs3_data_e[38]), .Y(exu_n20142));
XOR2X1 exu_ecc_chk_rs3_U143(.A(exu_n20144), .B(exu_n20143), .Y(exu_n20264));
XOR2X1 exu_ecc_chk_rs3_U142(.A(exu_spu_rs3_data_e[21]), .B(exu_spu_rs3_data_e[19]), .Y(exu_n20143));
XOR2X1 exu_ecc_chk_rs3_U141(.A(exu_spu_rs3_data_e[25]), .B(exu_spu_rs3_data_e[23]), .Y(exu_n20144));
XOR2X1 exu_ecc_chk_rs3_U140(.A(exu_n20146), .B(exu_n20145), .Y(exu_n20260));
XOR2X1 exu_ecc_chk_rs3_U139(.A(exu_n20148), .B(exu_n20147), .Y(exu_n20145));
XOR2X1 exu_ecc_chk_rs3_U138(.A(exu_n20264), .B(exu_n20149), .Y(exu_n20146));
XOR2X1 exu_ecc_chk_rs3_U137(.A(exu_n20262), .B(exu_n20266), .Y(exu_n20147));
XOR2X1 exu_ecc_chk_rs3_U136(.A(exu_spu_rs3_data_e[6]), .B(exu_spu_rs3_data_e[4]), .Y(exu_n20148));
XOR2X1 exu_ecc_chk_rs3_U135(.A(exu_spu_rs3_data_e[10]), .B(exu_spu_rs3_data_e[8]), .Y(exu_n20149));
XOR2X1 exu_ecc_chk_rs3_U134(.A(exu_n20151), .B(exu_n20150), .Y(exu_n20253));
XOR2X1 exu_ecc_chk_rs3_U133(.A(exu_spu_rs3_data_e[3]), .B(exu_n20152), .Y(exu_n20150));
XOR2X1 exu_ecc_chk_rs3_U132(.A(exu_spu_rs3_data_e[32]), .B(exu_spu_rs3_data_e[17]), .Y(exu_n20151));
XOR2X1 exu_ecc_chk_rs3_U131(.A(exu_spu_rs3_data_e[63]), .B(exu_spu_rs3_data_e[48]), .Y(exu_n20152));
XOR2X1 exu_ecc_chk_rs3_U130(.A(exu_n20154), .B(exu_n20153), .Y(exu_n20257));
XOR2X1 exu_ecc_chk_rs3_U129(.A(exu_spu_rs3_data_e[1]), .B(exu_n20155), .Y(exu_n20153));
XOR2X1 exu_ecc_chk_rs3_U128(.A(exu_spu_rs3_data_e[30]), .B(exu_spu_rs3_data_e[15]), .Y(exu_n20154));
XOR2X1 exu_ecc_chk_rs3_U127(.A(exu_spu_rs3_data_e[61]), .B(exu_spu_rs3_data_e[46]), .Y(exu_n20155));
XOR2X1 exu_ecc_chk_rs3_U126(.A(exu_n20157), .B(exu_n20156), .Y(exu_n20255));
XOR2X1 exu_ecc_chk_rs3_U125(.A(exu_spu_rs3_data_e[0]), .B(exu_n20158), .Y(exu_n20156));
XOR2X1 exu_ecc_chk_rs3_U124(.A(exu_spu_rs3_data_e[28]), .B(exu_spu_rs3_data_e[13]), .Y(exu_n20157));
XOR2X1 exu_ecc_chk_rs3_U123(.A(exu_spu_rs3_data_e[59]), .B(exu_spu_rs3_data_e[44]), .Y(exu_n20158));
XOR2X1 exu_ecc_chk_rs3_U122(.A(exu_n20160), .B(exu_n20159), .Y(ecc_rs3_err_e[0]));
XOR2X1 exu_ecc_chk_rs3_U121(.A(exu_n20162), .B(exu_n20161), .Y(exu_n20159));
XOR2X1 exu_ecc_chk_rs3_U120(.A(exu_n20164), .B(exu_n20163), .Y(exu_n20160));
XOR2X1 exu_ecc_chk_rs3_U119(.A(exu_n20255), .B(exu_n20165), .Y(exu_n20161));
XOR2X1 exu_ecc_chk_rs3_U118(.A(exu_n20253), .B(exu_n20257), .Y(exu_n20162));
XOR2X1 exu_ecc_chk_rs3_U117(.A(ecc_rs3_ecc_e[0]), .B(exu_n20260), .Y(exu_n20163));
XOR2X1 exu_ecc_chk_rs3_U116(.A(exu_spu_rs3_data_e[26]), .B(exu_spu_rs3_data_e[11]), .Y(exu_n20164));
XOR2X1 exu_ecc_chk_rs3_U115(.A(exu_spu_rs3_data_e[57]), .B(exu_spu_rs3_data_e[42]), .Y(exu_n20165));
XOR2X1 exu_ecc_chk_rs3_U114(.A(exu_n20167), .B(exu_n20166), .Y(exu_n20261));
XOR2X1 exu_ecc_chk_rs3_U113(.A(exu_spu_rs3_data_e[51]), .B(exu_spu_rs3_data_e[49]), .Y(exu_n20166));
XOR2X1 exu_ecc_chk_rs3_U112(.A(exu_spu_rs3_data_e[55]), .B(exu_spu_rs3_data_e[53]), .Y(exu_n20167));
XOR2X1 exu_ecc_chk_rs3_U111(.A(exu_n20169), .B(exu_n20168), .Y(exu_n20265));
XOR2X1 exu_ecc_chk_rs3_U110(.A(exu_spu_rs3_data_e[35]), .B(exu_spu_rs3_data_e[33]), .Y(exu_n20168));
XOR2X1 exu_ecc_chk_rs3_U109(.A(exu_spu_rs3_data_e[39]), .B(exu_spu_rs3_data_e[37]), .Y(exu_n20169));
XOR2X1 exu_ecc_chk_rs3_U108(.A(exu_n20171), .B(exu_n20170), .Y(exu_n20263));
XOR2X1 exu_ecc_chk_rs3_U107(.A(exu_spu_rs3_data_e[20]), .B(exu_spu_rs3_data_e[18]), .Y(exu_n20170));
XOR2X1 exu_ecc_chk_rs3_U106(.A(exu_spu_rs3_data_e[24]), .B(exu_spu_rs3_data_e[22]), .Y(exu_n20171));
XOR2X1 exu_ecc_chk_rs3_U105(.A(exu_n20173), .B(exu_n20172), .Y(exu_n20259));
XOR2X1 exu_ecc_chk_rs3_U104(.A(exu_n20175), .B(exu_n20174), .Y(exu_n20172));
XOR2X1 exu_ecc_chk_rs3_U103(.A(exu_n20263), .B(exu_n20176), .Y(exu_n20173));
XOR2X1 exu_ecc_chk_rs3_U102(.A(exu_n20261), .B(exu_n20265), .Y(exu_n20174));
XOR2X1 exu_ecc_chk_rs3_U101(.A(exu_spu_rs3_data_e[5]), .B(ecc_rs3_ecc_e[3]), .Y(exu_n20175));
XOR2X1 exu_ecc_chk_rs3_U100(.A(exu_spu_rs3_data_e[9]), .B(exu_spu_rs3_data_e[7]), .Y(exu_n20176));
XOR2X1 exu_ecc_chk_rs3_U99(.A(exu_n20178), .B(exu_n20177), .Y(exu_n20252));
XOR2X1 exu_ecc_chk_rs3_U98(.A(exu_spu_rs3_data_e[2]), .B(exu_n20179), .Y(exu_n20177));
XOR2X1 exu_ecc_chk_rs3_U97(.A(exu_spu_rs3_data_e[31]), .B(exu_spu_rs3_data_e[16]), .Y(exu_n20178));
XOR2X1 exu_ecc_chk_rs3_U96(.A(exu_spu_rs3_data_e[62]), .B(exu_spu_rs3_data_e[47]), .Y(exu_n20179));
XOR2X1 exu_ecc_chk_rs3_U95(.A(exu_n20181), .B(exu_n20180), .Y(exu_n20256));
XOR2X1 exu_ecc_chk_rs3_U94(.A(ecc_rs3_ecc_e[2]), .B(exu_n20182), .Y(exu_n20180));
XOR2X1 exu_ecc_chk_rs3_U93(.A(exu_spu_rs3_data_e[29]), .B(exu_spu_rs3_data_e[14]), .Y(exu_n20181));
XOR2X1 exu_ecc_chk_rs3_U92(.A(exu_spu_rs3_data_e[60]), .B(exu_spu_rs3_data_e[45]), .Y(exu_n20182));
XOR2X1 exu_ecc_chk_rs3_U91(.A(exu_n20184), .B(exu_n20183), .Y(exu_n20254));
XOR2X1 exu_ecc_chk_rs3_U90(.A(ecc_rs3_ecc_e[1]), .B(exu_n20185), .Y(exu_n20183));
XOR2X1 exu_ecc_chk_rs3_U89(.A(exu_spu_rs3_data_e[27]), .B(exu_spu_rs3_data_e[12]), .Y(exu_n20184));
XOR2X1 exu_ecc_chk_rs3_U88(.A(exu_spu_rs3_data_e[58]), .B(exu_spu_rs3_data_e[43]), .Y(exu_n20185));
XOR2X1 exu_ecc_chk_rs3_U87(.A(exu_n20187), .B(exu_n20186), .Y(ecc_chk_rs3_parity));
XOR2X1 exu_ecc_chk_rs3_U86(.A(exu_n20189), .B(exu_n20188), .Y(exu_n20186));
XOR2X1 exu_ecc_chk_rs3_U85(.A(exu_n20191), .B(exu_n20190), .Y(exu_n20187));
XOR2X1 exu_ecc_chk_rs3_U84(.A(exu_n20193), .B(exu_n20192), .Y(exu_n20188));
XOR2X1 exu_ecc_chk_rs3_U83(.A(exu_n20256), .B(exu_n20254), .Y(exu_n20189));
XOR2X1 exu_ecc_chk_rs3_U82(.A(exu_n20259), .B(exu_n20252), .Y(exu_n20190));
XOR2X1 exu_ecc_chk_rs3_U81(.A(ecc_rs3_ecc_e[4]), .B(ecc_rs3_err_e[0]), .Y(exu_n20191));
XOR2X1 exu_ecc_chk_rs3_U80(.A(ecc_rs3_ecc_e[6]), .B(ecc_rs3_ecc_e[5]), .Y(exu_n20192));
XOR2X1 exu_ecc_chk_rs3_U79(.A(exu_spu_rs3_data_e[41]), .B(ecc_rs3_ecc_e[7]), .Y(exu_n20193));
XOR2X1 exu_ecc_chk_rs3_U78(.A(exu_n20195), .B(exu_n20194), .Y(exu_n20258));
XOR2X1 exu_ecc_chk_rs3_U77(.A(exu_n20197), .B(exu_n20196), .Y(exu_n20194));
XOR2X1 exu_ecc_chk_rs3_U76(.A(exu_n20199), .B(exu_n20198), .Y(exu_n20195));
XOR2X1 exu_ecc_chk_rs3_U75(.A(exu_n20201), .B(exu_n20200), .Y(exu_n20196));
XOR2X1 exu_ecc_chk_rs3_U74(.A(exu_n20253), .B(exu_n20252), .Y(exu_n20197));
XOR2X1 exu_ecc_chk_rs3_U73(.A(exu_spu_rs3_data_e[10]), .B(exu_spu_rs3_data_e[9]), .Y(exu_n20198));
XOR2X1 exu_ecc_chk_rs3_U72(.A(exu_spu_rs3_data_e[25]), .B(exu_spu_rs3_data_e[24]), .Y(exu_n20199));
XOR2X1 exu_ecc_chk_rs3_U71(.A(exu_spu_rs3_data_e[40]), .B(exu_spu_rs3_data_e[39]), .Y(exu_n20200));
XOR2X1 exu_ecc_chk_rs3_U70(.A(exu_spu_rs3_data_e[56]), .B(exu_spu_rs3_data_e[55]), .Y(exu_n20201));
XOR2X1 exu_ecc_chk_rs3_U69(.A(exu_n20203), .B(exu_n20202), .Y(ecc_rs3_err_e[1]));
XOR2X1 exu_ecc_chk_rs3_U68(.A(exu_n20205), .B(exu_n20204), .Y(exu_n20202));
XOR2X1 exu_ecc_chk_rs3_U67(.A(exu_n20207), .B(exu_n20206), .Y(exu_n20203));
XOR2X1 exu_ecc_chk_rs3_U66(.A(exu_n20209), .B(exu_n20208), .Y(exu_n20204));
XOR2X1 exu_ecc_chk_rs3_U65(.A(exu_n20254), .B(exu_n20210), .Y(exu_n20205));
XOR2X1 exu_ecc_chk_rs3_U64(.A(exu_n20258), .B(exu_n20255), .Y(exu_n20206));
XOR2X1 exu_ecc_chk_rs3_U63(.A(exu_spu_rs3_data_e[6]), .B(exu_spu_rs3_data_e[5]), .Y(exu_n20207));
XOR2X1 exu_ecc_chk_rs3_U62(.A(exu_spu_rs3_data_e[21]), .B(exu_spu_rs3_data_e[20]), .Y(exu_n20208));
XOR2X1 exu_ecc_chk_rs3_U61(.A(exu_spu_rs3_data_e[36]), .B(exu_spu_rs3_data_e[35]), .Y(exu_n20209));
XOR2X1 exu_ecc_chk_rs3_U60(.A(exu_spu_rs3_data_e[52]), .B(exu_spu_rs3_data_e[51]), .Y(exu_n20210));
XOR2X1 exu_ecc_chk_rs3_U59(.A(exu_n20212), .B(exu_n20211), .Y(ecc_rs3_err_e[2]));
XOR2X1 exu_ecc_chk_rs3_U58(.A(exu_n20214), .B(exu_n20213), .Y(exu_n20211));
XOR2X1 exu_ecc_chk_rs3_U57(.A(exu_n20216), .B(exu_n20215), .Y(exu_n20212));
XOR2X1 exu_ecc_chk_rs3_U56(.A(exu_n20218), .B(exu_n20217), .Y(exu_n20213));
XOR2X1 exu_ecc_chk_rs3_U55(.A(exu_n20256), .B(exu_n20219), .Y(exu_n20214));
XOR2X1 exu_ecc_chk_rs3_U54(.A(exu_n20258), .B(exu_n20257), .Y(exu_n20215));
XOR2X1 exu_ecc_chk_rs3_U53(.A(exu_spu_rs3_data_e[8]), .B(exu_spu_rs3_data_e[7]), .Y(exu_n20216));
XOR2X1 exu_ecc_chk_rs3_U52(.A(exu_spu_rs3_data_e[23]), .B(exu_spu_rs3_data_e[22]), .Y(exu_n20217));
XOR2X1 exu_ecc_chk_rs3_U51(.A(exu_spu_rs3_data_e[38]), .B(exu_spu_rs3_data_e[37]), .Y(exu_n20218));
XOR2X1 exu_ecc_chk_rs3_U50(.A(exu_spu_rs3_data_e[54]), .B(exu_spu_rs3_data_e[53]), .Y(exu_n20219));
XOR2X1 exu_ecc_chk_rs3_U49(.A(exu_n20260), .B(exu_n20259), .Y(ecc_rs3_err_e[3]));
XOR2X1 exu_ecc_chk_rs3_U48(.A(exu_n20221), .B(exu_n20220), .Y(exu_n20267));
XOR2X1 exu_ecc_chk_rs3_U47(.A(exu_n20223), .B(exu_n20222), .Y(exu_n20220));
XOR2X1 exu_ecc_chk_rs3_U46(.A(exu_n20225), .B(exu_n20224), .Y(exu_n20221));
XOR2X1 exu_ecc_chk_rs3_U45(.A(exu_n20227), .B(exu_n20226), .Y(exu_n20222));
XOR2X1 exu_ecc_chk_rs3_U44(.A(exu_n20262), .B(exu_n20261), .Y(exu_n20223));
XOR2X1 exu_ecc_chk_rs3_U43(.A(exu_spu_rs3_data_e[42]), .B(exu_spu_rs3_data_e[41]), .Y(exu_n20224));
XOR2X1 exu_ecc_chk_rs3_U42(.A(exu_spu_rs3_data_e[44]), .B(exu_spu_rs3_data_e[43]), .Y(exu_n20225));
XOR2X1 exu_ecc_chk_rs3_U41(.A(exu_spu_rs3_data_e[46]), .B(exu_spu_rs3_data_e[45]), .Y(exu_n20226));
XOR2X1 exu_ecc_chk_rs3_U40(.A(exu_spu_rs3_data_e[48]), .B(exu_spu_rs3_data_e[47]), .Y(exu_n20227));
XOR2X1 exu_ecc_chk_rs3_U39(.A(exu_n20229), .B(exu_n20228), .Y(ecc_rs3_err_e[4]));
XOR2X1 exu_ecc_chk_rs3_U38(.A(exu_n20231), .B(exu_n20230), .Y(exu_n20228));
XOR2X1 exu_ecc_chk_rs3_U37(.A(exu_n20233), .B(exu_n20232), .Y(exu_n20229));
XOR2X1 exu_ecc_chk_rs3_U36(.A(exu_n20235), .B(exu_n20234), .Y(exu_n20230));
XOR2X1 exu_ecc_chk_rs3_U35(.A(exu_n20263), .B(exu_n20236), .Y(exu_n20231));
XOR2X1 exu_ecc_chk_rs3_U34(.A(exu_n20267), .B(exu_n20264), .Y(exu_n20232));
XOR2X1 exu_ecc_chk_rs3_U33(.A(exu_spu_rs3_data_e[11]), .B(ecc_rs3_ecc_e[4]), .Y(exu_n20233));
XOR2X1 exu_ecc_chk_rs3_U32(.A(exu_spu_rs3_data_e[13]), .B(exu_spu_rs3_data_e[12]), .Y(exu_n20234));
XOR2X1 exu_ecc_chk_rs3_U31(.A(exu_spu_rs3_data_e[15]), .B(exu_spu_rs3_data_e[14]), .Y(exu_n20235));
XOR2X1 exu_ecc_chk_rs3_U30(.A(exu_spu_rs3_data_e[17]), .B(exu_spu_rs3_data_e[16]), .Y(exu_n20236));
XOR2X1 exu_ecc_chk_rs3_U29(.A(exu_n20238), .B(exu_n20237), .Y(ecc_rs3_err_e[5]));
XOR2X1 exu_ecc_chk_rs3_U28(.A(exu_n20240), .B(exu_n20239), .Y(exu_n20237));
XOR2X1 exu_ecc_chk_rs3_U27(.A(exu_n20242), .B(exu_n20241), .Y(exu_n20238));
XOR2X1 exu_ecc_chk_rs3_U26(.A(exu_n20244), .B(exu_n20243), .Y(exu_n20239));
XOR2X1 exu_ecc_chk_rs3_U25(.A(exu_n20265), .B(exu_n20245), .Y(exu_n20240));
XOR2X1 exu_ecc_chk_rs3_U24(.A(exu_n20267), .B(exu_n20266), .Y(exu_n20241));
XOR2X1 exu_ecc_chk_rs3_U23(.A(exu_spu_rs3_data_e[26]), .B(ecc_rs3_ecc_e[5]), .Y(exu_n20242));
XOR2X1 exu_ecc_chk_rs3_U22(.A(exu_spu_rs3_data_e[28]), .B(exu_spu_rs3_data_e[27]), .Y(exu_n20243));
XOR2X1 exu_ecc_chk_rs3_U21(.A(exu_spu_rs3_data_e[30]), .B(exu_spu_rs3_data_e[29]), .Y(exu_n20244));
XOR2X1 exu_ecc_chk_rs3_U20(.A(exu_spu_rs3_data_e[32]), .B(exu_spu_rs3_data_e[31]), .Y(exu_n20245));
XOR2X1 exu_ecc_chk_rs3_U19(.A(exu_n20247), .B(exu_n20246), .Y(ecc_rs3_err_e[6]));
XOR2X1 exu_ecc_chk_rs3_U18(.A(exu_n20249), .B(exu_n20248), .Y(exu_n20246));
XOR2X1 exu_ecc_chk_rs3_U17(.A(exu_n20251), .B(exu_n20250), .Y(exu_n20247));
XOR2X1 exu_ecc_chk_rs3_U16(.A(exu_spu_rs3_data_e[57]), .B(ecc_rs3_ecc_e[6]), .Y(exu_n20248));
XOR2X1 exu_ecc_chk_rs3_U15(.A(exu_spu_rs3_data_e[59]), .B(exu_spu_rs3_data_e[58]), .Y(exu_n20249));
XOR2X1 exu_ecc_chk_rs3_U14(.A(exu_spu_rs3_data_e[61]), .B(exu_spu_rs3_data_e[60]), .Y(exu_n20250));
XOR2X1 exu_ecc_chk_rs3_U13(.A(exu_spu_rs3_data_e[63]), .B(exu_spu_rs3_data_e[62]), .Y(exu_n20251));
XOR2X1 exu_ecc_chk_rs2_U149(.A(exu_n20004), .B(exu_n20003), .Y(exu_n20126));
XOR2X1 exu_ecc_chk_rs2_U148(.A(div_input_data_e[116]), .B(div_input_data_e[114]), .Y(exu_n20003));
XOR2X1 exu_ecc_chk_rs2_U147(.A(div_input_data_e[120]), .B(div_input_data_e[118]), .Y(exu_n20004));
XOR2X1 exu_ecc_chk_rs2_U146(.A(exu_n20006), .B(exu_n20005), .Y(exu_n20130));
XOR2X1 exu_ecc_chk_rs2_U145(.A(div_input_data_e[100]), .B(div_input_data_e[98]), .Y(exu_n20005));
XOR2X1 exu_ecc_chk_rs2_U144(.A(div_input_data_e[104]), .B(div_input_data_e[102]), .Y(exu_n20006));
XOR2X1 exu_ecc_chk_rs2_U143(.A(exu_n20008), .B(exu_n20007), .Y(exu_n20128));
XOR2X1 exu_ecc_chk_rs2_U142(.A(div_input_data_e[85]), .B(div_input_data_e[83]), .Y(exu_n20007));
XOR2X1 exu_ecc_chk_rs2_U141(.A(div_input_data_e[89]), .B(div_input_data_e[87]), .Y(exu_n20008));
XOR2X1 exu_ecc_chk_rs2_U140(.A(exu_n20010), .B(exu_n20009), .Y(exu_n20124));
XOR2X1 exu_ecc_chk_rs2_U139(.A(exu_n20012), .B(exu_n20011), .Y(exu_n20009));
XOR2X1 exu_ecc_chk_rs2_U138(.A(exu_n20128), .B(exu_n20013), .Y(exu_n20010));
XOR2X1 exu_ecc_chk_rs2_U137(.A(exu_n20126), .B(exu_n20130), .Y(exu_n20011));
XOR2X1 exu_ecc_chk_rs2_U136(.A(div_input_data_e[70]), .B(div_input_data_e[68]), .Y(exu_n20012));
XOR2X1 exu_ecc_chk_rs2_U135(.A(div_input_data_e[74]), .B(div_input_data_e[72]), .Y(exu_n20013));
XOR2X1 exu_ecc_chk_rs2_U134(.A(exu_n20015), .B(exu_n20014), .Y(exu_n20117));
XOR2X1 exu_ecc_chk_rs2_U133(.A(div_input_data_e[67]), .B(exu_n20016), .Y(exu_n20014));
XOR2X1 exu_ecc_chk_rs2_U132(.A(div_input_data_e[96]), .B(div_input_data_e[81]), .Y(exu_n20015));
XOR2X1 exu_ecc_chk_rs2_U131(.A(div_input_data_e[127]), .B(div_input_data_e[112]), .Y(exu_n20016));
XOR2X1 exu_ecc_chk_rs2_U130(.A(exu_n20018), .B(exu_n20017), .Y(exu_n20121));
XOR2X1 exu_ecc_chk_rs2_U129(.A(div_input_data_e[65]), .B(exu_n20019), .Y(exu_n20017));
XOR2X1 exu_ecc_chk_rs2_U128(.A(div_input_data_e[94]), .B(div_input_data_e[79]), .Y(exu_n20018));
XOR2X1 exu_ecc_chk_rs2_U127(.A(div_input_data_e[125]), .B(div_input_data_e[110]), .Y(exu_n20019));
XOR2X1 exu_ecc_chk_rs2_U126(.A(exu_n20021), .B(exu_n20020), .Y(exu_n20119));
XOR2X1 exu_ecc_chk_rs2_U125(.A(div_input_data_e[64]), .B(exu_n20022), .Y(exu_n20020));
XOR2X1 exu_ecc_chk_rs2_U124(.A(div_input_data_e[92]), .B(div_input_data_e[77]), .Y(exu_n20021));
XOR2X1 exu_ecc_chk_rs2_U123(.A(div_input_data_e[123]), .B(div_input_data_e[108]), .Y(exu_n20022));
XOR2X1 exu_ecc_chk_rs2_U122(.A(exu_n20024), .B(exu_n20023), .Y(ecc_rs2_err_e[0]));
XOR2X1 exu_ecc_chk_rs2_U121(.A(exu_n20026), .B(exu_n20025), .Y(exu_n20023));
XOR2X1 exu_ecc_chk_rs2_U120(.A(exu_n20028), .B(exu_n20027), .Y(exu_n20024));
XOR2X1 exu_ecc_chk_rs2_U119(.A(exu_n20119), .B(exu_n20029), .Y(exu_n20025));
XOR2X1 exu_ecc_chk_rs2_U118(.A(exu_n20117), .B(exu_n20121), .Y(exu_n20026));
XOR2X1 exu_ecc_chk_rs2_U117(.A(ecc_rs2_ecc_e[0]), .B(exu_n20124), .Y(exu_n20027));
XOR2X1 exu_ecc_chk_rs2_U116(.A(div_input_data_e[90]), .B(div_input_data_e[75]), .Y(exu_n20028));
XOR2X1 exu_ecc_chk_rs2_U115(.A(div_input_data_e[121]), .B(div_input_data_e[106]), .Y(exu_n20029));
XOR2X1 exu_ecc_chk_rs2_U114(.A(exu_n20031), .B(exu_n20030), .Y(exu_n20125));
XOR2X1 exu_ecc_chk_rs2_U113(.A(div_input_data_e[115]), .B(div_input_data_e[113]), .Y(exu_n20030));
XOR2X1 exu_ecc_chk_rs2_U112(.A(div_input_data_e[119]), .B(div_input_data_e[117]), .Y(exu_n20031));
XOR2X1 exu_ecc_chk_rs2_U111(.A(exu_n20033), .B(exu_n20032), .Y(exu_n20129));
XOR2X1 exu_ecc_chk_rs2_U110(.A(div_input_data_e[99]), .B(div_input_data_e[97]), .Y(exu_n20032));
XOR2X1 exu_ecc_chk_rs2_U109(.A(div_input_data_e[103]), .B(div_input_data_e[101]), .Y(exu_n20033));
XOR2X1 exu_ecc_chk_rs2_U108(.A(exu_n20035), .B(exu_n20034), .Y(exu_n20127));
XOR2X1 exu_ecc_chk_rs2_U107(.A(div_input_data_e[84]), .B(div_input_data_e[82]), .Y(exu_n20034));
XOR2X1 exu_ecc_chk_rs2_U106(.A(div_input_data_e[88]), .B(div_input_data_e[86]), .Y(exu_n20035));
XOR2X1 exu_ecc_chk_rs2_U105(.A(exu_n20037), .B(exu_n20036), .Y(exu_n20123));
XOR2X1 exu_ecc_chk_rs2_U104(.A(exu_n20039), .B(exu_n20038), .Y(exu_n20036));
XOR2X1 exu_ecc_chk_rs2_U103(.A(exu_n20127), .B(exu_n20040), .Y(exu_n20037));
XOR2X1 exu_ecc_chk_rs2_U102(.A(exu_n20125), .B(exu_n20129), .Y(exu_n20038));
XOR2X1 exu_ecc_chk_rs2_U101(.A(div_input_data_e[69]), .B(ecc_rs2_ecc_e[3]), .Y(exu_n20039));
XOR2X1 exu_ecc_chk_rs2_U100(.A(div_input_data_e[73]), .B(div_input_data_e[71]), .Y(exu_n20040));
XOR2X1 exu_ecc_chk_rs2_U99(.A(exu_n20042), .B(exu_n20041), .Y(exu_n20116));
XOR2X1 exu_ecc_chk_rs2_U98(.A(div_input_data_e[66]), .B(exu_n20043), .Y(exu_n20041));
XOR2X1 exu_ecc_chk_rs2_U97(.A(div_input_data_e[95]), .B(div_input_data_e[80]), .Y(exu_n20042));
XOR2X1 exu_ecc_chk_rs2_U96(.A(div_input_data_e[126]), .B(div_input_data_e[111]), .Y(exu_n20043));
XOR2X1 exu_ecc_chk_rs2_U95(.A(exu_n20045), .B(exu_n20044), .Y(exu_n20120));
XOR2X1 exu_ecc_chk_rs2_U94(.A(ecc_rs2_ecc_e[2]), .B(exu_n20046), .Y(exu_n20044));
XOR2X1 exu_ecc_chk_rs2_U93(.A(div_input_data_e[93]), .B(div_input_data_e[78]), .Y(exu_n20045));
XOR2X1 exu_ecc_chk_rs2_U92(.A(div_input_data_e[124]), .B(div_input_data_e[109]), .Y(exu_n20046));
XOR2X1 exu_ecc_chk_rs2_U91(.A(exu_n20048), .B(exu_n20047), .Y(exu_n20118));
XOR2X1 exu_ecc_chk_rs2_U90(.A(ecc_rs2_ecc_e[1]), .B(exu_n20049), .Y(exu_n20047));
XOR2X1 exu_ecc_chk_rs2_U89(.A(div_input_data_e[91]), .B(div_input_data_e[76]), .Y(exu_n20048));
XOR2X1 exu_ecc_chk_rs2_U88(.A(div_input_data_e[122]), .B(div_input_data_e[107]), .Y(exu_n20049));
XOR2X1 exu_ecc_chk_rs2_U87(.A(exu_n20051), .B(exu_n20050), .Y(ecc_chk_rs2_parity));
XOR2X1 exu_ecc_chk_rs2_U86(.A(exu_n20053), .B(exu_n20052), .Y(exu_n20050));
XOR2X1 exu_ecc_chk_rs2_U85(.A(exu_n20055), .B(exu_n20054), .Y(exu_n20051));
XOR2X1 exu_ecc_chk_rs2_U84(.A(exu_n20057), .B(exu_n20056), .Y(exu_n20052));
XOR2X1 exu_ecc_chk_rs2_U83(.A(exu_n20120), .B(exu_n20118), .Y(exu_n20053));
XOR2X1 exu_ecc_chk_rs2_U82(.A(exu_n20123), .B(exu_n20116), .Y(exu_n20054));
XOR2X1 exu_ecc_chk_rs2_U81(.A(ecc_rs2_ecc_e[4]), .B(ecc_rs2_err_e[0]), .Y(exu_n20055));
XOR2X1 exu_ecc_chk_rs2_U80(.A(ecc_rs2_ecc_e[6]), .B(ecc_rs2_ecc_e[5]), .Y(exu_n20056));
XOR2X1 exu_ecc_chk_rs2_U79(.A(div_input_data_e[105]), .B(ecc_rs2_ecc_e[7]), .Y(exu_n20057));
XOR2X1 exu_ecc_chk_rs2_U78(.A(exu_n20059), .B(exu_n20058), .Y(exu_n20122));
XOR2X1 exu_ecc_chk_rs2_U77(.A(exu_n20061), .B(exu_n20060), .Y(exu_n20058));
XOR2X1 exu_ecc_chk_rs2_U76(.A(exu_n20063), .B(exu_n20062), .Y(exu_n20059));
XOR2X1 exu_ecc_chk_rs2_U75(.A(exu_n20065), .B(exu_n20064), .Y(exu_n20060));
XOR2X1 exu_ecc_chk_rs2_U74(.A(exu_n20117), .B(exu_n20116), .Y(exu_n20061));
XOR2X1 exu_ecc_chk_rs2_U73(.A(div_input_data_e[74]), .B(div_input_data_e[73]), .Y(exu_n20062));
XOR2X1 exu_ecc_chk_rs2_U72(.A(div_input_data_e[89]), .B(div_input_data_e[88]), .Y(exu_n20063));
XOR2X1 exu_ecc_chk_rs2_U71(.A(div_input_data_e[104]), .B(div_input_data_e[103]), .Y(exu_n20064));
XOR2X1 exu_ecc_chk_rs2_U70(.A(div_input_data_e[120]), .B(div_input_data_e[119]), .Y(exu_n20065));
XOR2X1 exu_ecc_chk_rs2_U69(.A(exu_n20067), .B(exu_n20066), .Y(ecc_rs2_err_e[1]));
XOR2X1 exu_ecc_chk_rs2_U68(.A(exu_n20069), .B(exu_n20068), .Y(exu_n20066));
XOR2X1 exu_ecc_chk_rs2_U67(.A(exu_n20071), .B(exu_n20070), .Y(exu_n20067));
XOR2X1 exu_ecc_chk_rs2_U66(.A(exu_n20073), .B(exu_n20072), .Y(exu_n20068));
XOR2X1 exu_ecc_chk_rs2_U65(.A(exu_n20118), .B(exu_n20074), .Y(exu_n20069));
XOR2X1 exu_ecc_chk_rs2_U64(.A(exu_n20122), .B(exu_n20119), .Y(exu_n20070));
XOR2X1 exu_ecc_chk_rs2_U63(.A(div_input_data_e[70]), .B(div_input_data_e[69]), .Y(exu_n20071));
XOR2X1 exu_ecc_chk_rs2_U62(.A(div_input_data_e[85]), .B(div_input_data_e[84]), .Y(exu_n20072));
XOR2X1 exu_ecc_chk_rs2_U61(.A(div_input_data_e[100]), .B(div_input_data_e[99]), .Y(exu_n20073));
XOR2X1 exu_ecc_chk_rs2_U60(.A(div_input_data_e[116]), .B(div_input_data_e[115]), .Y(exu_n20074));
XOR2X1 exu_ecc_chk_rs2_U59(.A(exu_n20076), .B(exu_n20075), .Y(ecc_rs2_err_e[2]));
XOR2X1 exu_ecc_chk_rs2_U58(.A(exu_n20078), .B(exu_n20077), .Y(exu_n20075));
XOR2X1 exu_ecc_chk_rs2_U57(.A(exu_n20080), .B(exu_n20079), .Y(exu_n20076));
XOR2X1 exu_ecc_chk_rs2_U56(.A(exu_n20082), .B(exu_n20081), .Y(exu_n20077));
XOR2X1 exu_ecc_chk_rs2_U55(.A(exu_n20120), .B(exu_n20083), .Y(exu_n20078));
XOR2X1 exu_ecc_chk_rs2_U54(.A(exu_n20122), .B(exu_n20121), .Y(exu_n20079));
XOR2X1 exu_ecc_chk_rs2_U53(.A(div_input_data_e[72]), .B(div_input_data_e[71]), .Y(exu_n20080));
XOR2X1 exu_ecc_chk_rs2_U52(.A(div_input_data_e[87]), .B(div_input_data_e[86]), .Y(exu_n20081));
XOR2X1 exu_ecc_chk_rs2_U51(.A(div_input_data_e[102]), .B(div_input_data_e[101]), .Y(exu_n20082));
XOR2X1 exu_ecc_chk_rs2_U50(.A(div_input_data_e[118]), .B(div_input_data_e[117]), .Y(exu_n20083));
XOR2X1 exu_ecc_chk_rs2_U49(.A(exu_n20124), .B(exu_n20123), .Y(ecc_rs2_err_e[3]));
XOR2X1 exu_ecc_chk_rs2_U48(.A(exu_n20085), .B(exu_n20084), .Y(exu_n20131));
XOR2X1 exu_ecc_chk_rs2_U47(.A(exu_n20087), .B(exu_n20086), .Y(exu_n20084));
XOR2X1 exu_ecc_chk_rs2_U46(.A(exu_n20089), .B(exu_n20088), .Y(exu_n20085));
XOR2X1 exu_ecc_chk_rs2_U45(.A(exu_n20091), .B(exu_n20090), .Y(exu_n20086));
XOR2X1 exu_ecc_chk_rs2_U44(.A(exu_n20126), .B(exu_n20125), .Y(exu_n20087));
XOR2X1 exu_ecc_chk_rs2_U43(.A(div_input_data_e[106]), .B(div_input_data_e[105]), .Y(exu_n20088));
XOR2X1 exu_ecc_chk_rs2_U42(.A(div_input_data_e[108]), .B(div_input_data_e[107]), .Y(exu_n20089));
XOR2X1 exu_ecc_chk_rs2_U41(.A(div_input_data_e[110]), .B(div_input_data_e[109]), .Y(exu_n20090));
XOR2X1 exu_ecc_chk_rs2_U40(.A(div_input_data_e[112]), .B(div_input_data_e[111]), .Y(exu_n20091));
XOR2X1 exu_ecc_chk_rs2_U39(.A(exu_n20093), .B(exu_n20092), .Y(ecc_rs2_err_e[4]));
XOR2X1 exu_ecc_chk_rs2_U38(.A(exu_n20095), .B(exu_n20094), .Y(exu_n20092));
XOR2X1 exu_ecc_chk_rs2_U37(.A(exu_n20097), .B(exu_n20096), .Y(exu_n20093));
XOR2X1 exu_ecc_chk_rs2_U36(.A(exu_n20099), .B(exu_n20098), .Y(exu_n20094));
XOR2X1 exu_ecc_chk_rs2_U35(.A(exu_n20127), .B(exu_n20100), .Y(exu_n20095));
XOR2X1 exu_ecc_chk_rs2_U34(.A(exu_n20131), .B(exu_n20128), .Y(exu_n20096));
XOR2X1 exu_ecc_chk_rs2_U33(.A(div_input_data_e[75]), .B(ecc_rs2_ecc_e[4]), .Y(exu_n20097));
XOR2X1 exu_ecc_chk_rs2_U32(.A(div_input_data_e[77]), .B(div_input_data_e[76]), .Y(exu_n20098));
XOR2X1 exu_ecc_chk_rs2_U31(.A(div_input_data_e[79]), .B(div_input_data_e[78]), .Y(exu_n20099));
XOR2X1 exu_ecc_chk_rs2_U30(.A(div_input_data_e[81]), .B(div_input_data_e[80]), .Y(exu_n20100));
XOR2X1 exu_ecc_chk_rs2_U29(.A(exu_n20102), .B(exu_n20101), .Y(ecc_rs2_err_e[5]));
XOR2X1 exu_ecc_chk_rs2_U28(.A(exu_n20104), .B(exu_n20103), .Y(exu_n20101));
XOR2X1 exu_ecc_chk_rs2_U27(.A(exu_n20106), .B(exu_n20105), .Y(exu_n20102));
XOR2X1 exu_ecc_chk_rs2_U26(.A(exu_n20108), .B(exu_n20107), .Y(exu_n20103));
XOR2X1 exu_ecc_chk_rs2_U25(.A(exu_n20129), .B(exu_n20109), .Y(exu_n20104));
XOR2X1 exu_ecc_chk_rs2_U24(.A(exu_n20131), .B(exu_n20130), .Y(exu_n20105));
XOR2X1 exu_ecc_chk_rs2_U23(.A(div_input_data_e[90]), .B(ecc_rs2_ecc_e[5]), .Y(exu_n20106));
XOR2X1 exu_ecc_chk_rs2_U22(.A(div_input_data_e[92]), .B(div_input_data_e[91]), .Y(exu_n20107));
XOR2X1 exu_ecc_chk_rs2_U21(.A(div_input_data_e[94]), .B(div_input_data_e[93]), .Y(exu_n20108));
XOR2X1 exu_ecc_chk_rs2_U20(.A(div_input_data_e[96]), .B(div_input_data_e[95]), .Y(exu_n20109));
XOR2X1 exu_ecc_chk_rs2_U19(.A(exu_n20111), .B(exu_n20110), .Y(ecc_rs2_err_e[6]));
XOR2X1 exu_ecc_chk_rs2_U18(.A(exu_n20113), .B(exu_n20112), .Y(exu_n20110));
XOR2X1 exu_ecc_chk_rs2_U17(.A(exu_n20115), .B(exu_n20114), .Y(exu_n20111));
XOR2X1 exu_ecc_chk_rs2_U16(.A(div_input_data_e[121]), .B(ecc_rs2_ecc_e[6]), .Y(exu_n20112));
XOR2X1 exu_ecc_chk_rs2_U15(.A(div_input_data_e[123]), .B(div_input_data_e[122]), .Y(exu_n20113));
XOR2X1 exu_ecc_chk_rs2_U14(.A(div_input_data_e[125]), .B(div_input_data_e[124]), .Y(exu_n20114));
XOR2X1 exu_ecc_chk_rs2_U13(.A(div_input_data_e[127]), .B(div_input_data_e[126]), .Y(exu_n20115));
DFFPOSX1 rml_cwp_spill_dff_q_reg[0](.D(exu_n19995), .CLK(rclk), .Q(exu_tlu_spill_wtype[0]));
DFFPOSX1 rml_cwp_spill_dff_q_reg[1](.D(exu_n19994), .CLK(rclk), .Q(exu_tlu_spill_wtype[1]));
DFFPOSX1 rml_cwp_spill_dff_q_reg[2](.D(exu_n19993), .CLK(rclk), .Q(exu_tlu_spill_wtype[2]));
DFFPOSX1 rml_cwp_spill_dff_q_reg[3](.D(exu_n19992), .CLK(rclk), .Q(exu_tlu_spill_other));
DFFPOSX1 rml_cwp_spill_dff_q_reg[4](.D(exu_n18420), .CLK(rclk), .Q(exu_tlu_spill_tid[0]));
DFFPOSX1 rml_cwp_spill_dff_q_reg[5](.D(exu_n18419), .CLK(rclk), .Q(exu_tlu_spill_tid[1]));
DFFPOSX1 rml_cwp_spill_dff_q_reg[6](.D(exu_n19991), .CLK(rclk), .Q(exu_tlu_spill));
DFFPOSX1 ecl_writeback_dff_sraddr_m2w_q_reg[0](.D(exu_n19989), .CLK(rclk), .Q(ecl_writeback_sraddr_w[0]));
DFFPOSX1 ecl_writeback_dff_sraddr_m2w_q_reg[1](.D(exu_n19988), .CLK(rclk), .Q(ecl_writeback_sraddr_w[1]));
DFFPOSX1 ecl_writeback_dff_sraddr_m2w_q_reg[2](.D(exu_n19987), .CLK(rclk), .Q(ecl_writeback_sraddr_w[2]));
DFFPOSX1 ecl_writeback_dff_sraddr_m2w_q_reg[3](.D(exu_n19986), .CLK(rclk), .Q(ecl_writeback_sraddr_w[3]));
DFFPOSX1 ecl_writeback_dff_sraddr_m2w_q_reg[4](.D(exu_n19985), .CLK(rclk), .Q(ecl_writeback_sraddr_w[4]));
DFFPOSX1 ecl_writeback_dff_sraddr_m2w_q_reg[5](.D(exu_n19984), .CLK(rclk), .Q(ecl_writeback_sraddr_w[5]));
DFFPOSX1 ecl_writeback_dff_sraddr_m2w_q_reg[6](.D(exu_n19983), .CLK(rclk), .Q(ecl_writeback_sraddr_w[6]));
DFFPOSX1 ecl_writeback_dff_sraddr_e2m_q_reg[0](.D(exu_n19981), .CLK(rclk), .Q(ecl_writeback_sraddr_m[0]));
DFFPOSX1 ecl_writeback_dff_sraddr_e2m_q_reg[1](.D(exu_n19980), .CLK(rclk), .Q(ecl_writeback_sraddr_m[1]));
DFFPOSX1 ecl_writeback_dff_sraddr_e2m_q_reg[2](.D(exu_n19979), .CLK(rclk), .Q(ecl_writeback_sraddr_m[2]));
DFFPOSX1 ecl_writeback_dff_sraddr_e2m_q_reg[3](.D(exu_n19978), .CLK(rclk), .Q(ecl_writeback_sraddr_m[3]));
DFFPOSX1 ecl_writeback_dff_sraddr_e2m_q_reg[4](.D(exu_n19977), .CLK(rclk), .Q(ecl_writeback_sraddr_m[4]));
DFFPOSX1 ecl_writeback_dff_sraddr_e2m_q_reg[5](.D(exu_n19976), .CLK(rclk), .Q(ecl_writeback_sraddr_m[5]));
DFFPOSX1 ecl_writeback_dff_sraddr_e2m_q_reg[6](.D(exu_n19975), .CLK(rclk), .Q(ecl_writeback_sraddr_m[6]));
DFFPOSX1 ecl_writeback_dff_sraddr_d2e_q_reg[0](.D(exu_n19973), .CLK(rclk), .Q(ecl_writeback_sraddr_e[0]));
DFFPOSX1 ecl_writeback_dff_sraddr_d2e_q_reg[1](.D(exu_n19972), .CLK(rclk), .Q(ecl_writeback_sraddr_e[1]));
DFFPOSX1 ecl_writeback_dff_sraddr_d2e_q_reg[2](.D(exu_n19971), .CLK(rclk), .Q(ecl_writeback_sraddr_e[2]));
DFFPOSX1 ecl_writeback_dff_sraddr_d2e_q_reg[3](.D(exu_n19970), .CLK(rclk), .Q(ecl_writeback_sraddr_e[3]));
DFFPOSX1 ecl_writeback_dff_sraddr_d2e_q_reg[4](.D(exu_n19969), .CLK(rclk), .Q(ecl_writeback_sraddr_e[4]));
DFFPOSX1 ecl_writeback_dff_sraddr_d2e_q_reg[5](.D(exu_n19968), .CLK(rclk), .Q(ecl_writeback_sraddr_e[5]));
DFFPOSX1 ecl_writeback_dff_sraddr_d2e_q_reg[6](.D(exu_n19967), .CLK(rclk), .Q(ecl_writeback_sraddr_e[6]));
DFFPOSX1 ecc_rs3o_err_e2m_q_reg[0](.D(exu_n19965), .CLK(rclk), .Q(ecc_rs3_err_m[0]));
DFFPOSX1 ecc_rs3o_err_e2m_q_reg[1](.D(exu_n19964), .CLK(rclk), .Q(ecc_rs3_err_m[1]));
DFFPOSX1 ecc_rs3o_err_e2m_q_reg[2](.D(exu_n19963), .CLK(rclk), .Q(ecc_rs3_err_m[2]));
DFFPOSX1 ecc_rs3o_err_e2m_q_reg[3](.D(exu_n19962), .CLK(rclk), .Q(ecc_rs3_err_m[3]));
DFFPOSX1 ecc_rs3o_err_e2m_q_reg[4](.D(exu_n19961), .CLK(rclk), .Q(ecc_rs3_err_m[4]));
DFFPOSX1 ecc_rs3o_err_e2m_q_reg[5](.D(exu_n19960), .CLK(rclk), .Q(ecc_rs3_err_m[5]));
DFFPOSX1 ecc_rs3o_err_e2m_q_reg[6](.D(exu_n19959), .CLK(rclk), .Q(ecc_rs3_err_m[6]));
DFFPOSX1 ecc_rs2_err_e2m_q_reg[0](.D(exu_n19957), .CLK(rclk), .Q(ecc_rs2_err_m[0]));
DFFPOSX1 ecc_rs2_err_e2m_q_reg[1](.D(exu_n19956), .CLK(rclk), .Q(ecc_rs2_err_m[1]));
DFFPOSX1 ecc_rs2_err_e2m_q_reg[2](.D(exu_n19955), .CLK(rclk), .Q(ecc_rs2_err_m[2]));
DFFPOSX1 ecc_rs2_err_e2m_q_reg[3](.D(exu_n19954), .CLK(rclk), .Q(ecc_rs2_err_m[3]));
DFFPOSX1 ecc_rs2_err_e2m_q_reg[4](.D(exu_n19953), .CLK(rclk), .Q(ecc_rs2_err_m[4]));
DFFPOSX1 ecc_rs2_err_e2m_q_reg[5](.D(exu_n19952), .CLK(rclk), .Q(ecc_rs2_err_m[5]));
DFFPOSX1 ecc_rs2_err_e2m_q_reg[6](.D(exu_n19951), .CLK(rclk), .Q(ecc_rs2_err_m[6]));
NAND2X1 exu_ecc_syn_log_mux_U32(.A(exu_n19946), .B(exu_n9998), .Y(exu_ifu_err_synd_m[0]));
NAND2X1 exu_ecc_syn_log_mux_U28(.A(exu_n19942), .B(exu_n9997), .Y(exu_ifu_err_synd_m[1]));
NAND2X1 exu_ecc_syn_log_mux_U24(.A(exu_n19938), .B(exu_n9996), .Y(exu_ifu_err_synd_m[2]));
NAND2X1 exu_ecc_syn_log_mux_U20(.A(exu_n19934), .B(exu_n9995), .Y(exu_ifu_err_synd_m[3]));
NAND2X1 exu_ecc_syn_log_mux_U16(.A(exu_n19930), .B(exu_n9994), .Y(exu_ifu_err_synd_m[4]));
NAND2X1 exu_ecc_syn_log_mux_U12(.A(exu_n19926), .B(exu_n9993), .Y(exu_ifu_err_synd_m[5]));
NAND2X1 exu_ecc_syn_log_mux_U8(.A(exu_n19922), .B(exu_n9992), .Y(exu_ifu_err_synd_m[6]));
DFFSR rml_rstff_q_reg[0](.D(exu_n19921), .CLK(rclk), .Q(rml_rml_reset_l));
DFFPOSX1 rml_cwp_tlu_data_dff_q_reg[0](.D(exu_n19919), .CLK(rclk), .Q(rml_cwp_tlu_swap_data[12]));
DFFPOSX1 rml_cwp_tlu_data_dff_q_reg[1](.D(exu_n19918), .CLK(rclk), .Q(rml_cwp_tlu_exu_cwp_w[0]));
DFFPOSX1 rml_cwp_tlu_data_dff_q_reg[2](.D(exu_n19917), .CLK(rclk), .Q(rml_cwp_tlu_exu_cwp_w[1]));
DFFPOSX1 rml_cwp_tlu_data_dff_q_reg[3](.D(exu_n19916), .CLK(rclk), .Q(rml_cwp_tlu_exu_cwp_w[2]));
DFFPOSX1 rml_cwp_tlu_data_dff_q_reg[4](.D(exu_n19915), .CLK(rclk), .Q(rml_cwp_cwpccr_update_w));
DFFPOSX1 ecl_divcntl_cc_sig_dff_q_reg[0](.D(exu_n19913), .CLK(rclk), .Q(ecl_divcntl_low32_nonzero_d1));
DFFPOSX1 ecl_divcntl_cc_sig_dff_q_reg[1](.D(exu_n19912), .CLK(rclk), .Q(ecl_divcntl_sel_div_d1));
DFFPOSX1 ecl_divcntl_cc_sig_dff_q_reg[2](.D(exu_n19911), .CLK(rclk), .Q(ecl_divcntl_gencc_in_31_d1));
DFFPOSX1 ecl_divcntl_cc_sig_dff_q_reg[3](.D(exu_n19910), .CLK(rclk), .Q(ecl_divcntl_gencc_in_msb_l_d1));
DFFPOSX1 ecl_divcntl_cc_sig_dff_q_reg[4](.D(exu_n19909), .CLK(rclk), .Q(ecl_divcntl_upper32_equal_d1));
DFFPOSX1 ecl_writeback_dff_rd_g2w2_q_reg[0](.D(exu_n19907), .CLK(rclk), .Q(ecl_wb_byplog_rd_w2[0]));
DFFPOSX1 ecl_writeback_dff_rd_g2w2_q_reg[1](.D(exu_n19906), .CLK(rclk), .Q(ecl_wb_byplog_rd_w2[1]));
DFFPOSX1 ecl_writeback_dff_rd_g2w2_q_reg[2](.D(exu_n19905), .CLK(rclk), .Q(ecl_wb_byplog_rd_w2[2]));
DFFPOSX1 ecl_writeback_dff_rd_g2w2_q_reg[3](.D(exu_n19904), .CLK(rclk), .Q(ecl_wb_byplog_rd_w2[3]));
DFFPOSX1 ecl_writeback_dff_rd_g2w2_q_reg[4](.D(exu_n19903), .CLK(rclk), .Q(ecl_wb_byplog_rd_w2[4]));
DFFPOSX1 ecl_writeback_dfill_rd_dff_q_reg[0](.D(exu_n19901), .CLK(rclk), .Q(ecl_wb_byplog_rd_g2[0]));
DFFPOSX1 ecl_writeback_dfill_rd_dff_q_reg[1](.D(exu_n19900), .CLK(rclk), .Q(ecl_wb_byplog_rd_g2[1]));
DFFPOSX1 ecl_writeback_dfill_rd_dff_q_reg[2](.D(exu_n19899), .CLK(rclk), .Q(ecl_wb_byplog_rd_g2[2]));
DFFPOSX1 ecl_writeback_dfill_rd_dff_q_reg[3](.D(exu_n19898), .CLK(rclk), .Q(ecl_wb_byplog_rd_g2[3]));
DFFPOSX1 ecl_writeback_dfill_rd_dff_q_reg[4](.D(exu_n19897), .CLK(rclk), .Q(ecl_wb_byplog_rd_g2[4]));
DFFPOSX1 ecl_dff_rd_m2w_q_reg[0](.D(exu_n19895), .CLK(rclk), .Q(ecl_ecl_irf_rd_w[0]));
DFFPOSX1 ecl_dff_rd_m2w_q_reg[1](.D(exu_n19894), .CLK(rclk), .Q(ecl_ecl_irf_rd_w[1]));
DFFPOSX1 ecl_dff_rd_m2w_q_reg[2](.D(exu_n19893), .CLK(rclk), .Q(ecl_ecl_irf_rd_w[2]));
DFFPOSX1 ecl_dff_rd_m2w_q_reg[3](.D(exu_n19892), .CLK(rclk), .Q(ecl_ecl_irf_rd_w[3]));
DFFPOSX1 ecl_dff_rd_m2w_q_reg[4](.D(exu_n19891), .CLK(rclk), .Q(ecl_ecl_irf_rd_w[4]));
DFFPOSX1 ecl_dff_rd_e2m_q_reg[0](.D(exu_n19889), .CLK(rclk), .Q(ecl_rd_m[0]));
DFFPOSX1 ecl_dff_rd_e2m_q_reg[1](.D(exu_n19888), .CLK(rclk), .Q(ecl_rd_m[1]));
DFFPOSX1 ecl_dff_rd_e2m_q_reg[2](.D(exu_n19887), .CLK(rclk), .Q(ecl_rd_m[2]));
DFFPOSX1 ecl_dff_rd_e2m_q_reg[3](.D(exu_n19886), .CLK(rclk), .Q(ecl_rd_m[3]));
DFFPOSX1 ecl_dff_rd_e2m_q_reg[4](.D(exu_n19885), .CLK(rclk), .Q(ecl_rd_m[4]));
DFFPOSX1 ecl_dff_rd_d2e_q_reg[0](.D(exu_n19883), .CLK(rclk), .Q(ecl_rd_e[0]));
DFFPOSX1 ecl_dff_rd_d2e_q_reg[1](.D(exu_n19882), .CLK(rclk), .Q(ecl_rd_e[1]));
DFFPOSX1 ecl_dff_rd_d2e_q_reg[2](.D(exu_n19881), .CLK(rclk), .Q(ecl_rd_e[2]));
DFFPOSX1 ecl_dff_rd_d2e_q_reg[3](.D(exu_n19880), .CLK(rclk), .Q(ecl_rd_e[3]));
DFFPOSX1 ecl_dff_rd_d2e_q_reg[4](.D(exu_n19879), .CLK(rclk), .Q(ecl_rd_e[4]));
DFFPOSX1 ecl_dff_ld_rd_m2g_q_reg[0](.D(exu_n19877), .CLK(rclk), .Q(ecl_ld_rd_g[0]));
DFFPOSX1 ecl_dff_ld_rd_m2g_q_reg[1](.D(exu_n19876), .CLK(rclk), .Q(ecl_ld_rd_g[1]));
DFFPOSX1 ecl_dff_ld_rd_m2g_q_reg[2](.D(exu_n19875), .CLK(rclk), .Q(ecl_ld_rd_g[2]));
DFFPOSX1 ecl_dff_ld_rd_m2g_q_reg[3](.D(exu_n19874), .CLK(rclk), .Q(ecl_ld_rd_g[3]));
DFFPOSX1 ecl_dff_ld_rd_m2g_q_reg[4](.D(exu_n19873), .CLK(rclk), .Q(ecl_ld_rd_g[4]));
DFFPOSX1 ecl_dff_rs3_e2m_q_reg[0](.D(exu_n19871), .CLK(rclk), .Q(ecl_ifu_exu_rs3_m[0]));
DFFPOSX1 ecl_dff_rs3_e2m_q_reg[1](.D(exu_n19870), .CLK(rclk), .Q(ecl_ifu_exu_rs3_m[1]));
DFFPOSX1 ecl_dff_rs3_e2m_q_reg[2](.D(exu_n19869), .CLK(rclk), .Q(ecl_ifu_exu_rs3_m[2]));
DFFPOSX1 ecl_dff_rs3_e2m_q_reg[3](.D(exu_n19868), .CLK(rclk), .Q(ecl_ifu_exu_rs3_m[3]));
DFFPOSX1 ecl_dff_rs3_e2m_q_reg[4](.D(exu_n19867), .CLK(rclk), .Q(ecl_ifu_exu_rs3_m[4]));
DFFPOSX1 ecl_dff_rs2_e2m_q_reg[0](.D(exu_n19865), .CLK(rclk), .Q(ecl_ifu_exu_rs2_m[0]));
DFFPOSX1 ecl_dff_rs2_e2m_q_reg[1](.D(exu_n19864), .CLK(rclk), .Q(ecl_ifu_exu_rs2_m[1]));
DFFPOSX1 ecl_dff_rs2_e2m_q_reg[2](.D(exu_n19863), .CLK(rclk), .Q(ecl_ifu_exu_rs2_m[2]));
DFFPOSX1 ecl_dff_rs2_e2m_q_reg[3](.D(exu_n19862), .CLK(rclk), .Q(ecl_ifu_exu_rs2_m[3]));
DFFPOSX1 ecl_dff_rs2_e2m_q_reg[4](.D(exu_n19861), .CLK(rclk), .Q(ecl_ifu_exu_rs2_m[4]));
DFFPOSX1 ecl_dff_rs1_e2m_q_reg[0](.D(exu_n19859), .CLK(rclk), .Q(ecl_ifu_exu_rs1_m[0]));
DFFPOSX1 ecl_dff_rs1_e2m_q_reg[1](.D(exu_n19858), .CLK(rclk), .Q(ecl_ifu_exu_rs1_m[1]));
DFFPOSX1 ecl_dff_rs1_e2m_q_reg[2](.D(exu_n19857), .CLK(rclk), .Q(ecl_ifu_exu_rs1_m[2]));
DFFPOSX1 ecl_dff_rs1_e2m_q_reg[3](.D(exu_n19856), .CLK(rclk), .Q(ecl_ifu_exu_rs1_m[3]));
DFFPOSX1 ecl_dff_rs1_e2m_q_reg[4](.D(exu_n19855), .CLK(rclk), .Q(ecl_ifu_exu_rs1_m[4]));
DFFPOSX1 ecl_dff_rs3_d2e_q_reg[0](.D(exu_n19853), .CLK(rclk), .Q(ecl_ifu_exu_rs3_e[0]));
DFFPOSX1 ecl_dff_rs3_d2e_q_reg[1](.D(exu_n19852), .CLK(rclk), .Q(ecl_ifu_exu_rs3_e[1]));
DFFPOSX1 ecl_dff_rs3_d2e_q_reg[2](.D(exu_n19851), .CLK(rclk), .Q(ecl_ifu_exu_rs3_e[2]));
DFFPOSX1 ecl_dff_rs3_d2e_q_reg[3](.D(exu_n19850), .CLK(rclk), .Q(ecl_ifu_exu_rs3_e[3]));
DFFPOSX1 ecl_dff_rs3_d2e_q_reg[4](.D(exu_n19849), .CLK(rclk), .Q(ecl_ifu_exu_rs3_e[4]));
DFFPOSX1 ecl_dff_rs2_d2e_q_reg[0](.D(exu_n19847), .CLK(rclk), .Q(ecl_ifu_exu_rs2_e[0]));
DFFPOSX1 ecl_dff_rs2_d2e_q_reg[1](.D(exu_n19846), .CLK(rclk), .Q(ecl_ifu_exu_rs2_e[1]));
DFFPOSX1 ecl_dff_rs2_d2e_q_reg[2](.D(exu_n19845), .CLK(rclk), .Q(ecl_ifu_exu_rs2_e[2]));
DFFPOSX1 ecl_dff_rs2_d2e_q_reg[3](.D(exu_n19844), .CLK(rclk), .Q(ecl_ifu_exu_rs2_e[3]));
DFFPOSX1 ecl_dff_rs2_d2e_q_reg[4](.D(exu_n19843), .CLK(rclk), .Q(ecl_ifu_exu_rs2_e[4]));
DFFPOSX1 ecl_dff_rs1_d2e_q_reg[0](.D(exu_n19841), .CLK(rclk), .Q(ecl_ifu_exu_rs1_e[0]));
DFFPOSX1 ecl_dff_rs1_d2e_q_reg[1](.D(exu_n19840), .CLK(rclk), .Q(ecl_ifu_exu_rs1_e[1]));
DFFPOSX1 ecl_dff_rs1_d2e_q_reg[2](.D(exu_n19839), .CLK(rclk), .Q(ecl_ifu_exu_rs1_e[2]));
DFFPOSX1 ecl_dff_rs1_d2e_q_reg[3](.D(exu_n19838), .CLK(rclk), .Q(ecl_ifu_exu_rs1_e[3]));
DFFPOSX1 ecl_dff_rs1_d2e_q_reg[4](.D(exu_n19837), .CLK(rclk), .Q(ecl_ifu_exu_rs1_e[4]));
DFFPOSX1 ecl_dff_rs3_s2d_q_reg[0](.D(exu_n19835), .CLK(rclk), .Q(ecl_ifu_exu_rs3_d[0]));
DFFPOSX1 ecl_dff_rs3_s2d_q_reg[1](.D(exu_n19834), .CLK(rclk), .Q(ecl_ifu_exu_rs3_d[1]));
DFFPOSX1 ecl_dff_rs3_s2d_q_reg[2](.D(exu_n19833), .CLK(rclk), .Q(ecl_ifu_exu_rs3_d[2]));
DFFPOSX1 ecl_dff_rs3_s2d_q_reg[3](.D(exu_n19832), .CLK(rclk), .Q(ecl_ifu_exu_rs3_d[3]));
DFFPOSX1 ecl_dff_rs3_s2d_q_reg[4](.D(exu_n19831), .CLK(rclk), .Q(ecl_ifu_exu_rs3_d[4]));
DFFPOSX1 ecl_dff_rs2_s2d_q_reg[0](.D(exu_n19829), .CLK(rclk), .Q(ecl_ifu_exu_rs2_d[0]));
DFFPOSX1 ecl_dff_rs2_s2d_q_reg[1](.D(exu_n19828), .CLK(rclk), .Q(ecl_ifu_exu_rs2_d[1]));
DFFPOSX1 ecl_dff_rs2_s2d_q_reg[2](.D(exu_n19827), .CLK(rclk), .Q(ecl_ifu_exu_rs2_d[2]));
DFFPOSX1 ecl_dff_rs2_s2d_q_reg[3](.D(exu_n19826), .CLK(rclk), .Q(ecl_ifu_exu_rs2_d[3]));
DFFPOSX1 ecl_dff_rs2_s2d_q_reg[4](.D(exu_n19825), .CLK(rclk), .Q(ecl_ifu_exu_rs2_d[4]));
DFFPOSX1 ecl_eccctl_gl_e2m_q_reg[0](.D(exu_n19823), .CLK(rclk), .Q(ecl_eccctl_gl_m[0]));
DFFPOSX1 ecl_eccctl_gl_e2m_q_reg[1](.D(exu_n19822), .CLK(rclk), .Q(ecl_eccctl_gl_m[1]));
DFFPOSX1 ecl_writeback_dff_thr_g2w2_q_reg[0](.D(exu_n19737), .CLK(rclk), .Q(ecl_wb_byplog_tid_w2[0]));
DFFPOSX1 ecl_writeback_dff_thr_g2w2_q_reg[1](.D(exu_n19736), .CLK(rclk), .Q(ecl_wb_byplog_tid_w2[1]));
DFFPOSX1 ecl_writeback_dfill_tid_dff_q_reg[0](.D(exu_n19820), .CLK(rclk), .Q(ecl_writeback_dfill_tid_g2[0]));
DFFPOSX1 ecl_writeback_dfill_tid_dff_q_reg[1](.D(exu_n19819), .CLK(rclk), .Q(ecl_writeback_dfill_tid_g2[1]));
DFFPOSX1 rml_dff_agp_thr3_q_reg[0](.D(exu_n19817), .CLK(rclk), .Q(rml_agp_thr3[0]));
DFFPOSX1 rml_dff_agp_thr3_q_reg[1](.D(exu_n19816), .CLK(rclk), .Q(rml_agp_thr3[1]));
DFFPOSX1 rml_dff_agp_thr2_q_reg[0](.D(exu_n19814), .CLK(rclk), .Q(rml_agp_thr2[0]));
DFFPOSX1 rml_dff_agp_thr2_q_reg[1](.D(exu_n19813), .CLK(rclk), .Q(rml_agp_thr2[1]));
DFFPOSX1 rml_dff_agp_thr1_q_reg[0](.D(exu_n19811), .CLK(rclk), .Q(rml_agp_thr1[0]));
DFFPOSX1 rml_dff_agp_thr1_q_reg[1](.D(exu_n19810), .CLK(rclk), .Q(rml_agp_thr1[1]));
DFFPOSX1 rml_dff_agp_thr0_q_reg[0](.D(exu_n19808), .CLK(rclk), .Q(rml_agp_thr0[0]));
DFFPOSX1 rml_dff_agp_thr0_q_reg[1](.D(exu_n19807), .CLK(rclk), .Q(rml_agp_thr0[1]));
DFFPOSX1 rml_tid_d2e_q_reg[0](.D(exu_n19805), .CLK(rclk), .Q(rml_tid_e[0]));
DFFPOSX1 rml_tid_d2e_q_reg[1](.D(exu_n19804), .CLK(rclk), .Q(rml_tid_e[1]));
DFFPOSX1 rml_tid_s2d_q_reg[0](.D(exu_n19790), .CLK(rclk), .Q(rml_tid_d[0]));
DFFPOSX1 rml_tid_s2d_q_reg[1](.D(exu_n19789), .CLK(rclk), .Q(rml_tid_d[1]));
DFFPOSX1 ecl_dff_irf_thr_m2w_q_reg[0](.D(exu_n19802), .CLK(rclk), .Q(ecl_ecl_irf_tid_w[0]));
DFFPOSX1 ecl_dff_irf_thr_m2w_q_reg[1](.D(exu_n19801), .CLK(rclk), .Q(ecl_ecl_irf_tid_w[1]));
DFFPOSX1 ecl_dff_tid_w2w1_q_reg[0](.D(exu_n19799), .CLK(rclk), .Q(ecl_tid_w1[0]));
DFFPOSX1 ecl_dff_tid_w2w1_q_reg[1](.D(exu_n19798), .CLK(rclk), .Q(ecl_tid_w1[1]));
DFFPOSX1 ecl_dff_tid_m2w_q_reg[0](.D(ecl_writeback_restore_tid_dff_n8), .CLK(rclk), .Q(ecl_tid_w[0]));
DFFPOSX1 ecl_dff_tid_m2w_q_reg[1](.D(ecl_writeback_restore_tid_dff_n13), .CLK(rclk), .Q(ecl_tid_w[1]));
DFFPOSX1 ecl_dff_thr_e2m_q_reg[0](.D(exu_n19796), .CLK(rclk), .Q(ecl_tid_m[0]));
DFFPOSX1 ecl_dff_thr_e2m_q_reg[1](.D(exu_n19795), .CLK(rclk), .Q(ecl_tid_m[1]));
DFFPOSX1 ecl_dff_tid_d2e_q_reg[0](.D(exu_n19793), .CLK(rclk), .Q(ecl_tid_e[0]));
DFFPOSX1 ecl_dff_tid_d2e_q_reg[1](.D(exu_n19792), .CLK(rclk), .Q(ecl_tid_e[1]));
DFFPOSX1 ecl_dff_thr_s2d_q_reg[0](.D(exu_n19790), .CLK(rclk), .Q(ecl_tid_d[0]));
DFFPOSX1 ecl_dff_thr_s2d_q_reg[1](.D(exu_n19789), .CLK(rclk), .Q(ecl_tid_d[1]));
DFFPOSX1 ecl_cc_d2e_q_reg[0](.D(exu_n19787), .CLK(rclk), .Q(ecl_cc_e_1));
DFFPOSX1 ecl_cc_d2e_q_reg[1](.D(exu_n19786), .CLK(rclk), .Q(ecl_cc_e_3));
DFFPOSX1 ecl_rsr_e2m_q_reg[0](.D(exu_n19784), .CLK(rclk), .Q(ecl_read_tlusr_m));
DFFPOSX1 ecl_rsr_e2m_q_reg[1](.D(exu_n19783), .CLK(rclk), .Q(ecl_byp_sel_ffusr_m));
DFFPOSX1 rml_cansave_reg_dff_reg_thr3_q_reg[0](.D(exu_n19781), .CLK(rclk), .Q(rml_cansave_reg_data_thr3[0]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr3_q_reg[1](.D(exu_n19780), .CLK(rclk), .Q(rml_cansave_reg_data_thr3[1]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr3_q_reg[2](.D(exu_n19779), .CLK(rclk), .Q(rml_cansave_reg_data_thr3[2]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr2_q_reg[0](.D(exu_n19777), .CLK(rclk), .Q(rml_cansave_reg_data_thr2[0]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr2_q_reg[1](.D(exu_n19776), .CLK(rclk), .Q(rml_cansave_reg_data_thr2[1]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr2_q_reg[2](.D(exu_n19775), .CLK(rclk), .Q(rml_cansave_reg_data_thr2[2]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr1_q_reg[0](.D(exu_n19773), .CLK(rclk), .Q(rml_cansave_reg_data_thr1[0]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr1_q_reg[1](.D(exu_n19772), .CLK(rclk), .Q(rml_cansave_reg_data_thr1[1]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr1_q_reg[2](.D(exu_n19771), .CLK(rclk), .Q(rml_cansave_reg_data_thr1[2]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr0_q_reg[0](.D(exu_n19769), .CLK(rclk), .Q(rml_cansave_reg_data_thr0[0]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr0_q_reg[1](.D(exu_n19768), .CLK(rclk), .Q(rml_cansave_reg_data_thr0[1]));
DFFPOSX1 rml_cansave_reg_dff_reg_thr0_q_reg[2](.D(exu_n19767), .CLK(rclk), .Q(rml_cansave_reg_data_thr0[2]));
DFFPOSX1 rml_cwp_dff_cwp_thr3_q_reg[0](.D(exu_n19765), .CLK(rclk), .Q(exu_tlu_cwp3_w[0]));
DFFPOSX1 rml_cwp_dff_cwp_thr3_q_reg[1](.D(exu_n19764), .CLK(rclk), .Q(exu_tlu_cwp3_w[1]));
DFFPOSX1 rml_cwp_dff_cwp_thr3_q_reg[2](.D(exu_n19763), .CLK(rclk), .Q(exu_tlu_cwp3_w[2]));
DFFPOSX1 rml_cwp_dff_cwp_thr2_q_reg[0](.D(exu_n19761), .CLK(rclk), .Q(exu_tlu_cwp2_w[0]));
DFFPOSX1 rml_cwp_dff_cwp_thr2_q_reg[1](.D(exu_n19760), .CLK(rclk), .Q(exu_tlu_cwp2_w[1]));
DFFPOSX1 rml_cwp_dff_cwp_thr2_q_reg[2](.D(exu_n19759), .CLK(rclk), .Q(exu_tlu_cwp2_w[2]));
DFFPOSX1 rml_cwp_dff_cwp_thr1_q_reg[0](.D(exu_n19757), .CLK(rclk), .Q(exu_tlu_cwp1_w[0]));
DFFPOSX1 rml_cwp_dff_cwp_thr1_q_reg[1](.D(exu_n19756), .CLK(rclk), .Q(exu_tlu_cwp1_w[1]));
DFFPOSX1 rml_cwp_dff_cwp_thr1_q_reg[2](.D(exu_n19755), .CLK(rclk), .Q(exu_tlu_cwp1_w[2]));
DFFPOSX1 rml_cwp_dff_cwp_thr0_q_reg[0](.D(exu_n19753), .CLK(rclk), .Q(exu_tlu_cwp0_w[0]));
DFFPOSX1 rml_cwp_dff_cwp_thr0_q_reg[1](.D(exu_n19752), .CLK(rclk), .Q(exu_tlu_cwp0_w[1]));
DFFPOSX1 rml_cwp_dff_cwp_thr0_q_reg[2](.D(exu_n19751), .CLK(rclk), .Q(exu_tlu_cwp0_w[2]));
DFFPOSX1 ecl_divcntl_muls_overlow_dff_q_reg[0](.D(exu_n19749), .CLK(rclk), .Q(ecl_divcntl_div_adder_out_31_w));
DFFPOSX1 ecl_divcntl_muls_overlow_dff_q_reg[1](.D(exu_n19748), .CLK(rclk), .Q(ecl_divcntl_rs2_data_31_w));
DFFPOSX1 ecl_divcntl_muls_overlow_dff_q_reg[2](.D(exu_n19747), .CLK(rclk), .Q(ecl_divcntl_muls_rs1_data_31_w));
DFFPOSX1 ecl_eccctl_cwp_e2m_q_reg[0](.D(exu_n19745), .CLK(rclk), .Q(ecl_eccctl_cwp_m[0]));
DFFPOSX1 ecl_eccctl_cwp_e2m_q_reg[1](.D(exu_n19744), .CLK(rclk), .Q(ecl_eccctl_cwp_m[1]));
DFFPOSX1 ecl_eccctl_cwp_e2m_q_reg[2](.D(exu_n19743), .CLK(rclk), .Q(ecl_eccctl_cwp_m[2]));
DFFPOSX1 ecl_eccctl_cwp_d2e_q_reg[0](.D(exu_n19741), .CLK(rclk), .Q(ecl_eccctl_cwp_e[0]));
DFFPOSX1 ecl_eccctl_cwp_d2e_q_reg[1](.D(exu_n19740), .CLK(rclk), .Q(ecl_eccctl_cwp_e[1]));
DFFPOSX1 ecl_eccctl_cwp_d2e_q_reg[2](.D(exu_n19739), .CLK(rclk), .Q(ecl_eccctl_cwp_e[2]));
DFFPOSX1 ecl_ccr_setcc_g2w2_q_reg[0](.D(exu_n19737), .CLK(rclk), .Q(ecl_ccr_thr_w2[0]));
DFFPOSX1 ecl_ccr_setcc_g2w2_q_reg[1](.D(exu_n19736), .CLK(rclk), .Q(ecl_ccr_thr_w2[1]));
DFFPOSX1 ecl_ccr_setcc_g2w2_q_reg[2](.D(exu_n19735), .CLK(rclk), .Q(ecl_ccr_setcc_w2));
DFFPOSX1 rml_cleanwin_d2e_q_reg[0](.D(exu_n19733), .CLK(rclk), .Q(rml_rml_ecl_cleanwin_e[0]));
DFFPOSX1 rml_cleanwin_d2e_q_reg[1](.D(exu_n19732), .CLK(rclk), .Q(rml_rml_ecl_cleanwin_e[1]));
DFFPOSX1 rml_cleanwin_d2e_q_reg[2](.D(exu_n19731), .CLK(rclk), .Q(rml_rml_ecl_cleanwin_e[2]));
DFFPOSX1 rml_otherwin_d2e_q_reg[0](.D(exu_n19729), .CLK(rclk), .Q(rml_rml_ecl_otherwin_e[0]));
DFFPOSX1 rml_otherwin_d2e_q_reg[1](.D(exu_n19728), .CLK(rclk), .Q(rml_rml_ecl_otherwin_e[1]));
DFFPOSX1 rml_otherwin_d2e_q_reg[2](.D(exu_n19727), .CLK(rclk), .Q(rml_rml_ecl_otherwin_e[2]));
DFFPOSX1 rml_canrestore_d2e_q_reg[0](.D(exu_n19725), .CLK(rclk), .Q(rml_rml_ecl_canrestore_e[0]));
DFFPOSX1 rml_canrestore_d2e_q_reg[1](.D(exu_n19724), .CLK(rclk), .Q(rml_rml_ecl_canrestore_e[1]));
DFFPOSX1 rml_canrestore_d2e_q_reg[2](.D(exu_n19723), .CLK(rclk), .Q(rml_rml_ecl_canrestore_e[2]));
DFFPOSX1 rml_cansave_d2e_q_reg[0](.D(exu_n19721), .CLK(rclk), .Q(rml_rml_ecl_cansave_e[0]));
DFFPOSX1 rml_cansave_d2e_q_reg[1](.D(exu_n19720), .CLK(rclk), .Q(rml_rml_ecl_cansave_e[1]));
DFFPOSX1 rml_cansave_d2e_q_reg[2](.D(exu_n19719), .CLK(rclk), .Q(rml_rml_ecl_cansave_e[2]));
DFFPOSX1 rml_next_cleanwin_m2w_q_reg[0](.D(exu_n19717), .CLK(rclk), .Q(rml_next_cleanwin_w[0]));
DFFPOSX1 rml_next_cleanwin_m2w_q_reg[1](.D(exu_n19716), .CLK(rclk), .Q(rml_next_cleanwin_w[1]));
DFFPOSX1 rml_next_cleanwin_m2w_q_reg[2](.D(exu_n19715), .CLK(rclk), .Q(rml_next_cleanwin_w[2]));
DFFPOSX1 rml_next_cleanwin_e2m_q_reg[0](.D(exu_n19713), .CLK(rclk), .Q(rml_next_cleanwin_m[0]));
DFFPOSX1 rml_next_cleanwin_e2m_q_reg[1](.D(exu_n19712), .CLK(rclk), .Q(rml_next_cleanwin_m[1]));
DFFPOSX1 rml_next_cleanwin_e2m_q_reg[2](.D(exu_n19711), .CLK(rclk), .Q(rml_next_cleanwin_m[2]));
DFFPOSX1 rml_next_otherwin_m2w_q_reg[0](.D(exu_n19709), .CLK(rclk), .Q(rml_next_otherwin_w[0]));
DFFPOSX1 rml_next_otherwin_m2w_q_reg[1](.D(exu_n19708), .CLK(rclk), .Q(rml_next_otherwin_w[1]));
DFFPOSX1 rml_next_otherwin_m2w_q_reg[2](.D(exu_n19707), .CLK(rclk), .Q(rml_next_otherwin_w[2]));
DFFPOSX1 rml_next_otherwin_e2m_q_reg[0](.D(exu_n19705), .CLK(rclk), .Q(rml_next_otherwin_m[0]));
DFFPOSX1 rml_next_otherwin_e2m_q_reg[1](.D(exu_n19704), .CLK(rclk), .Q(rml_next_otherwin_m[1]));
DFFPOSX1 rml_next_otherwin_e2m_q_reg[2](.D(exu_n19703), .CLK(rclk), .Q(rml_next_otherwin_m[2]));
DFFPOSX1 rml_next_canrestore_m2w_q_reg[0](.D(exu_n19701), .CLK(rclk), .Q(rml_next_canrestore_w[0]));
DFFPOSX1 rml_next_canrestore_m2w_q_reg[1](.D(exu_n19700), .CLK(rclk), .Q(rml_next_canrestore_w[1]));
DFFPOSX1 rml_next_canrestore_m2w_q_reg[2](.D(exu_n19699), .CLK(rclk), .Q(rml_next_canrestore_w[2]));
DFFPOSX1 rml_next_canrestore_e2m_q_reg[0](.D(exu_n19697), .CLK(rclk), .Q(rml_next_canrestore_m[0]));
DFFPOSX1 rml_next_canrestore_e2m_q_reg[1](.D(exu_n19696), .CLK(rclk), .Q(rml_next_canrestore_m[1]));
DFFPOSX1 rml_next_canrestore_e2m_q_reg[2](.D(exu_n19695), .CLK(rclk), .Q(rml_next_canrestore_m[2]));
DFFPOSX1 rml_next_cansave_m2w_q_reg[0](.D(exu_n19693), .CLK(rclk), .Q(rml_next_cansave_w[0]));
DFFPOSX1 rml_next_cansave_m2w_q_reg[1](.D(exu_n19692), .CLK(rclk), .Q(rml_next_cansave_w[1]));
DFFPOSX1 rml_next_cansave_m2w_q_reg[2](.D(exu_n19691), .CLK(rclk), .Q(rml_next_cansave_w[2]));
DFFPOSX1 rml_next_cansave_e2m_q_reg[0](.D(exu_n19689), .CLK(rclk), .Q(rml_next_cansave_m[0]));
DFFPOSX1 rml_next_cansave_e2m_q_reg[1](.D(exu_n19688), .CLK(rclk), .Q(rml_next_cansave_m[1]));
DFFPOSX1 rml_next_cansave_e2m_q_reg[2](.D(exu_n19687), .CLK(rclk), .Q(rml_next_cansave_m[2]));
DFFPOSX1 rml_next_cwp_m2w_q_reg[0](.D(exu_n19685), .CLK(rclk), .Q(rml_next_cwp_noreset_w[0]));
DFFPOSX1 rml_next_cwp_m2w_q_reg[1](.D(exu_n19684), .CLK(rclk), .Q(rml_next_cwp_noreset_w[1]));
DFFPOSX1 rml_next_cwp_m2w_q_reg[2](.D(exu_n19683), .CLK(rclk), .Q(rml_next_cwp_noreset_w[2]));
DFFPOSX1 rml_next_cwp_e2m_q_reg[0](.D(exu_n19681), .CLK(rclk), .Q(rml_next_cwp_m[0]));
DFFPOSX1 rml_next_cwp_e2m_q_reg[1](.D(exu_n19680), .CLK(rclk), .Q(rml_next_cwp_m[1]));
DFFPOSX1 rml_next_cwp_e2m_q_reg[2](.D(exu_n19679), .CLK(rclk), .Q(rml_next_cwp_m[2]));
DFFPOSX1 rml_wtype_d2e_q_reg[0](.D(exu_n19677), .CLK(rclk), .Q(rml_ecl_wtype_e[0]));
DFFPOSX1 rml_wtype_d2e_q_reg[1](.D(exu_n19676), .CLK(rclk), .Q(rml_ecl_wtype_e[1]));
DFFPOSX1 rml_wtype_d2e_q_reg[2](.D(exu_n19675), .CLK(rclk), .Q(rml_ecl_wtype_e[2]));
DFFPOSX1 ecl_dff_shiftop_d2e_q_reg[0](.D(exu_n19673), .CLK(rclk), .Q(ecl_shiftop_e_0));
DFFPOSX1 ecl_dff_shiftop_d2e_q_reg[1](.D(exu_n19672), .CLK(rclk), .Q(ecl_shft_lshift_e_l));
DFFPOSX1 ecl_dff_shiftop_d2e_q_reg[2](.D(exu_n19671), .CLK(rclk), .Q(ecl_shiftop_e[2]));
DFFPOSX1 rml_cwp_fastcmplt_dff_q_reg[0](.D(exu_n19669), .CLK(rclk), .Q(rml_cwp_cwp_fastcmplt_w));
DFFPOSX1 rml_cwp_full_swap_m2w_q_reg[0](.D(exu_n19668), .CLK(rclk), .Q(rml_cwp_full_swap_w));
DFFPOSX1 rml_cwp_full_swap_e2m_q_reg[0](.D(exu_n19667), .CLK(rclk), .Q(rml_cwp_full_swap_m));
DFFPOSX1 ecl_mdqctl_mulstate_dff_q_reg[0](.D(exu_n19666), .CLK(rclk), .Q(ecl_mdqctl_divcntl_muldone));
DFFPOSX1 ecl_mdqctl_dff_done_c32c4_q_reg[0](.D(exu_n19665), .CLK(rclk), .Q(ecl_div_mul_wen));
DFFPOSX1 ecl_mdqctl_dff_done_c22c3_q_reg[0](.D(exu_n19664), .CLK(rclk), .Q(ecl_mdqctl_mul_done_c3));
DFFPOSX1 ecl_mdqctl_dff_done_c1c2_q_reg[0](.D(exu_n19663), .CLK(rclk), .Q(ecl_mdqctl_mul_done_c2));
DFFPOSX1 ecl_mdqctl_dff_done_c02c1_q_reg[0](.D(exu_n19662), .CLK(rclk), .Q(ecl_mdqctl_mul_done_c1));
DFFPOSX1 ecl_mdqctl_dff_done_ack2c0_q_reg[0](.D(exu_n19661), .CLK(rclk), .Q(ecl_mdqctl_mul_done_c0));
DFFPOSX1 ecl_mdqctl_mul_ready_dff_q_reg[0](.D(exu_n19660), .CLK(rclk), .Q(exu_mul_input_vld));
DFFPOSX1 ecl_mdqctl_ismul_m2w_q_reg[0](.D(exu_n19659), .CLK(rclk), .Q(ecl_mdqctl_ismul_w));
DFFPOSX1 ecl_mdqctl_ismul_e2m_q_reg[0](.D(exu_n19658), .CLK(rclk), .Q(ecl_mdqctl_ismul_m));
DFFPOSX1 ecl_mdqctl_ismul_d2e_q_reg[0](.D(exu_n19657), .CLK(rclk), .Q(ecl_mdqctl_ismul_e));
DFFPOSX1 ecl_mdqctl_isdiv_m2w_q_reg[0](.D(exu_n19655), .CLK(rclk), .Q(ecl_mdqctl_isdiv_w));
DFFPOSX1 ecl_mdqctl_isdiv_e2m_q_reg[0](.D(exu_n19653), .CLK(rclk), .Q(ecl_mdqctl_isdiv_m));
DFFPOSX1 ecl_mdqctl_isdiv_d2e_q_reg[0](.D(exu_n19651), .CLK(rclk), .Q(ecl_div_ld_inputs));
DFFPOSX1 ecl_mdqctl_div_zero_e2m_q_reg[0](.D(exu_n19649), .CLK(rclk), .Q(ecl_mdqctl_div_zero_unqual_m));
DFFPOSX1 ecl_divcntl_muls_v_dff_q_reg[0](.D(exu_n19647), .CLK(rclk), .Q(ecl_divcntl_muls_v));
DFFPOSX1 ecl_divcntl_muls_c_dff_q_reg[0](.D(exu_n19645), .CLK(rclk), .Q(ecl_divcntl_muls_c));
DFFPOSX1 ecl_divcntl_last_cin_dff_q_reg[0](.D(exu_n19643), .CLK(rclk), .Q(ecl_divcntl_last_cin));
DFFPOSX1 ecl_divcntl_zero_rem_dff_q_reg[0](.D(exu_n19641), .CLK(rclk), .Q(ecl_divcntl_zero_rem_q));
DFFPOSX1 ecl_divcntl_sub_dff_q_reg[0](.D(exu_n19639), .CLK(rclk), .Q(ecl_divcntl_subtract));
DFFPOSX1 ecl_divcntl_q_dff_q_reg[0](.D(exu_n19638), .CLK(rclk), .Q(ecl_div_newq));
DFFPOSX1 ecl_eccctl_rs3_ue_e2m_q_reg[0](.D(exu_n19636), .CLK(rclk), .Q(ecl_eccctl_rs3_ue_m));
DFFPOSX1 ecl_eccctl_rs2_ce_e2m_q_reg[0](.D(exu_n19634), .CLK(rclk), .Q(ecl_eccctl_rs2_ce_m));
DFFPOSX1 ecl_eccctl_rs2_ue_e2m_q_reg[0](.D(exu_n19632), .CLK(rclk), .Q(ecl_eccctl_rs2_ue_m));
DFFPOSX1 ecl_eccctl_rs1_ce_e2m_q_reg[0](.D(exu_n19622), .CLK(rclk), .Q(ecl_eccctl_rs1_ce_m));
DFFPOSX1 ecl_eccctl_rs1_ue_e2m_q_reg[0](.D(exu_n19630), .CLK(rclk), .Q(ecl_eccctl_rs1_ue_m));
DFFPOSX1 ecl_eccctl_inj_irferr_m2w_q_reg[0](.D(exu_n19628), .CLK(rclk), .Q(exu_ifu_inj_ack));
DFFPOSX1 ecl_eccctl_ecc_sel_rs3_dff_q_reg[0](.D(exu_n19626), .CLK(rclk), .Q(ecl_eccctl_sel_rs3_m));
DFFPOSX1 ecl_eccctl_ecc_sel_rs2_dff_q_reg[0](.D(exu_n19624), .CLK(rclk), .Q(ecl_eccctl_sel_rs2_m));
DFFPOSX1 ecl_eccctl_ecc_sel_rs1_dff_q_reg[0](.D(exu_n19622), .CLK(rclk), .Q(ecl_eccctl_sel_rs1_m));
DFFPOSX1 ecl_eccctl_nceen_e2m_q_reg[0](.D(exu_n19620), .CLK(rclk), .Q(ecl_eccctl_nceen_m));
DFFPOSX1 ecl_eccctl_ecc_ue_e2m_q_reg[0](.D(exu_n19618), .CLK(rclk), .Q(exu_ifu_ecc_ue_m));
DFFPOSX1 ecl_eccctl_byp_sel_ecc_e2m_q_reg[0](.D(exu_n19616), .CLK(rclk), .Q(ecl_byp_sel_ecc_m));
DFFPOSX1 ecl_eccctl_rs3_rf_dff_q_reg[0](.D(exu_n19614), .CLK(rclk), .Q(ecl_eccctl_rs3_sel_rf_e));
DFFPOSX1 ecl_eccctl_rs2_rf_dff_q_reg[0](.D(exu_n19612), .CLK(rclk), .Q(ecl_eccctl_rs2_sel_rf_e));
DFFPOSX1 ecl_eccctl_rs1_rf_dff_q_reg[0](.D(exu_n19610), .CLK(rclk), .Q(ecl_eccctl_rs1_sel_rf_e));
DFFPOSX1 ecl_writeback_longop_done_e2m_q_reg[0](.D(exu_n19608), .CLK(rclk), .Q(ecl_writeback_short_longop_done_m));
DFFPOSX1 ecl_writeback_restore_ready_dff_q_reg[0](.D(exu_n19606), .CLK(rclk), .Q(ecl_writeback_restore_ready));
DFFPOSX1 ecl_writeback_restore_m2w_q_reg[0](.D(exu_n19604), .CLK(rclk), .Q(ecl_writeback_restore_w));
DFFPOSX1 ecl_writeback_restore_e2m_q_reg[0](.D(exu_n19602), .CLK(rclk), .Q(ecl_byp_restore_m));
DFFPOSX1 ecl_writeback_return_d2e_q_reg[0](.D(exu_n19600), .CLK(rclk), .Q(ecl_writeback_return_e));
DFFPOSX1 ecl_writeback_dff_yreg_wen_w2w1_q_reg[0](.D(exu_n19598), .CLK(rclk), .Q(ecl_writeback_yreg_wen_w1));
DFFPOSX1 ecl_writeback_dff_wrsr_m2w_q_reg[0](.D(exu_n19596), .CLK(rclk), .Q(ecl_writeback_wrsr_w));
DFFPOSX1 ecl_writeback_dff_wrsr_e2m_q_reg[0](.D(exu_n19594), .CLK(rclk), .Q(ecl_writeback_wrsr_m));
DFFPOSX1 ecl_writeback_dff_wrsr_d2e_q_reg[0](.D(exu_n19592), .CLK(rclk), .Q(exu_ffu_wsr_inst_e));
DFFPOSX1 ecl_writeback_dff_wb_e2m_q_reg[0](.D(exu_n19590), .CLK(rclk), .Q(ecl_bypass_m));
DFFPOSX1 ecl_writeback_dff_wb_d2e_q_reg[0](.D(exu_n19588), .CLK(rclk), .Q(ecl_wb_e));
DFFPOSX1 ecl_writeback_ecc_wen_m2w_q_reg[0](.D(exu_n19586), .CLK(rclk), .Q(ecl_writeback_inst_vld_noflush_wen_w));
DFFPOSX1 ecl_writeback_dff_lsu_wen_m2w_q_reg[0](.D(exu_n19584), .CLK(rclk), .Q(ecl_writeback_wen_no_inst_vld_w));
DFFPOSX1 ecl_writeback_wen_w2_dff_q_reg[0](.D(exu_n19582), .CLK(rclk), .Q(ecl_wb_byplog_wen_w2));
DFFPOSX1 ecl_writeback_dfill_vld_dff_q_reg[0](.D(exu_n19580), .CLK(rclk), .Q(ecl_wb_byplog_wen_g2));
DFFPOSX1 ecl_ccr_dff_setcc_m2w_q_reg[0](.D(exu_n19578), .CLK(rclk), .Q(ecl_ccr_setcc_w));
DFFPOSX1 ecl_ccr_dff_setcc_e2m_q_reg[0](.D(exu_n19576), .CLK(rclk), .Q(ecl_ccr_setcc_m));
DFFPOSX1 ecl_ccr_dff_setcc_d2e_q_reg[0](.D(exu_n19574), .CLK(rclk), .Q(ecl_ccr_setcc_e));
DFFPOSX1 bypass_w2_eccgen_Ip7ff_0__q_reg[0](.D(exu_n19572), .CLK(exu_n16179), .Q(bypass_w2_eccgen_p7_w[0]));
DFFPOSX1 bypass_w2_eccgen_Ip7ff_1__q_reg[0](.D(exu_n19570), .CLK(exu_n16179), .Q(bypass_w2_eccgen_p7_w[1]));
DFFPOSX1 bypass_w2_eccgen_Ip7ff_2__q_reg[0](.D(exu_n19568), .CLK(exu_n16179), .Q(bypass_w2_eccgen_p7_w[2]));
DFFPOSX1 bypass_w2_eccgen_Ip7ff_3__q_reg[0](.D(exu_n19566), .CLK(exu_n16179), .Q(bypass_w2_eccgen_p7_w[3]));
DFFPOSX1 bypass_w2_eccgen_Ip7ff_4__q_reg[0](.D(exu_n19564), .CLK(exu_n16179), .Q(bypass_w2_eccgen_p7_w[4]));
DFFPOSX1 bypass_w2_eccgen_Ip7ff_5__q_reg[0](.D(exu_n19562), .CLK(exu_n16179), .Q(bypass_w2_eccgen_p7_w[5]));
DFFPOSX1 bypass_w2_eccgen_Ip7ff_6__q_reg[0](.D(exu_n19560), .CLK(exu_n16179), .Q(bypass_w2_eccgen_p7_w[6]));
DFFPOSX1 bypass_w2_eccgen_Ip7ff_7__q_reg[0](.D(exu_n19558), .CLK(exu_n16179), .Q(bypass_w2_eccgen_p7_w[7]));
DFFPOSX1 bypass_w2_eccgen_Ip6ff_0__q_reg[0](.D(exu_n19556), .CLK(exu_n16179), .Q(bypass_w2_eccgen_p6_w[0]));
DFFPOSX1 bypass_w2_eccgen_Ip6ff_1__q_reg[0](.D(exu_n19554), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p6_w[1]));
DFFPOSX1 bypass_w2_eccgen_Ip5ff_0__q_reg[0](.D(exu_n19552), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p5_w[0]));
DFFPOSX1 bypass_w2_eccgen_Ip5ff_1__q_reg[0](.D(exu_n19550), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p5_w[1]));
DFFPOSX1 bypass_w2_eccgen_Ip4ff_0__q_reg[0](.D(exu_n19548), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p4_w[0]));
DFFPOSX1 bypass_w2_eccgen_Ip4ff_1__q_reg[0](.D(exu_n19546), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p4_w[1]));
DFFPOSX1 bypass_w2_eccgen_Ip4ff_2__q_reg[0](.D(exu_n19544), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p4_w[2]));
DFFPOSX1 bypass_w2_eccgen_Ip4ff_3__q_reg[0](.D(exu_n19542), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p4_w[3]));
DFFPOSX1 bypass_w2_eccgen_Ip3ff_0__q_reg[0](.D(exu_n19540), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p3_w[0]));
DFFPOSX1 bypass_w2_eccgen_Ip3ff_1__q_reg[0](.D(exu_n19538), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p3_w[1]));
DFFPOSX1 bypass_w2_eccgen_Ip3ff_2__q_reg[0](.D(exu_n19536), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p3_w[2]));
DFFPOSX1 bypass_w2_eccgen_Ip3ff_3__q_reg[0](.D(exu_n19534), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p3_w[3]));
DFFPOSX1 bypass_w2_eccgen_Ip3ff_4__q_reg[0](.D(exu_n19532), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p3_w[4]));
DFFPOSX1 bypass_w2_eccgen_Ip3ff_5__q_reg[0](.D(exu_n19530), .CLK(exu_n16178), .Q(bypass_w2_eccgen_p3_w[5]));
DFFPOSX1 bypass_w2_eccgen_Ip3ff_6__q_reg[0](.D(exu_n19528), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p3_w[6]));
DFFPOSX1 bypass_w2_eccgen_Ip3ff_7__q_reg[0](.D(exu_n19526), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p3_w[7]));
DFFPOSX1 bypass_w2_eccgen_Ip2ff_0__q_reg[0](.D(exu_n19524), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p2_w[0]));
DFFPOSX1 bypass_w2_eccgen_Ip2ff_1__q_reg[0](.D(exu_n19522), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p2_w[1]));
DFFPOSX1 bypass_w2_eccgen_Ip2ff_2__q_reg[0](.D(exu_n19520), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p2_w[2]));
DFFPOSX1 bypass_w2_eccgen_Ip2ff_3__q_reg[0](.D(exu_n19518), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p2_w[3]));
DFFPOSX1 bypass_w2_eccgen_Ip2ff_4__q_reg[0](.D(exu_n19516), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p2_w[4]));
DFFPOSX1 bypass_w2_eccgen_Ip2ff_5__q_reg[0](.D(exu_n19514), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p2_w[5]));
DFFPOSX1 bypass_w2_eccgen_Ip2ff_6__q_reg[0](.D(exu_n19512), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p2_w[6]));
DFFPOSX1 bypass_w2_eccgen_Ip2ff_7__q_reg[0](.D(exu_n19510), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p2_w[7]));
DFFPOSX1 bypass_w2_eccgen_Ip1ff_0__q_reg[0](.D(exu_n19508), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p1_w[0]));
DFFPOSX1 bypass_w2_eccgen_Ip1ff_1__q_reg[0](.D(exu_n19506), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p1_w[1]));
DFFPOSX1 bypass_w2_eccgen_Ip1ff_2__q_reg[0](.D(exu_n19504), .CLK(exu_n16177), .Q(bypass_w2_eccgen_p1_w[2]));
DFFPOSX1 bypass_w2_eccgen_Ip1ff_3__q_reg[0](.D(exu_n19502), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p1_w[3]));
DFFPOSX1 bypass_w2_eccgen_Ip1ff_4__q_reg[0](.D(exu_n19500), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p1_w[4]));
DFFPOSX1 bypass_w2_eccgen_Ip1ff_5__q_reg[0](.D(exu_n19498), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p1_w[5]));
DFFPOSX1 bypass_w2_eccgen_Ip1ff_6__q_reg[0](.D(exu_n19496), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p1_w[6]));
DFFPOSX1 bypass_w2_eccgen_Ip1ff_7__q_reg[0](.D(exu_n19494), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p1_w[7]));
DFFPOSX1 bypass_w2_eccgen_Ip0ff_0__q_reg[0](.D(exu_n19492), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p0_w[0]));
DFFPOSX1 bypass_w2_eccgen_Ip0ff_1__q_reg[0](.D(exu_n19490), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p0_w[1]));
DFFPOSX1 bypass_w2_eccgen_Ip0ff_2__q_reg[0](.D(exu_n19488), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p0_w[2]));
DFFPOSX1 bypass_w2_eccgen_Ip0ff_3__q_reg[0](.D(exu_n19486), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p0_w[3]));
DFFPOSX1 bypass_w2_eccgen_Ip0ff_4__q_reg[0](.D(exu_n19484), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p0_w[4]));
DFFPOSX1 bypass_w2_eccgen_Ip0ff_5__q_reg[0](.D(exu_n19482), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p0_w[5]));
DFFPOSX1 bypass_w2_eccgen_Ip0ff_6__q_reg[0](.D(exu_n19480), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p0_w[6]));
DFFPOSX1 bypass_w2_eccgen_Ip0ff_7__q_reg[0](.D(exu_n19478), .CLK(exu_n16176), .Q(bypass_w2_eccgen_p0_w[7]));
DFFPOSX1 bypass_w2_eccgen_Imsk_4__q_reg[0](.D(exu_n19380), .CLK(exu_n16175), .Q(bypass_w2_eccgen_msk_w4));
DFFPOSX1 bypass_w2_eccgen_Imsk_5__q_reg[0](.D(exu_n19378), .CLK(exu_n16175), .Q(bypass_w2_eccgen_msk_w5));
DFFPOSX1 bypass_w1_eccgen_Ip7ff_0__q_reg[0](.D(exu_n19476), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p7_w[0]));
DFFPOSX1 bypass_w1_eccgen_Ip7ff_1__q_reg[0](.D(exu_n19474), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p7_w[1]));
DFFPOSX1 bypass_w1_eccgen_Ip7ff_2__q_reg[0](.D(exu_n19472), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p7_w[2]));
DFFPOSX1 bypass_w1_eccgen_Ip7ff_3__q_reg[0](.D(exu_n19470), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p7_w[3]));
DFFPOSX1 bypass_w1_eccgen_Ip7ff_4__q_reg[0](.D(exu_n19468), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p7_w[4]));
DFFPOSX1 bypass_w1_eccgen_Ip7ff_5__q_reg[0](.D(exu_n19466), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p7_w[5]));
DFFPOSX1 bypass_w1_eccgen_Ip7ff_6__q_reg[0](.D(exu_n19464), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p7_w[6]));
DFFPOSX1 bypass_w1_eccgen_Ip7ff_7__q_reg[0](.D(exu_n19462), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p7_w[7]));
DFFPOSX1 bypass_w1_eccgen_Ip6ff_0__q_reg[0](.D(exu_n19460), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p6_w[0]));
DFFPOSX1 bypass_w1_eccgen_Ip6ff_1__q_reg[0](.D(exu_n19458), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p6_w[1]));
DFFPOSX1 bypass_w1_eccgen_Ip5ff_0__q_reg[0](.D(exu_n19456), .CLK(exu_n16175), .Q(bypass_w1_eccgen_p5_w[0]));
DFFPOSX1 bypass_w1_eccgen_Ip5ff_1__q_reg[0](.D(exu_n19454), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p5_w[1]));
DFFPOSX1 bypass_w1_eccgen_Ip4ff_0__q_reg[0](.D(exu_n19452), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p4_w[0]));
DFFPOSX1 bypass_w1_eccgen_Ip4ff_1__q_reg[0](.D(exu_n19450), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p4_w[1]));
DFFPOSX1 bypass_w1_eccgen_Ip4ff_2__q_reg[0](.D(exu_n19448), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p4_w[2]));
DFFPOSX1 bypass_w1_eccgen_Ip4ff_3__q_reg[0](.D(exu_n19446), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p4_w[3]));
DFFPOSX1 bypass_w1_eccgen_Ip3ff_0__q_reg[0](.D(exu_n19444), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p3_w[0]));
DFFPOSX1 bypass_w1_eccgen_Ip3ff_1__q_reg[0](.D(exu_n19442), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p3_w[1]));
DFFPOSX1 bypass_w1_eccgen_Ip3ff_2__q_reg[0](.D(exu_n19440), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p3_w[2]));
DFFPOSX1 bypass_w1_eccgen_Ip3ff_3__q_reg[0](.D(exu_n19438), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p3_w[3]));
DFFPOSX1 bypass_w1_eccgen_Ip3ff_4__q_reg[0](.D(exu_n19436), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p3_w[4]));
DFFPOSX1 bypass_w1_eccgen_Ip3ff_5__q_reg[0](.D(exu_n19434), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p3_w[5]));
DFFPOSX1 bypass_w1_eccgen_Ip3ff_6__q_reg[0](.D(exu_n19432), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p3_w[6]));
DFFPOSX1 bypass_w1_eccgen_Ip3ff_7__q_reg[0](.D(exu_n19430), .CLK(exu_n16174), .Q(bypass_w1_eccgen_p3_w[7]));
DFFPOSX1 bypass_w1_eccgen_Ip2ff_0__q_reg[0](.D(exu_n19428), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p2_w[0]));
DFFPOSX1 bypass_w1_eccgen_Ip2ff_1__q_reg[0](.D(exu_n19426), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p2_w[1]));
DFFPOSX1 bypass_w1_eccgen_Ip2ff_2__q_reg[0](.D(exu_n19424), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p2_w[2]));
DFFPOSX1 bypass_w1_eccgen_Ip2ff_3__q_reg[0](.D(exu_n19422), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p2_w[3]));
DFFPOSX1 bypass_w1_eccgen_Ip2ff_4__q_reg[0](.D(exu_n19420), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p2_w[4]));
DFFPOSX1 bypass_w1_eccgen_Ip2ff_5__q_reg[0](.D(exu_n19418), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p2_w[5]));
DFFPOSX1 bypass_w1_eccgen_Ip2ff_6__q_reg[0](.D(exu_n19416), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p2_w[6]));
DFFPOSX1 bypass_w1_eccgen_Ip2ff_7__q_reg[0](.D(exu_n19414), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p2_w[7]));
DFFPOSX1 bypass_w1_eccgen_Ip1ff_0__q_reg[0](.D(exu_n19412), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p1_w[0]));
DFFPOSX1 bypass_w1_eccgen_Ip1ff_1__q_reg[0](.D(exu_n19410), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p1_w[1]));
DFFPOSX1 bypass_w1_eccgen_Ip1ff_2__q_reg[0](.D(exu_n19408), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p1_w[2]));
DFFPOSX1 bypass_w1_eccgen_Ip1ff_3__q_reg[0](.D(exu_n19406), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p1_w[3]));
DFFPOSX1 bypass_w1_eccgen_Ip1ff_4__q_reg[0](.D(exu_n19404), .CLK(exu_n16173), .Q(bypass_w1_eccgen_p1_w[4]));
DFFPOSX1 bypass_w1_eccgen_Ip1ff_5__q_reg[0](.D(exu_n19402), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p1_w[5]));
DFFPOSX1 bypass_w1_eccgen_Ip1ff_6__q_reg[0](.D(exu_n19400), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p1_w[6]));
DFFPOSX1 bypass_w1_eccgen_Ip1ff_7__q_reg[0](.D(exu_n19398), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p1_w[7]));
DFFPOSX1 bypass_w1_eccgen_Ip0ff_0__q_reg[0](.D(exu_n19396), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p0_w[0]));
DFFPOSX1 bypass_w1_eccgen_Ip0ff_1__q_reg[0](.D(exu_n19394), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p0_w[1]));
DFFPOSX1 bypass_w1_eccgen_Ip0ff_2__q_reg[0](.D(exu_n19392), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p0_w[2]));
DFFPOSX1 bypass_w1_eccgen_Ip0ff_3__q_reg[0](.D(exu_n19390), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p0_w[3]));
DFFPOSX1 bypass_w1_eccgen_Ip0ff_4__q_reg[0](.D(exu_n19388), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p0_w[4]));
DFFPOSX1 bypass_w1_eccgen_Ip0ff_5__q_reg[0](.D(exu_n19386), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p0_w[5]));
DFFPOSX1 bypass_w1_eccgen_Ip0ff_6__q_reg[0](.D(exu_n19384), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p0_w[6]));
DFFPOSX1 bypass_w1_eccgen_Ip0ff_7__q_reg[0](.D(exu_n19382), .CLK(exu_n16172), .Q(bypass_w1_eccgen_p0_w[7]));
DFFPOSX1 bypass_w1_eccgen_Imsk_4__q_reg[0](.D(exu_n19380), .CLK(exu_n16172), .Q(bypass_w1_eccgen_msk_w4));
DFFPOSX1 bypass_w1_eccgen_Imsk_5__q_reg[0](.D(exu_n19378), .CLK(exu_n16172), .Q(bypass_w1_eccgen_msk_w5));
DFFPOSX1 rml_cleanwin_wen_m2w_q_reg[0](.D(exu_n19376), .CLK(rclk), .Q(rml_rml_cleanwin_wen_w));
DFFPOSX1 rml_cleanwin_wen_e2m_q_reg[0](.D(exu_n19374), .CLK(rclk), .Q(rml_cleanwin_wen_m));
DFFPOSX1 rml_otherwin_wen_m2w_q_reg[0](.D(exu_n19372), .CLK(rclk), .Q(rml_rml_otherwin_wen_w));
DFFPOSX1 rml_otherwin_wen_e2m_q_reg[0](.D(exu_n19370), .CLK(rclk), .Q(rml_otherwin_wen_m));
DFFPOSX1 rml_canrestore_wen_m2w_q_reg[0](.D(exu_n19368), .CLK(rclk), .Q(rml_rml_canrestore_wen_w));
DFFPOSX1 rml_canrestore_wen_e2m_q_reg[0](.D(exu_n19366), .CLK(rclk), .Q(rml_canrestore_wen_m));
DFFPOSX1 rml_cansave_wen_m2w_q_reg[0](.D(exu_n19364), .CLK(rclk), .Q(rml_rml_cansave_wen_w));
DFFPOSX1 rml_cansave_wen_e2m_q_reg[0](.D(exu_n19362), .CLK(rclk), .Q(rml_cansave_wen_m));
DFFPOSX1 rml_cwp_wen_m2w_q_reg[0](.D(exu_n19360), .CLK(rclk), .Q(rml_cwp_wen_nokill_w));
DFFPOSX1 rml_cwp_wen_e2m_q_reg[0](.D(exu_n19358), .CLK(rclk), .Q(rml_rml_cwp_wen_m));
DFFPOSX1 rml_dff_kill_restore_m2w_q_reg[0](.D(exu_n19356), .CLK(rclk), .Q(rml_kill_restore_w));
DFFPOSX1 rml_dff_did_restore_m2w_q_reg[0](.D(exu_n19354), .CLK(rclk), .Q(rml_did_restore_w));
DFFPOSX1 rml_dff_did_restore_e2m_q_reg[0](.D(exu_n19352), .CLK(rclk), .Q(rml_did_restore_m));
DFFPOSX1 rml_other_d2e_q_reg[0](.D(exu_n19350), .CLK(rclk), .Q(rml_ecl_other_e));
DFFPOSX1 rml_rml_kill_e2m_q_reg[0](.D(exu_n19348), .CLK(rclk), .Q(rml_ecl_kill_m));
DFFPOSX1 rml_spill_e2m_q_reg[0](.D(exu_n19346), .CLK(rclk), .Q(rml_spill_m));
DFFPOSX1 rml_win_trap_m2w_q_reg[0](.D(exu_n19344), .CLK(rclk), .Q(rml_win_trap_w));
DFFPOSX1 rml_win_trap_e2m_q_reg[0](.D(exu_n19342), .CLK(rclk), .Q(rml_win_trap_m));
DFFPOSX1 rml_restore_d2e_q_reg[0](.D(exu_n19294), .CLK(rclk), .Q(rml_restore_e));
DFFPOSX1 rml_save_e2m_q_reg[0](.D(exu_n19340), .CLK(rclk), .Q(rml_save_m));
DFFPOSX1 rml_save_d2e_q_reg[0](.D(exu_n19292), .CLK(rclk), .Q(rml_save_e));
DFFPOSX1 alu_invert_d2e_q_reg[0](.D(exu_n16321), .CLK(rclk), .Q(alu_invert_e));
DFFPOSX1 ecl_ld_thr_match_sg_dff_q_reg[0](.D(exu_n19336), .CLK(rclk), .Q(ecl_ld_thr_match_dg2));
DFFPOSX1 ecl_ld_thr_match_sm_dff_q_reg[0](.D(exu_n19334), .CLK(rclk), .Q(ecl_ld_thr_match_dg));
DFFPOSX1 ecl_thr_match_se_dff_q_reg[0](.D(exu_n19332), .CLK(rclk), .Q(ecl_thr_match_dm));
DFFPOSX1 ecl_thr_match_sd_dff_q_reg[0](.D(exu_n19330), .CLK(rclk), .Q(ecl_thr_match_de));
DFFPOSX1 ecl_fill_e2m_q_reg[0](.D(exu_n19328), .CLK(rclk), .Q(ecl_fill_trap_m));
DFFPOSX1 ecl_ttype_vld_e2m_q_reg[0](.D(exu_n19326), .CLK(rclk), .Q(ecl_early_ttype_vld_m));
DFFPOSX1 ecl_std_d2e_q_reg[0](.D(exu_n19324), .CLK(rclk), .Q(ecl_std_e));
DFFPOSX1 ecl_thr_match_ew_dff_q_reg[0](.D(exu_n19322), .CLK(rclk), .Q(ecl_thr_match_mw1));
DFFPOSX1 ecl_kill_rml_mw_q_reg[0](.D(exu_n19320), .CLK(rclk), .Q(ecl_kill_rml_w));
DFFPOSX1 ecl_flush_w_dff_q_reg[0](.D(exu_n19318), .CLK(rclk), .Q(ecl_flush_w1));
DFFPOSX1 ecl_flush_m2w_q_reg[0](.D(exu_n19316), .CLK(rclk), .Q(ecl_ifu_tlu_flush_w));
DFFPOSX1 ecl_early_flush_dff_q_reg[0](.D(exu_n19314), .CLK(rclk), .Q(ecl_part_early_flush_w));
DFFPOSX1 ecl_priv_trap_dff_q_reg[0](.D(exu_n19312), .CLK(rclk), .Q(ecl_tlu_priv_trap_w));
DFFPOSX1 ecl_inst_vld_ww1_q_reg[0](.D(exu_n19310), .CLK(rclk), .Q(ecl_inst_vld_w1));
DFFPOSX1 ecl_dff_range_check_other_e2m_q_reg[0](.D(exu_n19308), .CLK(rclk), .Q(ecl_ifu_exu_range_check_other_m));
DFFPOSX1 ecl_dff_range_check_other_d2e_q_reg[0](.D(exu_n19306), .CLK(rclk), .Q(ecl_ifu_exu_range_check_other_e));
DFFPOSX1 ecl_dff_range_check_jlret_e2m_q_reg[0](.D(exu_n19304), .CLK(rclk), .Q(ecl_ifu_exu_range_check_jlret_m));
DFFPOSX1 ecl_dff_range_check_jlret_d2e_q_reg[0](.D(exu_n19302), .CLK(rclk), .Q(ecl_ifu_exu_range_check_jlret_e));
DFFPOSX1 ecl_dff_misalign_addr_e2m_q_reg[0](.D(exu_n19300), .CLK(rclk), .Q(exu_tlu_misalign_addr_jmpl_rtn_m));
DFFPOSX1 ecl_dff_mem_invalid_e2m_q_reg[0](.D(exu_n19298), .CLK(rclk), .Q(ecl_alu_ecl_mem_addr_invalid_m_l));
DFFPOSX1 ecl_dff_addr_mask_d2e_q_reg[0](.D(exu_n19296), .CLK(rclk), .Q(ecl_addr_mask_e));
DFFPOSX1 ecl_restore_dff_q_reg[0](.D(exu_n19294), .CLK(rclk), .Q(ecl_restore_e));
DFFPOSX1 ecl_save_dff_q_reg[0](.D(exu_n19292), .CLK(rclk), .Q(ecl_save_e));
DFFPOSX1 ecl_rs2_31_e2m_q_reg[0](.D(exu_n19290), .CLK(rclk), .Q(ecl_rs2_data_31_m));
DFFPOSX1 ecl_mulsrs131_e2m_q_reg[0](.D(exu_n19288), .CLK(rclk), .Q(ecl_muls_rs1_31_m_l));
DFFPOSX1 ecl_zero_rs2_dff_q_reg[0](.D(exu_n19286), .CLK(rclk), .Q(ecl_div_zero_rs2_e));
DFFPOSX1 ecl_dff_muls_d2e_q_reg[0](.D(exu_n19284), .CLK(rclk), .Q(ecl_muls_e));
DFFPOSX1 ecl_c_used_dff_q_reg[0](.D(exu_n19282), .CLK(rclk), .Q(ecl_alu_cin_e));
DFFPOSX1 ecl_sub_dff_q_reg[0](.D(exu_n16320), .CLK(rclk), .Q(ecl_sub_e));
DFFPOSX1 ecl_dff_rs1_b0_m2w_q_reg[0](.D(exu_n19278), .CLK(rclk), .Q(ecl_div_yreg_data_31_g));
DFFPOSX1 ecl_casa_d2e_q_reg[0](.D(exu_n19276), .CLK(rclk), .Q(ecl_alu_casa_e));
DFFPOSX1 ecl_rs3_vld_d2e_q_reg[0](.D(exu_n19274), .CLK(rclk), .Q(ecl_rs3_vld_e));
DFFPOSX1 ecl_rs2_vld_d2e_q_reg[0](.D(exu_n19272), .CLK(rclk), .Q(ecl_rs2_vld_e));
DFFPOSX1 ecl_rs1_vld_d2e_q_reg[0](.D(exu_n19270), .CLK(rclk), .Q(ecl_rs1_vld_e));
DFFPOSX1 ecl_sethi_d2e_q_reg[0](.D(exu_n19268), .CLK(rclk), .Q(ecl_alu_sethi_inst_e));
DFFPOSX1 ecl_ldxa_dff_q_reg[0](.D(exu_n19266), .CLK(rclk), .Q(ecl_ldxa_g));
DFFPOSX1 ecl_dff_ialign_e2m_q_reg[0](.D(exu_n19264), .CLK(rclk), .Q(ecl_ialign_m));
DFFPOSX1 ecl_dff_ialign_d2e_q_reg[0](.D(exu_n19262), .CLK(rclk), .Q(ecl_ialign_e));
DFFPOSX1 ecl_dff_tagop_d2e_q_reg[0](.D(exu_n19260), .CLK(rclk), .Q(ecl_ifu_exu_tagop_e));
DFFPOSX1 ecl_dff_tv_d2e_q_reg[0](.D(exu_n19258), .CLK(rclk), .Q(ecl_ifu_exu_tv_e));
DFFPOSX1 ecl_dff_sel_sum_d2e_q_reg[0](.D(exu_n19256), .CLK(rclk), .Q(ecl_sel_sum_e));
DFFPOSX1 rml_cwp_cwp_output_queue_park_reg_q_reg[0](.D(exu_n19254), .CLK(rclk), .Q(rml_cwp_cwp_output_queue_pv[0]));
DFFPOSX1 rml_cwp_cwp_output_queue_park_reg_q_reg[1](.D(exu_n19253), .CLK(rclk), .Q(rml_cwp_cwp_output_queue_pv[1]));
DFFPOSX1 rml_cwp_cwp_output_queue_park_reg_q_reg[2](.D(exu_n19252), .CLK(rclk), .Q(rml_cwp_cwp_output_queue_pv[2]));
DFFPOSX1 rml_cwp_cwp_output_queue_park_reg_q_reg[3](.D(exu_n19251), .CLK(rclk), .Q(rml_cwp_cwp_output_queue_pv[3]));
DFFPOSX1 div_mul_data_dff_q_reg[0](.D(exu_n18551), .CLK(rclk), .Q(exu_mul_rs1_data[0]));
DFFPOSX1 div_mul_data_dff_q_reg[1](.D(exu_n18540), .CLK(rclk), .Q(exu_mul_rs1_data[1]));
DFFPOSX1 div_mul_data_dff_q_reg[2](.D(exu_n18529), .CLK(rclk), .Q(exu_mul_rs1_data[2]));
DFFPOSX1 div_mul_data_dff_q_reg[3](.D(exu_n18518), .CLK(rclk), .Q(exu_mul_rs1_data[3]));
DFFPOSX1 div_mul_data_dff_q_reg[4](.D(exu_n18507), .CLK(rclk), .Q(exu_mul_rs1_data[4]));
DFFPOSX1 div_mul_data_dff_q_reg[5](.D(exu_n18496), .CLK(rclk), .Q(exu_mul_rs1_data[5]));
DFFPOSX1 div_mul_data_dff_q_reg[6](.D(exu_n18485), .CLK(rclk), .Q(exu_mul_rs1_data[6]));
DFFPOSX1 div_mul_data_dff_q_reg[7](.D(exu_n18602), .CLK(rclk), .Q(exu_mul_rs1_data[7]));
DFFPOSX1 div_mul_data_dff_q_reg[8](.D(exu_n18591), .CLK(rclk), .Q(exu_mul_rs1_data[8]));
DFFPOSX1 div_mul_data_dff_q_reg[9](.D(exu_n18580), .CLK(rclk), .Q(exu_mul_rs1_data[9]));
DFFPOSX1 div_mul_data_dff_q_reg[10](.D(exu_n18569), .CLK(rclk), .Q(exu_mul_rs1_data[10]));
DFFPOSX1 div_mul_data_dff_q_reg[11](.D(exu_n18567), .CLK(rclk), .Q(exu_mul_rs1_data[11]));
DFFPOSX1 div_mul_data_dff_q_reg[12](.D(exu_n18566), .CLK(rclk), .Q(exu_mul_rs1_data[12]));
DFFPOSX1 div_mul_data_dff_q_reg[13](.D(exu_n18565), .CLK(rclk), .Q(exu_mul_rs1_data[13]));
DFFPOSX1 div_mul_data_dff_q_reg[14](.D(exu_n18564), .CLK(rclk), .Q(exu_mul_rs1_data[14]));
DFFPOSX1 div_mul_data_dff_q_reg[15](.D(exu_n18563), .CLK(rclk), .Q(exu_mul_rs1_data[15]));
DFFPOSX1 div_mul_data_dff_q_reg[16](.D(exu_n18562), .CLK(rclk), .Q(exu_mul_rs1_data[16]));
DFFPOSX1 div_mul_data_dff_q_reg[17](.D(exu_n18561), .CLK(rclk), .Q(exu_mul_rs1_data[17]));
DFFPOSX1 div_mul_data_dff_q_reg[18](.D(exu_n18560), .CLK(rclk), .Q(exu_mul_rs1_data[18]));
DFFPOSX1 div_mul_data_dff_q_reg[19](.D(exu_n18559), .CLK(rclk), .Q(exu_mul_rs1_data[19]));
DFFPOSX1 div_mul_data_dff_q_reg[20](.D(exu_n18558), .CLK(rclk), .Q(exu_mul_rs1_data[20]));
DFFPOSX1 div_mul_data_dff_q_reg[21](.D(exu_n18557), .CLK(rclk), .Q(exu_mul_rs1_data[21]));
DFFPOSX1 div_mul_data_dff_q_reg[22](.D(exu_n18556), .CLK(rclk), .Q(exu_mul_rs1_data[22]));
DFFPOSX1 div_mul_data_dff_q_reg[23](.D(exu_n18555), .CLK(rclk), .Q(exu_mul_rs1_data[23]));
DFFPOSX1 div_mul_data_dff_q_reg[24](.D(exu_n18554), .CLK(rclk), .Q(exu_mul_rs1_data[24]));
DFFPOSX1 div_mul_data_dff_q_reg[25](.D(exu_n18553), .CLK(rclk), .Q(exu_mul_rs1_data[25]));
DFFPOSX1 div_mul_data_dff_q_reg[26](.D(exu_n18552), .CLK(rclk), .Q(exu_mul_rs1_data[26]));
DFFPOSX1 div_mul_data_dff_q_reg[27](.D(exu_n18550), .CLK(rclk), .Q(exu_mul_rs1_data[27]));
DFFPOSX1 div_mul_data_dff_q_reg[28](.D(exu_n18549), .CLK(rclk), .Q(exu_mul_rs1_data[28]));
DFFPOSX1 div_mul_data_dff_q_reg[29](.D(exu_n18548), .CLK(rclk), .Q(exu_mul_rs1_data[29]));
DFFPOSX1 div_mul_data_dff_q_reg[30](.D(exu_n18547), .CLK(rclk), .Q(exu_mul_rs1_data[30]));
DFFPOSX1 div_mul_data_dff_q_reg[31](.D(exu_n18546), .CLK(rclk), .Q(exu_mul_rs1_data[31]));
DFFPOSX1 div_mul_data_dff_q_reg[32](.D(exu_n18545), .CLK(rclk), .Q(exu_mul_rs1_data[32]));
DFFPOSX1 div_mul_data_dff_q_reg[33](.D(exu_n18544), .CLK(rclk), .Q(exu_mul_rs1_data[33]));
DFFPOSX1 div_mul_data_dff_q_reg[34](.D(exu_n18543), .CLK(rclk), .Q(exu_mul_rs1_data[34]));
DFFPOSX1 div_mul_data_dff_q_reg[35](.D(exu_n18542), .CLK(rclk), .Q(exu_mul_rs1_data[35]));
DFFPOSX1 div_mul_data_dff_q_reg[36](.D(exu_n18541), .CLK(rclk), .Q(exu_mul_rs1_data[36]));
DFFPOSX1 div_mul_data_dff_q_reg[37](.D(exu_n18539), .CLK(rclk), .Q(exu_mul_rs1_data[37]));
DFFPOSX1 div_mul_data_dff_q_reg[38](.D(exu_n18538), .CLK(rclk), .Q(exu_mul_rs1_data[38]));
DFFPOSX1 div_mul_data_dff_q_reg[39](.D(exu_n18537), .CLK(rclk), .Q(exu_mul_rs1_data[39]));
DFFPOSX1 div_mul_data_dff_q_reg[40](.D(exu_n18536), .CLK(rclk), .Q(exu_mul_rs1_data[40]));
DFFPOSX1 div_mul_data_dff_q_reg[41](.D(exu_n18535), .CLK(rclk), .Q(exu_mul_rs1_data[41]));
DFFPOSX1 div_mul_data_dff_q_reg[42](.D(exu_n18534), .CLK(rclk), .Q(exu_mul_rs1_data[42]));
DFFPOSX1 div_mul_data_dff_q_reg[43](.D(exu_n18533), .CLK(rclk), .Q(exu_mul_rs1_data[43]));
DFFPOSX1 div_mul_data_dff_q_reg[44](.D(exu_n18532), .CLK(rclk), .Q(exu_mul_rs1_data[44]));
DFFPOSX1 div_mul_data_dff_q_reg[45](.D(exu_n18531), .CLK(rclk), .Q(exu_mul_rs1_data[45]));
DFFPOSX1 div_mul_data_dff_q_reg[46](.D(exu_n18530), .CLK(rclk), .Q(exu_mul_rs1_data[46]));
DFFPOSX1 div_mul_data_dff_q_reg[47](.D(exu_n18528), .CLK(rclk), .Q(exu_mul_rs1_data[47]));
DFFPOSX1 div_mul_data_dff_q_reg[48](.D(exu_n18527), .CLK(rclk), .Q(exu_mul_rs1_data[48]));
DFFPOSX1 div_mul_data_dff_q_reg[49](.D(exu_n18526), .CLK(rclk), .Q(exu_mul_rs1_data[49]));
DFFPOSX1 div_mul_data_dff_q_reg[50](.D(exu_n18525), .CLK(rclk), .Q(exu_mul_rs1_data[50]));
DFFPOSX1 div_mul_data_dff_q_reg[51](.D(exu_n18524), .CLK(rclk), .Q(exu_mul_rs1_data[51]));
DFFPOSX1 div_mul_data_dff_q_reg[52](.D(exu_n18523), .CLK(rclk), .Q(exu_mul_rs1_data[52]));
DFFPOSX1 div_mul_data_dff_q_reg[53](.D(exu_n18522), .CLK(rclk), .Q(exu_mul_rs1_data[53]));
DFFPOSX1 div_mul_data_dff_q_reg[54](.D(exu_n18521), .CLK(rclk), .Q(exu_mul_rs1_data[54]));
DFFPOSX1 div_mul_data_dff_q_reg[55](.D(exu_n18520), .CLK(rclk), .Q(exu_mul_rs1_data[55]));
DFFPOSX1 div_mul_data_dff_q_reg[56](.D(exu_n18519), .CLK(rclk), .Q(exu_mul_rs1_data[56]));
DFFPOSX1 div_mul_data_dff_q_reg[57](.D(exu_n18517), .CLK(rclk), .Q(exu_mul_rs1_data[57]));
DFFPOSX1 div_mul_data_dff_q_reg[58](.D(exu_n18516), .CLK(rclk), .Q(exu_mul_rs1_data[58]));
DFFPOSX1 div_mul_data_dff_q_reg[59](.D(exu_n18515), .CLK(rclk), .Q(exu_mul_rs1_data[59]));
DFFPOSX1 div_mul_data_dff_q_reg[60](.D(exu_n18514), .CLK(rclk), .Q(exu_mul_rs1_data[60]));
DFFPOSX1 div_mul_data_dff_q_reg[61](.D(exu_n18513), .CLK(rclk), .Q(exu_mul_rs1_data[61]));
DFFPOSX1 div_mul_data_dff_q_reg[62](.D(exu_n18512), .CLK(rclk), .Q(exu_mul_rs1_data[62]));
DFFPOSX1 div_mul_data_dff_q_reg[63](.D(exu_n18511), .CLK(rclk), .Q(exu_mul_rs1_data[63]));
DFFPOSX1 div_mul_data_dff_q_reg[64](.D(exu_n18510), .CLK(rclk), .Q(exu_mul_rs2_data[0]));
DFFPOSX1 div_mul_data_dff_q_reg[65](.D(exu_n18509), .CLK(rclk), .Q(exu_mul_rs2_data[1]));
DFFPOSX1 div_mul_data_dff_q_reg[66](.D(exu_n18508), .CLK(rclk), .Q(exu_mul_rs2_data[2]));
DFFPOSX1 div_mul_data_dff_q_reg[67](.D(exu_n18506), .CLK(rclk), .Q(exu_mul_rs2_data[3]));
DFFPOSX1 div_mul_data_dff_q_reg[68](.D(exu_n18505), .CLK(rclk), .Q(exu_mul_rs2_data[4]));
DFFPOSX1 div_mul_data_dff_q_reg[69](.D(exu_n18504), .CLK(rclk), .Q(exu_mul_rs2_data[5]));
DFFPOSX1 div_mul_data_dff_q_reg[70](.D(exu_n18503), .CLK(rclk), .Q(exu_mul_rs2_data[6]));
DFFPOSX1 div_mul_data_dff_q_reg[71](.D(exu_n18502), .CLK(rclk), .Q(exu_mul_rs2_data[7]));
DFFPOSX1 div_mul_data_dff_q_reg[72](.D(exu_n18501), .CLK(rclk), .Q(exu_mul_rs2_data[8]));
DFFPOSX1 div_mul_data_dff_q_reg[73](.D(exu_n18500), .CLK(rclk), .Q(exu_mul_rs2_data[9]));
DFFPOSX1 div_mul_data_dff_q_reg[74](.D(exu_n18499), .CLK(rclk), .Q(exu_mul_rs2_data[10]));
DFFPOSX1 div_mul_data_dff_q_reg[75](.D(exu_n18498), .CLK(rclk), .Q(exu_mul_rs2_data[11]));
DFFPOSX1 div_mul_data_dff_q_reg[76](.D(exu_n18497), .CLK(rclk), .Q(exu_mul_rs2_data[12]));
DFFPOSX1 div_mul_data_dff_q_reg[77](.D(exu_n18495), .CLK(rclk), .Q(exu_mul_rs2_data[13]));
DFFPOSX1 div_mul_data_dff_q_reg[78](.D(exu_n18494), .CLK(rclk), .Q(exu_mul_rs2_data[14]));
DFFPOSX1 div_mul_data_dff_q_reg[79](.D(exu_n18493), .CLK(rclk), .Q(exu_mul_rs2_data[15]));
DFFPOSX1 div_mul_data_dff_q_reg[80](.D(exu_n18492), .CLK(rclk), .Q(exu_mul_rs2_data[16]));
DFFPOSX1 div_mul_data_dff_q_reg[81](.D(exu_n18491), .CLK(rclk), .Q(exu_mul_rs2_data[17]));
DFFPOSX1 div_mul_data_dff_q_reg[82](.D(exu_n18490), .CLK(rclk), .Q(exu_mul_rs2_data[18]));
DFFPOSX1 div_mul_data_dff_q_reg[83](.D(exu_n18489), .CLK(rclk), .Q(exu_mul_rs2_data[19]));
DFFPOSX1 div_mul_data_dff_q_reg[84](.D(exu_n18488), .CLK(rclk), .Q(exu_mul_rs2_data[20]));
DFFPOSX1 div_mul_data_dff_q_reg[85](.D(exu_n18487), .CLK(rclk), .Q(exu_mul_rs2_data[21]));
DFFPOSX1 div_mul_data_dff_q_reg[86](.D(exu_n18486), .CLK(rclk), .Q(exu_mul_rs2_data[22]));
DFFPOSX1 div_mul_data_dff_q_reg[87](.D(exu_n18484), .CLK(rclk), .Q(exu_mul_rs2_data[23]));
DFFPOSX1 div_mul_data_dff_q_reg[88](.D(exu_n18483), .CLK(rclk), .Q(exu_mul_rs2_data[24]));
DFFPOSX1 div_mul_data_dff_q_reg[89](.D(exu_n18482), .CLK(rclk), .Q(exu_mul_rs2_data[25]));
DFFPOSX1 div_mul_data_dff_q_reg[90](.D(exu_n18481), .CLK(rclk), .Q(exu_mul_rs2_data[26]));
DFFPOSX1 div_mul_data_dff_q_reg[91](.D(exu_n18480), .CLK(rclk), .Q(exu_mul_rs2_data[27]));
DFFPOSX1 div_mul_data_dff_q_reg[92](.D(exu_n18479), .CLK(rclk), .Q(exu_mul_rs2_data[28]));
DFFPOSX1 div_mul_data_dff_q_reg[93](.D(exu_n18478), .CLK(rclk), .Q(exu_mul_rs2_data[29]));
DFFPOSX1 div_mul_data_dff_q_reg[94](.D(exu_n18477), .CLK(rclk), .Q(exu_mul_rs2_data[30]));
DFFPOSX1 div_mul_data_dff_q_reg[95](.D(exu_n18476), .CLK(rclk), .Q(exu_mul_rs2_data[31]));
DFFPOSX1 div_mul_data_dff_q_reg[96](.D(exu_n18475), .CLK(rclk), .Q(exu_mul_rs2_data[32]));
DFFPOSX1 div_mul_data_dff_q_reg[97](.D(exu_n18601), .CLK(rclk), .Q(exu_mul_rs2_data[33]));
DFFPOSX1 div_mul_data_dff_q_reg[98](.D(exu_n18600), .CLK(rclk), .Q(exu_mul_rs2_data[34]));
DFFPOSX1 div_mul_data_dff_q_reg[99](.D(exu_n18599), .CLK(rclk), .Q(exu_mul_rs2_data[35]));
DFFPOSX1 div_mul_data_dff_q_reg[100](.D(exu_n18598), .CLK(rclk), .Q(exu_mul_rs2_data[36]));
DFFPOSX1 div_mul_data_dff_q_reg[101](.D(exu_n18597), .CLK(rclk), .Q(exu_mul_rs2_data[37]));
DFFPOSX1 div_mul_data_dff_q_reg[102](.D(exu_n18596), .CLK(rclk), .Q(exu_mul_rs2_data[38]));
DFFPOSX1 div_mul_data_dff_q_reg[103](.D(exu_n18595), .CLK(rclk), .Q(exu_mul_rs2_data[39]));
DFFPOSX1 div_mul_data_dff_q_reg[104](.D(exu_n18594), .CLK(rclk), .Q(exu_mul_rs2_data[40]));
DFFPOSX1 div_mul_data_dff_q_reg[105](.D(exu_n18593), .CLK(rclk), .Q(exu_mul_rs2_data[41]));
DFFPOSX1 div_mul_data_dff_q_reg[106](.D(exu_n18592), .CLK(rclk), .Q(exu_mul_rs2_data[42]));
DFFPOSX1 div_mul_data_dff_q_reg[107](.D(exu_n18590), .CLK(rclk), .Q(exu_mul_rs2_data[43]));
DFFPOSX1 div_mul_data_dff_q_reg[108](.D(exu_n18589), .CLK(rclk), .Q(exu_mul_rs2_data[44]));
DFFPOSX1 div_mul_data_dff_q_reg[109](.D(exu_n18588), .CLK(rclk), .Q(exu_mul_rs2_data[45]));
DFFPOSX1 div_mul_data_dff_q_reg[110](.D(exu_n18587), .CLK(rclk), .Q(exu_mul_rs2_data[46]));
DFFPOSX1 div_mul_data_dff_q_reg[111](.D(exu_n18586), .CLK(rclk), .Q(exu_mul_rs2_data[47]));
DFFPOSX1 div_mul_data_dff_q_reg[112](.D(exu_n18585), .CLK(rclk), .Q(exu_mul_rs2_data[48]));
DFFPOSX1 div_mul_data_dff_q_reg[113](.D(exu_n18584), .CLK(rclk), .Q(exu_mul_rs2_data[49]));
DFFPOSX1 div_mul_data_dff_q_reg[114](.D(exu_n18583), .CLK(rclk), .Q(exu_mul_rs2_data[50]));
DFFPOSX1 div_mul_data_dff_q_reg[115](.D(exu_n18582), .CLK(rclk), .Q(exu_mul_rs2_data[51]));
DFFPOSX1 div_mul_data_dff_q_reg[116](.D(exu_n18581), .CLK(rclk), .Q(exu_mul_rs2_data[52]));
DFFPOSX1 div_mul_data_dff_q_reg[117](.D(exu_n18579), .CLK(rclk), .Q(exu_mul_rs2_data[53]));
DFFPOSX1 div_mul_data_dff_q_reg[118](.D(exu_n18578), .CLK(rclk), .Q(exu_mul_rs2_data[54]));
DFFPOSX1 div_mul_data_dff_q_reg[119](.D(exu_n18577), .CLK(rclk), .Q(exu_mul_rs2_data[55]));
DFFPOSX1 div_mul_data_dff_q_reg[120](.D(exu_n18576), .CLK(rclk), .Q(exu_mul_rs2_data[56]));
DFFPOSX1 div_mul_data_dff_q_reg[121](.D(exu_n18575), .CLK(rclk), .Q(exu_mul_rs2_data[57]));
DFFPOSX1 div_mul_data_dff_q_reg[122](.D(exu_n18574), .CLK(rclk), .Q(exu_mul_rs2_data[58]));
DFFPOSX1 div_mul_data_dff_q_reg[123](.D(exu_n18573), .CLK(rclk), .Q(exu_mul_rs2_data[59]));
DFFPOSX1 div_mul_data_dff_q_reg[124](.D(exu_n18572), .CLK(rclk), .Q(exu_mul_rs2_data[60]));
DFFPOSX1 div_mul_data_dff_q_reg[125](.D(exu_n18571), .CLK(rclk), .Q(exu_mul_rs2_data[61]));
DFFPOSX1 div_mul_data_dff_q_reg[126](.D(exu_n18570), .CLK(rclk), .Q(exu_mul_rs2_data[62]));
DFFPOSX1 div_mul_data_dff_q_reg[127](.D(exu_n18568), .CLK(rclk), .Q(exu_mul_rs2_data[63]));
XNOR2X1 exu_rml_canrestore_inc_U8(.A(exu_n16588), .B(rml_rml_ecl_canrestore_e[1]), .Y(exu_n18431));
XNOR2X1 exu_rml_canrestore_inc_U7(.A(exu_n15413), .B(exu_n18431), .Y(rml_rml_next_canrestore_e[1]));
XOR2X1 exu_rml_canrestore_inc_U3(.A(exu_n15074), .B(rml_rml_ecl_canrestore_e[2]), .Y(exu_n18427));
XOR2X1 exu_rml_canrestore_inc_U2(.A(rml_rml_next_canrestore_e[1]), .B(exu_n18427), .Y(rml_rml_next_canrestore_e[2]));
XNOR2X1 exu_rml_cansave_inc_U8(.A(exu_n16589), .B(rml_rml_ecl_cansave_e[1]), .Y(exu_n18426));
XNOR2X1 exu_rml_cansave_inc_U7(.A(exu_n15412), .B(exu_n18426), .Y(rml_rml_next_cansave_e[1]));
XOR2X1 exu_rml_cansave_inc_U3(.A(exu_n15073), .B(rml_rml_ecl_cansave_e[2]), .Y(exu_n18422));
XOR2X1 exu_rml_cansave_inc_U2(.A(rml_rml_next_cansave_e[1]), .B(exu_n18422), .Y(rml_rml_next_cansave_e[2]));
DFFPOSX1 rml_cwp_cwp_cmplt_dff_q_reg[0](.D(exu_n18421), .CLK(rclk), .Q(exu_tlu_cwp_retry));
DFFPOSX1 rml_cwp_cwp_cmplt_dff_q_reg[1](.D(exu_n18420), .CLK(rclk), .Q(exu_tlu_cwp_cmplt_tid[0]));
DFFPOSX1 rml_cwp_cwp_cmplt_dff_q_reg[2](.D(exu_n18419), .CLK(rclk), .Q(exu_tlu_cwp_cmplt_tid[1]));
DFFPOSX1 rml_cwp_cwp_cmplt_dff_q_reg[3](.D(exu_n18418), .CLK(rclk), .Q(exu_tlu_cwp_cmplt));
DFFPOSX1 rml_cwp_swap_done_dff_q_reg[0](.D(exu_n18416), .CLK(rclk), .Q(rml_ecl_swap_done[0]));
DFFPOSX1 rml_cwp_swap_done_dff_q_reg[1](.D(exu_n18415), .CLK(rclk), .Q(rml_ecl_swap_done[1]));
DFFPOSX1 rml_cwp_swap_done_dff_q_reg[2](.D(exu_n18414), .CLK(rclk), .Q(rml_ecl_swap_done[2]));
DFFPOSX1 rml_cwp_swap_done_dff_q_reg[3](.D(exu_n18413), .CLK(rclk), .Q(rml_ecl_swap_done[3]));
DFFPOSX1 rml_cwp_dff_swap_thr_q_reg[0](.D(exu_n18411), .CLK(rclk), .Q(rml_cwp_swap_thr[0]));
DFFPOSX1 rml_cwp_dff_swap_thr_q_reg[1](.D(exu_n18410), .CLK(rclk), .Q(rml_cwp_swap_thr[1]));
DFFPOSX1 rml_cwp_dff_swap_thr_q_reg[2](.D(exu_n18409), .CLK(rclk), .Q(rml_cwp_swap_thr[2]));
DFFPOSX1 rml_cwp_dff_swap_thr_q_reg[3](.D(exu_n18408), .CLK(rclk), .Q(rml_cwp_swap_thr[3]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr0_q_reg[2](.D(exu_n18381), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr0[2]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr0_q_reg[1](.D(exu_n18380), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr0[1]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr0_q_reg[0](.D(exu_n18379), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr0[0]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr1_q_reg[2](.D(exu_n18377), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr1[2]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr1_q_reg[1](.D(exu_n18376), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr1[1]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr1_q_reg[0](.D(exu_n18375), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr1[0]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr2_q_reg[2](.D(exu_n18373), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr2[2]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr2_q_reg[1](.D(exu_n18372), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr2[1]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr2_q_reg[0](.D(exu_n18371), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr2[0]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr3_q_reg[2](.D(exu_n18369), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr3[2]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr3_q_reg[1](.D(exu_n18368), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr3[1]));
DFFPOSX1 rml_lo_wstate_reg_dff_reg_thr3_q_reg[0](.D(exu_n18367), .CLK(rclk), .Q(rml_lo_wstate_reg_data_thr3[0]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr0_q_reg[2](.D(exu_n18341), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr0[2]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr0_q_reg[1](.D(exu_n18340), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr0[1]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr0_q_reg[0](.D(exu_n18339), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr0[0]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr1_q_reg[2](.D(exu_n18337), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr1[2]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr1_q_reg[1](.D(exu_n18336), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr1[1]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr1_q_reg[0](.D(exu_n18335), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr1[0]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr2_q_reg[2](.D(exu_n18333), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr2[2]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr2_q_reg[1](.D(exu_n18332), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr2[1]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr2_q_reg[0](.D(exu_n18331), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr2[0]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr3_q_reg[2](.D(exu_n18329), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr3[2]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr3_q_reg[1](.D(exu_n18328), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr3[1]));
DFFPOSX1 rml_hi_wstate_reg_dff_reg_thr3_q_reg[0](.D(exu_n18327), .CLK(rclk), .Q(rml_hi_wstate_reg_data_thr3[0]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr0_q_reg[2](.D(exu_n18297), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr0[2]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr0_q_reg[1](.D(exu_n18296), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr0[1]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr0_q_reg[0](.D(exu_n18295), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr0[0]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr1_q_reg[2](.D(exu_n18293), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr1[2]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr1_q_reg[1](.D(exu_n18292), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr1[1]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr1_q_reg[0](.D(exu_n18291), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr1[0]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr2_q_reg[2](.D(exu_n18289), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr2[2]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr2_q_reg[1](.D(exu_n18288), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr2[1]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr2_q_reg[0](.D(exu_n18287), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr2[0]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr3_q_reg[2](.D(exu_n18285), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr3[2]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr3_q_reg[1](.D(exu_n18284), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr3[1]));
DFFPOSX1 rml_cleanwin_reg_dff_reg_thr3_q_reg[0](.D(exu_n18283), .CLK(rclk), .Q(rml_cleanwin_reg_data_thr3[0]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr0_q_reg[2](.D(exu_n18253), .CLK(rclk), .Q(rml_otherwin_reg_data_thr0[2]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr0_q_reg[1](.D(exu_n18252), .CLK(rclk), .Q(rml_otherwin_reg_data_thr0[1]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr0_q_reg[0](.D(exu_n18251), .CLK(rclk), .Q(rml_otherwin_reg_data_thr0[0]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr1_q_reg[2](.D(exu_n18249), .CLK(rclk), .Q(rml_otherwin_reg_data_thr1[2]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr1_q_reg[1](.D(exu_n18248), .CLK(rclk), .Q(rml_otherwin_reg_data_thr1[1]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr1_q_reg[0](.D(exu_n18247), .CLK(rclk), .Q(rml_otherwin_reg_data_thr1[0]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr2_q_reg[2](.D(exu_n18245), .CLK(rclk), .Q(rml_otherwin_reg_data_thr2[2]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr2_q_reg[1](.D(exu_n18244), .CLK(rclk), .Q(rml_otherwin_reg_data_thr2[1]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr2_q_reg[0](.D(exu_n18243), .CLK(rclk), .Q(rml_otherwin_reg_data_thr2[0]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr3_q_reg[2](.D(exu_n18241), .CLK(rclk), .Q(rml_otherwin_reg_data_thr3[2]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr3_q_reg[1](.D(exu_n18240), .CLK(rclk), .Q(rml_otherwin_reg_data_thr3[1]));
DFFPOSX1 rml_otherwin_reg_dff_reg_thr3_q_reg[0](.D(exu_n18239), .CLK(rclk), .Q(rml_otherwin_reg_data_thr3[0]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr0_q_reg[2](.D(exu_n18209), .CLK(rclk), .Q(rml_canrestore_reg_data_thr0[2]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr0_q_reg[1](.D(exu_n18208), .CLK(rclk), .Q(rml_canrestore_reg_data_thr0[1]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr0_q_reg[0](.D(exu_n18207), .CLK(rclk), .Q(rml_canrestore_reg_data_thr0[0]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr1_q_reg[2](.D(exu_n18205), .CLK(rclk), .Q(rml_canrestore_reg_data_thr1[2]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr1_q_reg[1](.D(exu_n18204), .CLK(rclk), .Q(rml_canrestore_reg_data_thr1[1]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr1_q_reg[0](.D(exu_n18203), .CLK(rclk), .Q(rml_canrestore_reg_data_thr1[0]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr2_q_reg[2](.D(exu_n18201), .CLK(rclk), .Q(rml_canrestore_reg_data_thr2[2]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr2_q_reg[1](.D(exu_n18200), .CLK(rclk), .Q(rml_canrestore_reg_data_thr2[1]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr2_q_reg[0](.D(exu_n18199), .CLK(rclk), .Q(rml_canrestore_reg_data_thr2[0]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr3_q_reg[2](.D(exu_n18197), .CLK(rclk), .Q(rml_canrestore_reg_data_thr3[2]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr3_q_reg[1](.D(exu_n18196), .CLK(rclk), .Q(rml_canrestore_reg_data_thr3[1]));
DFFPOSX1 rml_canrestore_reg_dff_reg_thr3_q_reg[0](.D(exu_n18195), .CLK(rclk), .Q(rml_canrestore_reg_data_thr3[0]));
NAND2X1 exu_rml_cwp_irf_thr_mux_U5(.A(exu_n10783), .B(exu_n9775), .Y(rml_irf_cwpswap_tid_e[1]));
NAND2X1 exu_rml_cwp_irf_thr_mux_U4(.A(exu_n10782), .B(exu_n9774), .Y(rml_irf_cwpswap_tid_e[0]));
DFFPOSX1 rml_cwp_can_swap_flop_q_reg[0](.D(exu_n17980), .CLK(rclk), .Q(rml_cwp_just_swapped));
NAND2X1 exu_ecl_eccctl_ecc_rdlog_mux_U22(.A(exu_n17724), .B(exu_n9741), .Y(exu_ifu_err_reg_m[0]));
NAND2X1 exu_ecl_eccctl_ecc_rdlog_mux_U18(.A(exu_n17720), .B(exu_n9740), .Y(exu_ifu_err_reg_m[1]));
NAND2X1 exu_ecl_eccctl_ecc_rdlog_mux_U14(.A(exu_n17716), .B(exu_n9739), .Y(exu_ifu_err_reg_m[2]));
XOR2X1 exu_ecl_byplog_rs3h_w2_comp7_U13(.A(ecl_wb_byplog_rd_w2[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17704));
XNOR2X1 exu_ecl_byplog_rs3h_w2_comp7_U12(.A(ecl_wb_byplog_rd_w2[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17706));
XNOR2X1 exu_ecl_byplog_rs3h_w2_comp7_U11(.A(ecl_wb_byplog_tid_w2[0]), .B(ecl_tid_d[0]), .Y(exu_n17707));
XNOR2X1 exu_ecl_byplog_rs3h_w2_comp7_U7(.A(ecl_wb_byplog_tid_w2[1]), .B(ecl_tid_d[1]), .Y(exu_n17703));
XNOR2X1 exu_ecl_byplog_rs3h_w2_comp7_U5(.A(ecl_wb_byplog_rd_w2[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17701));
XNOR2X1 exu_ecl_byplog_rs3h_w2_comp7_U4(.A(ecl_wb_byplog_rd_w2[1]), .B(ecl_ifu_exu_rs3_d[1]), .Y(exu_n17702));
XOR2X1 exu_ecl_byplog_rs3h_w_comp7_U13(.A(ecl_ecl_irf_rd_w[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17693));
XNOR2X1 exu_ecl_byplog_rs3h_w_comp7_U12(.A(ecl_ecl_irf_rd_w[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17695));
XNOR2X1 exu_ecl_byplog_rs3h_w_comp7_U11(.A(ecl_ecl_irf_tid_w[0]), .B(ecl_tid_d[0]), .Y(exu_n17696));
XNOR2X1 exu_ecl_byplog_rs3h_w_comp7_U7(.A(ecl_ecl_irf_tid_w[1]), .B(ecl_tid_d[1]), .Y(exu_n17692));
XNOR2X1 exu_ecl_byplog_rs3h_w_comp7_U5(.A(ecl_ecl_irf_rd_w[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17690));
XNOR2X1 exu_ecl_byplog_rs3h_w_comp7_U4(.A(ecl_ecl_irf_rd_w[1]), .B(ecl_ifu_exu_rs3_d[1]), .Y(exu_n17691));
XOR2X1 exu_ecl_byplog_rs3_w2_comp7_U13(.A(ecl_wb_byplog_rd_w2[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17682));
XNOR2X1 exu_ecl_byplog_rs3_w2_comp7_U12(.A(ecl_wb_byplog_rd_w2[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17684));
XNOR2X1 exu_ecl_byplog_rs3_w2_comp7_U11(.A(ecl_wb_byplog_tid_w2[0]), .B(ecl_tid_d[0]), .Y(exu_n17685));
XNOR2X1 exu_ecl_byplog_rs3_w2_comp7_U8(.A(ecl_wb_byplog_rd_w2[0]), .B(ecl_ifu_exu_rs3_d[0]), .Y(exu_n17680));
XNOR2X1 exu_ecl_byplog_rs3_w2_comp7_U7(.A(ecl_wb_byplog_tid_w2[1]), .B(ecl_tid_d[1]), .Y(exu_n17681));
XNOR2X1 exu_ecl_byplog_rs3_w2_comp7_U5(.A(ecl_wb_byplog_rd_w2[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17678));
XNOR2X1 exu_ecl_byplog_rs3_w2_comp7_U4(.A(ecl_wb_byplog_rd_w2[1]), .B(ecl_ifu_exu_rs3_d[1]), .Y(exu_n17679));
XOR2X1 exu_ecl_byplog_rs3_w_comp7_U13(.A(ecl_ecl_irf_rd_w[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17670));
XNOR2X1 exu_ecl_byplog_rs3_w_comp7_U12(.A(ecl_ecl_irf_rd_w[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17672));
XNOR2X1 exu_ecl_byplog_rs3_w_comp7_U11(.A(ecl_ecl_irf_tid_w[0]), .B(ecl_tid_d[0]), .Y(exu_n17673));
XNOR2X1 exu_ecl_byplog_rs3_w_comp7_U8(.A(ecl_ecl_irf_rd_w[0]), .B(ecl_ifu_exu_rs3_d[0]), .Y(exu_n17668));
XNOR2X1 exu_ecl_byplog_rs3_w_comp7_U7(.A(ecl_ecl_irf_tid_w[1]), .B(ecl_tid_d[1]), .Y(exu_n17669));
XNOR2X1 exu_ecl_byplog_rs3_w_comp7_U5(.A(ecl_ecl_irf_rd_w[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17666));
XNOR2X1 exu_ecl_byplog_rs3_w_comp7_U4(.A(ecl_ecl_irf_rd_w[1]), .B(ecl_ifu_exu_rs3_d[1]), .Y(exu_n17667));
XOR2X1 exu_ecl_byplog_rs2_w2_comp7_U13(.A(ecl_wb_byplog_rd_w2[4]), .B(ecl_ifu_exu_rs2_d[4]), .Y(exu_n17658));
XNOR2X1 exu_ecl_byplog_rs2_w2_comp7_U12(.A(ecl_wb_byplog_rd_w2[3]), .B(ecl_ifu_exu_rs2_d[3]), .Y(exu_n17660));
XNOR2X1 exu_ecl_byplog_rs2_w2_comp7_U11(.A(ecl_wb_byplog_tid_w2[0]), .B(ecl_tid_d[0]), .Y(exu_n17661));
XNOR2X1 exu_ecl_byplog_rs2_w2_comp7_U8(.A(ecl_wb_byplog_rd_w2[0]), .B(ecl_ifu_exu_rs2_d[0]), .Y(exu_n17656));
XNOR2X1 exu_ecl_byplog_rs2_w2_comp7_U7(.A(ecl_wb_byplog_tid_w2[1]), .B(ecl_tid_d[1]), .Y(exu_n17657));
XNOR2X1 exu_ecl_byplog_rs2_w2_comp7_U5(.A(ecl_wb_byplog_rd_w2[2]), .B(ecl_ifu_exu_rs2_d[2]), .Y(exu_n17654));
XNOR2X1 exu_ecl_byplog_rs2_w2_comp7_U4(.A(ecl_wb_byplog_rd_w2[1]), .B(ecl_ifu_exu_rs2_d[1]), .Y(exu_n17655));
XOR2X1 exu_ecl_byplog_rs2_w_comp7_U13(.A(ecl_ecl_irf_rd_w[4]), .B(ecl_ifu_exu_rs2_d[4]), .Y(exu_n17646));
XNOR2X1 exu_ecl_byplog_rs2_w_comp7_U12(.A(ecl_ecl_irf_rd_w[3]), .B(ecl_ifu_exu_rs2_d[3]), .Y(exu_n17648));
XNOR2X1 exu_ecl_byplog_rs2_w_comp7_U11(.A(ecl_ecl_irf_tid_w[0]), .B(ecl_tid_d[0]), .Y(exu_n17649));
XNOR2X1 exu_ecl_byplog_rs2_w_comp7_U8(.A(ecl_ecl_irf_rd_w[0]), .B(ecl_ifu_exu_rs2_d[0]), .Y(exu_n17644));
XNOR2X1 exu_ecl_byplog_rs2_w_comp7_U7(.A(ecl_ecl_irf_tid_w[1]), .B(ecl_tid_d[1]), .Y(exu_n17645));
XNOR2X1 exu_ecl_byplog_rs2_w_comp7_U5(.A(ecl_ecl_irf_rd_w[2]), .B(ecl_ifu_exu_rs2_d[2]), .Y(exu_n17642));
XNOR2X1 exu_ecl_byplog_rs2_w_comp7_U4(.A(ecl_ecl_irf_rd_w[1]), .B(ecl_ifu_exu_rs2_d[1]), .Y(exu_n17643));
XOR2X1 exu_ecl_byplog_rs1_w2_comp7_U13(.A(ecl_wb_byplog_rd_w2[4]), .B(ecl_ifu_exu_rs1_d[4]), .Y(exu_n17634));
XNOR2X1 exu_ecl_byplog_rs1_w2_comp7_U12(.A(ecl_wb_byplog_rd_w2[3]), .B(ecl_ifu_exu_rs1_d[3]), .Y(exu_n17636));
XNOR2X1 exu_ecl_byplog_rs1_w2_comp7_U11(.A(ecl_wb_byplog_tid_w2[0]), .B(ecl_tid_d[0]), .Y(exu_n17637));
XNOR2X1 exu_ecl_byplog_rs1_w2_comp7_U8(.A(ecl_wb_byplog_rd_w2[0]), .B(ecl_ifu_exu_rs1_d[0]), .Y(exu_n17632));
XNOR2X1 exu_ecl_byplog_rs1_w2_comp7_U7(.A(ecl_wb_byplog_tid_w2[1]), .B(ecl_tid_d[1]), .Y(exu_n17633));
XNOR2X1 exu_ecl_byplog_rs1_w2_comp7_U5(.A(ecl_wb_byplog_rd_w2[2]), .B(ecl_ifu_exu_rs1_d[2]), .Y(exu_n17630));
XNOR2X1 exu_ecl_byplog_rs1_w2_comp7_U4(.A(ecl_wb_byplog_rd_w2[1]), .B(ecl_ifu_exu_rs1_d[1]), .Y(exu_n17631));
DFFPOSX1 ecl_divcntl_cnt6_cntr_dff_q_reg[0](.D(exu_n17625), .CLK(rclk), .Q(ecl_divcntl_cntr[0]));
DFFPOSX1 ecl_divcntl_cnt6_cntr_dff_q_reg[1](.D(exu_n17624), .CLK(rclk), .Q(ecl_divcntl_cntr[1]));
DFFPOSX1 ecl_divcntl_cnt6_cntr_dff_q_reg[2](.D(exu_n17623), .CLK(rclk), .Q(ecl_divcntl_cntr[2]));
DFFPOSX1 ecl_divcntl_cnt6_cntr_dff_q_reg[3](.D(exu_n17622), .CLK(rclk), .Q(ecl_divcntl_cntr[3]));
DFFPOSX1 ecl_divcntl_cnt6_cntr_dff_q_reg[4](.D(exu_n17621), .CLK(rclk), .Q(ecl_divcntl_cntr[4]));
DFFPOSX1 ecl_divcntl_cnt6_cntr_dff_q_reg[5](.D(exu_n17620), .CLK(rclk), .Q(ecl_divcntl_cntr[5]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[0](.D(exu_n17505), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[0]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[1](.D(exu_n17504), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[1]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[2](.D(exu_n17503), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[2]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[3](.D(exu_n17502), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[3]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[4](.D(exu_n17501), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[4]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[5](.D(exu_n17500), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[5]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[6](.D(exu_n17499), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[6]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[7](.D(exu_n17498), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[7]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[8](.D(exu_n17497), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[8]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[9](.D(exu_n17496), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[9]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[10](.D(exu_n17495), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[10]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[11](.D(exu_n17494), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[11]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[12](.D(exu_n17493), .CLK(rclk), .Q(rml_cwp_swap_slot3_data[12]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[13](.D(exu_n17492), .CLK(rclk), .Q(rml_cwp_swap_slot3_state_valid[0]));
DFFPOSX1 rml_cwp_slot3_data_dff_q_reg[14](.D(exu_n17491), .CLK(rclk), .Q(rml_cwp_swap_slot3_state[1]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[0](.D(exu_n17490), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[0]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[1](.D(exu_n17489), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[1]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[2](.D(exu_n17488), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[2]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[3](.D(exu_n17487), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[3]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[4](.D(exu_n17486), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[4]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[5](.D(exu_n17485), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[5]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[6](.D(exu_n17484), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[6]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[7](.D(exu_n17483), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[7]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[8](.D(exu_n17482), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[8]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[9](.D(exu_n17481), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[9]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[10](.D(exu_n17480), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[10]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[11](.D(exu_n17479), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[11]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[12](.D(exu_n17478), .CLK(rclk), .Q(rml_cwp_swap_slot2_data[12]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[13](.D(exu_n17477), .CLK(rclk), .Q(rml_cwp_swap_slot2_state_valid[0]));
DFFPOSX1 rml_cwp_slot2_data_dff_q_reg[14](.D(exu_n17475), .CLK(rclk), .Q(rml_cwp_swap_slot2_state[1]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[0](.D(exu_n17474), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[0]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[1](.D(exu_n17473), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[1]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[2](.D(exu_n17472), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[2]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[3](.D(exu_n17471), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[3]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[4](.D(exu_n17470), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[4]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[5](.D(exu_n17469), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[5]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[6](.D(exu_n17468), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[6]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[7](.D(exu_n17467), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[7]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[8](.D(exu_n17466), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[8]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[9](.D(exu_n17465), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[9]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[10](.D(exu_n17464), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[10]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[11](.D(exu_n17463), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[11]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[12](.D(exu_n17462), .CLK(rclk), .Q(rml_cwp_swap_slot1_data[12]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[13](.D(exu_n17461), .CLK(rclk), .Q(rml_cwp_swap_slot1_state_valid[0]));
DFFPOSX1 rml_cwp_slot1_data_dff_q_reg[14](.D(exu_n17460), .CLK(rclk), .Q(rml_cwp_swap_slot1_state[1]));
INVX1 exu_U1(.A(exu_n15351), .Y(exu_n15983));
INVX1 exu_U2(.A(ecl_shiftop_e[2]), .Y(exu_n16153));
INVX1 exu_U3(.A(exu_n15351), .Y(exu_n15984));
INVX1 exu_U4(.A(ecl_shiftop_e[2]), .Y(exu_n16152));
AND2X1 exu_U5(.A(alu_logic_rs1_data_bf1[63]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[63]));
AND2X1 exu_U6(.A(alu_logic_rs1_data_bf1[62]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[62]));
AND2X1 exu_U7(.A(alu_logic_rs1_data_bf1[61]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[61]));
AND2X1 exu_U8(.A(alu_logic_rs1_data_bf1[60]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[60]));
AND2X1 exu_U9(.A(alu_logic_rs1_data_bf1[59]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[59]));
AND2X1 exu_U10(.A(alu_logic_rs1_data_bf1[58]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[58]));
AND2X1 exu_U11(.A(alu_logic_rs1_data_bf1[57]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[57]));
AND2X1 exu_U12(.A(alu_logic_rs1_data_bf1[56]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[56]));
AND2X1 exu_U13(.A(alu_logic_rs1_data_bf1[55]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[55]));
AND2X1 exu_U14(.A(alu_logic_rs1_data_bf1[54]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[54]));
AND2X1 exu_U15(.A(alu_logic_rs1_data_bf1[53]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[53]));
AND2X1 exu_U16(.A(alu_logic_rs1_data_bf1[52]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[52]));
AND2X1 exu_U17(.A(alu_logic_rs1_data_bf1[51]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[51]));
AND2X1 exu_U18(.A(alu_logic_rs1_data_bf1[50]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[50]));
AND2X1 exu_U19(.A(alu_logic_rs1_data_bf1[49]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[49]));
AND2X1 exu_U20(.A(alu_logic_rs1_data_bf1[48]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[48]));
AND2X1 exu_U21(.A(alu_logic_rs1_data_bf1[47]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[47]));
AND2X1 exu_U22(.A(alu_logic_rs1_data_bf1[46]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[46]));
AND2X1 exu_U23(.A(alu_logic_rs1_data_bf1[45]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[45]));
AND2X1 exu_U24(.A(alu_logic_rs1_data_bf1[44]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[44]));
AND2X1 exu_U25(.A(alu_logic_rs1_data_bf1[43]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[43]));
AND2X1 exu_U26(.A(alu_logic_rs1_data_bf1[42]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[42]));
AND2X1 exu_U27(.A(alu_logic_rs1_data_bf1[41]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[41]));
AND2X1 exu_U28(.A(alu_logic_rs1_data_bf1[40]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[40]));
AND2X1 exu_U29(.A(alu_logic_rs1_data_bf1[39]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[39]));
AND2X1 exu_U30(.A(alu_logic_rs1_data_bf1[38]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[38]));
AND2X1 exu_U31(.A(alu_logic_rs1_data_bf1[37]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[37]));
AND2X1 exu_U32(.A(alu_logic_rs1_data_bf1[36]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[36]));
AND2X1 exu_U33(.A(alu_logic_rs1_data_bf1[35]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[35]));
AND2X1 exu_U34(.A(alu_logic_rs1_data_bf1[34]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[34]));
AND2X1 exu_U35(.A(alu_logic_rs1_data_bf1[33]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[33]));
AND2X1 exu_U36(.A(alu_logic_rs1_data_bf1[32]), .B(ecl_enshift_e), .Y(shft_shifter_input_b1[32]));
AND2X1 exu_U37(.A(alu_logic_rs1_data_bf1[31]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[31]));
AND2X1 exu_U38(.A(alu_logic_rs1_data_bf1[30]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[30]));
AND2X1 exu_U39(.A(alu_logic_rs1_data_bf1[29]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[29]));
AND2X1 exu_U40(.A(alu_logic_rs1_data_bf1[28]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[28]));
AND2X1 exu_U41(.A(alu_logic_rs1_data_bf1[27]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[27]));
AND2X1 exu_U42(.A(alu_logic_rs1_data_bf1[26]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[26]));
AND2X1 exu_U43(.A(alu_logic_rs1_data_bf1[24]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[24]));
AND2X1 exu_U44(.A(alu_logic_rs1_data_bf1[23]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[23]));
AND2X1 exu_U45(.A(alu_logic_rs1_data_bf1[22]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[22]));
AND2X1 exu_U46(.A(alu_logic_rs1_data_bf1[21]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[21]));
AND2X1 exu_U47(.A(alu_logic_rs1_data_bf1[20]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[20]));
AND2X1 exu_U48(.A(alu_logic_rs1_data_bf1[19]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[19]));
AND2X1 exu_U49(.A(alu_logic_rs1_data_bf1[18]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[18]));
AND2X1 exu_U50(.A(alu_logic_rs1_data_bf1[17]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[17]));
AND2X1 exu_U51(.A(alu_logic_rs1_data_bf1[16]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[16]));
INVX1 exu_U52(.A(ecl_shft_extendbit_e), .Y(exu_n16188));
INVX1 exu_U53(.A(ecl_shft_extendbit_e), .Y(exu_n16187));
AND2X1 exu_U54(.A(exu_n4434), .B(exu_n9288), .Y(shft_rshifterinput_b1[55]));
AND2X1 exu_U55(.A(exu_n4430), .B(exu_n9274), .Y(shft_rshifterinput_b1[39]));
AND2X1 exu_U56(.A(exu_n4456), .B(exu_n9289), .Y(shft_rshifterinput_b1[54]));
AND2X1 exu_U57(.A(exu_n4433), .B(exu_n9275), .Y(shft_rshifterinput_b1[38]));
AND2X1 exu_U58(.A(exu_n4455), .B(exu_n9290), .Y(shft_rshifterinput_b1[53]));
AND2X1 exu_U59(.A(exu_n4436), .B(exu_n9276), .Y(shft_rshifterinput_b1[37]));
AND2X1 exu_U60(.A(exu_n4449), .B(exu_n9291), .Y(shft_rshifterinput_b1[52]));
AND2X1 exu_U61(.A(exu_n4439), .B(exu_n9277), .Y(shft_rshifterinput_b1[36]));
AND2X1 exu_U62(.A(exu_n4454), .B(exu_n9282), .Y(shft_rshifterinput_b1[61]));
AND2X1 exu_U63(.A(exu_n4470), .B(exu_n9299), .Y(shft_rshifterinput_b1[45]));
AND2X1 exu_U64(.A(exu_n4458), .B(exu_n9286), .Y(shft_rshifterinput_b1[57]));
AND2X1 exu_U65(.A(exu_n4425), .B(exu_n9272), .Y(shft_rshifterinput_b1[41]));
AND2X1 exu_U66(.A(alu_logic_rs1_data_bf1[25]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[25]));
AND2X1 exu_U67(.A(exu_n4446), .B(exu_n9295), .Y(shft_rshifterinput_b1[49]));
AND2X1 exu_U68(.A(exu_n4461), .B(exu_n9292), .Y(shft_rshifterinput_b1[33]));
AND2X1 exu_U69(.A(exu_n4445), .B(exu_n9279), .Y(shft_rshifterinput_b1[63]));
AND2X1 exu_U70(.A(exu_n4464), .B(exu_n9297), .Y(shft_rshifterinput_b1[47]));
AND2X1 exu_U71(.A(exu_n4428), .B(exu_n9284), .Y(shft_rshifterinput_b1[59]));
AND2X1 exu_U72(.A(exu_n4476), .B(exu_n9301), .Y(shft_rshifterinput_b1[43]));
AND2X1 exu_U73(.A(exu_n4465), .B(exu_n9293), .Y(shft_rshifterinput_b1[51]));
AND2X1 exu_U74(.A(exu_n4442), .B(exu_n9278), .Y(shft_rshifterinput_b1[35]));
AND2X1 exu_U75(.A(exu_n4440), .B(exu_n9283), .Y(shft_rshifterinput_b1[60]));
AND2X1 exu_U76(.A(exu_n4473), .B(exu_n9300), .Y(shft_rshifterinput_b1[44]));
AND2X1 exu_U77(.A(exu_n4483), .B(exu_n9287), .Y(shft_rshifterinput_b1[56]));
AND2X1 exu_U78(.A(exu_n4427), .B(exu_n9273), .Y(shft_rshifterinput_b1[40]));
AND2X1 exu_U79(.A(exu_n4431), .B(exu_n9296), .Y(shft_rshifterinput_b1[48]));
AND2X1 exu_U80(.A(exu_n4482), .B(exu_n9303), .Y(shft_rshifterinput_b1[32]));
AND2X1 exu_U81(.A(exu_n4448), .B(exu_n9280), .Y(shft_rshifterinput_b1[62]));
AND2X1 exu_U82(.A(exu_n4467), .B(exu_n9298), .Y(shft_rshifterinput_b1[46]));
AND2X1 exu_U83(.A(exu_n4459), .B(exu_n9285), .Y(shft_rshifterinput_b1[58]));
AND2X1 exu_U84(.A(exu_n4479), .B(exu_n9302), .Y(shft_rshifterinput_b1[42]));
AND2X1 exu_U85(.A(exu_n4468), .B(exu_n9294), .Y(shft_rshifterinput_b1[50]));
AND2X1 exu_U86(.A(exu_n4451), .B(exu_n9281), .Y(shft_rshifterinput_b1[34]));
AND2X1 exu_U87(.A(exu_n3040), .B(exu_n8120), .Y(exu_n27759));
AND2X1 exu_U88(.A(exu_n16154), .B(alu_logic_rs1_data_bf1[31]), .Y(ecl_n105));
AND2X1 exu_U89(.A(exu_n3042), .B(exu_n8122), .Y(exu_n27765));
AND2X1 exu_U90(.A(exu_n3044), .B(exu_n8124), .Y(exu_n27771));
AND2X1 exu_U91(.A(exu_n3046), .B(exu_n8126), .Y(exu_n27777));
AND2X1 exu_U92(.A(exu_n3048), .B(exu_n8128), .Y(exu_n27784));
AND2X1 exu_U93(.A(exu_n3050), .B(exu_n8130), .Y(exu_n27790));
AND2X1 exu_U94(.A(exu_n3052), .B(exu_n8132), .Y(exu_n27796));
AND2X1 exu_U95(.A(exu_n3054), .B(exu_n8134), .Y(exu_n27802));
AND2X1 exu_U96(.A(exu_n3056), .B(exu_n8136), .Y(exu_n27808));
AND2X1 exu_U97(.A(exu_n3058), .B(exu_n8138), .Y(exu_n27814));
AND2X1 exu_U98(.A(exu_n3060), .B(exu_n8140), .Y(exu_n27820));
AND2X1 exu_U99(.A(exu_n3062), .B(exu_n8142), .Y(exu_n27826));
AND2X1 exu_U100(.A(exu_n3064), .B(exu_n8144), .Y(exu_n27832));
AND2X1 exu_U101(.A(exu_n3066), .B(exu_n8146), .Y(exu_n27838));
AND2X1 exu_U102(.A(exu_n2699), .B(exu_n7730), .Y(exu_n26753));
AND2X1 exu_U103(.A(exu_n3068), .B(exu_n8148), .Y(exu_n27845));
AND2X1 exu_U104(.A(exu_n2700), .B(exu_n7730), .Y(exu_n26757));
AND2X1 exu_U105(.A(exu_n3070), .B(exu_n8150), .Y(exu_n27851));
AND2X1 exu_U106(.A(exu_n2703), .B(exu_n7735), .Y(exu_n26761));
AND2X1 exu_U107(.A(exu_n2708), .B(exu_n7740), .Y(exu_n26764));
AND2X1 exu_U108(.A(exu_n2712), .B(exu_n7744), .Y(exu_n26772));
AND2X1 exu_U109(.A(exu_n2715), .B(exu_n7747), .Y(exu_n26776));
AND2X1 exu_U110(.A(exu_n2718), .B(exu_n7750), .Y(exu_n26780));
AND2X1 exu_U111(.A(exu_n2721), .B(exu_n7753), .Y(exu_n26784));
AND2X1 exu_U112(.A(exu_n2724), .B(exu_n7756), .Y(exu_n26788));
AND2X1 exu_U113(.A(exu_n2727), .B(exu_n7759), .Y(exu_n26792));
AND2X1 exu_U114(.A(exu_n2730), .B(exu_n7762), .Y(exu_n26796));
AND2X1 exu_U115(.A(exu_n2733), .B(exu_n7765), .Y(exu_n26800));
AND2X1 exu_U116(.A(exu_n2736), .B(exu_n7768), .Y(exu_n26804));
AND2X1 exu_U117(.A(exu_n2739), .B(exu_n7771), .Y(exu_n26808));
AND2X1 exu_U118(.A(exu_n2743), .B(exu_n7775), .Y(exu_n26816));
AND2X1 exu_U119(.A(exu_n2746), .B(exu_n7779), .Y(exu_n26820));
AND2X1 exu_U120(.A(exu_n2747), .B(exu_n7781), .Y(exu_n26826));
AND2X1 exu_U121(.A(exu_n2750), .B(exu_n7785), .Y(exu_n26831));
AND2X1 exu_U122(.A(exu_n2751), .B(exu_n7789), .Y(exu_n26836));
AND2X1 exu_U123(.A(exu_n2752), .B(exu_n7793), .Y(exu_n26841));
AND2X1 exu_U124(.A(exu_n2753), .B(exu_n7797), .Y(exu_n26846));
AND2X1 exu_U125(.A(exu_n2754), .B(exu_n7801), .Y(exu_n26851));
AND2X1 exu_U126(.A(exu_n2755), .B(exu_n7805), .Y(exu_n26856));
AND2X1 exu_U127(.A(exu_n2756), .B(exu_n7809), .Y(exu_n26861));
AND2X1 exu_U128(.A(exu_n2758), .B(exu_n7814), .Y(exu_n26870));
AND2X1 exu_U129(.A(exu_n2759), .B(exu_n7818), .Y(exu_n26875));
AND2X1 exu_U130(.A(exu_n2760), .B(exu_n7822), .Y(exu_n26880));
AND2X1 exu_U131(.A(exu_n2761), .B(exu_n7826), .Y(exu_n26885));
AND2X1 exu_U132(.A(exu_n2762), .B(exu_n7830), .Y(exu_n26890));
AND2X1 exu_U133(.A(exu_n2763), .B(exu_n7834), .Y(exu_n26895));
AND2X1 exu_U134(.A(exu_n2764), .B(exu_n7838), .Y(exu_n26900));
AND2X1 exu_U135(.A(exu_n2765), .B(exu_n7842), .Y(exu_n26905));
AND2X1 exu_U136(.A(exu_n3088), .B(exu_n7846), .Y(exu_n26911));
AND2X1 exu_U137(.A(exu_n3089), .B(exu_n7847), .Y(exu_n26915));
AND2X1 exu_U138(.A(exu_n3090), .B(exu_n7849), .Y(exu_n26923));
AND2X1 exu_U139(.A(alu_logic_rs1_data_bf1[15]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[15]));
AND2X1 exu_U140(.A(exu_n3091), .B(exu_n7850), .Y(exu_n26927));
AND2X1 exu_U141(.A(alu_logic_rs1_data_bf1[14]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[14]));
AND2X1 exu_U142(.A(exu_n3092), .B(exu_n7851), .Y(exu_n26931));
AND2X1 exu_U143(.A(alu_logic_rs1_data_bf1[13]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[13]));
AND2X1 exu_U144(.A(exu_n3093), .B(exu_n7852), .Y(exu_n26935));
AND2X1 exu_U145(.A(alu_logic_rs1_data_bf1[12]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[12]));
AND2X1 exu_U146(.A(exu_n3096), .B(exu_n7855), .Y(exu_n26947));
AND2X1 exu_U147(.A(exu_n3094), .B(exu_n7853), .Y(exu_n26939));
AND2X1 exu_U148(.A(alu_logic_rs1_data_bf1[11]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[11]));
AND2X1 exu_U149(.A(alu_logic_rs1_data_bf1[9]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[9]));
AND2X1 exu_U150(.A(exu_n3095), .B(exu_n7854), .Y(exu_n26943));
AND2X1 exu_U151(.A(alu_logic_rs1_data_bf1[10]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[10]));
AND2X1 exu_U152(.A(exu_n3097), .B(exu_n7856), .Y(exu_n26951));
AND2X1 exu_U153(.A(alu_logic_rs1_data_bf1[8]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[8]));
AND2X1 exu_U154(.A(exu_n3098), .B(exu_n7857), .Y(exu_n26955));
AND2X1 exu_U155(.A(alu_logic_rs1_data_bf1[7]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[7]));
AND2X1 exu_U156(.A(exu_n3099), .B(exu_n7858), .Y(exu_n26959));
AND2X1 exu_U157(.A(alu_logic_rs1_data_bf1[6]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[6]));
AND2X1 exu_U158(.A(exu_n3100), .B(exu_n7860), .Y(exu_n26967));
AND2X1 exu_U159(.A(exu_n15002), .B(exu_n8160), .Y(exu_n26745));
AND2X1 exu_U160(.A(alu_logic_rs1_data_bf1[5]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[5]));
AND2X1 exu_U161(.A(exu_n3101), .B(exu_n7863), .Y(exu_n26971));
AND2X1 exu_U162(.A(exu_n15003), .B(exu_n8161), .Y(exu_n26749));
INVX1 exu_U163(.A(div_input_data_e[66]), .Y(exu_n16517));
AND2X1 exu_U164(.A(alu_logic_rs1_data_bf1[4]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[4]));
AND2X1 exu_U165(.A(exu_n3102), .B(exu_n7866), .Y(exu_n26975));
AND2X1 exu_U166(.A(exu_n15004), .B(exu_n8162), .Y(exu_n26769));
AND2X1 exu_U167(.A(exu_n3103), .B(exu_n7869), .Y(exu_n26979));
AND2X1 exu_U168(.A(exu_n15005), .B(exu_n8163), .Y(exu_n26813));
AND2X1 exu_U169(.A(exu_n15008), .B(exu_n8154), .Y(exu_n26992));
AND2X1 exu_U170(.A(exu_n15000), .B(exu_n7721), .Y(exu_n26736));
AND2X1 exu_U171(.A(exu_n7), .B(exu_n8166), .Y(exu_n26963));
AND2X1 exu_U172(.A(exu_n15006), .B(exu_n8152), .Y(exu_n26984));
AND2X1 exu_U173(.A(exu_n15010), .B(exu_n8156), .Y(exu_n27000));
AND2X1 exu_U174(.A(exu_n5), .B(exu_n8164), .Y(exu_n26866));
AND2X1 exu_U175(.A(exu_n15009), .B(exu_n8155), .Y(exu_n26996));
AND2X1 exu_U176(.A(exu_n15001), .B(exu_n8159), .Y(exu_n26741));
AND2X1 exu_U177(.A(exu_n8), .B(exu_n8167), .Y(exu_n27008));
AND2X1 exu_U178(.A(exu_n15007), .B(exu_n8153), .Y(exu_n26988));
AND2X1 exu_U179(.A(exu_n15011), .B(exu_n8157), .Y(exu_n27004));
AND2X1 exu_U180(.A(exu_n6), .B(exu_n8165), .Y(exu_n26919));
INVX1 exu_U181(.A(div_input_data_e[68]), .Y(exu_n16519));
INVX1 exu_U182(.A(ecl_rd_m[0]), .Y(exu_n16561));
INVX1 exu_U183(.A(ecl_wb_byplog_rd_g2[0]), .Y(exu_n16559));
OR2X1 exu_U184(.A(div_adderin2[22]), .B(exu_n15907), .Y(div_spr_n97));
OR2X1 exu_U185(.A(exu_n13167), .B(exu_n14454), .Y(shft_lshift16_b1[63]));
AND2X1 exu_U186(.A(exu_n3041), .B(exu_n8121), .Y(exu_n27758));
OR2X1 exu_U187(.A(exu_n13168), .B(exu_n14455), .Y(shft_lshift16_b1[62]));
AND2X1 exu_U188(.A(exu_n3043), .B(exu_n8123), .Y(exu_n27764));
OR2X1 exu_U189(.A(exu_n13169), .B(exu_n14456), .Y(shft_lshift16_b1[61]));
AND2X1 exu_U190(.A(exu_n3045), .B(exu_n8125), .Y(exu_n27770));
OR2X1 exu_U191(.A(exu_n13170), .B(exu_n14457), .Y(shft_lshift16_b1[60]));
AND2X1 exu_U192(.A(exu_n3047), .B(exu_n8127), .Y(exu_n27776));
OR2X1 exu_U193(.A(exu_n13171), .B(exu_n14458), .Y(shft_lshift16_b1[59]));
AND2X1 exu_U194(.A(exu_n3049), .B(exu_n8129), .Y(exu_n27783));
OR2X1 exu_U195(.A(exu_n13172), .B(exu_n14459), .Y(shft_lshift16_b1[58]));
AND2X1 exu_U196(.A(exu_n3051), .B(exu_n8131), .Y(exu_n27789));
OR2X1 exu_U197(.A(exu_n13173), .B(exu_n14460), .Y(shft_lshift16_b1[57]));
AND2X1 exu_U198(.A(exu_n3053), .B(exu_n8133), .Y(exu_n27795));
OR2X1 exu_U199(.A(exu_n13174), .B(exu_n14461), .Y(shft_lshift16_b1[56]));
AND2X1 exu_U200(.A(exu_n3055), .B(exu_n8135), .Y(exu_n27801));
OR2X1 exu_U201(.A(exu_n13175), .B(exu_n14462), .Y(shft_lshift16_b1[55]));
AND2X1 exu_U202(.A(exu_n3057), .B(exu_n8137), .Y(exu_n27807));
OR2X1 exu_U203(.A(exu_n13176), .B(exu_n14463), .Y(shft_lshift16_b1[54]));
AND2X1 exu_U204(.A(exu_n3059), .B(exu_n8139), .Y(exu_n27813));
OR2X1 exu_U205(.A(exu_n13177), .B(exu_n14464), .Y(shft_lshift16_b1[53]));
AND2X1 exu_U206(.A(exu_n3061), .B(exu_n8141), .Y(exu_n27819));
OR2X1 exu_U207(.A(exu_n13178), .B(exu_n14465), .Y(shft_lshift16_b1[52]));
AND2X1 exu_U208(.A(exu_n3063), .B(exu_n8143), .Y(exu_n27825));
OR2X1 exu_U209(.A(exu_n13179), .B(exu_n14466), .Y(shft_lshift16_b1[51]));
AND2X1 exu_U210(.A(exu_n3065), .B(exu_n8145), .Y(exu_n27831));
OR2X1 exu_U211(.A(exu_n13180), .B(exu_n14467), .Y(shft_lshift16_b1[50]));
AND2X1 exu_U212(.A(exu_n3067), .B(exu_n8147), .Y(exu_n27837));
OR2X1 exu_U213(.A(exu_n12982), .B(exu_n14266), .Y(shft_rshift16_b1[63]));
AND2X1 exu_U214(.A(exu_n2702), .B(exu_n7727), .Y(exu_n26752));
OR2X1 exu_U215(.A(exu_n13181), .B(exu_n14468), .Y(shft_lshift16_b1[49]));
AND2X1 exu_U216(.A(exu_n3069), .B(exu_n8149), .Y(exu_n27844));
OR2X1 exu_U217(.A(exu_n12983), .B(exu_n14267), .Y(shft_rshift16_b1[62]));
AND2X1 exu_U218(.A(exu_n2702), .B(exu_n7732), .Y(exu_n26756));
OR2X1 exu_U219(.A(exu_n13182), .B(exu_n14469), .Y(shft_lshift16_b1[48]));
AND2X1 exu_U220(.A(exu_n3071), .B(exu_n8151), .Y(exu_n27850));
OR2X1 exu_U221(.A(exu_n12984), .B(exu_n14268), .Y(shft_rshift16_b1[61]));
AND2X1 exu_U222(.A(exu_n2705), .B(exu_n7737), .Y(exu_n26760));
OR2X1 exu_U223(.A(exu_n27859), .B(exu_n14470), .Y(shft_lshift16_b1[47]));
AND2X1 exu_U224(.A(exu_n3072), .B(exu_n8152), .Y(exu_n27856));
OR2X1 exu_U225(.A(exu_n12985), .B(exu_n14269), .Y(shft_rshift16_b1[60]));
AND2X1 exu_U226(.A(exu_n2706), .B(exu_n7777), .Y(exu_n26765));
OR2X1 exu_U227(.A(exu_n27863), .B(exu_n14471), .Y(shft_lshift16_b1[46]));
AND2X1 exu_U228(.A(exu_n3073), .B(exu_n8153), .Y(exu_n27860));
OR2X1 exu_U229(.A(exu_n12987), .B(exu_n14271), .Y(shft_rshift16_b1[59]));
AND2X1 exu_U230(.A(exu_n2710), .B(exu_n7777), .Y(exu_n26773));
OR2X1 exu_U231(.A(exu_n27867), .B(exu_n14472), .Y(shft_lshift16_b1[45]));
AND2X1 exu_U232(.A(exu_n3074), .B(exu_n8154), .Y(exu_n27864));
OR2X1 exu_U233(.A(exu_n12988), .B(exu_n14272), .Y(shft_rshift16_b1[58]));
AND2X1 exu_U234(.A(exu_n2713), .B(exu_n7777), .Y(exu_n26777));
OR2X1 exu_U235(.A(exu_n27871), .B(exu_n14473), .Y(shft_lshift16_b1[44]));
AND2X1 exu_U236(.A(exu_n3075), .B(exu_n8155), .Y(exu_n27868));
OR2X1 exu_U237(.A(exu_n12989), .B(exu_n14273), .Y(shft_rshift16_b1[57]));
AND2X1 exu_U238(.A(exu_n2716), .B(exu_n7777), .Y(exu_n26781));
OR2X1 exu_U239(.A(exu_n27875), .B(exu_n14474), .Y(shft_lshift16_b1[43]));
AND2X1 exu_U240(.A(exu_n3076), .B(exu_n8156), .Y(exu_n27872));
OR2X1 exu_U241(.A(exu_n12990), .B(exu_n14274), .Y(shft_rshift16_b1[56]));
AND2X1 exu_U242(.A(exu_n2719), .B(exu_n7777), .Y(exu_n26785));
OR2X1 exu_U243(.A(exu_n27879), .B(exu_n14475), .Y(shft_lshift16_b1[42]));
AND2X1 exu_U244(.A(exu_n3077), .B(exu_n8157), .Y(exu_n27876));
OR2X1 exu_U245(.A(exu_n12991), .B(exu_n14275), .Y(shft_rshift16_b1[55]));
AND2X1 exu_U246(.A(exu_n2722), .B(exu_n7777), .Y(exu_n26789));
OR2X1 exu_U247(.A(exu_n27883), .B(exu_n14476), .Y(shft_lshift16_b1[41]));
AND2X1 exu_U248(.A(exu_n3078), .B(exu_n8158), .Y(exu_n27880));
OR2X1 exu_U249(.A(exu_n12992), .B(exu_n14276), .Y(shft_rshift16_b1[54]));
AND2X1 exu_U250(.A(exu_n2725), .B(exu_n7777), .Y(exu_n26793));
OR2X1 exu_U251(.A(exu_n27887), .B(exu_n14477), .Y(shft_lshift16_b1[40]));
AND2X1 exu_U252(.A(exu_n3079), .B(exu_n8159), .Y(exu_n27884));
OR2X1 exu_U253(.A(exu_n12993), .B(exu_n14277), .Y(shft_rshift16_b1[53]));
AND2X1 exu_U254(.A(exu_n2728), .B(exu_n7777), .Y(exu_n26797));
OR2X1 exu_U255(.A(exu_n27892), .B(exu_n14478), .Y(shft_lshift16_b1[39]));
AND2X1 exu_U256(.A(exu_n3080), .B(exu_n8160), .Y(exu_n27889));
OR2X1 exu_U257(.A(exu_n12994), .B(exu_n14278), .Y(shft_rshift16_b1[52]));
AND2X1 exu_U258(.A(exu_n2731), .B(exu_n7777), .Y(exu_n26801));
OR2X1 exu_U259(.A(exu_n27896), .B(exu_n14479), .Y(shft_lshift16_b1[38]));
AND2X1 exu_U260(.A(exu_n3081), .B(exu_n8161), .Y(exu_n27893));
OR2X1 exu_U261(.A(exu_n12995), .B(exu_n14279), .Y(shft_rshift16_b1[51]));
AND2X1 exu_U262(.A(exu_n2734), .B(exu_n7777), .Y(exu_n26805));
OR2X1 exu_U263(.A(exu_n27900), .B(exu_n14480), .Y(shft_lshift16_b1[37]));
AND2X1 exu_U264(.A(exu_n3082), .B(exu_n8162), .Y(exu_n27897));
OR2X1 exu_U265(.A(exu_n12996), .B(exu_n14280), .Y(shft_rshift16_b1[50]));
AND2X1 exu_U266(.A(exu_n2737), .B(exu_n7777), .Y(exu_n26809));
OR2X1 exu_U267(.A(exu_n27904), .B(exu_n14481), .Y(shft_lshift16_b1[36]));
AND2X1 exu_U268(.A(exu_n3083), .B(exu_n8163), .Y(exu_n27901));
OR2X1 exu_U269(.A(exu_n12998), .B(exu_n14282), .Y(shft_rshift16_b1[49]));
AND2X1 exu_U270(.A(exu_n2741), .B(exu_n7777), .Y(exu_n26817));
OR2X1 exu_U271(.A(exu_n27908), .B(exu_n14482), .Y(shft_lshift16_b1[35]));
AND2X1 exu_U272(.A(exu_n3084), .B(exu_n8164), .Y(exu_n27905));
OR2X1 exu_U273(.A(exu_n12999), .B(exu_n14283), .Y(shft_rshift16_b1[48]));
AND2X1 exu_U274(.A(exu_n2744), .B(exu_n7777), .Y(exu_n26821));
OR2X1 exu_U275(.A(exu_n27912), .B(exu_n14483), .Y(shft_lshift16_b1[34]));
AND2X1 exu_U276(.A(exu_n3085), .B(exu_n8165), .Y(exu_n27909));
OR2X1 exu_U277(.A(exu_n13000), .B(exu_n14284), .Y(shft_rshift16_b1[47]));
AND2X1 exu_U278(.A(exu_n2749), .B(exu_n7783), .Y(exu_n26825));
OR2X1 exu_U279(.A(exu_n27916), .B(exu_n14484), .Y(shft_lshift16_b1[33]));
AND2X1 exu_U280(.A(exu_n3086), .B(exu_n8166), .Y(exu_n27913));
OR2X1 exu_U281(.A(exu_n13001), .B(exu_n14285), .Y(shft_rshift16_b1[46]));
AND2X1 exu_U282(.A(exu_n2766), .B(exu_n7787), .Y(exu_n26830));
OR2X1 exu_U283(.A(exu_n27920), .B(exu_n14485), .Y(shft_lshift16_b1[32]));
AND2X1 exu_U284(.A(exu_n3087), .B(exu_n8167), .Y(exu_n27917));
OR2X1 exu_U285(.A(exu_n13002), .B(exu_n14286), .Y(shft_rshift16_b1[45]));
AND2X1 exu_U286(.A(exu_n2766), .B(exu_n7791), .Y(exu_n26835));
AND2X1 exu_U287(.A(exu_n3088), .B(exu_n8168), .Y(exu_n27921));
OR2X1 exu_U288(.A(exu_n13003), .B(exu_n14287), .Y(shft_rshift16_b1[44]));
AND2X1 exu_U289(.A(exu_n2766), .B(exu_n7795), .Y(exu_n26840));
AND2X1 exu_U290(.A(exu_n3089), .B(exu_n8169), .Y(exu_n27924));
OR2X1 exu_U291(.A(exu_n13004), .B(exu_n14288), .Y(shft_rshift16_b1[43]));
AND2X1 exu_U292(.A(exu_n2766), .B(exu_n7799), .Y(exu_n26845));
AND2X1 exu_U293(.A(exu_n3090), .B(exu_n8170), .Y(exu_n27928));
OR2X1 exu_U294(.A(exu_n13005), .B(exu_n14289), .Y(shft_rshift16_b1[42]));
AND2X1 exu_U295(.A(exu_n2766), .B(exu_n7803), .Y(exu_n26850));
AND2X1 exu_U296(.A(exu_n3091), .B(exu_n8171), .Y(exu_n27931));
OR2X1 exu_U297(.A(exu_n13006), .B(exu_n14290), .Y(shft_rshift16_b1[41]));
AND2X1 exu_U298(.A(exu_n2766), .B(exu_n7807), .Y(exu_n26855));
AND2X1 exu_U299(.A(exu_n3092), .B(exu_n8172), .Y(exu_n27934));
OR2X1 exu_U300(.A(exu_n13007), .B(exu_n14291), .Y(shft_rshift16_b1[40]));
AND2X1 exu_U301(.A(exu_n2766), .B(exu_n7811), .Y(exu_n26860));
AND2X1 exu_U302(.A(exu_n3093), .B(exu_n8173), .Y(exu_n27937));
OR2X1 exu_U303(.A(exu_n13009), .B(exu_n14293), .Y(shft_rshift16_b1[39]));
AND2X1 exu_U304(.A(exu_n2766), .B(exu_n7816), .Y(exu_n26869));
AND2X1 exu_U305(.A(exu_n3094), .B(exu_n8174), .Y(exu_n27940));
OR2X1 exu_U306(.A(exu_n13010), .B(exu_n14294), .Y(shft_rshift16_b1[38]));
AND2X1 exu_U307(.A(exu_n2766), .B(exu_n7820), .Y(exu_n26874));
AND2X1 exu_U308(.A(exu_n3095), .B(exu_n8175), .Y(exu_n27943));
OR2X1 exu_U309(.A(exu_n13011), .B(exu_n14295), .Y(shft_rshift16_b1[37]));
AND2X1 exu_U310(.A(exu_n2766), .B(exu_n7824), .Y(exu_n26879));
AND2X1 exu_U311(.A(exu_n3096), .B(exu_n8176), .Y(exu_n27946));
OR2X1 exu_U312(.A(exu_n13012), .B(exu_n14296), .Y(shft_rshift16_b1[36]));
AND2X1 exu_U313(.A(exu_n2766), .B(exu_n7828), .Y(exu_n26884));
AND2X1 exu_U314(.A(exu_n3097), .B(exu_n8177), .Y(exu_n27949));
OR2X1 exu_U315(.A(exu_n13013), .B(exu_n14297), .Y(shft_rshift16_b1[35]));
AND2X1 exu_U316(.A(exu_n2766), .B(exu_n7832), .Y(exu_n26889));
AND2X1 exu_U317(.A(exu_n3098), .B(exu_n8178), .Y(exu_n27952));
OR2X1 exu_U318(.A(exu_n13014), .B(exu_n14298), .Y(shft_rshift16_b1[34]));
AND2X1 exu_U319(.A(exu_n2766), .B(exu_n7836), .Y(exu_n26894));
AND2X1 exu_U320(.A(exu_n3099), .B(exu_n8179), .Y(exu_n27955));
OR2X1 exu_U321(.A(exu_n13015), .B(exu_n14299), .Y(shft_rshift16_b1[33]));
AND2X1 exu_U322(.A(exu_n2766), .B(exu_n7840), .Y(exu_n26899));
AND2X1 exu_U323(.A(exu_n3100), .B(exu_n8180), .Y(exu_n27959));
OR2X1 exu_U324(.A(exu_n13016), .B(exu_n14300), .Y(shft_rshift16_b1[32]));
AND2X1 exu_U325(.A(exu_n2766), .B(exu_n7844), .Y(exu_n26904));
AND2X1 exu_U326(.A(exu_n3101), .B(exu_n8181), .Y(exu_n27962));
OR2X1 exu_U327(.A(exu_n13017), .B(exu_n14301), .Y(shft_rshift16_b1[31]));
AND2X1 exu_U328(.A(exu_n2767), .B(exu_n7817), .Y(exu_n26910));
AND2X1 exu_U329(.A(exu_n3102), .B(exu_n8182), .Y(exu_n27965));
OR2X1 exu_U330(.A(exu_n13018), .B(exu_n14302), .Y(shft_rshift16_b1[30]));
AND2X1 exu_U331(.A(exu_n2768), .B(exu_n7821), .Y(exu_n26914));
AND2X1 exu_U332(.A(exu_n3103), .B(exu_n8183), .Y(exu_n27968));
OR2X1 exu_U333(.A(exu_n13020), .B(exu_n14304), .Y(shft_rshift16_b1[29]));
AND2X1 exu_U334(.A(exu_n2770), .B(exu_n7825), .Y(exu_n26922));
OR2X1 exu_U335(.A(exu_n13021), .B(exu_n14305), .Y(shft_rshift16_b1[28]));
AND2X1 exu_U336(.A(exu_n2771), .B(exu_n7769), .Y(exu_n26926));
OR2X1 exu_U337(.A(exu_n13022), .B(exu_n14306), .Y(shft_rshift16_b1[27]));
AND2X1 exu_U338(.A(exu_n2772), .B(exu_n7780), .Y(exu_n26930));
OR2X1 exu_U339(.A(exu_n13023), .B(exu_n14307), .Y(shft_rshift16_b1[26]));
AND2X1 exu_U340(.A(exu_n2773), .B(exu_n7792), .Y(exu_n26934));
OR2X1 exu_U341(.A(exu_n13026), .B(exu_n14310), .Y(shft_rshift16_b1[23]));
AND2X1 exu_U342(.A(exu_n2776), .B(exu_n7728), .Y(exu_n26946));
OR2X1 exu_U343(.A(exu_n13024), .B(exu_n14308), .Y(shft_rshift16_b1[25]));
AND2X1 exu_U344(.A(exu_n2774), .B(exu_n7808), .Y(exu_n26938));
OR2X1 exu_U345(.A(exu_n13025), .B(exu_n14309), .Y(shft_rshift16_b1[24]));
AND2X1 exu_U346(.A(exu_n2775), .B(exu_n7804), .Y(exu_n26942));
OR2X1 exu_U347(.A(exu_n13027), .B(exu_n14311), .Y(shft_rshift16_b1[22]));
AND2X1 exu_U348(.A(exu_n2777), .B(exu_n7733), .Y(exu_n26950));
INVX1 exu_U349(.A(div_input_data_e[67]), .Y(exu_n16518));
OR2X1 exu_U350(.A(exu_n13028), .B(exu_n14312), .Y(shft_rshift16_b1[21]));
AND2X1 exu_U351(.A(exu_n2778), .B(exu_n7738), .Y(exu_n26954));
OR2X1 exu_U352(.A(exu_n13029), .B(exu_n14313), .Y(shft_rshift16_b1[20]));
AND2X1 exu_U353(.A(exu_n2779), .B(exu_n7741), .Y(exu_n26958));
OR2X1 exu_U354(.A(exu_n13031), .B(exu_n14315), .Y(shft_rshift16_b1[19]));
AND2X1 exu_U355(.A(exu_n2781), .B(exu_n7862), .Y(exu_n26966));
OR2X1 exu_U356(.A(exu_n12980), .B(exu_n14264), .Y(shft_rshift16_b1[7]));
AND2X1 exu_U357(.A(exu_n2697), .B(exu_n7724), .Y(exu_n26744));
OR2X1 exu_U358(.A(exu_n13032), .B(exu_n14316), .Y(shft_rshift16_b1[18]));
AND2X1 exu_U359(.A(exu_n2782), .B(exu_n7865), .Y(exu_n26970));
OR2X1 exu_U360(.A(exu_n12981), .B(exu_n14265), .Y(shft_rshift16_b1[6]));
AND2X1 exu_U361(.A(exu_n2698), .B(exu_n7725), .Y(exu_n26748));
OR2X1 exu_U362(.A(exu_n13033), .B(exu_n14317), .Y(shft_rshift16_b1[17]));
AND2X1 exu_U363(.A(exu_n2783), .B(exu_n7868), .Y(exu_n26974));
OR2X1 exu_U364(.A(exu_n12986), .B(exu_n14270), .Y(shft_rshift16_b1[5]));
AND2X1 exu_U365(.A(exu_n2709), .B(exu_n7742), .Y(exu_n26768));
AND2X1 exu_U366(.A(alu_logic_rs1_data_bf1[3]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[3]));
OR2X1 exu_U367(.A(exu_n13034), .B(exu_n14318), .Y(shft_rshift16_b1[16]));
AND2X1 exu_U368(.A(exu_n2784), .B(exu_n7870), .Y(exu_n26978));
OR2X1 exu_U369(.A(exu_n12997), .B(exu_n14281), .Y(shft_rshift16_b1[4]));
AND2X1 exu_U370(.A(exu_n2740), .B(exu_n7773), .Y(exu_n26812));
AND2X1 exu_U371(.A(alu_logic_rs1_data_bf1[2]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[2]));
OR2X1 exu_U372(.A(exu_n13037), .B(exu_n14321), .Y(shft_rshift16_b1[13]));
AND2X1 exu_U373(.A(exu_n2787), .B(exu_n7873), .Y(exu_n26991));
OR2X1 exu_U374(.A(exu_n12978), .B(exu_n14262), .Y(shft_rshift16_b1[9]));
AND2X1 exu_U375(.A(exu_n2695), .B(exu_n7722), .Y(exu_n26735));
OR2X1 exu_U376(.A(exu_n13030), .B(exu_n14314), .Y(shft_rshift16_b1[1]));
AND2X1 exu_U377(.A(exu_n2780), .B(exu_n7859), .Y(exu_n26962));
OR2X1 exu_U378(.A(exu_n13035), .B(exu_n14319), .Y(shft_rshift16_b1[15]));
AND2X1 exu_U379(.A(exu_n2785), .B(exu_n7871), .Y(exu_n26983));
OR2X1 exu_U380(.A(exu_n13039), .B(exu_n14323), .Y(shft_rshift16_b1[11]));
AND2X1 exu_U381(.A(exu_n2789), .B(exu_n7875), .Y(exu_n26999));
OR2X1 exu_U382(.A(exu_n13008), .B(exu_n14292), .Y(shft_rshift16_b1[3]));
AND2X1 exu_U383(.A(exu_n2757), .B(exu_n7813), .Y(exu_n26865));
AND2X1 exu_U384(.A(alu_logic_rs1_data_bf1[1]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[1]));
OR2X1 exu_U385(.A(exu_n13038), .B(exu_n14322), .Y(shft_rshift16_b1[12]));
AND2X1 exu_U386(.A(exu_n2788), .B(exu_n7874), .Y(exu_n26995));
OR2X1 exu_U387(.A(exu_n12979), .B(exu_n14263), .Y(shft_rshift16_b1[8]));
AND2X1 exu_U388(.A(exu_n2696), .B(exu_n7723), .Y(exu_n26740));
OR2X1 exu_U389(.A(exu_n13041), .B(exu_n14325), .Y(shft_rshift16_b1[0]));
AND2X1 exu_U390(.A(exu_n2791), .B(exu_n7877), .Y(exu_n27007));
OR2X1 exu_U391(.A(exu_n13036), .B(exu_n14320), .Y(shft_rshift16_b1[14]));
AND2X1 exu_U392(.A(exu_n2786), .B(exu_n7872), .Y(exu_n26987));
OR2X1 exu_U393(.A(exu_n13040), .B(exu_n14324), .Y(shft_rshift16_b1[10]));
AND2X1 exu_U394(.A(exu_n2790), .B(exu_n7876), .Y(exu_n27003));
OR2X1 exu_U395(.A(exu_n13019), .B(exu_n14303), .Y(shft_rshift16_b1[2]));
AND2X1 exu_U396(.A(exu_n2769), .B(exu_n7848), .Y(exu_n26918));
OR2X1 exu_U397(.A(exu_n16561), .B(ecl_ifu_exu_rs1_d[0]), .Y(exu_n16655));
OR2X1 exu_U398(.A(exu_n16559), .B(ecl_ifu_exu_rs2_d[0]), .Y(exu_n16683));
OR2X1 exu_U399(.A(exu_n16561), .B(ecl_ifu_exu_rs2_d[0]), .Y(exu_n16711));
OR2X1 exu_U400(.A(exu_n16559), .B(ecl_ifu_exu_rs1_d[0]), .Y(exu_n16627));
INVX1 exu_U401(.A(ecl_ifu_exu_rs1_d[1]), .Y(exu_n16399));
OR2X1 exu_U402(.A(exu_n16561), .B(ecl_ifu_exu_rs3_d[0]), .Y(exu_n17431));
INVX1 exu_U403(.A(ecl_rd_m[1]), .Y(exu_n16562));
OR2X1 exu_U404(.A(exu_n16559), .B(ecl_ifu_exu_rs3_d[0]), .Y(exu_n17403));
INVX1 exu_U405(.A(ecl_wb_byplog_rd_g2[1]), .Y(exu_n16560));
OR2X1 exu_U406(.A(div_adderin2[46]), .B(exu_n15882), .Y(div_spr_n45));
OR2X1 exu_U407(.A(div_adderin2[38]), .B(exu_n15891), .Y(div_spr_n63));
OR2X1 exu_U408(.A(div_adderin2[62]), .B(exu_n15864), .Y(div_spr_n9));
OR2X1 exu_U409(.A(div_adderin2[54]), .B(exu_n15873), .Y(div_spr_n27));
OR2X1 exu_U410(.A(div_adderin2[8]), .B(exu_n15861), .Y(div_spr_n1));
OR2X1 exu_U411(.A(div_adderin2[4]), .B(exu_n15878), .Y(div_spr_n17));
OR2X1 exu_U412(.A(div_adderin2[29]), .B(exu_n15900), .Y(div_spr_n81));
OR2X1 exu_U413(.A(div_adderin2[26]), .B(exu_n15903), .Y(div_spr_n89));
OR2X1 exu_U414(.A(div_adderin2[15]), .B(exu_n15915), .Y(div_spr_n113));
OR2X1 exu_U415(.A(div_adderin2[13]), .B(exu_n15917), .Y(div_spr_n117));
OR2X1 exu_U416(.A(div_adderin2[11]), .B(exu_n15919), .Y(div_spr_n121));
OR2X1 exu_U417(.A(div_adderin2[9]), .B(exu_n15860), .Y(div_spr_n125));
OR2X1 exu_U418(.A(div_adderin2[0]), .B(exu_n15859), .Y(div_spr_n105));
OR2X1 exu_U419(.A(div_adderin2[18]), .B(exu_n15912), .Y(div_spr_n107));
OR2X1 exu_U420(.A(div_adderin2[17]), .B(exu_n15913), .Y(div_spr_n109));
OR2X1 exu_U421(.A(div_adderin2[16]), .B(exu_n15914), .Y(div_spr_n111));
OR2X1 exu_U422(.A(div_adderin2[20]), .B(exu_n15909), .Y(div_spr_n101));
OR2X1 exu_U423(.A(div_adderin2[19]), .B(exu_n15911), .Y(div_spr_n103));
OR2X1 exu_U424(.A(div_adderin2[21]), .B(exu_n15908), .Y(div_spr_n99));
AND2X1 exu_U425(.A(exu_n3883), .B(exu_n8962), .Y(div_z_in[23]));
AND2X1 exu_U426(.A(exu_n3108), .B(exu_n8188), .Y(exu_n27993));
AND2X1 exu_U427(.A(ecl_shiftop_e_0), .B(ecl_shiftop_e[2]), .Y(ecl_n104));
AND2X1 exu_U428(.A(exu_n3110), .B(exu_n8190), .Y(exu_n27999));
INVX1 exu_U429(.A(div_input_data_e[126]), .Y(exu_n16550));
AND2X1 exu_U430(.A(exu_n3112), .B(exu_n8192), .Y(exu_n28005));
INVX1 exu_U431(.A(div_input_data_e[125]), .Y(exu_n16549));
AND2X1 exu_U432(.A(exu_n2801), .B(exu_n7886), .Y(exu_n27038));
AND2X1 exu_U433(.A(exu_n3114), .B(exu_n8194), .Y(exu_n28011));
INVX1 exu_U434(.A(div_input_data_e[124]), .Y(exu_n16548));
AND2X1 exu_U435(.A(exu_n3117), .B(exu_n8197), .Y(exu_n28020));
INVX1 exu_U436(.A(div_input_data_e[123]), .Y(exu_n16547));
AND2X1 exu_U437(.A(exu_n2803), .B(exu_n7886), .Y(exu_n27044));
AND2X1 exu_U438(.A(exu_n3119), .B(exu_n8199), .Y(exu_n28026));
INVX1 exu_U439(.A(div_input_data_e[122]), .Y(exu_n16546));
AND2X1 exu_U440(.A(exu_n2806), .B(exu_n7890), .Y(exu_n27055));
AND2X1 exu_U441(.A(exu_n3121), .B(exu_n8201), .Y(exu_n28032));
INVX1 exu_U442(.A(div_input_data_e[121]), .Y(exu_n16545));
AND2X1 exu_U443(.A(exu_n2807), .B(exu_n7892), .Y(exu_n27060));
AND2X1 exu_U444(.A(exu_n3123), .B(exu_n8203), .Y(exu_n28038));
INVX1 exu_U445(.A(div_input_data_e[120]), .Y(exu_n16544));
AND2X1 exu_U446(.A(exu_n2810), .B(exu_n7891), .Y(exu_n27040));
AND2X1 exu_U447(.A(exu_n3125), .B(exu_n8205), .Y(exu_n28044));
INVX1 exu_U448(.A(div_input_data_e[119]), .Y(exu_n16543));
AND2X1 exu_U449(.A(exu_n2809), .B(exu_n7895), .Y(exu_n27068));
AND2X1 exu_U450(.A(exu_n3127), .B(exu_n8207), .Y(exu_n28050));
INVX1 exu_U451(.A(div_input_data_e[118]), .Y(exu_n16542));
AND2X1 exu_U452(.A(exu_n2811), .B(exu_n7896), .Y(exu_n27073));
AND2X1 exu_U453(.A(exu_n3129), .B(exu_n8209), .Y(exu_n28056));
INVX1 exu_U454(.A(div_input_data_e[117]), .Y(exu_n16541));
AND2X1 exu_U455(.A(exu_n2813), .B(exu_n7897), .Y(exu_n27078));
AND2X1 exu_U456(.A(exu_n3131), .B(exu_n8211), .Y(exu_n28062));
INVX1 exu_U457(.A(div_input_data_e[116]), .Y(exu_n16540));
AND2X1 exu_U458(.A(exu_n2815), .B(exu_n7898), .Y(exu_n27083));
AND2X1 exu_U459(.A(exu_n3133), .B(exu_n8213), .Y(exu_n28068));
INVX1 exu_U460(.A(div_input_data_e[115]), .Y(exu_n16539));
AND2X1 exu_U461(.A(exu_n2817), .B(exu_n7899), .Y(exu_n27088));
AND2X1 exu_U462(.A(exu_n3135), .B(exu_n8215), .Y(exu_n28074));
INVX1 exu_U463(.A(div_input_data_e[114]), .Y(exu_n16538));
AND2X1 exu_U464(.A(exu_n2819), .B(exu_n7900), .Y(exu_n27093));
AND2X1 exu_U465(.A(exu_n3138), .B(exu_n8218), .Y(exu_n28083));
INVX1 exu_U466(.A(div_input_data_e[113]), .Y(exu_n16537));
AND2X1 exu_U467(.A(exu_n2821), .B(exu_n7902), .Y(exu_n27099));
AND2X1 exu_U468(.A(exu_n3140), .B(exu_n8220), .Y(exu_n28089));
INVX1 exu_U469(.A(div_input_data_e[112]), .Y(exu_n16536));
AND2X1 exu_U470(.A(exu_n2825), .B(exu_n7906), .Y(exu_n27111));
AND2X1 exu_U471(.A(exu_n3142), .B(exu_n8222), .Y(exu_n28095));
INVX1 exu_U472(.A(div_input_data_e[111]), .Y(exu_n16535));
AND2X1 exu_U473(.A(exu_n2827), .B(exu_n7908), .Y(exu_n27117));
AND2X1 exu_U474(.A(exu_n3144), .B(exu_n8224), .Y(exu_n28101));
INVX1 exu_U475(.A(div_input_data_e[110]), .Y(exu_n16534));
AND2X1 exu_U476(.A(exu_n2829), .B(exu_n7910), .Y(exu_n27123));
AND2X1 exu_U477(.A(exu_n3146), .B(exu_n8226), .Y(exu_n28107));
INVX1 exu_U478(.A(div_input_data_e[109]), .Y(exu_n16533));
AND2X1 exu_U479(.A(exu_n2831), .B(exu_n7912), .Y(exu_n27129));
AND2X1 exu_U480(.A(exu_n3148), .B(exu_n8228), .Y(exu_n28113));
INVX1 exu_U481(.A(div_input_data_e[108]), .Y(exu_n16532));
AND2X1 exu_U482(.A(exu_n2833), .B(exu_n7914), .Y(exu_n27135));
AND2X1 exu_U483(.A(exu_n3150), .B(exu_n8230), .Y(exu_n28119));
INVX1 exu_U484(.A(div_input_data_e[107]), .Y(exu_n16531));
AND2X1 exu_U485(.A(exu_n2835), .B(exu_n7916), .Y(exu_n27141));
AND2X1 exu_U486(.A(exu_n3152), .B(exu_n8232), .Y(exu_n28125));
INVX1 exu_U487(.A(div_input_data_e[106]), .Y(exu_n16530));
AND2X1 exu_U488(.A(exu_n2837), .B(exu_n7918), .Y(exu_n27147));
AND2X1 exu_U489(.A(exu_n3154), .B(exu_n8234), .Y(exu_n28131));
INVX1 exu_U490(.A(div_input_data_e[105]), .Y(exu_n16529));
AND2X1 exu_U491(.A(exu_n2839), .B(exu_n7920), .Y(exu_n27153));
AND2X1 exu_U492(.A(exu_n3156), .B(exu_n8236), .Y(exu_n28137));
INVX1 exu_U493(.A(div_input_data_e[104]), .Y(exu_n16528));
AND2X1 exu_U494(.A(exu_n2841), .B(exu_n7922), .Y(exu_n27159));
AND2X1 exu_U495(.A(exu_n3158), .B(exu_n8238), .Y(exu_n28144));
INVX1 exu_U496(.A(div_input_data_e[103]), .Y(exu_n16527));
AND2X1 exu_U497(.A(exu_n2843), .B(exu_n7924), .Y(exu_n27165));
AND2X1 exu_U498(.A(exu_n3160), .B(exu_n8240), .Y(exu_n28150));
INVX1 exu_U499(.A(div_input_data_e[102]), .Y(exu_n16526));
AND2X1 exu_U500(.A(exu_n2847), .B(exu_n7928), .Y(exu_n27177));
AND2X1 exu_U501(.A(exu_n3162), .B(exu_n8242), .Y(exu_n28156));
INVX1 exu_U502(.A(div_input_data_e[101]), .Y(exu_n16525));
AND2X1 exu_U503(.A(exu_n2849), .B(exu_n7930), .Y(exu_n27183));
AND2X1 exu_U504(.A(exu_n3164), .B(exu_n8244), .Y(exu_n28162));
INVX1 exu_U505(.A(div_input_data_e[100]), .Y(exu_n16524));
AND2X1 exu_U506(.A(exu_n2851), .B(exu_n7932), .Y(exu_n27189));
AND2X1 exu_U507(.A(exu_n3166), .B(exu_n8246), .Y(exu_n28168));
INVX1 exu_U508(.A(div_input_data_e[99]), .Y(exu_n16523));
AND2X1 exu_U509(.A(exu_n2853), .B(exu_n7934), .Y(exu_n27195));
AND2X1 exu_U510(.A(exu_n3168), .B(exu_n8248), .Y(exu_n28174));
INVX1 exu_U511(.A(div_input_data_e[98]), .Y(exu_n16522));
AND2X1 exu_U512(.A(exu_n2855), .B(exu_n7936), .Y(exu_n27201));
AND2X1 exu_U513(.A(exu_n3170), .B(exu_n8250), .Y(exu_n28180));
INVX1 exu_U514(.A(div_input_data_e[97]), .Y(exu_n16521));
AND2X1 exu_U515(.A(exu_n2857), .B(exu_n7938), .Y(exu_n27207));
AND2X1 exu_U516(.A(exu_n3172), .B(exu_n8252), .Y(exu_n28186));
INVX1 exu_U517(.A(div_input_data_e[96]), .Y(exu_n16520));
AND2X1 exu_U518(.A(exu_n2859), .B(exu_n7940), .Y(exu_n27213));
AND2X1 exu_U519(.A(exu_n3174), .B(exu_n8254), .Y(exu_n28192));
AND2X1 exu_U520(.A(exu_n2861), .B(exu_n7942), .Y(exu_n27219));
AND2X1 exu_U521(.A(exu_n3176), .B(exu_n8256), .Y(exu_n28198));
AND2X1 exu_U522(.A(exu_n2863), .B(exu_n7944), .Y(exu_n27225));
AND2X1 exu_U523(.A(exu_n3178), .B(exu_n8258), .Y(exu_n28205));
AND2X1 exu_U524(.A(exu_n2865), .B(exu_n7946), .Y(exu_n27231));
AND2X1 exu_U525(.A(exu_n3180), .B(exu_n8260), .Y(exu_n28211));
AND2X1 exu_U526(.A(exu_n2869), .B(exu_n7950), .Y(exu_n27243));
AND2X1 exu_U527(.A(exu_n3182), .B(exu_n8262), .Y(exu_n28217));
AND2X1 exu_U528(.A(exu_n2871), .B(exu_n7952), .Y(exu_n27249));
AND2X1 exu_U529(.A(exu_n3184), .B(exu_n8264), .Y(exu_n28223));
AND2X1 exu_U530(.A(exu_n2873), .B(exu_n7954), .Y(exu_n27255));
AND2X1 exu_U531(.A(exu_n3186), .B(exu_n8266), .Y(exu_n28229));
AND2X1 exu_U532(.A(exu_n2875), .B(exu_n7956), .Y(exu_n27261));
AND2X1 exu_U533(.A(exu_n3188), .B(exu_n8268), .Y(exu_n28235));
AND2X1 exu_U534(.A(exu_n2877), .B(exu_n7958), .Y(exu_n27267));
AND2X1 exu_U535(.A(exu_n3190), .B(exu_n8270), .Y(exu_n28241));
AND2X1 exu_U536(.A(exu_n2879), .B(exu_n7960), .Y(exu_n27273));
AND2X1 exu_U537(.A(exu_n3192), .B(exu_n8272), .Y(exu_n28247));
AND2X1 exu_U538(.A(exu_n2881), .B(exu_n7962), .Y(exu_n27279));
AND2X1 exu_U539(.A(exu_n3194), .B(exu_n8274), .Y(exu_n28253));
AND2X1 exu_U540(.A(exu_n2883), .B(exu_n7964), .Y(exu_n27285));
AND2X1 exu_U541(.A(exu_n3196), .B(exu_n8276), .Y(exu_n28259));
AND2X1 exu_U542(.A(exu_n2885), .B(exu_n7966), .Y(exu_n27291));
AND2X1 exu_U543(.A(exu_n3198), .B(exu_n8278), .Y(exu_n28266));
AND2X1 exu_U544(.A(exu_n2887), .B(exu_n7968), .Y(exu_n27297));
AND2X1 exu_U545(.A(exu_n3200), .B(exu_n8280), .Y(exu_n28272));
AND2X1 exu_U546(.A(exu_n2891), .B(exu_n7972), .Y(exu_n27309));
AND2X1 exu_U547(.A(exu_n3202), .B(exu_n8282), .Y(exu_n28278));
AND2X1 exu_U548(.A(exu_n2893), .B(exu_n7974), .Y(exu_n27315));
AND2X1 exu_U549(.A(exu_n3204), .B(exu_n8284), .Y(exu_n28284));
AND2X1 exu_U550(.A(exu_n2895), .B(exu_n7976), .Y(exu_n27321));
AND2X1 exu_U551(.A(exu_n3206), .B(exu_n8286), .Y(exu_n28290));
AND2X1 exu_U552(.A(exu_n2897), .B(exu_n7978), .Y(exu_n27327));
AND2X1 exu_U553(.A(exu_n3208), .B(exu_n8288), .Y(exu_n28296));
AND2X1 exu_U554(.A(exu_n2899), .B(exu_n7980), .Y(exu_n27333));
AND2X1 exu_U555(.A(exu_n3210), .B(exu_n8290), .Y(exu_n28302));
AND2X1 exu_U556(.A(exu_n2901), .B(exu_n7982), .Y(exu_n27339));
AND2X1 exu_U557(.A(exu_n3212), .B(exu_n8292), .Y(exu_n28308));
AND2X1 exu_U558(.A(exu_n2907), .B(exu_n7988), .Y(exu_n27357));
AND2X1 exu_U559(.A(exu_n2903), .B(exu_n7984), .Y(exu_n27345));
AND2X1 exu_U560(.A(exu_n2905), .B(exu_n7986), .Y(exu_n27351));
AND2X1 exu_U561(.A(exu_n2909), .B(exu_n7990), .Y(exu_n27363));
AND2X1 exu_U562(.A(exu_n2792), .B(exu_n7878), .Y(exu_n27012));
AND2X1 exu_U563(.A(exu_n2794), .B(exu_n7880), .Y(exu_n27018));
AND2X1 exu_U564(.A(exu_n2796), .B(exu_n7882), .Y(exu_n27024));
AND2X1 exu_U565(.A(exu_n2798), .B(exu_n7884), .Y(exu_n27030));
AND2X1 exu_U566(.A(exu_n2804), .B(exu_n7888), .Y(exu_n27049));
AND2X1 exu_U567(.A(exu_n2823), .B(exu_n7904), .Y(exu_n27105));
AND2X1 exu_U568(.A(exu_n2889), .B(exu_n7970), .Y(exu_n27303));
AND2X1 exu_U569(.A(exu_n2845), .B(exu_n7926), .Y(exu_n27171));
INVX1 exu_U570(.A(div_input_data_e[64]), .Y(exu_n16514));
AND2X1 exu_U571(.A(exu_n2911), .B(exu_n7992), .Y(exu_n27369));
AND2X1 exu_U572(.A(exu_n2867), .B(exu_n7948), .Y(exu_n27237));
AND2X1 exu_U573(.A(alu_logic_rs1_data_bf1[0]), .B(ecl_enshift_e), .Y(shft_rshifterinput_b1[0]));
INVX1 exu_U574(.A(ecl_rd_e[0]), .Y(exu_n16563));
INVX1 exu_U575(.A(ecl_ifu_exu_rs2_d[1]), .Y(exu_n16568));
INVX1 exu_U576(.A(ecl_ld_rd_g[0]), .Y(exu_n16565));
INVX1 exu_U577(.A(ecl_ifu_exu_rs3_d[1]), .Y(exu_n16567));
OR2X1 exu_U578(.A(exu_n16563), .B(ecl_ifu_exu_rs3_d[0]), .Y(exu_n17445));
OR2X1 exu_U579(.A(exu_n16563), .B(ecl_ifu_exu_rs1_d[0]), .Y(exu_n16669));
OR2X1 exu_U580(.A(exu_n16565), .B(ecl_ifu_exu_rs1_d[0]), .Y(exu_n16641));
OR2X1 exu_U581(.A(div_adderin2[42]), .B(exu_n15886), .Y(div_spr_n53));
OR2X1 exu_U582(.A(div_adderin2[41]), .B(exu_n15887), .Y(div_spr_n55));
OR2X1 exu_U583(.A(div_adderin2[40]), .B(exu_n15888), .Y(div_spr_n57));
OR2X1 exu_U584(.A(div_adderin2[39]), .B(exu_n15890), .Y(div_spr_n59));
OR2X1 exu_U585(.A(div_adderin2[44]), .B(exu_n15884), .Y(div_spr_n49));
OR2X1 exu_U586(.A(div_adderin2[43]), .B(exu_n15885), .Y(div_spr_n51));
OR2X1 exu_U587(.A(div_adderin2[45]), .B(exu_n15883), .Y(div_spr_n47));
AND2X1 exu_U588(.A(exu_n3857), .B(exu_n8936), .Y(div_z_in[47]));
OR2X1 exu_U589(.A(div_adderin2[34]), .B(exu_n15895), .Y(div_spr_n71));
OR2X1 exu_U590(.A(div_adderin2[33]), .B(exu_n15896), .Y(div_spr_n73));
OR2X1 exu_U591(.A(div_adderin2[32]), .B(exu_n15858), .Y(div_spr_n75));
OR2X1 exu_U592(.A(div_adderin2[31]), .B(exu_n15897), .Y(div_spr_n77));
OR2X1 exu_U593(.A(div_adderin2[36]), .B(exu_n15893), .Y(div_spr_n67));
OR2X1 exu_U594(.A(div_adderin2[35]), .B(exu_n15894), .Y(div_spr_n69));
OR2X1 exu_U595(.A(div_adderin2[37]), .B(exu_n15892), .Y(div_spr_n65));
AND2X1 exu_U596(.A(exu_n3866), .B(exu_n8945), .Y(div_z_in[39]));
OR2X1 exu_U597(.A(div_adderin2[58]), .B(exu_n15869), .Y(div_spr_n19));
OR2X1 exu_U598(.A(div_adderin2[57]), .B(exu_n15870), .Y(div_spr_n21));
OR2X1 exu_U599(.A(div_adderin2[56]), .B(exu_n15871), .Y(div_spr_n23));
OR2X1 exu_U600(.A(div_adderin2[55]), .B(exu_n15872), .Y(div_spr_n25));
OR2X1 exu_U601(.A(div_adderin2[60]), .B(exu_n15866), .Y(div_spr_n13));
OR2X1 exu_U602(.A(div_adderin2[59]), .B(exu_n15868), .Y(div_spr_n15));
OR2X1 exu_U603(.A(div_adderin2[61]), .B(exu_n15865), .Y(div_spr_n11));
AND2X1 exu_U604(.A(exu_n3839), .B(exu_n8918), .Y(div_z_in[63]));
OR2X1 exu_U605(.A(div_adderin2[50]), .B(exu_n15877), .Y(div_spr_n35));
OR2X1 exu_U606(.A(div_adderin2[49]), .B(exu_n15879), .Y(div_spr_n37));
OR2X1 exu_U607(.A(div_adderin2[48]), .B(exu_n15880), .Y(div_spr_n41));
OR2X1 exu_U608(.A(div_adderin2[47]), .B(exu_n15881), .Y(div_spr_n43));
OR2X1 exu_U609(.A(div_adderin2[52]), .B(exu_n15875), .Y(div_spr_n31));
OR2X1 exu_U610(.A(div_adderin2[51]), .B(exu_n15876), .Y(div_spr_n33));
OR2X1 exu_U611(.A(div_adderin2[53]), .B(exu_n15874), .Y(div_spr_n29));
AND2X1 exu_U612(.A(exu_n3848), .B(exu_n8927), .Y(div_z_in[55]));
OR2X1 exu_U613(.A(div_adderin2[6]), .B(exu_n15863), .Y(div_spr_n5));
OR2X1 exu_U614(.A(div_adderin2[5]), .B(exu_n15867), .Y(div_spr_n7));
OR2X1 exu_U615(.A(div_adderin2[7]), .B(exu_n15862), .Y(div_spr_n3));
AND2X1 exu_U616(.A(exu_n3835), .B(exu_n8914), .Y(div_z_in[9]));
OR2X1 exu_U617(.A(div_adderin2[2]), .B(exu_n15899), .Y(div_spr_n61));
OR2X1 exu_U618(.A(div_adderin2[30]), .B(exu_n15898), .Y(div_spr_n79));
OR2X1 exu_U619(.A(div_adderin2[3]), .B(exu_n15889), .Y(div_spr_n39));
AND2X1 exu_U620(.A(exu_n3843), .B(exu_n8922), .Y(div_z_in[5]));
OR2X1 exu_U621(.A(div_adderin2[28]), .B(exu_n15901), .Y(div_spr_n85));
OR2X1 exu_U622(.A(div_adderin2[27]), .B(exu_n15902), .Y(div_spr_n87));
OR2X1 exu_U623(.A(div_adderin2[1]), .B(exu_n15910), .Y(div_spr_n83));
AND2X1 exu_U624(.A(exu_n3875), .B(exu_n8954), .Y(div_z_in[30]));
OR2X1 exu_U625(.A(div_adderin2[24]), .B(exu_n15905), .Y(div_spr_n93));
OR2X1 exu_U626(.A(div_adderin2[23]), .B(exu_n15906), .Y(div_spr_n95));
OR2X1 exu_U627(.A(div_adderin2[25]), .B(exu_n15904), .Y(div_spr_n91));
AND2X1 exu_U628(.A(exu_n3879), .B(exu_n8958), .Y(div_z_in[27]));
OR2X1 exu_U629(.A(div_adderin2[14]), .B(exu_n15916), .Y(div_spr_n115));
AND2X1 exu_U630(.A(exu_n3891), .B(exu_n8970), .Y(div_z_in[16]));
OR2X1 exu_U631(.A(div_adderin2[12]), .B(exu_n15918), .Y(div_spr_n119));
AND2X1 exu_U632(.A(exu_n3893), .B(exu_n8972), .Y(div_z_in[14]));
OR2X1 exu_U633(.A(div_adderin2[10]), .B(exu_n15920), .Y(div_spr_n123));
AND2X1 exu_U634(.A(exu_n3895), .B(exu_n8974), .Y(div_z_in[12]));
AND2X1 exu_U635(.A(exu_n3897), .B(exu_n8976), .Y(div_z_in[10]));
AND2X1 exu_U636(.A(exu_n3887), .B(exu_n8966), .Y(div_z_in[1]));
AND2X1 exu_U637(.A(exu_n3888), .B(exu_n8967), .Y(div_z_in[19]));
AND2X1 exu_U638(.A(exu_n3889), .B(exu_n8968), .Y(div_z_in[18]));
AND2X1 exu_U639(.A(exu_n3890), .B(exu_n8969), .Y(div_z_in[17]));
AND2X1 exu_U640(.A(exu_n3885), .B(exu_n8964), .Y(div_z_in[21]));
AND2X1 exu_U641(.A(exu_n3886), .B(exu_n8965), .Y(div_z_in[20]));
AND2X1 exu_U642(.A(exu_n3884), .B(exu_n8963), .Y(div_z_in[22]));
OR2X1 exu_U643(.A(alu_addsub_rs2_data[46]), .B(alu_logic_rs1_data_bf1[46]), .Y(exu_n31533));
OR2X1 exu_U644(.A(alu_addsub_rs2_data[62]), .B(alu_logic_rs1_data_bf1[62]), .Y(exu_n31497));
OR2X1 exu_U645(.A(alu_addsub_rs2_data[54]), .B(alu_logic_rs1_data_bf1[54]), .Y(exu_n31515));
OR2X1 exu_U646(.A(alu_addsub_rs2_data_22), .B(alu_logic_rs1_data_bf1[22]), .Y(exu_n31585));
OR2X1 exu_U647(.A(alu_addsub_rs2_data_8), .B(alu_logic_rs1_data_bf1[8]), .Y(exu_n31489));
OR2X1 exu_U648(.A(exu_n13183), .B(exu_n14488), .Y(shft_lshift4_b1[63]));
AND2X1 exu_U649(.A(exu_n3109), .B(exu_n8189), .Y(exu_n27992));
OR2X1 exu_U650(.A(exu_n13184), .B(exu_n14489), .Y(shft_lshift4_b1[62]));
AND2X1 exu_U651(.A(exu_n3111), .B(exu_n8191), .Y(exu_n27998));
OR2X1 exu_U652(.A(exu_n13047), .B(exu_n14330), .Y(shft_rshift4_b1[63]));
AND2X1 exu_U653(.A(exu_n2800), .B(exu_n7886), .Y(exu_n27035));
OR2X1 exu_U654(.A(exu_n13185), .B(exu_n14490), .Y(shft_lshift4_b1[61]));
AND2X1 exu_U655(.A(exu_n3113), .B(exu_n8193), .Y(exu_n28004));
OR2X1 exu_U656(.A(exu_n13046), .B(exu_n14331), .Y(shft_rshift4_b1[62]));
AND2X1 exu_U657(.A(exu_n2810), .B(exu_n7887), .Y(exu_n27037));
OR2X1 exu_U658(.A(exu_n13186), .B(exu_n14491), .Y(shft_lshift4_b1[60]));
AND2X1 exu_U659(.A(exu_n3115), .B(exu_n8195), .Y(exu_n28010));
OR2X1 exu_U660(.A(exu_n13047), .B(exu_n14332), .Y(shft_rshift4_b1[61]));
AND2X1 exu_U661(.A(exu_n2802), .B(exu_n7886), .Y(exu_n27041));
OR2X1 exu_U662(.A(exu_n13187), .B(exu_n14492), .Y(shft_lshift4_b1[59]));
AND2X1 exu_U663(.A(exu_n3118), .B(exu_n8198), .Y(exu_n28019));
OR2X1 exu_U664(.A(exu_n13048), .B(exu_n14333), .Y(shft_rshift4_b1[60]));
AND2X1 exu_U665(.A(exu_n2810), .B(exu_n7887), .Y(exu_n27043));
OR2X1 exu_U666(.A(exu_n13188), .B(exu_n14493), .Y(shft_lshift4_b1[58]));
AND2X1 exu_U667(.A(exu_n3120), .B(exu_n8200), .Y(exu_n28025));
OR2X1 exu_U668(.A(exu_n13050), .B(exu_n14335), .Y(shft_rshift4_b1[59]));
AND2X1 exu_U669(.A(exu_n2810), .B(exu_n7891), .Y(exu_n27054));
OR2X1 exu_U670(.A(exu_n13189), .B(exu_n14494), .Y(shft_lshift4_b1[57]));
AND2X1 exu_U671(.A(exu_n3122), .B(exu_n8202), .Y(exu_n28031));
OR2X1 exu_U672(.A(exu_n13051), .B(exu_n14336), .Y(shft_rshift4_b1[58]));
AND2X1 exu_U673(.A(exu_n2810), .B(exu_n7893), .Y(exu_n27059));
OR2X1 exu_U674(.A(exu_n13190), .B(exu_n14495), .Y(shft_lshift4_b1[56]));
AND2X1 exu_U675(.A(exu_n3124), .B(exu_n8204), .Y(exu_n28037));
OR2X1 exu_U676(.A(exu_n13047), .B(exu_n14337), .Y(shft_rshift4_b1[57]));
AND2X1 exu_U677(.A(exu_n2808), .B(exu_n7894), .Y(exu_n27064));
OR2X1 exu_U678(.A(exu_n13191), .B(exu_n14496), .Y(shft_lshift4_b1[55]));
AND2X1 exu_U679(.A(exu_n3126), .B(exu_n8206), .Y(exu_n28043));
OR2X1 exu_U680(.A(exu_n13052), .B(exu_n14338), .Y(shft_rshift4_b1[56]));
AND2X1 exu_U681(.A(exu_n2810), .B(exu_n7893), .Y(exu_n27067));
OR2X1 exu_U682(.A(exu_n13192), .B(exu_n14497), .Y(shft_lshift4_b1[54]));
AND2X1 exu_U683(.A(exu_n3128), .B(exu_n8208), .Y(exu_n28049));
OR2X1 exu_U684(.A(exu_n13053), .B(exu_n14339), .Y(shft_rshift4_b1[55]));
AND2X1 exu_U685(.A(exu_n2812), .B(exu_n7891), .Y(exu_n27072));
OR2X1 exu_U686(.A(exu_n13193), .B(exu_n14498), .Y(shft_lshift4_b1[53]));
AND2X1 exu_U687(.A(exu_n3130), .B(exu_n8210), .Y(exu_n28055));
OR2X1 exu_U688(.A(exu_n13054), .B(exu_n14340), .Y(shft_rshift4_b1[54]));
AND2X1 exu_U689(.A(exu_n2814), .B(exu_n7887), .Y(exu_n27077));
OR2X1 exu_U690(.A(exu_n13194), .B(exu_n14499), .Y(shft_lshift4_b1[52]));
AND2X1 exu_U691(.A(exu_n3132), .B(exu_n8212), .Y(exu_n28061));
OR2X1 exu_U692(.A(exu_n13055), .B(exu_n14341), .Y(shft_rshift4_b1[53]));
AND2X1 exu_U693(.A(exu_n2816), .B(exu_n7893), .Y(exu_n27082));
OR2X1 exu_U694(.A(exu_n13195), .B(exu_n14500), .Y(shft_lshift4_b1[51]));
AND2X1 exu_U695(.A(exu_n3134), .B(exu_n8214), .Y(exu_n28067));
OR2X1 exu_U696(.A(exu_n13056), .B(exu_n14342), .Y(shft_rshift4_b1[52]));
AND2X1 exu_U697(.A(exu_n2818), .B(exu_n7887), .Y(exu_n27087));
OR2X1 exu_U698(.A(exu_n13196), .B(exu_n14501), .Y(shft_lshift4_b1[50]));
AND2X1 exu_U699(.A(exu_n3136), .B(exu_n8216), .Y(exu_n28073));
OR2X1 exu_U700(.A(exu_n13057), .B(exu_n14343), .Y(shft_rshift4_b1[51]));
AND2X1 exu_U701(.A(exu_n2820), .B(exu_n7901), .Y(exu_n27092));
OR2X1 exu_U702(.A(exu_n13197), .B(exu_n14502), .Y(shft_lshift4_b1[49]));
AND2X1 exu_U703(.A(exu_n3139), .B(exu_n8219), .Y(exu_n28082));
OR2X1 exu_U704(.A(exu_n13058), .B(exu_n14344), .Y(shft_rshift4_b1[50]));
AND2X1 exu_U705(.A(exu_n2822), .B(exu_n7903), .Y(exu_n27098));
OR2X1 exu_U706(.A(exu_n13198), .B(exu_n14503), .Y(shft_lshift4_b1[48]));
AND2X1 exu_U707(.A(exu_n3141), .B(exu_n8221), .Y(exu_n28088));
OR2X1 exu_U708(.A(exu_n13060), .B(exu_n14346), .Y(shft_rshift4_b1[49]));
AND2X1 exu_U709(.A(exu_n2826), .B(exu_n7907), .Y(exu_n27110));
OR2X1 exu_U710(.A(exu_n13199), .B(exu_n14504), .Y(shft_lshift4_b1[47]));
AND2X1 exu_U711(.A(exu_n3143), .B(exu_n8223), .Y(exu_n28094));
OR2X1 exu_U712(.A(exu_n13061), .B(exu_n14347), .Y(shft_rshift4_b1[48]));
AND2X1 exu_U713(.A(exu_n2828), .B(exu_n7909), .Y(exu_n27116));
OR2X1 exu_U714(.A(exu_n13200), .B(exu_n14505), .Y(shft_lshift4_b1[46]));
AND2X1 exu_U715(.A(exu_n3145), .B(exu_n8225), .Y(exu_n28100));
OR2X1 exu_U716(.A(exu_n13062), .B(exu_n14348), .Y(shft_rshift4_b1[47]));
AND2X1 exu_U717(.A(exu_n2830), .B(exu_n7911), .Y(exu_n27122));
OR2X1 exu_U718(.A(exu_n13201), .B(exu_n14506), .Y(shft_lshift4_b1[45]));
AND2X1 exu_U719(.A(exu_n3147), .B(exu_n8227), .Y(exu_n28106));
OR2X1 exu_U720(.A(exu_n13063), .B(exu_n14349), .Y(shft_rshift4_b1[46]));
AND2X1 exu_U721(.A(exu_n2832), .B(exu_n7913), .Y(exu_n27128));
OR2X1 exu_U722(.A(exu_n13202), .B(exu_n14507), .Y(shft_lshift4_b1[44]));
AND2X1 exu_U723(.A(exu_n3149), .B(exu_n8229), .Y(exu_n28112));
OR2X1 exu_U724(.A(exu_n13064), .B(exu_n14350), .Y(shft_rshift4_b1[45]));
AND2X1 exu_U725(.A(exu_n2834), .B(exu_n7915), .Y(exu_n27134));
OR2X1 exu_U726(.A(exu_n13203), .B(exu_n14508), .Y(shft_lshift4_b1[43]));
AND2X1 exu_U727(.A(exu_n3151), .B(exu_n8231), .Y(exu_n28118));
OR2X1 exu_U728(.A(exu_n13065), .B(exu_n14351), .Y(shft_rshift4_b1[44]));
AND2X1 exu_U729(.A(exu_n2836), .B(exu_n7917), .Y(exu_n27140));
OR2X1 exu_U730(.A(exu_n13204), .B(exu_n14509), .Y(shft_lshift4_b1[42]));
AND2X1 exu_U731(.A(exu_n3153), .B(exu_n8233), .Y(exu_n28124));
OR2X1 exu_U732(.A(exu_n13066), .B(exu_n14352), .Y(shft_rshift4_b1[43]));
AND2X1 exu_U733(.A(exu_n2838), .B(exu_n7919), .Y(exu_n27146));
OR2X1 exu_U734(.A(exu_n13205), .B(exu_n14510), .Y(shft_lshift4_b1[41]));
AND2X1 exu_U735(.A(exu_n3155), .B(exu_n8235), .Y(exu_n28130));
OR2X1 exu_U736(.A(exu_n13067), .B(exu_n14353), .Y(shft_rshift4_b1[42]));
AND2X1 exu_U737(.A(exu_n2840), .B(exu_n7921), .Y(exu_n27152));
OR2X1 exu_U738(.A(exu_n13206), .B(exu_n14511), .Y(shft_lshift4_b1[40]));
AND2X1 exu_U739(.A(exu_n3157), .B(exu_n8237), .Y(exu_n28136));
OR2X1 exu_U740(.A(exu_n13068), .B(exu_n14354), .Y(shft_rshift4_b1[41]));
AND2X1 exu_U741(.A(exu_n2842), .B(exu_n7923), .Y(exu_n27158));
OR2X1 exu_U742(.A(exu_n13207), .B(exu_n14512), .Y(shft_lshift4_b1[39]));
AND2X1 exu_U743(.A(exu_n3159), .B(exu_n8239), .Y(exu_n28143));
OR2X1 exu_U744(.A(exu_n13069), .B(exu_n14355), .Y(shft_rshift4_b1[40]));
AND2X1 exu_U745(.A(exu_n2844), .B(exu_n7925), .Y(exu_n27164));
OR2X1 exu_U746(.A(exu_n13208), .B(exu_n14513), .Y(shft_lshift4_b1[38]));
AND2X1 exu_U747(.A(exu_n3161), .B(exu_n8241), .Y(exu_n28149));
OR2X1 exu_U748(.A(exu_n13071), .B(exu_n14357), .Y(shft_rshift4_b1[39]));
AND2X1 exu_U749(.A(exu_n2848), .B(exu_n7929), .Y(exu_n27176));
OR2X1 exu_U750(.A(exu_n13209), .B(exu_n14514), .Y(shft_lshift4_b1[37]));
AND2X1 exu_U751(.A(exu_n3163), .B(exu_n8243), .Y(exu_n28155));
OR2X1 exu_U752(.A(exu_n13072), .B(exu_n14358), .Y(shft_rshift4_b1[38]));
AND2X1 exu_U753(.A(exu_n2850), .B(exu_n7931), .Y(exu_n27182));
OR2X1 exu_U754(.A(exu_n13210), .B(exu_n14515), .Y(shft_lshift4_b1[36]));
AND2X1 exu_U755(.A(exu_n3165), .B(exu_n8245), .Y(exu_n28161));
OR2X1 exu_U756(.A(exu_n13073), .B(exu_n14359), .Y(shft_rshift4_b1[37]));
AND2X1 exu_U757(.A(exu_n2852), .B(exu_n7933), .Y(exu_n27188));
OR2X1 exu_U758(.A(exu_n13211), .B(exu_n14516), .Y(shft_lshift4_b1[35]));
AND2X1 exu_U759(.A(exu_n3167), .B(exu_n8247), .Y(exu_n28167));
OR2X1 exu_U760(.A(exu_n13074), .B(exu_n14360), .Y(shft_rshift4_b1[36]));
AND2X1 exu_U761(.A(exu_n2854), .B(exu_n7935), .Y(exu_n27194));
OR2X1 exu_U762(.A(exu_n13212), .B(exu_n14517), .Y(shft_lshift4_b1[34]));
AND2X1 exu_U763(.A(exu_n3169), .B(exu_n8249), .Y(exu_n28173));
OR2X1 exu_U764(.A(exu_n13075), .B(exu_n14361), .Y(shft_rshift4_b1[35]));
AND2X1 exu_U765(.A(exu_n2856), .B(exu_n7937), .Y(exu_n27200));
OR2X1 exu_U766(.A(exu_n13213), .B(exu_n14518), .Y(shft_lshift4_b1[33]));
AND2X1 exu_U767(.A(exu_n3171), .B(exu_n8251), .Y(exu_n28179));
OR2X1 exu_U768(.A(exu_n13076), .B(exu_n14362), .Y(shft_rshift4_b1[34]));
AND2X1 exu_U769(.A(exu_n2858), .B(exu_n7939), .Y(exu_n27206));
OR2X1 exu_U770(.A(exu_n13214), .B(exu_n14519), .Y(shft_lshift4_b1[32]));
AND2X1 exu_U771(.A(exu_n3173), .B(exu_n8253), .Y(exu_n28185));
OR2X1 exu_U772(.A(exu_n13077), .B(exu_n14363), .Y(shft_rshift4_b1[33]));
AND2X1 exu_U773(.A(exu_n2860), .B(exu_n7941), .Y(exu_n27212));
OR2X1 exu_U774(.A(exu_n13215), .B(exu_n14520), .Y(shft_lshift4_b1[31]));
AND2X1 exu_U775(.A(exu_n3175), .B(exu_n8255), .Y(exu_n28191));
OR2X1 exu_U776(.A(exu_n13078), .B(exu_n14364), .Y(shft_rshift4_b1[32]));
AND2X1 exu_U777(.A(exu_n2862), .B(exu_n7943), .Y(exu_n27218));
OR2X1 exu_U778(.A(exu_n13216), .B(exu_n14521), .Y(shft_lshift4_b1[30]));
AND2X1 exu_U779(.A(exu_n3177), .B(exu_n8257), .Y(exu_n28197));
OR2X1 exu_U780(.A(exu_n13079), .B(exu_n14365), .Y(shft_rshift4_b1[31]));
AND2X1 exu_U781(.A(exu_n2864), .B(exu_n7945), .Y(exu_n27224));
OR2X1 exu_U782(.A(exu_n13217), .B(exu_n14522), .Y(shft_lshift4_b1[29]));
AND2X1 exu_U783(.A(exu_n3179), .B(exu_n8259), .Y(exu_n28204));
OR2X1 exu_U784(.A(exu_n13080), .B(exu_n14366), .Y(shft_rshift4_b1[30]));
AND2X1 exu_U785(.A(exu_n2866), .B(exu_n7947), .Y(exu_n27230));
OR2X1 exu_U786(.A(exu_n13218), .B(exu_n14523), .Y(shft_lshift4_b1[28]));
AND2X1 exu_U787(.A(exu_n3181), .B(exu_n8261), .Y(exu_n28210));
OR2X1 exu_U788(.A(exu_n13082), .B(exu_n14368), .Y(shft_rshift4_b1[29]));
AND2X1 exu_U789(.A(exu_n2870), .B(exu_n7951), .Y(exu_n27242));
OR2X1 exu_U790(.A(exu_n13219), .B(exu_n14524), .Y(shft_lshift4_b1[27]));
AND2X1 exu_U791(.A(exu_n3183), .B(exu_n8263), .Y(exu_n28216));
OR2X1 exu_U792(.A(exu_n13083), .B(exu_n14369), .Y(shft_rshift4_b1[28]));
AND2X1 exu_U793(.A(exu_n2872), .B(exu_n7953), .Y(exu_n27248));
OR2X1 exu_U794(.A(exu_n13220), .B(exu_n14525), .Y(shft_lshift4_b1[26]));
AND2X1 exu_U795(.A(exu_n3185), .B(exu_n8265), .Y(exu_n28222));
OR2X1 exu_U796(.A(exu_n13084), .B(exu_n14370), .Y(shft_rshift4_b1[27]));
AND2X1 exu_U797(.A(exu_n2874), .B(exu_n7955), .Y(exu_n27254));
OR2X1 exu_U798(.A(exu_n13221), .B(exu_n14526), .Y(shft_lshift4_b1[25]));
AND2X1 exu_U799(.A(exu_n3187), .B(exu_n8267), .Y(exu_n28228));
OR2X1 exu_U800(.A(exu_n13085), .B(exu_n14371), .Y(shft_rshift4_b1[26]));
AND2X1 exu_U801(.A(exu_n2876), .B(exu_n7957), .Y(exu_n27260));
OR2X1 exu_U802(.A(exu_n13222), .B(exu_n14527), .Y(shft_lshift4_b1[24]));
AND2X1 exu_U803(.A(exu_n3189), .B(exu_n8269), .Y(exu_n28234));
OR2X1 exu_U804(.A(exu_n13086), .B(exu_n14372), .Y(shft_rshift4_b1[25]));
AND2X1 exu_U805(.A(exu_n2878), .B(exu_n7959), .Y(exu_n27266));
OR2X1 exu_U806(.A(exu_n13223), .B(exu_n14528), .Y(shft_lshift4_b1[23]));
AND2X1 exu_U807(.A(exu_n3191), .B(exu_n8271), .Y(exu_n28240));
OR2X1 exu_U808(.A(exu_n13087), .B(exu_n14373), .Y(shft_rshift4_b1[24]));
AND2X1 exu_U809(.A(exu_n2880), .B(exu_n7961), .Y(exu_n27272));
OR2X1 exu_U810(.A(exu_n13224), .B(exu_n14529), .Y(shft_lshift4_b1[22]));
AND2X1 exu_U811(.A(exu_n3193), .B(exu_n8273), .Y(exu_n28246));
OR2X1 exu_U812(.A(exu_n13088), .B(exu_n14374), .Y(shft_rshift4_b1[23]));
AND2X1 exu_U813(.A(exu_n2882), .B(exu_n7963), .Y(exu_n27278));
OR2X1 exu_U814(.A(exu_n13225), .B(exu_n14530), .Y(shft_lshift4_b1[21]));
AND2X1 exu_U815(.A(exu_n3195), .B(exu_n8275), .Y(exu_n28252));
OR2X1 exu_U816(.A(exu_n13089), .B(exu_n14375), .Y(shft_rshift4_b1[22]));
AND2X1 exu_U817(.A(exu_n2884), .B(exu_n7965), .Y(exu_n27284));
OR2X1 exu_U818(.A(exu_n13226), .B(exu_n14531), .Y(shft_lshift4_b1[20]));
AND2X1 exu_U819(.A(exu_n3197), .B(exu_n8277), .Y(exu_n28258));
OR2X1 exu_U820(.A(exu_n13090), .B(exu_n14376), .Y(shft_rshift4_b1[21]));
AND2X1 exu_U821(.A(exu_n2886), .B(exu_n7967), .Y(exu_n27290));
OR2X1 exu_U822(.A(exu_n13227), .B(exu_n14532), .Y(shft_lshift4_b1[19]));
AND2X1 exu_U823(.A(exu_n3199), .B(exu_n8279), .Y(exu_n28265));
OR2X1 exu_U824(.A(exu_n13091), .B(exu_n14377), .Y(shft_rshift4_b1[20]));
AND2X1 exu_U825(.A(exu_n2888), .B(exu_n7969), .Y(exu_n27296));
OR2X1 exu_U826(.A(exu_n13228), .B(exu_n14533), .Y(shft_lshift4_b1[18]));
AND2X1 exu_U827(.A(exu_n3201), .B(exu_n8281), .Y(exu_n28271));
OR2X1 exu_U828(.A(exu_n13093), .B(exu_n14379), .Y(shft_rshift4_b1[19]));
AND2X1 exu_U829(.A(exu_n2892), .B(exu_n7973), .Y(exu_n27308));
OR2X1 exu_U830(.A(exu_n13229), .B(exu_n14534), .Y(shft_lshift4_b1[17]));
AND2X1 exu_U831(.A(exu_n3203), .B(exu_n8283), .Y(exu_n28277));
OR2X1 exu_U832(.A(exu_n13094), .B(exu_n14380), .Y(shft_rshift4_b1[18]));
AND2X1 exu_U833(.A(exu_n2894), .B(exu_n7975), .Y(exu_n27314));
OR2X1 exu_U834(.A(exu_n13230), .B(exu_n14535), .Y(shft_lshift4_b1[16]));
AND2X1 exu_U835(.A(exu_n3205), .B(exu_n8285), .Y(exu_n28283));
OR2X1 exu_U836(.A(exu_n13095), .B(exu_n14381), .Y(shft_rshift4_b1[17]));
AND2X1 exu_U837(.A(exu_n2896), .B(exu_n7977), .Y(exu_n27320));
OR2X1 exu_U838(.A(exu_n13231), .B(exu_n14536), .Y(shft_lshift4_b1[15]));
AND2X1 exu_U839(.A(exu_n3207), .B(exu_n8287), .Y(exu_n28289));
OR2X1 exu_U840(.A(exu_n13096), .B(exu_n14382), .Y(shft_rshift4_b1[16]));
AND2X1 exu_U841(.A(exu_n2898), .B(exu_n7979), .Y(exu_n27326));
OR2X1 exu_U842(.A(exu_n13232), .B(exu_n14537), .Y(shft_lshift4_b1[14]));
AND2X1 exu_U843(.A(exu_n3209), .B(exu_n8289), .Y(exu_n28295));
OR2X1 exu_U844(.A(exu_n13097), .B(exu_n14383), .Y(shft_rshift4_b1[15]));
AND2X1 exu_U845(.A(exu_n2900), .B(exu_n7981), .Y(exu_n27332));
OR2X1 exu_U846(.A(exu_n13233), .B(exu_n14538), .Y(shft_lshift4_b1[13]));
AND2X1 exu_U847(.A(exu_n3211), .B(exu_n8291), .Y(exu_n28301));
OR2X1 exu_U848(.A(exu_n13098), .B(exu_n14384), .Y(shft_rshift4_b1[14]));
AND2X1 exu_U849(.A(exu_n2902), .B(exu_n7983), .Y(exu_n27338));
OR2X1 exu_U850(.A(exu_n13234), .B(exu_n14539), .Y(shft_lshift4_b1[12]));
AND2X1 exu_U851(.A(exu_n3213), .B(exu_n8293), .Y(exu_n28307));
OR2X1 exu_U852(.A(exu_n13101), .B(exu_n14387), .Y(shft_rshift4_b1[11]));
AND2X1 exu_U853(.A(exu_n2908), .B(exu_n7989), .Y(exu_n27356));
OR2X1 exu_U854(.A(exu_n13099), .B(exu_n14385), .Y(shft_rshift4_b1[13]));
AND2X1 exu_U855(.A(exu_n2904), .B(exu_n7985), .Y(exu_n27344));
OR2X1 exu_U856(.A(exu_n28316), .B(exu_n14540), .Y(shft_lshift4_b1[11]));
AND2X1 exu_U857(.A(exu_n3214), .B(exu_n8294), .Y(exu_n28313));
OR2X1 exu_U858(.A(exu_n27981), .B(exu_n14486), .Y(shft_lshift4_b1[9]));
AND2X1 exu_U859(.A(exu_n3104), .B(exu_n8184), .Y(exu_n27978));
OR2X1 exu_U860(.A(exu_n13100), .B(exu_n14386), .Y(shft_rshift4_b1[12]));
AND2X1 exu_U861(.A(exu_n2906), .B(exu_n7987), .Y(exu_n27350));
OR2X1 exu_U862(.A(exu_n28320), .B(exu_n14541), .Y(shft_lshift4_b1[10]));
AND2X1 exu_U863(.A(exu_n3215), .B(exu_n8295), .Y(exu_n28317));
OR2X1 exu_U864(.A(exu_n13102), .B(exu_n14388), .Y(shft_rshift4_b1[10]));
AND2X1 exu_U865(.A(exu_n2910), .B(exu_n7991), .Y(exu_n27362));
OR2X1 exu_U866(.A(exu_n27985), .B(exu_n14487), .Y(shft_lshift4_b1[8]));
AND2X1 exu_U867(.A(exu_n3105), .B(exu_n8185), .Y(exu_n27982));
OR2X1 exu_U868(.A(exu_n13042), .B(exu_n14326), .Y(shft_rshift4_b1[9]));
AND2X1 exu_U869(.A(exu_n2793), .B(exu_n7879), .Y(exu_n27011));
AND2X1 exu_U870(.A(exu_n3106), .B(exu_n8186), .Y(exu_n27986));
OR2X1 exu_U871(.A(exu_n13043), .B(exu_n14327), .Y(shft_rshift4_b1[8]));
AND2X1 exu_U872(.A(exu_n2795), .B(exu_n7881), .Y(exu_n27017));
AND2X1 exu_U873(.A(exu_n3107), .B(exu_n8187), .Y(exu_n27989));
OR2X1 exu_U874(.A(exu_n13044), .B(exu_n14328), .Y(shft_rshift4_b1[7]));
AND2X1 exu_U875(.A(exu_n2797), .B(exu_n7883), .Y(exu_n27023));
AND2X1 exu_U876(.A(exu_n3116), .B(exu_n8196), .Y(exu_n28016));
OR2X1 exu_U877(.A(exu_n13045), .B(exu_n14329), .Y(shft_rshift4_b1[6]));
AND2X1 exu_U878(.A(exu_n2799), .B(exu_n7885), .Y(exu_n27029));
AND2X1 exu_U879(.A(exu_n3137), .B(exu_n8217), .Y(exu_n28079));
OR2X1 exu_U880(.A(exu_n13049), .B(exu_n14334), .Y(shft_rshift4_b1[5]));
AND2X1 exu_U881(.A(exu_n2805), .B(exu_n7889), .Y(exu_n27048));
OR2X1 exu_U882(.A(exu_n13059), .B(exu_n14345), .Y(shft_rshift4_b1[4]));
AND2X1 exu_U883(.A(exu_n2824), .B(exu_n7905), .Y(exu_n27104));
INVX1 exu_U884(.A(div_input_data_e[65]), .Y(exu_n16516));
OR2X1 exu_U885(.A(exu_n13092), .B(exu_n14378), .Y(shft_rshift4_b1[1]));
AND2X1 exu_U886(.A(exu_n2890), .B(exu_n7971), .Y(exu_n27302));
OR2X1 exu_U887(.A(exu_n13070), .B(exu_n14356), .Y(shft_rshift4_b1[3]));
AND2X1 exu_U888(.A(exu_n2846), .B(exu_n7927), .Y(exu_n27170));
OR2X1 exu_U889(.A(exu_n13103), .B(exu_n14389), .Y(shft_rshift4_b1[0]));
AND2X1 exu_U890(.A(exu_n2912), .B(exu_n7993), .Y(exu_n27368));
OR2X1 exu_U891(.A(exu_n13081), .B(exu_n14367), .Y(shft_rshift4_b1[2]));
AND2X1 exu_U892(.A(exu_n2868), .B(exu_n7949), .Y(exu_n27236));
AND2X1 exu_U893(.A(ecc_syn_mux_n1), .B(exu_n9360), .Y(ecc_err_m[6]));
AND2X1 exu_U894(.A(exu_n4580), .B(exu_n9361), .Y(ecc_syn_mux_n1));
AND2X1 exu_U895(.A(exu_n4581), .B(exu_n9363), .Y(ecc_syn_mux_n5));
AND2X1 exu_U896(.A(exu_n12), .B(exu_n4982), .Y(exu_n16664));
OR2X1 exu_U897(.A(exu_n16565), .B(ecl_ifu_exu_rs2_d[0]), .Y(exu_n16697));
AND2X1 exu_U898(.A(exu_n16), .B(exu_n4984), .Y(exu_n16692));
OR2X1 exu_U899(.A(exu_n16563), .B(ecl_ifu_exu_rs2_d[0]), .Y(exu_n16725));
INVX1 exu_U900(.A(ecl_rd_e[1]), .Y(exu_n16564));
AND2X1 exu_U901(.A(exu_n18), .B(exu_n4987), .Y(exu_n16720));
OR2X1 exu_U902(.A(exu_n16565), .B(ecl_ifu_exu_rs3_d[0]), .Y(exu_n17417));
INVX1 exu_U903(.A(ecl_ld_rd_g[1]), .Y(exu_n16566));
AND2X1 exu_U904(.A(exu_n10), .B(exu_n4979), .Y(exu_n16636));
AND2X1 exu_U905(.A(exu_n2913), .B(exu_n7994), .Y(exu_n27375));
AND2X1 exu_U906(.A(exu_n2914), .B(exu_n7995), .Y(exu_n27374));
AND2X1 exu_U907(.A(exu_n3217), .B(exu_n8297), .Y(exu_n28322));
AND2X1 exu_U908(.A(exu_n3216), .B(exu_n8296), .Y(exu_n28323));
AND2X1 exu_U909(.A(exu_n17375), .B(ecl_wb_byplog_rd_g2[0]), .Y(exu_n17377));
AND2X1 exu_U910(.A(exu_n17389), .B(ecl_rd_m[0]), .Y(exu_n17391));
INVX1 exu_U911(.A(tlu_exu_pic_onebelow_m), .Y(exu_n16318));
AND2X1 exu_U912(.A(exu_n154), .B(exu_n5121), .Y(exu_n17440));
AND2X1 exu_U913(.A(exu_n152), .B(exu_n5118), .Y(exu_n17412));
AND2X1 exu_U914(.A(exu_n3861), .B(exu_n8940), .Y(div_z_in[43]));
AND2X1 exu_U915(.A(exu_n3862), .B(exu_n8941), .Y(div_z_in[42]));
AND2X1 exu_U916(.A(exu_n3863), .B(exu_n8942), .Y(div_z_in[41]));
AND2X1 exu_U917(.A(exu_n3864), .B(exu_n8943), .Y(div_z_in[40]));
AND2X1 exu_U918(.A(exu_n3859), .B(exu_n8938), .Y(div_z_in[45]));
AND2X1 exu_U919(.A(exu_n3860), .B(exu_n8939), .Y(div_z_in[44]));
AND2X1 exu_U920(.A(exu_n3858), .B(exu_n8937), .Y(div_z_in[46]));
AND2X1 exu_U921(.A(exu_n3870), .B(exu_n8949), .Y(div_z_in[35]));
AND2X1 exu_U922(.A(exu_n3871), .B(exu_n8950), .Y(div_z_in[34]));
AND2X1 exu_U923(.A(exu_n3872), .B(exu_n8951), .Y(div_z_in[33]));
AND2X1 exu_U924(.A(exu_n3873), .B(exu_n8952), .Y(div_z_in[32]));
AND2X1 exu_U925(.A(exu_n3868), .B(exu_n8947), .Y(div_z_in[37]));
AND2X1 exu_U926(.A(exu_n3869), .B(exu_n8948), .Y(div_z_in[36]));
AND2X1 exu_U927(.A(exu_n3867), .B(exu_n8946), .Y(div_z_in[38]));
AND2X1 exu_U928(.A(exu_n3844), .B(exu_n8923), .Y(div_z_in[59]));
AND2X1 exu_U929(.A(exu_n3845), .B(exu_n8924), .Y(div_z_in[58]));
AND2X1 exu_U930(.A(exu_n3846), .B(exu_n8925), .Y(div_z_in[57]));
AND2X1 exu_U931(.A(exu_n3847), .B(exu_n8926), .Y(div_z_in[56]));
AND2X1 exu_U932(.A(exu_n3841), .B(exu_n8920), .Y(div_z_in[61]));
AND2X1 exu_U933(.A(exu_n3842), .B(exu_n8921), .Y(div_z_in[60]));
AND2X1 exu_U934(.A(exu_n3840), .B(exu_n8919), .Y(div_z_in[62]));
AND2X1 exu_U935(.A(exu_n3852), .B(exu_n8931), .Y(div_z_in[51]));
AND2X1 exu_U936(.A(exu_n3853), .B(exu_n8932), .Y(div_z_in[50]));
AND2X1 exu_U937(.A(exu_n3855), .B(exu_n8934), .Y(div_z_in[49]));
AND2X1 exu_U938(.A(exu_n3856), .B(exu_n8935), .Y(div_z_in[48]));
AND2X1 exu_U939(.A(exu_n3850), .B(exu_n8929), .Y(div_z_in[53]));
AND2X1 exu_U940(.A(exu_n3851), .B(exu_n8930), .Y(div_z_in[52]));
AND2X1 exu_U941(.A(exu_n3849), .B(exu_n8928), .Y(div_z_in[54]));
AND2X1 exu_U942(.A(exu_n3837), .B(exu_n8916), .Y(div_z_in[7]));
AND2X1 exu_U943(.A(exu_n3838), .B(exu_n8917), .Y(div_z_in[6]));
AND2X1 exu_U944(.A(exu_n3836), .B(exu_n8915), .Y(div_z_in[8]));
AND2X1 exu_U945(.A(exu_n3865), .B(exu_n8944), .Y(div_z_in[3]));
AND2X1 exu_U946(.A(exu_n3874), .B(exu_n8953), .Y(div_z_in[31]));
AND2X1 exu_U947(.A(exu_n3854), .B(exu_n8933), .Y(div_z_in[4]));
AND2X1 exu_U948(.A(exu_n3877), .B(exu_n8956), .Y(div_z_in[29]));
AND2X1 exu_U949(.A(exu_n3878), .B(exu_n8957), .Y(div_z_in[28]));
AND2X1 exu_U950(.A(exu_n3876), .B(exu_n8955), .Y(div_z_in[2]));
AND2X1 exu_U951(.A(exu_n3881), .B(exu_n8960), .Y(div_z_in[25]));
AND2X1 exu_U952(.A(exu_n3882), .B(exu_n8961), .Y(div_z_in[24]));
AND2X1 exu_U953(.A(exu_n3880), .B(exu_n8959), .Y(div_z_in[26]));
AND2X1 exu_U954(.A(exu_n3892), .B(exu_n8971), .Y(div_z_in[15]));
AND2X1 exu_U955(.A(exu_n3894), .B(exu_n8973), .Y(div_z_in[13]));
AND2X1 exu_U956(.A(exu_n3896), .B(exu_n8975), .Y(div_z_in[11]));
AND2X1 exu_U957(.A(exu_n3898), .B(exu_n8977), .Y(div_z_in[0]));
AND2X1 exu_U958(.A(exu_n4908), .B(exu_n9622), .Y(div_n41));
INVX1 exu_U959(.A(div_input_data_e[127]), .Y(exu_n16551));
OR2X1 exu_U960(.A(alu_addsub_rs2_data[38]), .B(alu_logic_rs1_data_bf1[38]), .Y(exu_n31551));
OR2X1 exu_U961(.A(alu_addsub_rs2_data[36]), .B(alu_logic_rs1_data_bf1[36]), .Y(exu_n31555));
OR2X1 exu_U962(.A(alu_addsub_rs2_data[34]), .B(alu_logic_rs1_data_bf1[34]), .Y(exu_n31559));
OR2X1 exu_U963(.A(alu_addsub_rs2_data[32]), .B(alu_logic_rs1_data_bf1[32]), .Y(exu_n31563));
OR2X1 exu_U964(.A(alu_addsub_rs2_data[42]), .B(alu_logic_rs1_data_bf1[42]), .Y(exu_n31541));
OR2X1 exu_U965(.A(alu_addsub_rs2_data[41]), .B(alu_logic_rs1_data_bf1[41]), .Y(exu_n31543));
OR2X1 exu_U966(.A(alu_addsub_rs2_data[40]), .B(alu_logic_rs1_data_bf1[40]), .Y(exu_n31545));
OR2X1 exu_U967(.A(alu_addsub_rs2_data[39]), .B(alu_logic_rs1_data_bf1[39]), .Y(exu_n31547));
OR2X1 exu_U968(.A(alu_addsub_rs2_data[44]), .B(alu_logic_rs1_data_bf1[44]), .Y(exu_n31537));
OR2X1 exu_U969(.A(alu_addsub_rs2_data[43]), .B(alu_logic_rs1_data_bf1[43]), .Y(exu_n31539));
OR2X1 exu_U970(.A(alu_addsub_rs2_data[45]), .B(alu_logic_rs1_data_bf1[45]), .Y(exu_n31535));
AND2X1 exu_U971(.A(exu_n3665), .B(exu_n8682), .Y(alu_zcomp_in[47]));
OR2X1 exu_U972(.A(alu_addsub_rs2_data[58]), .B(alu_logic_rs1_data_bf1[58]), .Y(exu_n31507));
OR2X1 exu_U973(.A(alu_addsub_rs2_data[57]), .B(alu_logic_rs1_data_bf1[57]), .Y(exu_n31509));
OR2X1 exu_U974(.A(alu_addsub_rs2_data[56]), .B(alu_logic_rs1_data_bf1[56]), .Y(exu_n31511));
OR2X1 exu_U975(.A(alu_addsub_rs2_data[55]), .B(alu_logic_rs1_data_bf1[55]), .Y(exu_n31513));
OR2X1 exu_U976(.A(alu_addsub_rs2_data[60]), .B(alu_logic_rs1_data_bf1[60]), .Y(exu_n31501));
OR2X1 exu_U977(.A(alu_addsub_rs2_data[59]), .B(alu_logic_rs1_data_bf1[59]), .Y(exu_n31503));
OR2X1 exu_U978(.A(alu_addsub_rs2_data[61]), .B(alu_logic_rs1_data_bf1[61]), .Y(exu_n31499));
AND2X1 exu_U979(.A(exu_n3647), .B(exu_n8664), .Y(alu_zcomp_in[63]));
OR2X1 exu_U980(.A(alu_addsub_rs2_data[50]), .B(alu_logic_rs1_data_bf1[50]), .Y(exu_n31523));
OR2X1 exu_U981(.A(alu_addsub_rs2_data[49]), .B(alu_logic_rs1_data_bf1[49]), .Y(exu_n31525));
OR2X1 exu_U982(.A(alu_addsub_rs2_data[48]), .B(alu_logic_rs1_data_bf1[48]), .Y(exu_n31529));
OR2X1 exu_U983(.A(alu_addsub_rs2_data[47]), .B(alu_logic_rs1_data_bf1[47]), .Y(exu_n31531));
OR2X1 exu_U984(.A(alu_addsub_rs2_data[52]), .B(alu_logic_rs1_data_bf1[52]), .Y(exu_n31519));
OR2X1 exu_U985(.A(alu_addsub_rs2_data[51]), .B(alu_logic_rs1_data_bf1[51]), .Y(exu_n31521));
OR2X1 exu_U986(.A(alu_addsub_rs2_data[53]), .B(alu_logic_rs1_data_bf1[53]), .Y(exu_n31517));
AND2X1 exu_U987(.A(exu_n3656), .B(exu_n8673), .Y(alu_zcomp_in[55]));
INVX1 exu_U988(.A(ecl_ifu_exu_aluop_e[2]), .Y(exu_n16402));
INVX1 exu_U989(.A(ecl_ifu_exu_aluop_e[1]), .Y(exu_n16401));
OR2X1 exu_U990(.A(alu_addsub_rs2_data_15), .B(alu_logic_rs1_data_bf1[15]), .Y(exu_n31601));
OR2X1 exu_U991(.A(alu_addsub_rs2_data_13), .B(alu_logic_rs1_data_bf1[13]), .Y(exu_n31605));
OR2X1 exu_U992(.A(alu_addsub_rs2_data_11), .B(alu_logic_rs1_data_bf1[11]), .Y(exu_n31609));
OR2X1 exu_U993(.A(alu_addsub_rs2_data_9), .B(alu_logic_rs1_data_bf1[9]), .Y(exu_n31613));
OR2X1 exu_U994(.A(alu_addsub_rs2_data_0), .B(alu_logic_rs1_data_bf1[0]), .Y(exu_n31593));
OR2X1 exu_U995(.A(alu_addsub_rs2_data_18), .B(alu_logic_rs1_data_bf1[18]), .Y(exu_n31595));
OR2X1 exu_U996(.A(alu_addsub_rs2_data_17), .B(alu_logic_rs1_data_bf1[17]), .Y(exu_n31597));
OR2X1 exu_U997(.A(alu_addsub_rs2_data_16), .B(alu_logic_rs1_data_bf1[16]), .Y(exu_n31599));
OR2X1 exu_U998(.A(alu_addsub_rs2_data_20), .B(alu_logic_rs1_data_bf1[20]), .Y(exu_n31589));
OR2X1 exu_U999(.A(alu_addsub_rs2_data_19), .B(alu_logic_rs1_data_bf1[19]), .Y(exu_n31591));
OR2X1 exu_U1000(.A(alu_addsub_rs2_data_21), .B(alu_logic_rs1_data_bf1[21]), .Y(exu_n31587));
AND2X1 exu_U1001(.A(exu_n3691), .B(exu_n8708), .Y(alu_zcomp_in[23]));
OR2X1 exu_U1002(.A(alu_addsub_rs2_data_29), .B(alu_logic_rs1_data_bf1[29]), .Y(exu_n31569));
OR2X1 exu_U1003(.A(alu_addsub_rs2_data_28), .B(alu_logic_rs1_data_bf1[28]), .Y(exu_n31573));
OR2X1 exu_U1004(.A(alu_addsub_rs2_data_26), .B(alu_logic_rs1_data_bf1[26]), .Y(exu_n31577));
OR2X1 exu_U1005(.A(alu_addsub_rs2_data_24), .B(alu_logic_rs1_data_bf1[24]), .Y(exu_n31581));
OR2X1 exu_U1006(.A(alu_addsub_rs2_data_4), .B(alu_logic_rs1_data_bf1[4]), .Y(exu_n31505));
OR2X1 exu_U1007(.A(alu_addsub_rs2_data_3), .B(alu_logic_rs1_data_bf1[3]), .Y(exu_n31527));
OR2X1 exu_U1008(.A(alu_addsub_rs2_data_2), .B(alu_logic_rs1_data_bf1[2]), .Y(exu_n31549));
OR2X1 exu_U1009(.A(alu_addsub_rs2_data_30), .B(alu_logic_rs1_data_bf1[30]), .Y(exu_n31567));
OR2X1 exu_U1010(.A(alu_addsub_rs2_data_6), .B(alu_logic_rs1_data_bf1[6]), .Y(exu_n31493));
OR2X1 exu_U1011(.A(alu_addsub_rs2_data_5), .B(alu_logic_rs1_data_bf1[5]), .Y(exu_n31495));
OR2X1 exu_U1012(.A(alu_addsub_rs2_data_7), .B(alu_logic_rs1_data_bf1[7]), .Y(exu_n31491));
AND2X1 exu_U1013(.A(exu_n3643), .B(exu_n8660), .Y(alu_zcomp_in[9]));
AND2X1 exu_U1014(.A(exu_n3224), .B(exu_n8304), .Y(exu_n28347));
AND2X1 exu_U1015(.A(exu_n3225), .B(exu_n8305), .Y(exu_n28346));
OR2X1 exu_U1016(.A(exu_n15680), .B(alu_logic_rs1_data_bf1[61]), .Y(exu_n17348));
AND2X1 exu_U1017(.A(exu_n2923), .B(exu_n8004), .Y(exu_n27398));
AND2X1 exu_U1018(.A(exu_n3226), .B(exu_n8306), .Y(exu_n28353));
AND2X1 exu_U1019(.A(exu_n3227), .B(exu_n8307), .Y(exu_n28352));
AND2X1 exu_U1020(.A(alu_logic_rs1_data_bf1[62]), .B(alu_logic_n102), .Y(alu_logic_result_and[62]));
OR2X1 exu_U1021(.A(alu_logic_n102), .B(alu_logic_rs1_data_bf1[62]), .Y(alu_logic_result_or[62]));
AND2X1 exu_U1022(.A(exu_n3412), .B(exu_n8493), .Y(exu_n28948));
OR2X1 exu_U1023(.A(exu_n15679), .B(alu_logic_rs1_data_bf1[60]), .Y(exu_n17341));
AND2X1 exu_U1024(.A(exu_n2924), .B(exu_n8005), .Y(exu_n27408));
AND2X1 exu_U1025(.A(exu_n2925), .B(exu_n8004), .Y(exu_n27407));
AND2X1 exu_U1026(.A(exu_n3228), .B(exu_n8308), .Y(exu_n28359));
AND2X1 exu_U1027(.A(exu_n3229), .B(exu_n8309), .Y(exu_n28358));
AND2X1 exu_U1028(.A(alu_logic_rs1_data_bf1[61]), .B(alu_logic_n103), .Y(alu_logic_result_and[61]));
OR2X1 exu_U1029(.A(alu_logic_n103), .B(alu_logic_rs1_data_bf1[61]), .Y(alu_logic_result_or[61]));
AND2X1 exu_U1030(.A(exu_n3414), .B(exu_n8495), .Y(exu_n28954));
OR2X1 exu_U1031(.A(exu_n15678), .B(alu_logic_rs1_data_bf1[59]), .Y(exu_n17336));
AND2X1 exu_U1032(.A(exu_n2926), .B(exu_n8006), .Y(exu_n27413));
AND2X1 exu_U1033(.A(exu_n2927), .B(exu_n8007), .Y(exu_n27412));
AND2X1 exu_U1034(.A(exu_n3230), .B(exu_n8310), .Y(exu_n28365));
AND2X1 exu_U1035(.A(exu_n3231), .B(exu_n8311), .Y(exu_n28364));
AND2X1 exu_U1036(.A(alu_logic_rs1_data_bf1[60]), .B(alu_logic_n104), .Y(alu_logic_result_and[60]));
OR2X1 exu_U1037(.A(alu_logic_n104), .B(alu_logic_rs1_data_bf1[60]), .Y(alu_logic_result_or[60]));
AND2X1 exu_U1038(.A(exu_n3416), .B(exu_n8497), .Y(exu_n28960));
OR2X1 exu_U1039(.A(exu_n15677), .B(alu_logic_rs1_data_bf1[58]), .Y(exu_n17331));
AND2X1 exu_U1040(.A(exu_n2930), .B(exu_n8010), .Y(exu_n27425));
AND2X1 exu_U1041(.A(exu_n2931), .B(exu_n8011), .Y(exu_n27424));
AND2X1 exu_U1042(.A(exu_n3234), .B(exu_n8314), .Y(exu_n28377));
AND2X1 exu_U1043(.A(exu_n3235), .B(exu_n8315), .Y(exu_n28376));
AND2X1 exu_U1044(.A(alu_logic_rs1_data_bf1[59]), .B(alu_logic_n106), .Y(alu_logic_result_and[59]));
OR2X1 exu_U1045(.A(alu_logic_n106), .B(alu_logic_rs1_data_bf1[59]), .Y(alu_logic_result_or[59]));
AND2X1 exu_U1046(.A(exu_n3420), .B(exu_n8501), .Y(exu_n28972));
OR2X1 exu_U1047(.A(exu_n15676), .B(alu_logic_rs1_data_bf1[57]), .Y(exu_n17326));
AND2X1 exu_U1048(.A(exu_n2932), .B(exu_n8012), .Y(exu_n27431));
AND2X1 exu_U1049(.A(exu_n2933), .B(exu_n8013), .Y(exu_n27430));
AND2X1 exu_U1050(.A(exu_n3236), .B(exu_n8316), .Y(exu_n28383));
AND2X1 exu_U1051(.A(exu_n3237), .B(exu_n8317), .Y(exu_n28382));
AND2X1 exu_U1052(.A(alu_logic_rs1_data_bf1[58]), .B(alu_logic_n107), .Y(alu_logic_result_and[58]));
OR2X1 exu_U1053(.A(alu_logic_n107), .B(alu_logic_rs1_data_bf1[58]), .Y(alu_logic_result_or[58]));
AND2X1 exu_U1054(.A(exu_n3422), .B(exu_n8503), .Y(exu_n28978));
OR2X1 exu_U1055(.A(exu_n15675), .B(alu_logic_rs1_data_bf1[56]), .Y(exu_n17321));
AND2X1 exu_U1056(.A(exu_n2934), .B(exu_n8014), .Y(exu_n27437));
AND2X1 exu_U1057(.A(exu_n2935), .B(exu_n8015), .Y(exu_n27436));
AND2X1 exu_U1058(.A(exu_n3238), .B(exu_n8318), .Y(exu_n28389));
AND2X1 exu_U1059(.A(exu_n3239), .B(exu_n8319), .Y(exu_n28388));
AND2X1 exu_U1060(.A(alu_logic_rs1_data_bf1[57]), .B(alu_logic_n108), .Y(alu_logic_result_and[57]));
OR2X1 exu_U1061(.A(alu_logic_n108), .B(alu_logic_rs1_data_bf1[57]), .Y(alu_logic_result_or[57]));
AND2X1 exu_U1062(.A(exu_n3424), .B(exu_n8505), .Y(exu_n28984));
OR2X1 exu_U1063(.A(exu_n15674), .B(alu_logic_rs1_data_bf1[55]), .Y(exu_n17316));
AND2X1 exu_U1064(.A(exu_n2936), .B(exu_n8016), .Y(exu_n27443));
AND2X1 exu_U1065(.A(exu_n2937), .B(exu_n8017), .Y(exu_n27442));
AND2X1 exu_U1066(.A(exu_n3240), .B(exu_n8320), .Y(exu_n28395));
AND2X1 exu_U1067(.A(exu_n3241), .B(exu_n8321), .Y(exu_n28394));
AND2X1 exu_U1068(.A(alu_logic_rs1_data_bf1[56]), .B(alu_logic_n109), .Y(alu_logic_result_and[56]));
OR2X1 exu_U1069(.A(alu_logic_n109), .B(alu_logic_rs1_data_bf1[56]), .Y(alu_logic_result_or[56]));
AND2X1 exu_U1070(.A(exu_n3426), .B(exu_n8507), .Y(exu_n28990));
OR2X1 exu_U1071(.A(exu_n15673), .B(alu_logic_rs1_data_bf1[54]), .Y(exu_n17311));
AND2X1 exu_U1072(.A(exu_n2938), .B(exu_n8018), .Y(exu_n27449));
AND2X1 exu_U1073(.A(exu_n2939), .B(exu_n8019), .Y(exu_n27448));
AND2X1 exu_U1074(.A(exu_n3242), .B(exu_n8322), .Y(exu_n28401));
AND2X1 exu_U1075(.A(exu_n3243), .B(exu_n8323), .Y(exu_n28400));
AND2X1 exu_U1076(.A(alu_logic_rs1_data_bf1[55]), .B(alu_logic_n110), .Y(alu_logic_result_and[55]));
OR2X1 exu_U1077(.A(alu_logic_n110), .B(alu_logic_rs1_data_bf1[55]), .Y(alu_logic_result_or[55]));
AND2X1 exu_U1078(.A(exu_n3428), .B(exu_n8509), .Y(exu_n28996));
OR2X1 exu_U1079(.A(exu_n15672), .B(alu_logic_rs1_data_bf1[53]), .Y(exu_n17306));
AND2X1 exu_U1080(.A(exu_n2940), .B(exu_n8020), .Y(exu_n27455));
AND2X1 exu_U1081(.A(exu_n2941), .B(exu_n8021), .Y(exu_n27454));
AND2X1 exu_U1082(.A(exu_n3244), .B(exu_n8324), .Y(exu_n28407));
AND2X1 exu_U1083(.A(exu_n3245), .B(exu_n8325), .Y(exu_n28406));
AND2X1 exu_U1084(.A(alu_logic_rs1_data_bf1[54]), .B(alu_logic_n111), .Y(alu_logic_result_and[54]));
OR2X1 exu_U1085(.A(alu_logic_n111), .B(alu_logic_rs1_data_bf1[54]), .Y(alu_logic_result_or[54]));
AND2X1 exu_U1086(.A(exu_n3430), .B(exu_n8511), .Y(exu_n29002));
OR2X1 exu_U1087(.A(exu_n15671), .B(alu_logic_rs1_data_bf1[52]), .Y(exu_n17301));
AND2X1 exu_U1088(.A(exu_n2942), .B(exu_n8022), .Y(exu_n27461));
AND2X1 exu_U1089(.A(exu_n2943), .B(exu_n8023), .Y(exu_n27460));
AND2X1 exu_U1090(.A(exu_n3246), .B(exu_n8326), .Y(exu_n28413));
AND2X1 exu_U1091(.A(exu_n3247), .B(exu_n8327), .Y(exu_n28412));
AND2X1 exu_U1092(.A(alu_logic_rs1_data_bf1[53]), .B(alu_logic_n112), .Y(alu_logic_result_and[53]));
OR2X1 exu_U1093(.A(alu_logic_n112), .B(alu_logic_rs1_data_bf1[53]), .Y(alu_logic_result_or[53]));
AND2X1 exu_U1094(.A(exu_n3432), .B(exu_n8513), .Y(exu_n29008));
OR2X1 exu_U1095(.A(exu_n15670), .B(alu_logic_rs1_data_bf1[51]), .Y(exu_n17296));
AND2X1 exu_U1096(.A(exu_n2944), .B(exu_n8024), .Y(exu_n27467));
AND2X1 exu_U1097(.A(exu_n2945), .B(exu_n8025), .Y(exu_n27466));
AND2X1 exu_U1098(.A(exu_n3248), .B(exu_n8328), .Y(exu_n28419));
AND2X1 exu_U1099(.A(exu_n3249), .B(exu_n8329), .Y(exu_n28418));
AND2X1 exu_U1100(.A(alu_logic_rs1_data_bf1[52]), .B(alu_logic_n113), .Y(alu_logic_result_and[52]));
OR2X1 exu_U1101(.A(alu_logic_n113), .B(alu_logic_rs1_data_bf1[52]), .Y(alu_logic_result_or[52]));
AND2X1 exu_U1102(.A(exu_n3434), .B(exu_n8515), .Y(exu_n29014));
OR2X1 exu_U1103(.A(exu_n15669), .B(alu_logic_rs1_data_bf1[50]), .Y(exu_n17289));
AND2X1 exu_U1104(.A(exu_n2946), .B(exu_n8026), .Y(exu_n27473));
AND2X1 exu_U1105(.A(exu_n2947), .B(exu_n8027), .Y(exu_n27472));
AND2X1 exu_U1106(.A(exu_n3250), .B(exu_n8330), .Y(exu_n28425));
AND2X1 exu_U1107(.A(exu_n3251), .B(exu_n8331), .Y(exu_n28424));
AND2X1 exu_U1108(.A(alu_logic_rs1_data_bf1[51]), .B(alu_logic_n114), .Y(alu_logic_result_and[51]));
OR2X1 exu_U1109(.A(alu_logic_n114), .B(alu_logic_rs1_data_bf1[51]), .Y(alu_logic_result_or[51]));
AND2X1 exu_U1110(.A(exu_n3436), .B(exu_n8517), .Y(exu_n29020));
OR2X1 exu_U1111(.A(exu_n15668), .B(alu_logic_rs1_data_bf1[49]), .Y(exu_n17284));
AND2X1 exu_U1112(.A(exu_n2948), .B(exu_n8028), .Y(exu_n27479));
AND2X1 exu_U1113(.A(exu_n2949), .B(exu_n8029), .Y(exu_n27478));
AND2X1 exu_U1114(.A(exu_n3252), .B(exu_n8332), .Y(exu_n28431));
AND2X1 exu_U1115(.A(exu_n3253), .B(exu_n8333), .Y(exu_n28430));
AND2X1 exu_U1116(.A(alu_logic_rs1_data_bf1[50]), .B(alu_logic_n115), .Y(alu_logic_result_and[50]));
OR2X1 exu_U1117(.A(alu_logic_n115), .B(alu_logic_rs1_data_bf1[50]), .Y(alu_logic_result_or[50]));
AND2X1 exu_U1118(.A(exu_n3438), .B(exu_n8519), .Y(exu_n29026));
OR2X1 exu_U1119(.A(exu_n15667), .B(alu_logic_rs1_data_bf1[48]), .Y(exu_n17279));
AND2X1 exu_U1120(.A(exu_n2952), .B(exu_n8032), .Y(exu_n27491));
AND2X1 exu_U1121(.A(exu_n2953), .B(exu_n8033), .Y(exu_n27490));
AND2X1 exu_U1122(.A(exu_n3256), .B(exu_n8336), .Y(exu_n28443));
AND2X1 exu_U1123(.A(exu_n3257), .B(exu_n8337), .Y(exu_n28442));
AND2X1 exu_U1124(.A(alu_logic_rs1_data_bf1[49]), .B(alu_logic_n117), .Y(alu_logic_result_and[49]));
OR2X1 exu_U1125(.A(alu_logic_n117), .B(alu_logic_rs1_data_bf1[49]), .Y(alu_logic_result_or[49]));
AND2X1 exu_U1126(.A(exu_n3442), .B(exu_n8523), .Y(exu_n29038));
OR2X1 exu_U1127(.A(exu_n15666), .B(alu_logic_rs1_data_bf1[47]), .Y(exu_n17274));
AND2X1 exu_U1128(.A(exu_n2954), .B(exu_n8034), .Y(exu_n27497));
AND2X1 exu_U1129(.A(exu_n2955), .B(exu_n8035), .Y(exu_n27496));
AND2X1 exu_U1130(.A(exu_n3258), .B(exu_n8338), .Y(exu_n28449));
AND2X1 exu_U1131(.A(exu_n3259), .B(exu_n8339), .Y(exu_n28448));
AND2X1 exu_U1132(.A(alu_logic_rs1_data_bf1[48]), .B(alu_logic_n118), .Y(alu_logic_result_and[48]));
OR2X1 exu_U1133(.A(alu_logic_n118), .B(alu_logic_rs1_data_bf1[48]), .Y(alu_logic_result_or[48]));
AND2X1 exu_U1134(.A(exu_n3444), .B(exu_n8525), .Y(exu_n29044));
AND2X1 exu_U1135(.A(exu_n2956), .B(exu_n8036), .Y(exu_n27503));
AND2X1 exu_U1136(.A(exu_n2957), .B(exu_n8037), .Y(exu_n27502));
AND2X1 exu_U1137(.A(exu_n3260), .B(exu_n8340), .Y(exu_n28455));
AND2X1 exu_U1138(.A(exu_n3261), .B(exu_n8341), .Y(exu_n28454));
AND2X1 exu_U1139(.A(alu_logic_rs1_data_bf1[47]), .B(alu_logic_n119), .Y(alu_logic_result_and[47]));
OR2X1 exu_U1140(.A(alu_logic_n119), .B(alu_logic_rs1_data_bf1[47]), .Y(alu_logic_result_or[47]));
AND2X1 exu_U1141(.A(exu_n3446), .B(exu_n8527), .Y(exu_n29050));
AND2X1 exu_U1142(.A(exu_n2958), .B(exu_n8038), .Y(exu_n27509));
AND2X1 exu_U1143(.A(exu_n2959), .B(exu_n8039), .Y(exu_n27508));
AND2X1 exu_U1144(.A(exu_n3262), .B(exu_n8342), .Y(exu_n28461));
AND2X1 exu_U1145(.A(exu_n3263), .B(exu_n8343), .Y(exu_n28460));
AND2X1 exu_U1146(.A(alu_logic_rs1_data_bf1[46]), .B(alu_logic_n120), .Y(alu_logic_result_and[46]));
OR2X1 exu_U1147(.A(alu_logic_n120), .B(alu_logic_rs1_data_bf1[46]), .Y(alu_logic_result_or[46]));
AND2X1 exu_U1148(.A(exu_n3448), .B(exu_n8529), .Y(exu_n29056));
AND2X1 exu_U1149(.A(exu_n2960), .B(exu_n8040), .Y(exu_n27515));
AND2X1 exu_U1150(.A(exu_n2961), .B(exu_n8041), .Y(exu_n27514));
AND2X1 exu_U1151(.A(exu_n3264), .B(exu_n8344), .Y(exu_n28467));
AND2X1 exu_U1152(.A(exu_n3265), .B(exu_n8345), .Y(exu_n28466));
AND2X1 exu_U1153(.A(alu_logic_rs1_data_bf1[45]), .B(alu_logic_n121), .Y(alu_logic_result_and[45]));
OR2X1 exu_U1154(.A(alu_logic_n121), .B(alu_logic_rs1_data_bf1[45]), .Y(alu_logic_result_or[45]));
AND2X1 exu_U1155(.A(exu_n3450), .B(exu_n8531), .Y(exu_n29062));
AND2X1 exu_U1156(.A(exu_n2962), .B(exu_n8042), .Y(exu_n27521));
AND2X1 exu_U1157(.A(exu_n2963), .B(exu_n8043), .Y(exu_n27520));
AND2X1 exu_U1158(.A(exu_n3266), .B(exu_n8346), .Y(exu_n28473));
AND2X1 exu_U1159(.A(exu_n3267), .B(exu_n8347), .Y(exu_n28472));
AND2X1 exu_U1160(.A(alu_logic_rs1_data_bf1[44]), .B(alu_logic_n122), .Y(alu_logic_result_and[44]));
OR2X1 exu_U1161(.A(alu_logic_n122), .B(alu_logic_rs1_data_bf1[44]), .Y(alu_logic_result_or[44]));
AND2X1 exu_U1162(.A(exu_n3452), .B(exu_n8533), .Y(exu_n29068));
AND2X1 exu_U1163(.A(exu_n2964), .B(exu_n8044), .Y(exu_n27527));
AND2X1 exu_U1164(.A(exu_n2965), .B(exu_n8045), .Y(exu_n27526));
AND2X1 exu_U1165(.A(exu_n3268), .B(exu_n8348), .Y(exu_n28479));
AND2X1 exu_U1166(.A(exu_n3269), .B(exu_n8349), .Y(exu_n28478));
AND2X1 exu_U1167(.A(alu_logic_rs1_data_bf1[43]), .B(alu_logic_n123), .Y(alu_logic_result_and[43]));
OR2X1 exu_U1168(.A(alu_logic_n123), .B(alu_logic_rs1_data_bf1[43]), .Y(alu_logic_result_or[43]));
AND2X1 exu_U1169(.A(exu_n3454), .B(exu_n8535), .Y(exu_n29074));
AND2X1 exu_U1170(.A(exu_n2966), .B(exu_n8046), .Y(exu_n27533));
AND2X1 exu_U1171(.A(exu_n2967), .B(exu_n8047), .Y(exu_n27532));
AND2X1 exu_U1172(.A(exu_n3270), .B(exu_n8350), .Y(exu_n28485));
AND2X1 exu_U1173(.A(exu_n3271), .B(exu_n8351), .Y(exu_n28484));
AND2X1 exu_U1174(.A(alu_logic_rs1_data_bf1[42]), .B(alu_logic_n124), .Y(alu_logic_result_and[42]));
OR2X1 exu_U1175(.A(alu_logic_n124), .B(alu_logic_rs1_data_bf1[42]), .Y(alu_logic_result_or[42]));
AND2X1 exu_U1176(.A(exu_n3456), .B(exu_n8537), .Y(exu_n29080));
AND2X1 exu_U1177(.A(exu_n2968), .B(exu_n8048), .Y(exu_n27539));
AND2X1 exu_U1178(.A(exu_n2969), .B(exu_n8049), .Y(exu_n27538));
AND2X1 exu_U1179(.A(exu_n3272), .B(exu_n8352), .Y(exu_n28491));
AND2X1 exu_U1180(.A(exu_n3273), .B(exu_n8353), .Y(exu_n28490));
AND2X1 exu_U1181(.A(alu_logic_rs1_data_bf1[41]), .B(alu_logic_n125), .Y(alu_logic_result_and[41]));
OR2X1 exu_U1182(.A(alu_logic_n125), .B(alu_logic_rs1_data_bf1[41]), .Y(alu_logic_result_or[41]));
AND2X1 exu_U1183(.A(exu_n3458), .B(exu_n8539), .Y(exu_n29086));
AND2X1 exu_U1184(.A(exu_n2970), .B(exu_n8050), .Y(exu_n27545));
AND2X1 exu_U1185(.A(exu_n2971), .B(exu_n8051), .Y(exu_n27544));
AND2X1 exu_U1186(.A(exu_n3274), .B(exu_n8354), .Y(exu_n28497));
AND2X1 exu_U1187(.A(exu_n3275), .B(exu_n8355), .Y(exu_n28496));
AND2X1 exu_U1188(.A(alu_logic_rs1_data_bf1[40]), .B(alu_logic_n126), .Y(alu_logic_result_and[40]));
OR2X1 exu_U1189(.A(alu_logic_n126), .B(alu_logic_rs1_data_bf1[40]), .Y(alu_logic_result_or[40]));
AND2X1 exu_U1190(.A(exu_n3460), .B(exu_n8541), .Y(exu_n29092));
AND2X1 exu_U1191(.A(exu_n2974), .B(exu_n8054), .Y(exu_n27557));
AND2X1 exu_U1192(.A(exu_n2975), .B(exu_n8055), .Y(exu_n27556));
AND2X1 exu_U1193(.A(exu_n3278), .B(exu_n8358), .Y(exu_n28509));
AND2X1 exu_U1194(.A(exu_n3279), .B(exu_n8359), .Y(exu_n28508));
AND2X1 exu_U1195(.A(alu_logic_rs1_data_bf1[39]), .B(alu_logic_n128), .Y(alu_logic_result_and[39]));
OR2X1 exu_U1196(.A(alu_logic_n128), .B(alu_logic_rs1_data_bf1[39]), .Y(alu_logic_result_or[39]));
AND2X1 exu_U1197(.A(exu_n3464), .B(exu_n8545), .Y(exu_n29104));
AND2X1 exu_U1198(.A(exu_n2976), .B(exu_n8056), .Y(exu_n27563));
AND2X1 exu_U1199(.A(exu_n2977), .B(exu_n8057), .Y(exu_n27562));
AND2X1 exu_U1200(.A(exu_n3280), .B(exu_n8360), .Y(exu_n28515));
AND2X1 exu_U1201(.A(exu_n3281), .B(exu_n8361), .Y(exu_n28514));
AND2X1 exu_U1202(.A(alu_logic_rs1_data_bf1[38]), .B(alu_logic_n129), .Y(alu_logic_result_and[38]));
OR2X1 exu_U1203(.A(alu_logic_n129), .B(alu_logic_rs1_data_bf1[38]), .Y(alu_logic_result_or[38]));
AND2X1 exu_U1204(.A(exu_n3466), .B(exu_n8547), .Y(exu_n29110));
AND2X1 exu_U1205(.A(exu_n2978), .B(exu_n8058), .Y(exu_n27569));
AND2X1 exu_U1206(.A(exu_n2979), .B(exu_n8059), .Y(exu_n27568));
AND2X1 exu_U1207(.A(exu_n3282), .B(exu_n8362), .Y(exu_n28521));
AND2X1 exu_U1208(.A(exu_n3283), .B(exu_n8363), .Y(exu_n28520));
AND2X1 exu_U1209(.A(alu_logic_rs1_data_bf1[37]), .B(alu_logic_n130), .Y(alu_logic_result_and[37]));
OR2X1 exu_U1210(.A(alu_logic_n130), .B(alu_logic_rs1_data_bf1[37]), .Y(alu_logic_result_or[37]));
AND2X1 exu_U1211(.A(exu_n3468), .B(exu_n8549), .Y(exu_n29116));
AND2X1 exu_U1212(.A(exu_n2980), .B(exu_n8060), .Y(exu_n27575));
AND2X1 exu_U1213(.A(exu_n2981), .B(exu_n8061), .Y(exu_n27574));
AND2X1 exu_U1214(.A(exu_n3284), .B(exu_n8364), .Y(exu_n28527));
AND2X1 exu_U1215(.A(exu_n3285), .B(exu_n8365), .Y(exu_n28526));
AND2X1 exu_U1216(.A(alu_logic_rs1_data_bf1[36]), .B(alu_logic_n131), .Y(alu_logic_result_and[36]));
OR2X1 exu_U1217(.A(alu_logic_n131), .B(alu_logic_rs1_data_bf1[36]), .Y(alu_logic_result_or[36]));
AND2X1 exu_U1218(.A(exu_n3470), .B(exu_n8551), .Y(exu_n29122));
AND2X1 exu_U1219(.A(exu_n2982), .B(exu_n8062), .Y(exu_n27581));
AND2X1 exu_U1220(.A(exu_n2983), .B(exu_n8063), .Y(exu_n27580));
AND2X1 exu_U1221(.A(exu_n3286), .B(exu_n8366), .Y(exu_n28533));
AND2X1 exu_U1222(.A(exu_n3287), .B(exu_n8367), .Y(exu_n28532));
AND2X1 exu_U1223(.A(alu_logic_rs1_data_bf1[35]), .B(alu_logic_n132), .Y(alu_logic_result_and[35]));
OR2X1 exu_U1224(.A(alu_logic_n132), .B(alu_logic_rs1_data_bf1[35]), .Y(alu_logic_result_or[35]));
AND2X1 exu_U1225(.A(exu_n3472), .B(exu_n8553), .Y(exu_n29128));
AND2X1 exu_U1226(.A(exu_n2984), .B(exu_n8064), .Y(exu_n27587));
AND2X1 exu_U1227(.A(exu_n2985), .B(exu_n8065), .Y(exu_n27586));
AND2X1 exu_U1228(.A(exu_n3288), .B(exu_n8368), .Y(exu_n28539));
AND2X1 exu_U1229(.A(exu_n3289), .B(exu_n8369), .Y(exu_n28538));
AND2X1 exu_U1230(.A(alu_logic_rs1_data_bf1[34]), .B(alu_logic_n133), .Y(alu_logic_result_and[34]));
OR2X1 exu_U1231(.A(alu_logic_n133), .B(alu_logic_rs1_data_bf1[34]), .Y(alu_logic_result_or[34]));
AND2X1 exu_U1232(.A(exu_n3474), .B(exu_n8555), .Y(exu_n29134));
AND2X1 exu_U1233(.A(exu_n2986), .B(exu_n8066), .Y(exu_n27593));
AND2X1 exu_U1234(.A(exu_n2987), .B(exu_n8067), .Y(exu_n27592));
AND2X1 exu_U1235(.A(exu_n3290), .B(exu_n8370), .Y(exu_n28545));
AND2X1 exu_U1236(.A(exu_n3291), .B(exu_n8371), .Y(exu_n28544));
AND2X1 exu_U1237(.A(alu_logic_rs1_data_bf1[33]), .B(alu_logic_n134), .Y(alu_logic_result_and[33]));
OR2X1 exu_U1238(.A(alu_logic_n134), .B(alu_logic_rs1_data_bf1[33]), .Y(alu_logic_result_or[33]));
AND2X1 exu_U1239(.A(exu_n3476), .B(exu_n8557), .Y(exu_n29140));
AND2X1 exu_U1240(.A(exu_n2988), .B(exu_n8068), .Y(exu_n27599));
AND2X1 exu_U1241(.A(exu_n2989), .B(exu_n8069), .Y(exu_n27598));
AND2X1 exu_U1242(.A(exu_n3292), .B(exu_n8372), .Y(exu_n28551));
AND2X1 exu_U1243(.A(exu_n3293), .B(exu_n8373), .Y(exu_n28550));
AND2X1 exu_U1244(.A(alu_logic_rs1_data_bf1[32]), .B(alu_logic_n135), .Y(alu_logic_result_and[32]));
OR2X1 exu_U1245(.A(alu_logic_n135), .B(alu_logic_rs1_data_bf1[32]), .Y(alu_logic_result_or[32]));
AND2X1 exu_U1246(.A(exu_n3478), .B(exu_n8559), .Y(exu_n29146));
AND2X1 exu_U1247(.A(exu_n2990), .B(exu_n8070), .Y(exu_n27605));
AND2X1 exu_U1248(.A(exu_n2991), .B(exu_n8071), .Y(exu_n27604));
AND2X1 exu_U1249(.A(exu_n3294), .B(exu_n8374), .Y(exu_n28557));
AND2X1 exu_U1250(.A(exu_n3295), .B(exu_n8375), .Y(exu_n28556));
AND2X1 exu_U1251(.A(exu_n2992), .B(exu_n8072), .Y(exu_n27611));
AND2X1 exu_U1252(.A(exu_n2993), .B(exu_n8073), .Y(exu_n27610));
AND2X1 exu_U1253(.A(exu_n3296), .B(exu_n8376), .Y(exu_n28563));
AND2X1 exu_U1254(.A(exu_n3297), .B(exu_n8377), .Y(exu_n28562));
AND2X1 exu_U1255(.A(alu_logic_rs1_data_bf1[30]), .B(alu_logic_n137), .Y(alu_logic_result_and[30]));
OR2X1 exu_U1256(.A(alu_logic_n137), .B(alu_logic_rs1_data_bf1[30]), .Y(alu_logic_result_or[30]));
AND2X1 exu_U1257(.A(exu_n3482), .B(exu_n8563), .Y(exu_n29158));
AND2X1 exu_U1258(.A(exu_n2996), .B(exu_n8076), .Y(exu_n27623));
AND2X1 exu_U1259(.A(exu_n2997), .B(exu_n8077), .Y(exu_n27622));
AND2X1 exu_U1260(.A(exu_n3299), .B(exu_n8379), .Y(exu_n28573));
AND2X1 exu_U1261(.A(exu_n3300), .B(exu_n8380), .Y(exu_n28572));
AND2X1 exu_U1262(.A(alu_logic_rs1_data_bf1[29]), .B(alu_logic_n139), .Y(alu_logic_result_and[29]));
OR2X1 exu_U1263(.A(alu_logic_n139), .B(alu_logic_rs1_data_bf1[29]), .Y(alu_logic_result_or[29]));
AND2X1 exu_U1264(.A(exu_n3486), .B(exu_n8567), .Y(exu_n29170));
AND2X1 exu_U1265(.A(exu_n2998), .B(exu_n8078), .Y(exu_n27629));
AND2X1 exu_U1266(.A(exu_n2999), .B(exu_n8079), .Y(exu_n27628));
AND2X1 exu_U1267(.A(exu_n3301), .B(exu_n8381), .Y(exu_n28579));
AND2X1 exu_U1268(.A(exu_n3302), .B(exu_n8382), .Y(exu_n28578));
AND2X1 exu_U1269(.A(alu_logic_rs1_data_bf1[28]), .B(alu_logic_n140), .Y(alu_logic_result_and[28]));
OR2X1 exu_U1270(.A(alu_logic_n140), .B(alu_logic_rs1_data_bf1[28]), .Y(alu_logic_result_or[28]));
AND2X1 exu_U1271(.A(exu_n3488), .B(exu_n8569), .Y(exu_n29176));
AND2X1 exu_U1272(.A(exu_n3000), .B(exu_n8080), .Y(exu_n27635));
AND2X1 exu_U1273(.A(exu_n3001), .B(exu_n8081), .Y(exu_n27634));
AND2X1 exu_U1274(.A(exu_n3303), .B(exu_n8383), .Y(exu_n28585));
AND2X1 exu_U1275(.A(exu_n3304), .B(exu_n8384), .Y(exu_n28584));
AND2X1 exu_U1276(.A(alu_logic_rs1_data_bf1[27]), .B(alu_logic_n141), .Y(alu_logic_result_and[27]));
OR2X1 exu_U1277(.A(alu_logic_n141), .B(alu_logic_rs1_data_bf1[27]), .Y(alu_logic_result_or[27]));
AND2X1 exu_U1278(.A(exu_n3490), .B(exu_n8571), .Y(exu_n29182));
AND2X1 exu_U1279(.A(exu_n3002), .B(exu_n8082), .Y(exu_n27641));
AND2X1 exu_U1280(.A(exu_n3003), .B(exu_n8083), .Y(exu_n27640));
AND2X1 exu_U1281(.A(exu_n3305), .B(exu_n8385), .Y(exu_n28591));
AND2X1 exu_U1282(.A(exu_n3306), .B(exu_n8386), .Y(exu_n28590));
AND2X1 exu_U1283(.A(alu_logic_rs1_data_bf1[26]), .B(alu_logic_n142), .Y(alu_logic_result_and[26]));
OR2X1 exu_U1284(.A(alu_logic_n142), .B(alu_logic_rs1_data_bf1[26]), .Y(alu_logic_result_or[26]));
AND2X1 exu_U1285(.A(exu_n3492), .B(exu_n8573), .Y(exu_n29188));
AND2X1 exu_U1286(.A(exu_n3004), .B(exu_n8084), .Y(exu_n27647));
AND2X1 exu_U1287(.A(exu_n3005), .B(exu_n8085), .Y(exu_n27646));
AND2X1 exu_U1288(.A(exu_n3307), .B(exu_n8387), .Y(exu_n28597));
AND2X1 exu_U1289(.A(exu_n3308), .B(exu_n8388), .Y(exu_n28596));
AND2X1 exu_U1290(.A(alu_logic_rs1_data_bf1[25]), .B(alu_logic_n143), .Y(alu_logic_result_and[25]));
OR2X1 exu_U1291(.A(alu_logic_n143), .B(alu_logic_rs1_data_bf1[25]), .Y(alu_logic_result_or[25]));
AND2X1 exu_U1292(.A(exu_n3494), .B(exu_n8575), .Y(exu_n29194));
AND2X1 exu_U1293(.A(exu_n3006), .B(exu_n8086), .Y(exu_n27653));
AND2X1 exu_U1294(.A(exu_n3007), .B(exu_n8087), .Y(exu_n27652));
AND2X1 exu_U1295(.A(exu_n3309), .B(exu_n8389), .Y(exu_n28603));
AND2X1 exu_U1296(.A(exu_n3310), .B(exu_n8390), .Y(exu_n28602));
AND2X1 exu_U1297(.A(alu_logic_rs1_data_bf1[24]), .B(alu_logic_n144), .Y(alu_logic_result_and[24]));
OR2X1 exu_U1298(.A(alu_logic_n144), .B(alu_logic_rs1_data_bf1[24]), .Y(alu_logic_result_or[24]));
AND2X1 exu_U1299(.A(exu_n3496), .B(exu_n8577), .Y(exu_n29200));
AND2X1 exu_U1300(.A(exu_n3008), .B(exu_n8088), .Y(exu_n27659));
AND2X1 exu_U1301(.A(exu_n3009), .B(exu_n8089), .Y(exu_n27658));
AND2X1 exu_U1302(.A(exu_n3311), .B(exu_n8391), .Y(exu_n28609));
AND2X1 exu_U1303(.A(exu_n3312), .B(exu_n8392), .Y(exu_n28608));
AND2X1 exu_U1304(.A(alu_logic_rs1_data_bf1[23]), .B(alu_logic_n145), .Y(alu_logic_result_and[23]));
OR2X1 exu_U1305(.A(alu_logic_n145), .B(alu_logic_rs1_data_bf1[23]), .Y(alu_logic_result_or[23]));
AND2X1 exu_U1306(.A(exu_n3498), .B(exu_n8579), .Y(exu_n29206));
AND2X1 exu_U1307(.A(exu_n3010), .B(exu_n8090), .Y(exu_n27665));
AND2X1 exu_U1308(.A(exu_n3011), .B(exu_n8091), .Y(exu_n27664));
AND2X1 exu_U1309(.A(exu_n3313), .B(exu_n8393), .Y(exu_n28615));
AND2X1 exu_U1310(.A(exu_n3314), .B(exu_n8394), .Y(exu_n28614));
AND2X1 exu_U1311(.A(alu_logic_rs1_data_bf1[22]), .B(alu_logic_n146), .Y(alu_logic_result_and[22]));
OR2X1 exu_U1312(.A(alu_logic_n146), .B(alu_logic_rs1_data_bf1[22]), .Y(alu_logic_result_or[22]));
AND2X1 exu_U1313(.A(exu_n3500), .B(exu_n8581), .Y(exu_n29212));
AND2X1 exu_U1314(.A(exu_n3012), .B(exu_n8092), .Y(exu_n27671));
AND2X1 exu_U1315(.A(exu_n3013), .B(exu_n8093), .Y(exu_n27670));
AND2X1 exu_U1316(.A(exu_n3315), .B(exu_n8395), .Y(exu_n28621));
AND2X1 exu_U1317(.A(exu_n3316), .B(exu_n8396), .Y(exu_n28620));
AND2X1 exu_U1318(.A(alu_logic_rs1_data_bf1[21]), .B(alu_logic_n147), .Y(alu_logic_result_and[21]));
OR2X1 exu_U1319(.A(alu_logic_n147), .B(alu_logic_rs1_data_bf1[21]), .Y(alu_logic_result_or[21]));
AND2X1 exu_U1320(.A(exu_n3502), .B(exu_n8583), .Y(exu_n29218));
AND2X1 exu_U1321(.A(exu_n3014), .B(exu_n8094), .Y(exu_n27677));
AND2X1 exu_U1322(.A(exu_n3015), .B(exu_n8095), .Y(exu_n27676));
AND2X1 exu_U1323(.A(exu_n3317), .B(exu_n8397), .Y(exu_n28627));
AND2X1 exu_U1324(.A(exu_n3318), .B(exu_n8398), .Y(exu_n28626));
AND2X1 exu_U1325(.A(alu_logic_rs1_data_bf1[20]), .B(alu_logic_n148), .Y(alu_logic_result_and[20]));
OR2X1 exu_U1326(.A(alu_logic_n148), .B(alu_logic_rs1_data_bf1[20]), .Y(alu_logic_result_or[20]));
AND2X1 exu_U1327(.A(exu_n3504), .B(exu_n8585), .Y(exu_n29224));
AND2X1 exu_U1328(.A(exu_n3018), .B(exu_n8098), .Y(exu_n27689));
AND2X1 exu_U1329(.A(exu_n3019), .B(exu_n8099), .Y(exu_n27688));
AND2X1 exu_U1330(.A(exu_n3319), .B(exu_n8400), .Y(exu_n28636));
AND2X1 exu_U1331(.A(exu_n3320), .B(exu_n8401), .Y(exu_n28635));
AND2X1 exu_U1332(.A(alu_logic_rs1_data_bf1[19]), .B(alu_logic_n150), .Y(alu_logic_result_and[19]));
OR2X1 exu_U1333(.A(alu_logic_n150), .B(alu_logic_rs1_data_bf1[19]), .Y(alu_logic_result_or[19]));
AND2X1 exu_U1334(.A(exu_n3508), .B(exu_n8589), .Y(exu_n29236));
AND2X1 exu_U1335(.A(exu_n3020), .B(exu_n8100), .Y(exu_n27695));
AND2X1 exu_U1336(.A(exu_n3021), .B(exu_n8101), .Y(exu_n27694));
AND2X1 exu_U1337(.A(exu_n3321), .B(exu_n8402), .Y(exu_n28642));
AND2X1 exu_U1338(.A(exu_n3322), .B(exu_n8403), .Y(exu_n28641));
AND2X1 exu_U1339(.A(alu_logic_rs1_data_bf1[18]), .B(alu_logic_n151), .Y(alu_logic_result_and[18]));
OR2X1 exu_U1340(.A(alu_logic_n151), .B(alu_logic_rs1_data_bf1[18]), .Y(alu_logic_result_or[18]));
AND2X1 exu_U1341(.A(exu_n3510), .B(exu_n8591), .Y(exu_n29242));
AND2X1 exu_U1342(.A(exu_n3022), .B(exu_n8102), .Y(exu_n27701));
AND2X1 exu_U1343(.A(exu_n3023), .B(exu_n8103), .Y(exu_n27700));
AND2X1 exu_U1344(.A(exu_n3323), .B(exu_n8404), .Y(exu_n28648));
AND2X1 exu_U1345(.A(exu_n3324), .B(exu_n8405), .Y(exu_n28647));
AND2X1 exu_U1346(.A(alu_logic_rs1_data_bf1[17]), .B(alu_logic_n152), .Y(alu_logic_result_and[17]));
OR2X1 exu_U1347(.A(alu_logic_n152), .B(alu_logic_rs1_data_bf1[17]), .Y(alu_logic_result_or[17]));
AND2X1 exu_U1348(.A(exu_n3512), .B(exu_n8593), .Y(exu_n29248));
AND2X1 exu_U1349(.A(exu_n3024), .B(exu_n8104), .Y(exu_n27707));
AND2X1 exu_U1350(.A(exu_n3025), .B(exu_n8105), .Y(exu_n27706));
AND2X1 exu_U1351(.A(exu_n3325), .B(exu_n8406), .Y(exu_n28654));
AND2X1 exu_U1352(.A(exu_n3326), .B(exu_n8407), .Y(exu_n28653));
AND2X1 exu_U1353(.A(alu_logic_rs1_data_bf1[16]), .B(alu_logic_n153), .Y(alu_logic_result_and[16]));
OR2X1 exu_U1354(.A(alu_logic_n153), .B(alu_logic_rs1_data_bf1[16]), .Y(alu_logic_result_or[16]));
AND2X1 exu_U1355(.A(exu_n3514), .B(exu_n8595), .Y(exu_n29254));
AND2X1 exu_U1356(.A(exu_n3026), .B(exu_n8106), .Y(exu_n27713));
AND2X1 exu_U1357(.A(exu_n3027), .B(exu_n8107), .Y(exu_n27712));
AND2X1 exu_U1358(.A(exu_n3327), .B(exu_n8408), .Y(exu_n28660));
AND2X1 exu_U1359(.A(exu_n3328), .B(exu_n8409), .Y(exu_n28659));
AND2X1 exu_U1360(.A(alu_logic_rs1_data_bf1[15]), .B(alu_logic_n154), .Y(alu_logic_result_and[15]));
OR2X1 exu_U1361(.A(alu_logic_n154), .B(alu_logic_rs1_data_bf1[15]), .Y(alu_logic_result_or[15]));
AND2X1 exu_U1362(.A(exu_n3516), .B(exu_n8597), .Y(exu_n29260));
AND2X1 exu_U1363(.A(exu_n3028), .B(exu_n8108), .Y(exu_n27719));
AND2X1 exu_U1364(.A(exu_n3029), .B(exu_n8109), .Y(exu_n27718));
AND2X1 exu_U1365(.A(exu_n3329), .B(exu_n8410), .Y(exu_n28666));
AND2X1 exu_U1366(.A(exu_n3330), .B(exu_n8411), .Y(exu_n28665));
AND2X1 exu_U1367(.A(alu_logic_rs1_data_bf1[14]), .B(alu_logic_n155), .Y(alu_logic_result_and[14]));
OR2X1 exu_U1368(.A(alu_logic_n155), .B(alu_logic_rs1_data_bf1[14]), .Y(alu_logic_result_or[14]));
AND2X1 exu_U1369(.A(exu_n3518), .B(exu_n8599), .Y(exu_n29266));
AND2X1 exu_U1370(.A(exu_n3030), .B(exu_n8110), .Y(exu_n27725));
AND2X1 exu_U1371(.A(exu_n3031), .B(exu_n8111), .Y(exu_n27724));
AND2X1 exu_U1372(.A(exu_n3331), .B(exu_n8412), .Y(exu_n28672));
AND2X1 exu_U1373(.A(exu_n3332), .B(exu_n8413), .Y(exu_n28671));
AND2X1 exu_U1374(.A(alu_logic_rs1_data_bf1[13]), .B(alu_logic_n156), .Y(alu_logic_result_and[13]));
OR2X1 exu_U1375(.A(alu_logic_n156), .B(alu_logic_rs1_data_bf1[13]), .Y(alu_logic_result_or[13]));
AND2X1 exu_U1376(.A(exu_n3520), .B(exu_n8601), .Y(exu_n29272));
AND2X1 exu_U1377(.A(exu_n3032), .B(exu_n8112), .Y(exu_n27731));
AND2X1 exu_U1378(.A(exu_n3033), .B(exu_n8113), .Y(exu_n27730));
AND2X1 exu_U1379(.A(exu_n3333), .B(exu_n8414), .Y(exu_n28678));
AND2X1 exu_U1380(.A(exu_n3334), .B(exu_n8415), .Y(exu_n28677));
AND2X1 exu_U1381(.A(alu_logic_rs1_data_bf1[12]), .B(alu_logic_n157), .Y(alu_logic_result_and[12]));
OR2X1 exu_U1382(.A(alu_logic_n157), .B(alu_logic_rs1_data_bf1[12]), .Y(alu_logic_result_or[12]));
AND2X1 exu_U1383(.A(exu_n3522), .B(exu_n8603), .Y(exu_n29278));
AND2X1 exu_U1384(.A(exu_n3034), .B(exu_n8114), .Y(exu_n27737));
AND2X1 exu_U1385(.A(exu_n3035), .B(exu_n8115), .Y(exu_n27736));
AND2X1 exu_U1386(.A(exu_n3335), .B(exu_n8416), .Y(exu_n28684));
AND2X1 exu_U1387(.A(exu_n3336), .B(exu_n8417), .Y(exu_n28683));
AND2X1 exu_U1388(.A(alu_logic_rs1_data_bf1[11]), .B(alu_logic_n158), .Y(alu_logic_result_and[11]));
OR2X1 exu_U1389(.A(alu_logic_n158), .B(alu_logic_rs1_data_bf1[11]), .Y(alu_logic_result_or[11]));
AND2X1 exu_U1390(.A(exu_n3524), .B(exu_n8605), .Y(exu_n29284));
AND2X1 exu_U1391(.A(exu_n3036), .B(exu_n8116), .Y(exu_n27743));
AND2X1 exu_U1392(.A(exu_n3037), .B(exu_n8117), .Y(exu_n27742));
AND2X1 exu_U1393(.A(exu_n3337), .B(exu_n8418), .Y(exu_n28690));
AND2X1 exu_U1394(.A(exu_n3338), .B(exu_n8419), .Y(exu_n28689));
AND2X1 exu_U1395(.A(alu_logic_rs1_data_bf1[10]), .B(alu_logic_n159), .Y(alu_logic_result_and[10]));
OR2X1 exu_U1396(.A(alu_logic_n159), .B(alu_logic_rs1_data_bf1[10]), .Y(alu_logic_result_or[10]));
AND2X1 exu_U1397(.A(exu_n3526), .B(exu_n8607), .Y(exu_n29290));
AND2X1 exu_U1398(.A(exu_n2915), .B(exu_n7996), .Y(exu_n27381));
AND2X1 exu_U1399(.A(exu_n2916), .B(exu_n7997), .Y(exu_n27380));
AND2X1 exu_U1400(.A(exu_n3218), .B(exu_n8298), .Y(exu_n28329));
AND2X1 exu_U1401(.A(exu_n3219), .B(exu_n8299), .Y(exu_n28328));
AND2X1 exu_U1402(.A(alu_logic_rs1_data_bf1[8]), .B(alu_logic_n98), .Y(alu_logic_result_and[8]));
OR2X1 exu_U1403(.A(alu_logic_n98), .B(alu_logic_rs1_data_bf1[8]), .Y(alu_logic_result_or[8]));
AND2X1 exu_U1404(.A(exu_n3404), .B(exu_n8485), .Y(exu_n28924));
AND2X1 exu_U1405(.A(exu_n2917), .B(exu_n7998), .Y(exu_n27387));
AND2X1 exu_U1406(.A(exu_n2918), .B(exu_n7999), .Y(exu_n27386));
AND2X1 exu_U1407(.A(exu_n3220), .B(exu_n8300), .Y(exu_n28335));
AND2X1 exu_U1408(.A(exu_n3221), .B(exu_n8301), .Y(exu_n28334));
AND2X1 exu_U1409(.A(alu_logic_rs1_data_bf1[7]), .B(alu_logic_n99), .Y(alu_logic_result_and[7]));
OR2X1 exu_U1410(.A(alu_logic_n99), .B(alu_logic_rs1_data_bf1[7]), .Y(alu_logic_result_or[7]));
AND2X1 exu_U1411(.A(exu_n3406), .B(exu_n8487), .Y(exu_n28930));
AND2X1 exu_U1412(.A(exu_n2919), .B(exu_n8000), .Y(exu_n27393));
AND2X1 exu_U1413(.A(exu_n2920), .B(exu_n8001), .Y(exu_n27392));
AND2X1 exu_U1414(.A(exu_n3222), .B(exu_n8302), .Y(exu_n28341));
AND2X1 exu_U1415(.A(exu_n3223), .B(exu_n8303), .Y(exu_n28340));
AND2X1 exu_U1416(.A(alu_logic_rs1_data_bf1[6]), .B(alu_logic_n100), .Y(alu_logic_result_and[6]));
OR2X1 exu_U1417(.A(alu_logic_n100), .B(alu_logic_rs1_data_bf1[6]), .Y(alu_logic_result_or[6]));
AND2X1 exu_U1418(.A(exu_n3408), .B(exu_n8489), .Y(exu_n28936));
AND2X1 exu_U1419(.A(exu_n2928), .B(exu_n8008), .Y(exu_n27419));
AND2X1 exu_U1420(.A(exu_n2929), .B(exu_n8009), .Y(exu_n27418));
AND2X1 exu_U1421(.A(exu_n3232), .B(exu_n8312), .Y(exu_n28371));
AND2X1 exu_U1422(.A(exu_n3233), .B(exu_n8313), .Y(exu_n28370));
AND2X1 exu_U1423(.A(alu_logic_rs1_data_bf1[5]), .B(alu_logic_n105), .Y(alu_logic_result_and[5]));
OR2X1 exu_U1424(.A(alu_logic_n105), .B(alu_logic_rs1_data_bf1[5]), .Y(alu_logic_result_or[5]));
AND2X1 exu_U1425(.A(exu_n3418), .B(exu_n8499), .Y(exu_n28966));
AND2X1 exu_U1426(.A(exu_n2950), .B(exu_n8030), .Y(exu_n27485));
AND2X1 exu_U1427(.A(exu_n2951), .B(exu_n8031), .Y(exu_n27484));
AND2X1 exu_U1428(.A(exu_n3254), .B(exu_n8334), .Y(exu_n28437));
AND2X1 exu_U1429(.A(exu_n3255), .B(exu_n8335), .Y(exu_n28436));
AND2X1 exu_U1430(.A(alu_logic_rs1_data_bf1[4]), .B(alu_logic_n116), .Y(alu_logic_result_and[4]));
OR2X1 exu_U1431(.A(alu_logic_n116), .B(alu_logic_rs1_data_bf1[4]), .Y(alu_logic_result_or[4]));
AND2X1 exu_U1432(.A(exu_n3440), .B(exu_n8521), .Y(exu_n29032));
AND2X1 exu_U1433(.A(exu_n2972), .B(exu_n8052), .Y(exu_n27551));
AND2X1 exu_U1434(.A(exu_n2973), .B(exu_n8053), .Y(exu_n27550));
AND2X1 exu_U1435(.A(exu_n3276), .B(exu_n8356), .Y(exu_n28503));
AND2X1 exu_U1436(.A(exu_n3277), .B(exu_n8357), .Y(exu_n28502));
AND2X1 exu_U1437(.A(alu_logic_rs1_data_bf1[3]), .B(alu_logic_n127), .Y(alu_logic_result_and[3]));
OR2X1 exu_U1438(.A(alu_logic_n127), .B(alu_logic_rs1_data_bf1[3]), .Y(alu_logic_result_or[3]));
AND2X1 exu_U1439(.A(exu_n3462), .B(exu_n8543), .Y(exu_n29098));
AND2X1 exu_U1440(.A(exu_n2994), .B(exu_n8074), .Y(exu_n27617));
AND2X1 exu_U1441(.A(exu_n2995), .B(exu_n8075), .Y(exu_n27616));
AND2X1 exu_U1442(.A(exu_n3298), .B(exu_n8378), .Y(exu_n28568));
AND2X1 exu_U1443(.A(alu_logic_rs1_data_bf1[2]), .B(alu_logic_n138), .Y(alu_logic_result_and[2]));
OR2X1 exu_U1444(.A(alu_logic_n138), .B(alu_logic_rs1_data_bf1[2]), .Y(alu_logic_result_or[2]));
AND2X1 exu_U1445(.A(exu_n3484), .B(exu_n8565), .Y(exu_n29164));
AND2X1 exu_U1446(.A(exu_n3016), .B(exu_n8096), .Y(exu_n27683));
AND2X1 exu_U1447(.A(exu_n3017), .B(exu_n8097), .Y(exu_n27682));
AND2X1 exu_U1448(.A(alu_logic_rs1_data_bf1[1]), .B(alu_logic_n149), .Y(alu_logic_result_and[1]));
OR2X1 exu_U1449(.A(alu_logic_n149), .B(alu_logic_rs1_data_bf1[1]), .Y(alu_logic_result_or[1]));
AND2X1 exu_U1450(.A(exu_n3506), .B(exu_n8587), .Y(exu_n29230));
AND2X1 exu_U1451(.A(exu_n3038), .B(exu_n8118), .Y(exu_n27749));
AND2X1 exu_U1452(.A(exu_n3039), .B(exu_n8119), .Y(exu_n27748));
AND2X1 exu_U1453(.A(alu_logic_rs1_data_bf1[0]), .B(alu_logic_n160), .Y(alu_logic_result_and[0]));
OR2X1 exu_U1454(.A(alu_logic_n160), .B(alu_logic_rs1_data_bf1[0]), .Y(alu_logic_result_or[0]));
AND2X1 exu_U1455(.A(exu_n3528), .B(exu_n8609), .Y(exu_n29296));
OR2X1 exu_U1456(.A(exu_n13454), .B(exu_n14774), .Y(ecc_decode_n23));
AND2X1 exu_U1457(.A(exu_n15459), .B(exu_n15202), .Y(ecc_decode_n37));
AND2X1 exu_U1458(.A(exu_n15202), .B(ecc_err_m[4]), .Y(ecc_decode_n43));
AND2X1 exu_U1459(.A(exu_n4585), .B(exu_n9371), .Y(ecc_syn_mux_n21));
AND2X1 exu_U1460(.A(exu_n4582), .B(exu_n9365), .Y(ecc_syn_mux_n9));
AND2X1 exu_U1461(.A(exu_n4584), .B(exu_n9369), .Y(ecc_syn_mux_n17));
AND2X1 exu_U1462(.A(exu_n156), .B(exu_n5122), .Y(exu_n17454));
AND2X1 exu_U1463(.A(exu_n14), .B(exu_n4983), .Y(exu_n16678));
AND2X1 exu_U1464(.A(alu_logic_rs1_data_bf1[9]), .B(alu_logic_n97), .Y(alu_logic_result_and[9]));
OR2X1 exu_U1465(.A(alu_logic_n97), .B(alu_logic_rs1_data_bf1[9]), .Y(alu_logic_result_or[9]));
AND2X1 exu_U1466(.A(exu_n3402), .B(exu_n8483), .Y(exu_n28918));
OR2X1 exu_U1467(.A(exu_n13104), .B(exu_n14390), .Y(shft_rshift1[9]));
OR2X1 exu_U1468(.A(exu_n13235), .B(exu_n14542), .Y(shft_lshift1[9]));
AND2X1 exu_U1469(.A(exu_n17396), .B(ecl_rd_e[0]), .Y(exu_n17398));
INVX1 exu_U1470(.A(lsu_exu_st_dtlb_perr_g), .Y(exu_n16372));
AND2X1 exu_U1471(.A(exu_n11), .B(exu_n4981), .Y(exu_n16650));
INVX1 exu_U1472(.A(ecl_ifu_exu_aluop_e[0]), .Y(exu_n16400));
AND2X1 exu_U1473(.A(exu_n4918), .B(exu_n9632), .Y(div_n71));
AND2X1 exu_U1474(.A(exu_n4921), .B(exu_n9634), .Y(div_n77));
AND2X1 exu_U1475(.A(exu_n4923), .B(exu_n9637), .Y(div_n85));
AND2X1 exu_U1476(.A(exu_n4926), .B(exu_n9639), .Y(div_n91));
AND2X1 exu_U1477(.A(exu_n4913), .B(exu_n9627), .Y(div_n55));
AND2X1 exu_U1478(.A(exu_n4912), .B(exu_n9626), .Y(div_n56));
AND2X1 exu_U1479(.A(exu_n4916), .B(exu_n9629), .Y(div_n61));
AND2X1 exu_U1480(.A(exu_n4915), .B(exu_n9628), .Y(div_n62));
AND2X1 exu_U1481(.A(exu_n4911), .B(exu_n9624), .Y(div_n47));
AND2X1 exu_U1482(.A(exu_n4910), .B(exu_n9623), .Y(div_n48));
AND2X1 exu_U1483(.A(exu_n4907), .B(exu_n9621), .Y(div_n42));
INVX1 exu_U1484(.A(ecl_writeback_sraddr_w[2]), .Y(exu_n16555));
AND2X1 exu_U1485(.A(ecl_writeback_n58), .B(ecl_writeback_sraddr_w[3]), .Y(ecl_writeback_n144));
AND2X1 exu_U1486(.A(exu_n3718), .B(exu_n8797), .Y(div_gencc_in[57]));
AND2X1 exu_U1487(.A(exu_n3720), .B(exu_n8799), .Y(div_gencc_in[55]));
AND2X1 exu_U1488(.A(exu_n3719), .B(exu_n8798), .Y(div_gencc_in[56]));
AND2X1 exu_U1489(.A(exu_n3733), .B(exu_n8812), .Y(div_gencc_in[43]));
AND2X1 exu_U1490(.A(exu_n3735), .B(exu_n8814), .Y(div_gencc_in[41]));
AND2X1 exu_U1491(.A(exu_n3734), .B(exu_n8813), .Y(div_gencc_in[42]));
AND2X1 exu_U1492(.A(exu_n3725), .B(exu_n8804), .Y(div_gencc_in[50]));
AND2X1 exu_U1493(.A(exu_n3728), .B(exu_n8807), .Y(div_gencc_in[48]));
AND2X1 exu_U1494(.A(exu_n3727), .B(exu_n8806), .Y(div_gencc_in[49]));
AND2X1 exu_U1495(.A(exu_n3755), .B(exu_n8834), .Y(div_gencc_in_23));
AND2X1 exu_U1496(.A(exu_n3707), .B(exu_n10243), .Y(div_gencc_in_9));
OR2X1 exu_U1497(.A(alu_addsub_rs2_data[37]), .B(alu_logic_rs1_data_bf1[37]), .Y(exu_n31553));
AND2X1 exu_U1498(.A(exu_n3674), .B(exu_n8691), .Y(alu_zcomp_in[39]));
OR2X1 exu_U1499(.A(alu_addsub_rs2_data[35]), .B(alu_logic_rs1_data_bf1[35]), .Y(exu_n31557));
AND2X1 exu_U1500(.A(exu_n3676), .B(exu_n8693), .Y(alu_zcomp_in[37]));
OR2X1 exu_U1501(.A(alu_addsub_rs2_data[33]), .B(alu_logic_rs1_data_bf1[33]), .Y(exu_n31561));
AND2X1 exu_U1502(.A(exu_n3678), .B(exu_n8695), .Y(alu_zcomp_in[35]));
OR2X1 exu_U1503(.A(alu_ecl_adderin2_31_e), .B(alu_logic_rs1_data_bf1[31]), .Y(exu_n31565));
AND2X1 exu_U1504(.A(exu_n3680), .B(exu_n8697), .Y(alu_zcomp_in[33]));
AND2X1 exu_U1505(.A(exu_n3669), .B(exu_n8686), .Y(alu_zcomp_in[43]));
AND2X1 exu_U1506(.A(exu_n3670), .B(exu_n8687), .Y(alu_zcomp_in[42]));
AND2X1 exu_U1507(.A(exu_n3671), .B(exu_n8688), .Y(alu_zcomp_in[41]));
AND2X1 exu_U1508(.A(exu_n3672), .B(exu_n8689), .Y(alu_zcomp_in[40]));
AND2X1 exu_U1509(.A(exu_n3667), .B(exu_n8684), .Y(alu_zcomp_in[45]));
AND2X1 exu_U1510(.A(exu_n3668), .B(exu_n8685), .Y(alu_zcomp_in[44]));
AND2X1 exu_U1511(.A(exu_n3666), .B(exu_n8683), .Y(alu_zcomp_in[46]));
AND2X1 exu_U1512(.A(exu_n3652), .B(exu_n8669), .Y(alu_zcomp_in[59]));
AND2X1 exu_U1513(.A(exu_n3653), .B(exu_n8670), .Y(alu_zcomp_in[58]));
AND2X1 exu_U1514(.A(exu_n3654), .B(exu_n8671), .Y(alu_zcomp_in[57]));
AND2X1 exu_U1515(.A(exu_n3655), .B(exu_n8672), .Y(alu_zcomp_in[56]));
AND2X1 exu_U1516(.A(exu_n3649), .B(exu_n8666), .Y(alu_zcomp_in[61]));
AND2X1 exu_U1517(.A(exu_n3650), .B(exu_n8667), .Y(alu_zcomp_in[60]));
AND2X1 exu_U1518(.A(exu_n3648), .B(exu_n8665), .Y(alu_zcomp_in[62]));
AND2X1 exu_U1519(.A(exu_n3660), .B(exu_n8677), .Y(alu_zcomp_in[51]));
AND2X1 exu_U1520(.A(exu_n3661), .B(exu_n8678), .Y(alu_zcomp_in[50]));
AND2X1 exu_U1521(.A(exu_n3663), .B(exu_n8680), .Y(alu_zcomp_in[49]));
AND2X1 exu_U1522(.A(exu_n3664), .B(exu_n8681), .Y(alu_zcomp_in[48]));
AND2X1 exu_U1523(.A(exu_n3658), .B(exu_n8675), .Y(alu_zcomp_in[53]));
AND2X1 exu_U1524(.A(exu_n3659), .B(exu_n8676), .Y(alu_zcomp_in[52]));
AND2X1 exu_U1525(.A(exu_n3657), .B(exu_n8674), .Y(alu_zcomp_in[54]));
OR2X1 exu_U1526(.A(alu_addsub_rs2_data_14), .B(alu_logic_rs1_data_bf1[14]), .Y(exu_n31603));
AND2X1 exu_U1527(.A(exu_n3699), .B(exu_n8716), .Y(alu_zcomp_in[16]));
OR2X1 exu_U1528(.A(alu_addsub_rs2_data_12), .B(alu_logic_rs1_data_bf1[12]), .Y(exu_n31607));
AND2X1 exu_U1529(.A(exu_n3701), .B(exu_n8718), .Y(alu_zcomp_in[14]));
OR2X1 exu_U1530(.A(alu_addsub_rs2_data_10), .B(alu_logic_rs1_data_bf1[10]), .Y(exu_n31611));
AND2X1 exu_U1531(.A(exu_n3703), .B(exu_n8720), .Y(alu_zcomp_in[12]));
AND2X1 exu_U1532(.A(exu_n3705), .B(exu_n8722), .Y(alu_zcomp_in[10]));
AND2X1 exu_U1533(.A(exu_n3695), .B(exu_n8712), .Y(alu_zcomp_in[1]));
AND2X1 exu_U1534(.A(exu_n3696), .B(exu_n8713), .Y(alu_zcomp_in[19]));
AND2X1 exu_U1535(.A(exu_n3697), .B(exu_n8714), .Y(alu_zcomp_in[18]));
AND2X1 exu_U1536(.A(exu_n3698), .B(exu_n8715), .Y(alu_zcomp_in[17]));
AND2X1 exu_U1537(.A(exu_n3693), .B(exu_n8710), .Y(alu_zcomp_in[21]));
AND2X1 exu_U1538(.A(exu_n3694), .B(exu_n8711), .Y(alu_zcomp_in[20]));
AND2X1 exu_U1539(.A(exu_n3692), .B(exu_n8709), .Y(alu_zcomp_in[22]));
OR2X1 exu_U1540(.A(alu_addsub_rs2_data_1), .B(alu_logic_rs1_data_bf1[1]), .Y(exu_n31571));
AND2X1 exu_U1541(.A(exu_n3683), .B(exu_n8700), .Y(alu_zcomp_in[30]));
OR2X1 exu_U1542(.A(alu_addsub_rs2_data_27), .B(alu_logic_rs1_data_bf1[27]), .Y(exu_n31575));
AND2X1 exu_U1543(.A(exu_n3685), .B(exu_n8702), .Y(alu_zcomp_in[29]));
OR2X1 exu_U1544(.A(alu_addsub_rs2_data_25), .B(alu_logic_rs1_data_bf1[25]), .Y(exu_n31579));
AND2X1 exu_U1545(.A(exu_n3687), .B(exu_n8704), .Y(alu_zcomp_in[27]));
OR2X1 exu_U1546(.A(alu_addsub_rs2_data_23), .B(alu_logic_rs1_data_bf1[23]), .Y(exu_n31583));
AND2X1 exu_U1547(.A(exu_n3689), .B(exu_n8706), .Y(alu_zcomp_in[25]));
AND2X1 exu_U1548(.A(exu_n3651), .B(exu_n8668), .Y(alu_zcomp_in[5]));
AND2X1 exu_U1549(.A(exu_n3662), .B(exu_n8679), .Y(alu_zcomp_in[4]));
AND2X1 exu_U1550(.A(exu_n3673), .B(exu_n8690), .Y(alu_zcomp_in[3]));
AND2X1 exu_U1551(.A(exu_n3682), .B(exu_n8699), .Y(alu_zcomp_in[31]));
AND2X1 exu_U1552(.A(exu_n3645), .B(exu_n8662), .Y(alu_zcomp_in[7]));
AND2X1 exu_U1553(.A(exu_n3646), .B(exu_n8663), .Y(alu_zcomp_in[6]));
AND2X1 exu_U1554(.A(exu_n3644), .B(exu_n8661), .Y(alu_zcomp_in[8]));
INVX1 exu_U1555(.A(ecl_writeback_sraddr_w[1]), .Y(exu_n16554));
INVX1 exu_U1556(.A(ecl_tid_w1[0]), .Y(exu_n16575));
OR2X1 exu_U1557(.A(exu_n13108), .B(exu_n14394), .Y(shft_rshift1[63]));
AND2X1 exu_U1558(.A(exu_n2921), .B(exu_n8002), .Y(exu_n27399));
OR2X1 exu_U1559(.A(exu_n13239), .B(exu_n14546), .Y(shft_lshift1[63]));
AND2X1 exu_U1560(.A(exu_n147), .B(exu_n5114), .Y(exu_n17352));
OR2X1 exu_U1561(.A(exu_n13108), .B(exu_n14395), .Y(shft_rshift1[62]));
AND2X1 exu_U1562(.A(exu_n2922), .B(exu_n8003), .Y(exu_n27402));
OR2X1 exu_U1563(.A(exu_n13240), .B(exu_n14547), .Y(shft_lshift1[62]));
OR2X1 exu_U1564(.A(exu_n13333), .B(exu_n14640), .Y(alu_logic_out[62]));
AND2X1 exu_U1565(.A(exu_n3413), .B(exu_n8494), .Y(exu_n28947));
AND2X1 exu_U1566(.A(exu_n146), .B(exu_n5113), .Y(exu_n17347));
OR2X1 exu_U1567(.A(exu_n13109), .B(exu_n14396), .Y(shft_rshift1[61]));
OR2X1 exu_U1568(.A(exu_n13241), .B(exu_n14548), .Y(shft_lshift1[61]));
OR2X1 exu_U1569(.A(exu_n13334), .B(exu_n14641), .Y(alu_logic_out[61]));
AND2X1 exu_U1570(.A(exu_n3415), .B(exu_n8496), .Y(exu_n28953));
AND2X1 exu_U1571(.A(exu_n145), .B(exu_n5112), .Y(exu_n17340));
OR2X1 exu_U1572(.A(exu_n13110), .B(exu_n14397), .Y(shft_rshift1[60]));
OR2X1 exu_U1573(.A(exu_n13242), .B(exu_n14549), .Y(shft_lshift1[60]));
OR2X1 exu_U1574(.A(exu_n13335), .B(exu_n14642), .Y(alu_logic_out[60]));
AND2X1 exu_U1575(.A(exu_n3417), .B(exu_n8498), .Y(exu_n28959));
AND2X1 exu_U1576(.A(exu_n144), .B(exu_n5111), .Y(exu_n17335));
OR2X1 exu_U1577(.A(exu_n13112), .B(exu_n14399), .Y(shft_rshift1[59]));
OR2X1 exu_U1578(.A(exu_n13244), .B(exu_n14551), .Y(shft_lshift1[59]));
OR2X1 exu_U1579(.A(exu_n13337), .B(exu_n14644), .Y(alu_logic_out[59]));
AND2X1 exu_U1580(.A(exu_n3421), .B(exu_n8502), .Y(exu_n28971));
AND2X1 exu_U1581(.A(exu_n143), .B(exu_n5110), .Y(exu_n17330));
OR2X1 exu_U1582(.A(exu_n13113), .B(exu_n14400), .Y(shft_rshift1[58]));
OR2X1 exu_U1583(.A(exu_n13245), .B(exu_n14552), .Y(shft_lshift1[58]));
OR2X1 exu_U1584(.A(exu_n13338), .B(exu_n14645), .Y(alu_logic_out[58]));
AND2X1 exu_U1585(.A(exu_n3423), .B(exu_n8504), .Y(exu_n28977));
AND2X1 exu_U1586(.A(exu_n142), .B(exu_n5109), .Y(exu_n17325));
OR2X1 exu_U1587(.A(exu_n13114), .B(exu_n14401), .Y(shft_rshift1[57]));
OR2X1 exu_U1588(.A(exu_n13246), .B(exu_n14553), .Y(shft_lshift1[57]));
OR2X1 exu_U1589(.A(exu_n13339), .B(exu_n14646), .Y(alu_logic_out[57]));
AND2X1 exu_U1590(.A(exu_n3425), .B(exu_n8506), .Y(exu_n28983));
AND2X1 exu_U1591(.A(exu_n141), .B(exu_n5108), .Y(exu_n17320));
OR2X1 exu_U1592(.A(exu_n13115), .B(exu_n14402), .Y(shft_rshift1[56]));
OR2X1 exu_U1593(.A(exu_n13247), .B(exu_n14554), .Y(shft_lshift1[56]));
OR2X1 exu_U1594(.A(exu_n13340), .B(exu_n14647), .Y(alu_logic_out[56]));
AND2X1 exu_U1595(.A(exu_n3427), .B(exu_n8508), .Y(exu_n28989));
AND2X1 exu_U1596(.A(exu_n140), .B(exu_n5107), .Y(exu_n17315));
OR2X1 exu_U1597(.A(exu_n13116), .B(exu_n14403), .Y(shft_rshift1[55]));
OR2X1 exu_U1598(.A(exu_n13248), .B(exu_n14555), .Y(shft_lshift1[55]));
OR2X1 exu_U1599(.A(exu_n13341), .B(exu_n14648), .Y(alu_logic_out[55]));
AND2X1 exu_U1600(.A(exu_n3429), .B(exu_n8510), .Y(exu_n28995));
AND2X1 exu_U1601(.A(exu_n139), .B(exu_n5106), .Y(exu_n17310));
OR2X1 exu_U1602(.A(exu_n13117), .B(exu_n14404), .Y(shft_rshift1[54]));
OR2X1 exu_U1603(.A(exu_n13249), .B(exu_n14556), .Y(shft_lshift1[54]));
OR2X1 exu_U1604(.A(exu_n13342), .B(exu_n14649), .Y(alu_logic_out[54]));
AND2X1 exu_U1605(.A(exu_n3431), .B(exu_n8512), .Y(exu_n29001));
AND2X1 exu_U1606(.A(exu_n138), .B(exu_n5105), .Y(exu_n17305));
OR2X1 exu_U1607(.A(exu_n13118), .B(exu_n14405), .Y(shft_rshift1[53]));
OR2X1 exu_U1608(.A(exu_n13250), .B(exu_n14557), .Y(shft_lshift1[53]));
OR2X1 exu_U1609(.A(exu_n13343), .B(exu_n14650), .Y(alu_logic_out[53]));
AND2X1 exu_U1610(.A(exu_n3433), .B(exu_n8514), .Y(exu_n29007));
AND2X1 exu_U1611(.A(exu_n137), .B(exu_n5104), .Y(exu_n17300));
OR2X1 exu_U1612(.A(exu_n13119), .B(exu_n14406), .Y(shft_rshift1[52]));
OR2X1 exu_U1613(.A(exu_n13251), .B(exu_n14558), .Y(shft_lshift1[52]));
OR2X1 exu_U1614(.A(exu_n13344), .B(exu_n14651), .Y(alu_logic_out[52]));
AND2X1 exu_U1615(.A(exu_n3435), .B(exu_n8516), .Y(exu_n29013));
AND2X1 exu_U1616(.A(exu_n136), .B(exu_n5103), .Y(exu_n17295));
OR2X1 exu_U1617(.A(exu_n13120), .B(exu_n14407), .Y(shft_rshift1[51]));
OR2X1 exu_U1618(.A(exu_n13252), .B(exu_n14559), .Y(shft_lshift1[51]));
OR2X1 exu_U1619(.A(exu_n13345), .B(exu_n14652), .Y(alu_logic_out[51]));
AND2X1 exu_U1620(.A(exu_n3437), .B(exu_n8518), .Y(exu_n29019));
AND2X1 exu_U1621(.A(exu_n135), .B(exu_n5102), .Y(exu_n17288));
OR2X1 exu_U1622(.A(exu_n13121), .B(exu_n14408), .Y(shft_rshift1[50]));
OR2X1 exu_U1623(.A(exu_n13253), .B(exu_n14560), .Y(shft_lshift1[50]));
OR2X1 exu_U1624(.A(exu_n13346), .B(exu_n14653), .Y(alu_logic_out[50]));
AND2X1 exu_U1625(.A(exu_n3439), .B(exu_n8520), .Y(exu_n29025));
AND2X1 exu_U1626(.A(exu_n134), .B(exu_n5101), .Y(exu_n17283));
OR2X1 exu_U1627(.A(exu_n13123), .B(exu_n14410), .Y(shft_rshift1[49]));
OR2X1 exu_U1628(.A(exu_n13255), .B(exu_n14562), .Y(shft_lshift1[49]));
OR2X1 exu_U1629(.A(exu_n13348), .B(exu_n14655), .Y(alu_logic_out[49]));
AND2X1 exu_U1630(.A(exu_n3443), .B(exu_n8524), .Y(exu_n29037));
AND2X1 exu_U1631(.A(exu_n133), .B(exu_n5100), .Y(exu_n17278));
OR2X1 exu_U1632(.A(exu_n13124), .B(exu_n14411), .Y(shft_rshift1[48]));
OR2X1 exu_U1633(.A(exu_n13256), .B(exu_n14563), .Y(shft_lshift1[48]));
OR2X1 exu_U1634(.A(exu_n13349), .B(exu_n14656), .Y(alu_logic_out[48]));
AND2X1 exu_U1635(.A(exu_n3445), .B(exu_n8526), .Y(exu_n29043));
OR2X1 exu_U1636(.A(exu_n13125), .B(exu_n14412), .Y(shft_rshift1[47]));
OR2X1 exu_U1637(.A(exu_n13257), .B(exu_n14564), .Y(shft_lshift1[47]));
OR2X1 exu_U1638(.A(exu_n13350), .B(exu_n14657), .Y(alu_logic_out[47]));
AND2X1 exu_U1639(.A(exu_n3447), .B(exu_n8528), .Y(exu_n29049));
OR2X1 exu_U1640(.A(exu_n13126), .B(exu_n14413), .Y(shft_rshift1[46]));
OR2X1 exu_U1641(.A(exu_n13258), .B(exu_n14565), .Y(shft_lshift1[46]));
OR2X1 exu_U1642(.A(exu_n13351), .B(exu_n14658), .Y(alu_logic_out[46]));
AND2X1 exu_U1643(.A(exu_n3449), .B(exu_n8530), .Y(exu_n29055));
OR2X1 exu_U1644(.A(exu_n13127), .B(exu_n14414), .Y(shft_rshift1[45]));
OR2X1 exu_U1645(.A(exu_n13259), .B(exu_n14566), .Y(shft_lshift1[45]));
OR2X1 exu_U1646(.A(exu_n13352), .B(exu_n14659), .Y(alu_logic_out[45]));
AND2X1 exu_U1647(.A(exu_n3451), .B(exu_n8532), .Y(exu_n29061));
OR2X1 exu_U1648(.A(exu_n13128), .B(exu_n14415), .Y(shft_rshift1[44]));
OR2X1 exu_U1649(.A(exu_n13260), .B(exu_n14567), .Y(shft_lshift1[44]));
OR2X1 exu_U1650(.A(exu_n13353), .B(exu_n14660), .Y(alu_logic_out[44]));
AND2X1 exu_U1651(.A(exu_n3453), .B(exu_n8534), .Y(exu_n29067));
OR2X1 exu_U1652(.A(exu_n13129), .B(exu_n14416), .Y(shft_rshift1[43]));
OR2X1 exu_U1653(.A(exu_n13261), .B(exu_n14568), .Y(shft_lshift1[43]));
OR2X1 exu_U1654(.A(exu_n13354), .B(exu_n14661), .Y(alu_logic_out[43]));
AND2X1 exu_U1655(.A(exu_n3455), .B(exu_n8536), .Y(exu_n29073));
OR2X1 exu_U1656(.A(exu_n13130), .B(exu_n14417), .Y(shft_rshift1[42]));
OR2X1 exu_U1657(.A(exu_n13262), .B(exu_n14569), .Y(shft_lshift1[42]));
OR2X1 exu_U1658(.A(exu_n13355), .B(exu_n14662), .Y(alu_logic_out[42]));
AND2X1 exu_U1659(.A(exu_n3457), .B(exu_n8538), .Y(exu_n29079));
OR2X1 exu_U1660(.A(exu_n13131), .B(exu_n14418), .Y(shft_rshift1[41]));
OR2X1 exu_U1661(.A(exu_n13263), .B(exu_n14570), .Y(shft_lshift1[41]));
OR2X1 exu_U1662(.A(exu_n13356), .B(exu_n14663), .Y(alu_logic_out[41]));
AND2X1 exu_U1663(.A(exu_n3459), .B(exu_n8540), .Y(exu_n29085));
OR2X1 exu_U1664(.A(exu_n13132), .B(exu_n14419), .Y(shft_rshift1[40]));
OR2X1 exu_U1665(.A(exu_n13264), .B(exu_n14571), .Y(shft_lshift1[40]));
OR2X1 exu_U1666(.A(exu_n13357), .B(exu_n14664), .Y(alu_logic_out[40]));
AND2X1 exu_U1667(.A(exu_n3461), .B(exu_n8542), .Y(exu_n29091));
OR2X1 exu_U1668(.A(exu_n13134), .B(exu_n14421), .Y(shft_rshift1[39]));
OR2X1 exu_U1669(.A(exu_n13266), .B(exu_n14573), .Y(shft_lshift1[39]));
OR2X1 exu_U1670(.A(exu_n13359), .B(exu_n14666), .Y(alu_logic_out[39]));
AND2X1 exu_U1671(.A(exu_n3465), .B(exu_n8546), .Y(exu_n29103));
OR2X1 exu_U1672(.A(exu_n13135), .B(exu_n14422), .Y(shft_rshift1[38]));
OR2X1 exu_U1673(.A(exu_n13267), .B(exu_n14574), .Y(shft_lshift1[38]));
OR2X1 exu_U1674(.A(exu_n13360), .B(exu_n14667), .Y(alu_logic_out[38]));
AND2X1 exu_U1675(.A(exu_n3467), .B(exu_n8548), .Y(exu_n29109));
OR2X1 exu_U1676(.A(exu_n13136), .B(exu_n14423), .Y(shft_rshift1[37]));
OR2X1 exu_U1677(.A(exu_n13268), .B(exu_n14575), .Y(shft_lshift1[37]));
OR2X1 exu_U1678(.A(exu_n13361), .B(exu_n14668), .Y(alu_logic_out[37]));
AND2X1 exu_U1679(.A(exu_n3469), .B(exu_n8550), .Y(exu_n29115));
OR2X1 exu_U1680(.A(exu_n13137), .B(exu_n14424), .Y(shft_rshift1[36]));
OR2X1 exu_U1681(.A(exu_n13269), .B(exu_n14576), .Y(shft_lshift1[36]));
OR2X1 exu_U1682(.A(exu_n13362), .B(exu_n14669), .Y(alu_logic_out[36]));
AND2X1 exu_U1683(.A(exu_n3471), .B(exu_n8552), .Y(exu_n29121));
OR2X1 exu_U1684(.A(exu_n13138), .B(exu_n14425), .Y(shft_rshift1[35]));
OR2X1 exu_U1685(.A(exu_n13270), .B(exu_n14577), .Y(shft_lshift1[35]));
OR2X1 exu_U1686(.A(exu_n13363), .B(exu_n14670), .Y(alu_logic_out[35]));
AND2X1 exu_U1687(.A(exu_n3473), .B(exu_n8554), .Y(exu_n29127));
OR2X1 exu_U1688(.A(exu_n13139), .B(exu_n14426), .Y(shft_rshift1[34]));
OR2X1 exu_U1689(.A(exu_n13271), .B(exu_n14578), .Y(shft_lshift1[34]));
OR2X1 exu_U1690(.A(exu_n13364), .B(exu_n14671), .Y(alu_logic_out[34]));
AND2X1 exu_U1691(.A(exu_n3475), .B(exu_n8556), .Y(exu_n29133));
OR2X1 exu_U1692(.A(exu_n13140), .B(exu_n14427), .Y(shft_rshift1[33]));
OR2X1 exu_U1693(.A(exu_n13272), .B(exu_n14579), .Y(shft_lshift1[33]));
OR2X1 exu_U1694(.A(exu_n13365), .B(exu_n14672), .Y(alu_logic_out[33]));
AND2X1 exu_U1695(.A(exu_n3477), .B(exu_n8558), .Y(exu_n29139));
OR2X1 exu_U1696(.A(exu_n13141), .B(exu_n14428), .Y(shft_rshift1[32]));
OR2X1 exu_U1697(.A(exu_n13273), .B(exu_n14580), .Y(shft_lshift1[32]));
OR2X1 exu_U1698(.A(exu_n13366), .B(exu_n14673), .Y(alu_logic_out[32]));
AND2X1 exu_U1699(.A(exu_n3479), .B(exu_n8560), .Y(exu_n29145));
OR2X1 exu_U1700(.A(exu_n13142), .B(exu_n14429), .Y(shft_rshift1[31]));
OR2X1 exu_U1701(.A(exu_n13274), .B(exu_n14581), .Y(shft_lshift1[31]));
OR2X1 exu_U1702(.A(exu_n13143), .B(exu_n14430), .Y(shft_rshift1[30]));
OR2X1 exu_U1703(.A(exu_n13275), .B(exu_n14582), .Y(shft_lshift1[30]));
OR2X1 exu_U1704(.A(exu_n13368), .B(exu_n14675), .Y(alu_logic_out_30));
AND2X1 exu_U1705(.A(exu_n3483), .B(exu_n8564), .Y(exu_n29157));
OR2X1 exu_U1706(.A(exu_n13145), .B(exu_n14432), .Y(shft_rshift1[29]));
OR2X1 exu_U1707(.A(exu_n13276), .B(exu_n14584), .Y(shft_lshift1[29]));
OR2X1 exu_U1708(.A(exu_n13370), .B(exu_n14677), .Y(alu_logic_out_29));
AND2X1 exu_U1709(.A(exu_n3487), .B(exu_n8568), .Y(exu_n29169));
OR2X1 exu_U1710(.A(exu_n13146), .B(exu_n14433), .Y(shft_rshift1[28]));
OR2X1 exu_U1711(.A(exu_n13277), .B(exu_n14585), .Y(shft_lshift1[28]));
OR2X1 exu_U1712(.A(exu_n13371), .B(exu_n14678), .Y(alu_logic_out_28));
AND2X1 exu_U1713(.A(exu_n3489), .B(exu_n8570), .Y(exu_n29175));
OR2X1 exu_U1714(.A(exu_n13147), .B(exu_n14434), .Y(shft_rshift1[27]));
OR2X1 exu_U1715(.A(exu_n13278), .B(exu_n14586), .Y(shft_lshift1[27]));
OR2X1 exu_U1716(.A(exu_n13372), .B(exu_n14679), .Y(alu_logic_out_27));
AND2X1 exu_U1717(.A(exu_n3491), .B(exu_n8572), .Y(exu_n29181));
OR2X1 exu_U1718(.A(exu_n13148), .B(exu_n14435), .Y(shft_rshift1[26]));
OR2X1 exu_U1719(.A(exu_n13279), .B(exu_n14587), .Y(shft_lshift1[26]));
OR2X1 exu_U1720(.A(exu_n13373), .B(exu_n14680), .Y(alu_logic_out_26));
AND2X1 exu_U1721(.A(exu_n3493), .B(exu_n8574), .Y(exu_n29187));
OR2X1 exu_U1722(.A(exu_n13149), .B(exu_n14436), .Y(shft_rshift1[25]));
OR2X1 exu_U1723(.A(exu_n13280), .B(exu_n14588), .Y(shft_lshift1[25]));
OR2X1 exu_U1724(.A(exu_n13374), .B(exu_n14681), .Y(alu_logic_out_25));
AND2X1 exu_U1725(.A(exu_n3495), .B(exu_n8576), .Y(exu_n29193));
OR2X1 exu_U1726(.A(exu_n13150), .B(exu_n14437), .Y(shft_rshift1[24]));
OR2X1 exu_U1727(.A(exu_n13281), .B(exu_n14589), .Y(shft_lshift1[24]));
OR2X1 exu_U1728(.A(exu_n13375), .B(exu_n14682), .Y(alu_logic_out_24));
AND2X1 exu_U1729(.A(exu_n3497), .B(exu_n8578), .Y(exu_n29199));
OR2X1 exu_U1730(.A(exu_n13151), .B(exu_n14438), .Y(shft_rshift1[23]));
OR2X1 exu_U1731(.A(exu_n13282), .B(exu_n14590), .Y(shft_lshift1[23]));
OR2X1 exu_U1732(.A(exu_n13376), .B(exu_n14683), .Y(alu_logic_out_23));
AND2X1 exu_U1733(.A(exu_n3499), .B(exu_n8580), .Y(exu_n29205));
OR2X1 exu_U1734(.A(exu_n13152), .B(exu_n14439), .Y(shft_rshift1[22]));
OR2X1 exu_U1735(.A(exu_n13283), .B(exu_n14591), .Y(shft_lshift1[22]));
OR2X1 exu_U1736(.A(exu_n13377), .B(exu_n14684), .Y(alu_logic_out_22));
AND2X1 exu_U1737(.A(exu_n3501), .B(exu_n8582), .Y(exu_n29211));
OR2X1 exu_U1738(.A(exu_n13153), .B(exu_n14440), .Y(shft_rshift1[21]));
OR2X1 exu_U1739(.A(exu_n13284), .B(exu_n14592), .Y(shft_lshift1[21]));
OR2X1 exu_U1740(.A(exu_n13378), .B(exu_n14685), .Y(alu_logic_out_21));
AND2X1 exu_U1741(.A(exu_n3503), .B(exu_n8584), .Y(exu_n29217));
OR2X1 exu_U1742(.A(exu_n13154), .B(exu_n14441), .Y(shft_rshift1[20]));
OR2X1 exu_U1743(.A(exu_n13285), .B(exu_n14593), .Y(shft_lshift1[20]));
OR2X1 exu_U1744(.A(exu_n13379), .B(exu_n14686), .Y(alu_logic_out_20));
AND2X1 exu_U1745(.A(exu_n3505), .B(exu_n8586), .Y(exu_n29223));
OR2X1 exu_U1746(.A(exu_n13156), .B(exu_n14443), .Y(shft_rshift1[19]));
OR2X1 exu_U1747(.A(exu_n13286), .B(exu_n14594), .Y(shft_lshift1[19]));
OR2X1 exu_U1748(.A(exu_n13381), .B(exu_n14688), .Y(alu_logic_out_19));
AND2X1 exu_U1749(.A(exu_n3509), .B(exu_n8590), .Y(exu_n29235));
OR2X1 exu_U1750(.A(exu_n13157), .B(exu_n14444), .Y(shft_rshift1[18]));
OR2X1 exu_U1751(.A(exu_n13287), .B(exu_n14595), .Y(shft_lshift1[18]));
OR2X1 exu_U1752(.A(exu_n13382), .B(exu_n14689), .Y(alu_logic_out_18));
AND2X1 exu_U1753(.A(exu_n3511), .B(exu_n8592), .Y(exu_n29241));
OR2X1 exu_U1754(.A(exu_n13158), .B(exu_n14445), .Y(shft_rshift1[17]));
OR2X1 exu_U1755(.A(exu_n13288), .B(exu_n14596), .Y(shft_lshift1[17]));
OR2X1 exu_U1756(.A(exu_n13383), .B(exu_n14690), .Y(alu_logic_out_17));
AND2X1 exu_U1757(.A(exu_n3513), .B(exu_n8594), .Y(exu_n29247));
OR2X1 exu_U1758(.A(exu_n13159), .B(exu_n14446), .Y(shft_rshift1[16]));
OR2X1 exu_U1759(.A(exu_n13289), .B(exu_n14597), .Y(shft_lshift1[16]));
OR2X1 exu_U1760(.A(exu_n13384), .B(exu_n14691), .Y(alu_logic_out_16));
AND2X1 exu_U1761(.A(exu_n3515), .B(exu_n8596), .Y(exu_n29253));
OR2X1 exu_U1762(.A(exu_n13160), .B(exu_n14447), .Y(shft_rshift1[15]));
OR2X1 exu_U1763(.A(exu_n13290), .B(exu_n14598), .Y(shft_lshift1[15]));
OR2X1 exu_U1764(.A(exu_n13385), .B(exu_n14692), .Y(alu_logic_out_15));
AND2X1 exu_U1765(.A(exu_n3517), .B(exu_n8598), .Y(exu_n29259));
OR2X1 exu_U1766(.A(exu_n13161), .B(exu_n14448), .Y(shft_rshift1[14]));
OR2X1 exu_U1767(.A(exu_n13291), .B(exu_n14599), .Y(shft_lshift1[14]));
OR2X1 exu_U1768(.A(exu_n13386), .B(exu_n14693), .Y(alu_logic_out_14));
AND2X1 exu_U1769(.A(exu_n3519), .B(exu_n8600), .Y(exu_n29265));
OR2X1 exu_U1770(.A(exu_n13162), .B(exu_n14449), .Y(shft_rshift1[13]));
OR2X1 exu_U1771(.A(exu_n13292), .B(exu_n14600), .Y(shft_lshift1[13]));
OR2X1 exu_U1772(.A(exu_n13387), .B(exu_n14694), .Y(alu_logic_out_13));
AND2X1 exu_U1773(.A(exu_n3521), .B(exu_n8602), .Y(exu_n29271));
OR2X1 exu_U1774(.A(exu_n13163), .B(exu_n14450), .Y(shft_rshift1[12]));
OR2X1 exu_U1775(.A(exu_n13293), .B(exu_n14601), .Y(shft_lshift1[12]));
OR2X1 exu_U1776(.A(exu_n13388), .B(exu_n14695), .Y(alu_logic_out_12));
AND2X1 exu_U1777(.A(exu_n3523), .B(exu_n8604), .Y(exu_n29277));
OR2X1 exu_U1778(.A(exu_n13164), .B(exu_n14451), .Y(shft_rshift1[11]));
OR2X1 exu_U1779(.A(exu_n13294), .B(exu_n14602), .Y(shft_lshift1[11]));
OR2X1 exu_U1780(.A(exu_n13389), .B(exu_n14696), .Y(alu_logic_out_11));
AND2X1 exu_U1781(.A(exu_n3525), .B(exu_n8606), .Y(exu_n29283));
OR2X1 exu_U1782(.A(exu_n13165), .B(exu_n14452), .Y(shft_rshift1[10]));
OR2X1 exu_U1783(.A(exu_n13295), .B(exu_n14603), .Y(shft_lshift1[10]));
OR2X1 exu_U1784(.A(exu_n13390), .B(exu_n14697), .Y(alu_logic_out_10));
AND2X1 exu_U1785(.A(exu_n3527), .B(exu_n8608), .Y(exu_n29289));
OR2X1 exu_U1786(.A(exu_n13105), .B(exu_n14391), .Y(shft_rshift1[8]));
OR2X1 exu_U1787(.A(exu_n13236), .B(exu_n14543), .Y(shft_lshift1[8]));
OR2X1 exu_U1788(.A(exu_n13329), .B(exu_n14636), .Y(alu_logic_out_8));
AND2X1 exu_U1789(.A(exu_n3405), .B(exu_n8486), .Y(exu_n28923));
OR2X1 exu_U1790(.A(exu_n13106), .B(exu_n14392), .Y(shft_rshift1[7]));
OR2X1 exu_U1791(.A(exu_n13237), .B(exu_n14544), .Y(shft_lshift1[7]));
OR2X1 exu_U1792(.A(exu_n13330), .B(exu_n14637), .Y(alu_logic_out_7));
AND2X1 exu_U1793(.A(exu_n3407), .B(exu_n8488), .Y(exu_n28929));
OR2X1 exu_U1794(.A(exu_n13107), .B(exu_n14393), .Y(shft_rshift1[6]));
OR2X1 exu_U1795(.A(exu_n13238), .B(exu_n14545), .Y(shft_lshift1[6]));
OR2X1 exu_U1796(.A(exu_n13331), .B(exu_n14638), .Y(alu_logic_out_6));
AND2X1 exu_U1797(.A(exu_n3409), .B(exu_n8490), .Y(exu_n28935));
OR2X1 exu_U1798(.A(exu_n13111), .B(exu_n14398), .Y(shft_rshift1[5]));
OR2X1 exu_U1799(.A(exu_n13243), .B(exu_n14550), .Y(shft_lshift1[5]));
OR2X1 exu_U1800(.A(exu_n13336), .B(exu_n14643), .Y(alu_logic_out_5));
AND2X1 exu_U1801(.A(exu_n3419), .B(exu_n8500), .Y(exu_n28965));
OR2X1 exu_U1802(.A(exu_n13122), .B(exu_n14409), .Y(shft_rshift1[4]));
OR2X1 exu_U1803(.A(exu_n13254), .B(exu_n14561), .Y(shft_lshift1[4]));
OR2X1 exu_U1804(.A(exu_n13347), .B(exu_n14654), .Y(alu_logic_out_4));
AND2X1 exu_U1805(.A(exu_n3441), .B(exu_n8522), .Y(exu_n29031));
OR2X1 exu_U1806(.A(exu_n13133), .B(exu_n14420), .Y(shft_rshift1[3]));
OR2X1 exu_U1807(.A(exu_n13265), .B(exu_n14572), .Y(shft_lshift1[3]));
OR2X1 exu_U1808(.A(exu_n13358), .B(exu_n14665), .Y(alu_logic_out_3));
AND2X1 exu_U1809(.A(exu_n3463), .B(exu_n8544), .Y(exu_n29097));
OR2X1 exu_U1810(.A(exu_n13144), .B(exu_n14431), .Y(shft_rshift1[2]));
OR2X1 exu_U1811(.A(exu_n28571), .B(exu_n14583), .Y(shft_lshift1[2]));
OR2X1 exu_U1812(.A(exu_n13369), .B(exu_n14676), .Y(alu_logic_out_2));
AND2X1 exu_U1813(.A(exu_n3485), .B(exu_n8566), .Y(exu_n29163));
OR2X1 exu_U1814(.A(exu_n13155), .B(exu_n14442), .Y(shft_rshift1[1]));
AND2X1 exu_U1815(.A(exu_n11058), .B(exu_n8399), .Y(exu_n28632));
OR2X1 exu_U1816(.A(exu_n13380), .B(exu_n14687), .Y(alu_logic_out_1));
AND2X1 exu_U1817(.A(exu_n3507), .B(exu_n8588), .Y(exu_n29229));
OR2X1 exu_U1818(.A(exu_n13166), .B(exu_n14453), .Y(shft_rshift1[0]));
OR2X1 exu_U1819(.A(exu_n13391), .B(exu_n14698), .Y(alu_logic_out_0));
AND2X1 exu_U1820(.A(exu_n3529), .B(exu_n8610), .Y(exu_n29295));
AND2X1 exu_U1821(.A(exu_n15199), .B(ecc_err_m[0]), .Y(ecc_decode_n20));
AND2X1 exu_U1822(.A(exu_n15199), .B(exu_n15689), .Y(ecc_decode_n19));
AND2X1 exu_U1823(.A(exu_n15200), .B(exu_n15459), .Y(ecc_decode_n48));
AND2X1 exu_U1824(.A(exu_n4586), .B(exu_n9373), .Y(ecc_syn_mux_n25));
INVX1 exu_U1825(.A(ecl_ialign_m), .Y(exu_n16615));
AND2X1 exu_U1826(.A(exu_n15200), .B(ecc_err_m[4]), .Y(ecc_decode_n34));
AND2X1 exu_U1827(.A(exu_n4583), .B(exu_n9367), .Y(ecc_syn_mux_n13));
OR2X1 exu_U1828(.A(exu_n13440), .B(exu_n14759), .Y(ecl_byplog_rs1_n32));
AND2X1 exu_U1829(.A(exu_n13), .B(ecl_byplog_rs1_n17), .Y(ecl_byplog_rs1_n47));
AND2X1 exu_U1830(.A(exu_n17), .B(exu_n4986), .Y(exu_n16706));
AND2X1 exu_U1831(.A(exu_n218), .B(exu_n5143), .Y(ecl_byplog_rs2_match_w2));
AND2X1 exu_U1832(.A(ecl_ld_thr_match_dg2), .B(exu_n4985), .Y(ecl_byplog_rs2_n41));
AND2X1 exu_U1833(.A(exu_n20), .B(exu_n4988), .Y(exu_n16734));
OR2X1 exu_U1834(.A(exu_n13436), .B(exu_n14759), .Y(ecl_byplog_rs2_n32));
AND2X1 exu_U1835(.A(exu_n19), .B(ecl_byplog_rs2_n15), .Y(ecl_byplog_rs2_n42));
AND2X1 exu_U1836(.A(exu_n15423), .B(exu_n15820), .Y(ecl_byplog_rs2_n33));
AND2X1 exu_U1837(.A(exu_n153), .B(exu_n5120), .Y(exu_n17426));
AND2X1 exu_U1838(.A(exu_n15421), .B(exu_n15818), .Y(exu_n19203));
AND2X1 exu_U1839(.A(ecl_byp_ldxa_g), .B(exu_n15207), .Y(ecl_byplog_rs1_n46));
AND2X1 exu_U1840(.A(exu_n216), .B(exu_n5141), .Y(ecl_byplog_rs1_match_w2));
AND2X1 exu_U1841(.A(ecl_ld_thr_match_dg2), .B(exu_n4980), .Y(ecl_byplog_rs1_n45));
AND2X1 exu_U1842(.A(ecl_byplog_rs1_n32), .B(ecl_byplog_rs1_n17), .Y(ecl_byplog_rs1_n35));
OR2X1 exu_U1843(.A(exu_n13328), .B(exu_n14635), .Y(alu_logic_out_9));
AND2X1 exu_U1844(.A(exu_n3403), .B(exu_n8484), .Y(exu_n28917));
AND2X1 exu_U1845(.A(exu_n17382), .B(ecl_ld_rd_g[0]), .Y(exu_n17384));
AND2X1 exu_U1846(.A(exu_n222), .B(exu_n5147), .Y(ecl_byplog_rs3h_match_w2));
AND2X1 exu_U1847(.A(ecl_ld_thr_match_dg2), .B(exu_n5117), .Y(exu_n19247));
AND2X1 exu_U1848(.A(ecl_byp_ldxa_g), .B(exu_n15209), .Y(exu_n19250));
AND2X1 exu_U1849(.A(exu_n15422), .B(exu_n15819), .Y(exu_n19239));
OR2X1 exu_U1850(.A(exu_n12144), .B(exu_n14759), .Y(exu_n19238));
AND2X1 exu_U1851(.A(exu_n150), .B(exu_n19222), .Y(exu_n19248));
INVX1 exu_U1852(.A(ecl_ccr_setcc_w), .Y(exu_n16601));
AND2X1 exu_U1853(.A(exu_n3987), .B(exu_n9003), .Y(exu_n31664));
AND2X1 exu_U1854(.A(exu_n3972), .B(exu_n8988), .Y(exu_n31620));
AND2X1 exu_U1855(.A(exu_n3975), .B(exu_n8990), .Y(exu_n31626));
AND2X1 exu_U1856(.A(exu_n3977), .B(exu_n8993), .Y(exu_n31634));
AND2X1 exu_U1857(.A(exu_n3980), .B(exu_n8995), .Y(exu_n31640));
AND2X1 exu_U1858(.A(exu_n3982), .B(exu_n8998), .Y(exu_n31650));
AND2X1 exu_U1859(.A(exu_n3985), .B(exu_n9000), .Y(exu_n31656));
OR2X1 exu_U1860(.A(ecl_part_early_flush_w), .B(ecl_tlu_priv_trap_w), .Y(ecl_rml_early_flush_w));
OR2X1 exu_U1861(.A(ecl_writeback_n131), .B(ecl_writeback_sraddr_w[1]), .Y(ecl_writeback_n133));
OR2X1 exu_U1862(.A(exu_n16555), .B(exu_n15361), .Y(ecl_writeback_n131));
AND2X1 exu_U1863(.A(exu_n3638), .B(exu_n8655), .Y(alu_va_e[51]));
AND2X1 exu_U1864(.A(exu_n3636), .B(exu_n8653), .Y(alu_va_e[53]));
AND2X1 exu_U1865(.A(exu_n3637), .B(exu_n8654), .Y(alu_va_e[52]));
AND2X1 exu_U1866(.A(exu_n3640), .B(exu_n8657), .Y(alu_va_e[49]));
AND2X1 exu_U1867(.A(exu_n3639), .B(exu_n8656), .Y(alu_va_e[50]));
AND2X1 exu_U1868(.A(exu_n3641), .B(exu_n8658), .Y(alu_va_e[48]));
AND2X1 exu_U1869(.A(exu_n3630), .B(exu_n8647), .Y(alu_va_e[59]));
AND2X1 exu_U1870(.A(exu_n3628), .B(exu_n8645), .Y(alu_va_e[61]));
AND2X1 exu_U1871(.A(exu_n3627), .B(exu_n8644), .Y(alu_va_e[62]));
AND2X1 exu_U1872(.A(exu_n3629), .B(exu_n8646), .Y(alu_va_e[60]));
AND2X1 exu_U1873(.A(exu_n3635), .B(exu_n8652), .Y(alu_va_e[54]));
AND2X1 exu_U1874(.A(exu_n3634), .B(exu_n8651), .Y(alu_va_e[55]));
AND2X1 exu_U1875(.A(exu_n3632), .B(exu_n8649), .Y(alu_va_e[57]));
AND2X1 exu_U1876(.A(exu_n3631), .B(exu_n8648), .Y(alu_va_e[58]));
AND2X1 exu_U1877(.A(exu_n3633), .B(exu_n8650), .Y(alu_va_e[56]));
AND2X1 exu_U1878(.A(ecl_n93), .B(exu_n9665), .Y(ecl_n92));
AND2X1 exu_U1879(.A(ecl_thr_match_mw1), .B(ecl_inst_vld_w1), .Y(ecl_n98));
INVX1 exu_U1880(.A(rml_rml_ecl_cansave_e[1]), .Y(exu_n16590));
OR2X1 exu_U1881(.A(exu_n12086), .B(exu_n13502), .Y(ecl_byplog_rs1_N2));
AND2X1 exu_U1882(.A(ecl_byp_ldxa_g), .B(exu_n15208), .Y(ecl_byplog_rs2_n46));
AND2X1 exu_U1883(.A(ecl_byp_ldxa_g), .B(exu_n15210), .Y(exu_n19214));
OR2X1 exu_U1884(.A(exu_n12141), .B(exu_n14759), .Y(exu_n19202));
AND2X1 exu_U1885(.A(exu_n155), .B(exu_n19186), .Y(exu_n19212));
AND2X1 exu_U1886(.A(exu_n4550), .B(exu_n16599), .Y(ecl_bypass_w));
INVX1 exu_U1887(.A(ecl_writeback_inst_vld_noflush_wen_w), .Y(exu_n16599));
AND2X1 exu_U1888(.A(exu_n220), .B(exu_n5145), .Y(ecl_byplog_rs3_match_w2));
AND2X1 exu_U1889(.A(ecl_ld_thr_match_dg2), .B(exu_n5119), .Y(exu_n19211));
AND2X1 exu_U1890(.A(exu_n4968), .B(exu_n9672), .Y(ecl_n69));
AND2X1 exu_U1891(.A(exu_n4967), .B(exu_n16400), .Y(ecl_n68));
AND2X1 exu_U1892(.A(exu_n4917), .B(exu_n9631), .Y(div_n72));
AND2X1 exu_U1893(.A(exu_n4920), .B(exu_n9633), .Y(div_n78));
AND2X1 exu_U1894(.A(exu_n4922), .B(exu_n9636), .Y(div_n86));
AND2X1 exu_U1895(.A(exu_n4925), .B(exu_n9638), .Y(div_n92));
AND2X1 exu_U1896(.A(exu_n4909), .B(exu_n9620), .Y(div_n38));
OR2X1 exu_U1897(.A(exu_n15361), .B(exu_n14767), .Y(ecl_writeback_n142));
AND2X1 exu_U1898(.A(exu_n3742), .B(exu_n8821), .Y(div_gencc_in[35]));
AND2X1 exu_U1899(.A(exu_n3743), .B(exu_n8822), .Y(div_gencc_in[34]));
AND2X1 exu_U1900(.A(exu_n3740), .B(exu_n8819), .Y(div_gencc_in[37]));
AND2X1 exu_U1901(.A(exu_n3741), .B(exu_n8820), .Y(div_gencc_in[36]));
AND2X1 exu_U1902(.A(exu_n3738), .B(exu_n8817), .Y(div_gencc_in[39]));
AND2X1 exu_U1903(.A(exu_n3739), .B(exu_n8818), .Y(div_gencc_in[38]));
AND2X1 exu_U1904(.A(exu_n3736), .B(exu_n8815), .Y(div_gencc_in[40]));
AND2X1 exu_U1905(.A(exu_n3717), .B(exu_n8796), .Y(div_gencc_in[58]));
AND2X1 exu_U1906(.A(exu_n3716), .B(exu_n8795), .Y(div_gencc_in[59]));
AND2X1 exu_U1907(.A(exu_n3745), .B(exu_n8824), .Y(div_gencc_in[32]));
AND2X1 exu_U1908(.A(exu_n3714), .B(exu_n8793), .Y(div_gencc_in[60]));
AND2X1 exu_U1909(.A(exu_n3744), .B(exu_n8823), .Y(div_gencc_in[33]));
AND2X1 exu_U1910(.A(exu_n3713), .B(exu_n8792), .Y(div_gencc_in[61]));
AND2X1 exu_U1911(.A(exu_n3732), .B(exu_n8811), .Y(div_gencc_in[44]));
AND2X1 exu_U1912(.A(exu_n3712), .B(exu_n8791), .Y(div_gencc_in[62]));
AND2X1 exu_U1913(.A(exu_n3731), .B(exu_n8810), .Y(div_gencc_in[45]));
AND2X1 exu_U1914(.A(exu_n3730), .B(exu_n8809), .Y(div_gencc_in[46]));
AND2X1 exu_U1915(.A(exu_n3729), .B(exu_n8808), .Y(div_gencc_in[47]));
AND2X1 exu_U1916(.A(exu_n3721), .B(exu_n8800), .Y(div_gencc_in[54]));
AND2X1 exu_U1917(.A(exu_n3724), .B(exu_n8803), .Y(div_gencc_in[51]));
AND2X1 exu_U1918(.A(exu_n3723), .B(exu_n8802), .Y(div_gencc_in[52]));
AND2X1 exu_U1919(.A(exu_n3722), .B(exu_n8801), .Y(div_gencc_in[53]));
AND2X1 exu_U1920(.A(exu_n3763), .B(exu_n8842), .Y(div_gencc_in_16));
AND2X1 exu_U1921(.A(exu_n3765), .B(exu_n8844), .Y(div_gencc_in_14));
AND2X1 exu_U1922(.A(exu_n3767), .B(exu_n8846), .Y(div_gencc_in_12));
AND2X1 exu_U1923(.A(exu_n3769), .B(exu_n8848), .Y(div_gencc_in_10));
AND2X1 exu_U1924(.A(exu_n3759), .B(exu_n8838), .Y(div_gencc_in_1));
AND2X1 exu_U1925(.A(exu_n3760), .B(exu_n8839), .Y(div_gencc_in_19));
AND2X1 exu_U1926(.A(exu_n3761), .B(exu_n8840), .Y(div_gencc_in_18));
AND2X1 exu_U1927(.A(exu_n3762), .B(exu_n8841), .Y(div_gencc_in_17));
AND2X1 exu_U1928(.A(exu_n3757), .B(exu_n8836), .Y(div_gencc_in_21));
AND2X1 exu_U1929(.A(exu_n3758), .B(exu_n8837), .Y(div_gencc_in_20));
AND2X1 exu_U1930(.A(exu_n3756), .B(exu_n8835), .Y(div_gencc_in_22));
AND2X1 exu_U1931(.A(exu_n3747), .B(exu_n8826), .Y(div_gencc_in_30));
AND2X1 exu_U1932(.A(exu_n3749), .B(exu_n8828), .Y(div_gencc_in_29));
AND2X1 exu_U1933(.A(exu_n3751), .B(exu_n8830), .Y(div_gencc_in_27));
AND2X1 exu_U1934(.A(exu_n3753), .B(exu_n8832), .Y(div_gencc_in_25));
AND2X1 exu_U1935(.A(exu_n3715), .B(exu_n8794), .Y(div_gencc_in_5));
AND2X1 exu_U1936(.A(exu_n3726), .B(exu_n8805), .Y(div_gencc_in_4));
AND2X1 exu_U1937(.A(exu_n3709), .B(exu_n8788), .Y(div_gencc_in_7));
AND2X1 exu_U1938(.A(exu_n3710), .B(exu_n8789), .Y(div_gencc_in_6));
AND2X1 exu_U1939(.A(exu_n3708), .B(exu_n8787), .Y(div_gencc_in_8));
AND2X1 exu_U1940(.A(alu_logic_rs1_data_bf1[63]), .B(alu_logic_n101), .Y(alu_logic_result_and[63]));
OR2X1 exu_U1941(.A(alu_logic_n101), .B(alu_logic_rs1_data_bf1[63]), .Y(alu_logic_result_or[63]));
AND2X1 exu_U1942(.A(exu_n3410), .B(exu_n8491), .Y(exu_n28942));
AND2X1 exu_U1943(.A(exu_n3675), .B(exu_n8692), .Y(alu_zcomp_in[38]));
AND2X1 exu_U1944(.A(exu_n3677), .B(exu_n8694), .Y(alu_zcomp_in[36]));
AND2X1 exu_U1945(.A(exu_n3679), .B(exu_n8696), .Y(alu_zcomp_in[34]));
AND2X1 exu_U1946(.A(exu_n3681), .B(exu_n8698), .Y(alu_zcomp_in[32]));
AND2X1 exu_U1947(.A(exu_n4938), .B(exu_n9653), .Y(alu_n103));
AND2X1 exu_U1948(.A(exu_n4943), .B(exu_n9658), .Y(alu_n117));
AND2X1 exu_U1949(.A(exu_n4946), .B(exu_n9660), .Y(alu_n123));
OR2X1 exu_U1950(.A(exu_n15681), .B(alu_logic_rs1_data_bf1[62]), .Y(exu_n17353));
AND2X1 exu_U1951(.A(alu_logic_rs1_data_bf1[31]), .B(alu_logic_n136), .Y(alu_logic_result_and[31]));
OR2X1 exu_U1952(.A(alu_logic_n136), .B(alu_logic_rs1_data_bf1[31]), .Y(alu_logic_result_or[31]));
AND2X1 exu_U1953(.A(exu_n3480), .B(exu_n8561), .Y(exu_n29152));
AND2X1 exu_U1954(.A(exu_n3700), .B(exu_n8717), .Y(alu_zcomp_in[15]));
AND2X1 exu_U1955(.A(exu_n3702), .B(exu_n8719), .Y(alu_zcomp_in[13]));
AND2X1 exu_U1956(.A(exu_n3704), .B(exu_n8721), .Y(alu_zcomp_in[11]));
AND2X1 exu_U1957(.A(exu_n3706), .B(exu_n8723), .Y(alu_zcomp_in[0]));
AND2X1 exu_U1958(.A(exu_n4928), .B(exu_n9642), .Y(alu_n73));
AND2X1 exu_U1959(.A(exu_n3684), .B(exu_n8701), .Y(alu_zcomp_in[2]));
AND2X1 exu_U1960(.A(exu_n3686), .B(exu_n8703), .Y(alu_zcomp_in[28]));
AND2X1 exu_U1961(.A(exu_n3688), .B(exu_n8705), .Y(alu_zcomp_in[26]));
AND2X1 exu_U1962(.A(exu_n3690), .B(exu_n8707), .Y(alu_zcomp_in[24]));
AND2X1 exu_U1963(.A(exu_n4933), .B(exu_n9647), .Y(alu_n87));
INVX1 exu_U1964(.A(exu_ifu_brpc_e[31]), .Y(exu_n16512));
AND2X1 exu_U1965(.A(exu_n4545), .B(ecl_writeback_n176), .Y(ecl_writeback_n86));
INVX1 exu_U1966(.A(ecl_mdqctl_wb_multhr_g[1]), .Y(exu_n16510));
OR2X1 exu_U1967(.A(exu_n16575), .B(ecl_tid_w1[1]), .Y(ecl_writeback_n181));
INVX1 exu_U1968(.A(ecl_mdqctl_wb_multhr_g[0]), .Y(exu_n16509));
OR2X1 exu_U1969(.A(exu_n15775), .B(exu_n14769), .Y(ecl_writeback_n78));
OR2X1 exu_U1970(.A(exu_n15775), .B(exu_n14768), .Y(ecl_writeback_n74));
AND2X1 exu_U1971(.A(exu_n11242), .B(exu_n8727), .Y(shft_alu_shift_out_e[63]));
AND2X1 exu_U1972(.A(exu_n11244), .B(exu_n8728), .Y(shft_alu_shift_out_e[62]));
AND2X1 exu_U1973(.A(exu_n11246), .B(exu_n8729), .Y(shft_alu_shift_out_e[61]));
AND2X1 exu_U1974(.A(exu_n11248), .B(exu_n8730), .Y(shft_alu_shift_out_e[60]));
AND2X1 exu_U1975(.A(exu_n11252), .B(exu_n8732), .Y(shft_alu_shift_out_e[59]));
AND2X1 exu_U1976(.A(exu_n11254), .B(exu_n8733), .Y(shft_alu_shift_out_e[58]));
AND2X1 exu_U1977(.A(exu_n11256), .B(exu_n8734), .Y(shft_alu_shift_out_e[57]));
AND2X1 exu_U1978(.A(exu_n11258), .B(exu_n8735), .Y(shft_alu_shift_out_e[56]));
AND2X1 exu_U1979(.A(exu_n11260), .B(exu_n8736), .Y(shft_alu_shift_out_e[55]));
AND2X1 exu_U1980(.A(exu_n11262), .B(exu_n8737), .Y(shft_alu_shift_out_e[54]));
AND2X1 exu_U1981(.A(exu_n11264), .B(exu_n8738), .Y(shft_alu_shift_out_e[53]));
AND2X1 exu_U1982(.A(exu_n11266), .B(exu_n8739), .Y(shft_alu_shift_out_e[52]));
AND2X1 exu_U1983(.A(exu_n11268), .B(exu_n8740), .Y(shft_alu_shift_out_e[51]));
AND2X1 exu_U1984(.A(exu_n11270), .B(exu_n8741), .Y(shft_alu_shift_out_e[50]));
AND2X1 exu_U1985(.A(exu_n11274), .B(exu_n8743), .Y(shft_alu_shift_out_e[49]));
AND2X1 exu_U1986(.A(exu_n11276), .B(exu_n8744), .Y(shft_alu_shift_out_e[48]));
AND2X1 exu_U1987(.A(exu_n11278), .B(exu_n8745), .Y(shft_alu_shift_out_e[47]));
AND2X1 exu_U1988(.A(exu_n11280), .B(exu_n8746), .Y(shft_alu_shift_out_e[46]));
AND2X1 exu_U1989(.A(exu_n11282), .B(exu_n8747), .Y(shft_alu_shift_out_e[45]));
AND2X1 exu_U1990(.A(exu_n11284), .B(exu_n8748), .Y(shft_alu_shift_out_e[44]));
AND2X1 exu_U1991(.A(exu_n11286), .B(exu_n8749), .Y(shft_alu_shift_out_e[43]));
AND2X1 exu_U1992(.A(exu_n11288), .B(exu_n8750), .Y(shft_alu_shift_out_e[42]));
AND2X1 exu_U1993(.A(exu_n11290), .B(exu_n8751), .Y(shft_alu_shift_out_e[41]));
AND2X1 exu_U1994(.A(exu_n11292), .B(exu_n8752), .Y(shft_alu_shift_out_e[40]));
AND2X1 exu_U1995(.A(exu_n11296), .B(exu_n8754), .Y(shft_alu_shift_out_e[39]));
AND2X1 exu_U1996(.A(exu_n11298), .B(exu_n8755), .Y(shft_alu_shift_out_e[38]));
AND2X1 exu_U1997(.A(exu_n11300), .B(exu_n8756), .Y(shft_alu_shift_out_e[37]));
AND2X1 exu_U1998(.A(exu_n11302), .B(exu_n8757), .Y(shft_alu_shift_out_e[36]));
AND2X1 exu_U1999(.A(exu_n11304), .B(exu_n8758), .Y(shft_alu_shift_out_e[35]));
AND2X1 exu_U2000(.A(exu_n11306), .B(exu_n8759), .Y(shft_alu_shift_out_e[34]));
AND2X1 exu_U2001(.A(exu_n11308), .B(exu_n8760), .Y(shft_alu_shift_out_e[33]));
AND2X1 exu_U2002(.A(exu_n11310), .B(exu_n8761), .Y(shft_alu_shift_out_e[32]));
AND2X1 exu_U2003(.A(exu_n11312), .B(exu_n8762), .Y(shft_alu_shift_out_e[31]));
AND2X1 exu_U2004(.A(exu_n11314), .B(exu_n8763), .Y(shft_alu_shift_out_e[30]));
AND2X1 exu_U2005(.A(exu_n11318), .B(exu_n8765), .Y(shft_alu_shift_out_e[29]));
AND2X1 exu_U2006(.A(exu_n11320), .B(exu_n8766), .Y(shft_alu_shift_out_e[28]));
AND2X1 exu_U2007(.A(exu_n11322), .B(exu_n8767), .Y(shft_alu_shift_out_e[27]));
AND2X1 exu_U2008(.A(exu_n11324), .B(exu_n8768), .Y(shft_alu_shift_out_e[26]));
AND2X1 exu_U2009(.A(exu_n11326), .B(exu_n8769), .Y(shft_alu_shift_out_e[25]));
AND2X1 exu_U2010(.A(exu_n11328), .B(exu_n8770), .Y(shft_alu_shift_out_e[24]));
AND2X1 exu_U2011(.A(exu_n11330), .B(exu_n8771), .Y(shft_alu_shift_out_e[23]));
AND2X1 exu_U2012(.A(exu_n11332), .B(exu_n8772), .Y(shft_alu_shift_out_e[22]));
AND2X1 exu_U2013(.A(exu_n11334), .B(exu_n8773), .Y(shft_alu_shift_out_e[21]));
AND2X1 exu_U2014(.A(exu_n11336), .B(exu_n8774), .Y(shft_alu_shift_out_e[20]));
AND2X1 exu_U2015(.A(exu_n11340), .B(exu_n8776), .Y(shft_alu_shift_out_e[19]));
AND2X1 exu_U2016(.A(exu_n11342), .B(exu_n8777), .Y(shft_alu_shift_out_e[18]));
AND2X1 exu_U2017(.A(exu_n11344), .B(exu_n8778), .Y(shft_alu_shift_out_e[17]));
AND2X1 exu_U2018(.A(exu_n11346), .B(exu_n8779), .Y(shft_alu_shift_out_e[16]));
AND2X1 exu_U2019(.A(exu_n11348), .B(exu_n8780), .Y(shft_alu_shift_out_e[15]));
AND2X1 exu_U2020(.A(exu_n11350), .B(exu_n8781), .Y(shft_alu_shift_out_e[14]));
AND2X1 exu_U2021(.A(exu_n11352), .B(exu_n8782), .Y(shft_alu_shift_out_e[13]));
AND2X1 exu_U2022(.A(exu_n11354), .B(exu_n8783), .Y(shft_alu_shift_out_e[12]));
AND2X1 exu_U2023(.A(exu_n11356), .B(exu_n8784), .Y(shft_alu_shift_out_e[11]));
AND2X1 exu_U2024(.A(exu_n11358), .B(exu_n8785), .Y(shft_alu_shift_out_e[10]));
INVX1 exu_U2025(.A(ecl_tid_e[1]), .Y(exu_n16580));
AND2X1 exu_U2026(.A(exu_n11236), .B(exu_n8724), .Y(shft_alu_shift_out_e[8]));
AND2X1 exu_U2027(.A(exu_n11238), .B(exu_n8725), .Y(shft_alu_shift_out_e[7]));
AND2X1 exu_U2028(.A(exu_n11240), .B(exu_n8726), .Y(shft_alu_shift_out_e[6]));
AND2X1 exu_U2029(.A(exu_n11250), .B(exu_n8731), .Y(shft_alu_shift_out_e[5]));
INVX1 exu_U2030(.A(exu_n16159), .Y(exu_n16158));
AND2X1 exu_U2031(.A(exu_n11272), .B(exu_n8742), .Y(shft_alu_shift_out_e[4]));
AND2X1 exu_U2032(.A(exu_n11294), .B(exu_n8753), .Y(shft_alu_shift_out_e[3]));
AND2X1 exu_U2033(.A(exu_n11316), .B(exu_n8764), .Y(shft_alu_shift_out_e[2]));
AND2X1 exu_U2034(.A(exu_n11338), .B(exu_n8775), .Y(shft_alu_shift_out_e[1]));
AND2X1 exu_U2035(.A(exu_n11360), .B(exu_n8786), .Y(shft_alu_shift_out_e[0]));
AND2X1 exu_U2036(.A(exu_n22833), .B(exu_n6387), .Y(ecc_ecc_datain_m[63]));
AND2X1 exu_U2037(.A(exu_n1493), .B(exu_n6388), .Y(exu_n22833));
AND2X1 exu_U2038(.A(exu_n22837), .B(exu_n6389), .Y(ecc_ecc_datain_m[62]));
AND2X1 exu_U2039(.A(exu_n1494), .B(exu_n6390), .Y(exu_n22837));
AND2X1 exu_U2040(.A(exu_n22841), .B(exu_n6391), .Y(ecc_ecc_datain_m[61]));
AND2X1 exu_U2041(.A(exu_n1495), .B(exu_n6392), .Y(exu_n22841));
AND2X1 exu_U2042(.A(exu_n22845), .B(exu_n6393), .Y(ecc_ecc_datain_m[60]));
AND2X1 exu_U2043(.A(exu_n1496), .B(exu_n6394), .Y(exu_n22845));
AND2X1 exu_U2044(.A(exu_n22853), .B(exu_n6397), .Y(ecc_ecc_datain_m[59]));
AND2X1 exu_U2045(.A(exu_n1498), .B(exu_n6398), .Y(exu_n22853));
AND2X1 exu_U2046(.A(exu_n22857), .B(exu_n6399), .Y(ecc_ecc_datain_m[58]));
AND2X1 exu_U2047(.A(exu_n1499), .B(exu_n6400), .Y(exu_n22857));
AND2X1 exu_U2048(.A(exu_n22861), .B(exu_n6401), .Y(ecc_ecc_datain_m[57]));
AND2X1 exu_U2049(.A(exu_n1500), .B(exu_n6402), .Y(exu_n22861));
AND2X1 exu_U2050(.A(exu_n22865), .B(exu_n6403), .Y(ecc_ecc_datain_m[56]));
AND2X1 exu_U2051(.A(exu_n1501), .B(exu_n6404), .Y(exu_n22865));
AND2X1 exu_U2052(.A(exu_n22869), .B(exu_n6405), .Y(ecc_ecc_datain_m[55]));
AND2X1 exu_U2053(.A(exu_n1502), .B(exu_n6406), .Y(exu_n22869));
AND2X1 exu_U2054(.A(exu_n22873), .B(exu_n6407), .Y(ecc_ecc_datain_m[54]));
AND2X1 exu_U2055(.A(exu_n1503), .B(exu_n6408), .Y(exu_n22873));
AND2X1 exu_U2056(.A(exu_n22877), .B(exu_n6409), .Y(ecc_ecc_datain_m[53]));
AND2X1 exu_U2057(.A(exu_n1504), .B(exu_n6410), .Y(exu_n22877));
AND2X1 exu_U2058(.A(exu_n22881), .B(exu_n6411), .Y(ecc_ecc_datain_m[52]));
AND2X1 exu_U2059(.A(exu_n1505), .B(exu_n6412), .Y(exu_n22881));
AND2X1 exu_U2060(.A(exu_n22885), .B(exu_n6413), .Y(ecc_ecc_datain_m[51]));
AND2X1 exu_U2061(.A(exu_n1506), .B(exu_n6414), .Y(exu_n22885));
AND2X1 exu_U2062(.A(exu_n22889), .B(exu_n6415), .Y(ecc_ecc_datain_m[50]));
AND2X1 exu_U2063(.A(exu_n1507), .B(exu_n6416), .Y(exu_n22889));
AND2X1 exu_U2064(.A(exu_n22897), .B(exu_n6419), .Y(ecc_ecc_datain_m[49]));
AND2X1 exu_U2065(.A(exu_n1509), .B(exu_n6420), .Y(exu_n22897));
AND2X1 exu_U2066(.A(exu_n22901), .B(exu_n6421), .Y(ecc_ecc_datain_m[48]));
AND2X1 exu_U2067(.A(exu_n1510), .B(exu_n6422), .Y(exu_n22901));
AND2X1 exu_U2068(.A(exu_n22905), .B(exu_n6423), .Y(ecc_ecc_datain_m[47]));
AND2X1 exu_U2069(.A(exu_n1511), .B(exu_n6424), .Y(exu_n22905));
AND2X1 exu_U2070(.A(exu_n22909), .B(exu_n6425), .Y(ecc_ecc_datain_m[46]));
AND2X1 exu_U2071(.A(exu_n1512), .B(exu_n6426), .Y(exu_n22909));
AND2X1 exu_U2072(.A(exu_n22913), .B(exu_n6427), .Y(ecc_ecc_datain_m[45]));
AND2X1 exu_U2073(.A(exu_n1513), .B(exu_n6428), .Y(exu_n22913));
AND2X1 exu_U2074(.A(exu_n22917), .B(exu_n6429), .Y(ecc_ecc_datain_m[44]));
AND2X1 exu_U2075(.A(exu_n1514), .B(exu_n6430), .Y(exu_n22917));
AND2X1 exu_U2076(.A(exu_n22921), .B(exu_n6431), .Y(ecc_ecc_datain_m[43]));
AND2X1 exu_U2077(.A(exu_n1515), .B(exu_n6432), .Y(exu_n22921));
AND2X1 exu_U2078(.A(exu_n22925), .B(exu_n6433), .Y(ecc_ecc_datain_m[42]));
AND2X1 exu_U2079(.A(exu_n1516), .B(exu_n6434), .Y(exu_n22925));
AND2X1 exu_U2080(.A(exu_n22929), .B(exu_n6435), .Y(ecc_ecc_datain_m[41]));
AND2X1 exu_U2081(.A(exu_n1517), .B(exu_n6436), .Y(exu_n22929));
AND2X1 exu_U2082(.A(exu_n22933), .B(exu_n6437), .Y(ecc_ecc_datain_m[40]));
AND2X1 exu_U2083(.A(exu_n1518), .B(exu_n6438), .Y(exu_n22933));
AND2X1 exu_U2084(.A(exu_n22941), .B(exu_n6441), .Y(ecc_ecc_datain_m[39]));
AND2X1 exu_U2085(.A(exu_n1520), .B(exu_n6442), .Y(exu_n22941));
AND2X1 exu_U2086(.A(exu_n22945), .B(exu_n6443), .Y(ecc_ecc_datain_m[38]));
AND2X1 exu_U2087(.A(exu_n1521), .B(exu_n6444), .Y(exu_n22945));
AND2X1 exu_U2088(.A(exu_n22949), .B(exu_n6445), .Y(ecc_ecc_datain_m[37]));
AND2X1 exu_U2089(.A(exu_n1522), .B(exu_n6446), .Y(exu_n22949));
AND2X1 exu_U2090(.A(exu_n22953), .B(exu_n6447), .Y(ecc_ecc_datain_m[36]));
AND2X1 exu_U2091(.A(exu_n1523), .B(exu_n6448), .Y(exu_n22953));
AND2X1 exu_U2092(.A(exu_n22957), .B(exu_n6449), .Y(ecc_ecc_datain_m[35]));
AND2X1 exu_U2093(.A(exu_n1524), .B(exu_n6450), .Y(exu_n22957));
AND2X1 exu_U2094(.A(exu_n22961), .B(exu_n6451), .Y(ecc_ecc_datain_m[34]));
AND2X1 exu_U2095(.A(exu_n1525), .B(exu_n6452), .Y(exu_n22961));
AND2X1 exu_U2096(.A(exu_n22965), .B(exu_n6453), .Y(ecc_ecc_datain_m[33]));
AND2X1 exu_U2097(.A(exu_n1526), .B(exu_n6454), .Y(exu_n22965));
AND2X1 exu_U2098(.A(exu_n22969), .B(exu_n6455), .Y(ecc_ecc_datain_m[32]));
AND2X1 exu_U2099(.A(exu_n1527), .B(exu_n6456), .Y(exu_n22969));
AND2X1 exu_U2100(.A(exu_n22973), .B(exu_n6457), .Y(ecc_ecc_datain_m[31]));
AND2X1 exu_U2101(.A(exu_n1528), .B(exu_n6458), .Y(exu_n22973));
AND2X1 exu_U2102(.A(exu_n22977), .B(exu_n6459), .Y(ecc_ecc_datain_m[30]));
AND2X1 exu_U2103(.A(exu_n1529), .B(exu_n6460), .Y(exu_n22977));
AND2X1 exu_U2104(.A(exu_n22985), .B(exu_n6463), .Y(ecc_ecc_datain_m[29]));
AND2X1 exu_U2105(.A(exu_n1531), .B(exu_n6464), .Y(exu_n22985));
AND2X1 exu_U2106(.A(exu_n22989), .B(exu_n6465), .Y(ecc_ecc_datain_m[28]));
AND2X1 exu_U2107(.A(exu_n1532), .B(exu_n6466), .Y(exu_n22989));
AND2X1 exu_U2108(.A(exu_n22993), .B(exu_n6467), .Y(ecc_ecc_datain_m[27]));
AND2X1 exu_U2109(.A(exu_n1533), .B(exu_n6468), .Y(exu_n22993));
AND2X1 exu_U2110(.A(exu_n22997), .B(exu_n6469), .Y(ecc_ecc_datain_m[26]));
AND2X1 exu_U2111(.A(exu_n1534), .B(exu_n6470), .Y(exu_n22997));
AND2X1 exu_U2112(.A(exu_n23001), .B(exu_n6471), .Y(ecc_ecc_datain_m[25]));
AND2X1 exu_U2113(.A(exu_n1535), .B(exu_n6472), .Y(exu_n23001));
AND2X1 exu_U2114(.A(exu_n23005), .B(exu_n6473), .Y(ecc_ecc_datain_m[24]));
AND2X1 exu_U2115(.A(exu_n1536), .B(exu_n6474), .Y(exu_n23005));
AND2X1 exu_U2116(.A(exu_n23009), .B(exu_n6475), .Y(ecc_ecc_datain_m[23]));
AND2X1 exu_U2117(.A(exu_n1537), .B(exu_n6476), .Y(exu_n23009));
AND2X1 exu_U2118(.A(exu_n23013), .B(exu_n6477), .Y(ecc_ecc_datain_m[22]));
AND2X1 exu_U2119(.A(exu_n1538), .B(exu_n6478), .Y(exu_n23013));
AND2X1 exu_U2120(.A(exu_n23017), .B(exu_n6479), .Y(ecc_ecc_datain_m[21]));
AND2X1 exu_U2121(.A(exu_n1539), .B(exu_n6480), .Y(exu_n23017));
AND2X1 exu_U2122(.A(exu_n23021), .B(exu_n6481), .Y(ecc_ecc_datain_m[20]));
AND2X1 exu_U2123(.A(exu_n1540), .B(exu_n6482), .Y(exu_n23021));
AND2X1 exu_U2124(.A(exu_n23029), .B(exu_n6485), .Y(ecc_ecc_datain_m[19]));
AND2X1 exu_U2125(.A(exu_n1542), .B(exu_n6486), .Y(exu_n23029));
AND2X1 exu_U2126(.A(exu_n23033), .B(exu_n6487), .Y(ecc_ecc_datain_m[18]));
AND2X1 exu_U2127(.A(exu_n1543), .B(exu_n6488), .Y(exu_n23033));
AND2X1 exu_U2128(.A(exu_n23037), .B(exu_n6489), .Y(ecc_ecc_datain_m[17]));
AND2X1 exu_U2129(.A(exu_n1544), .B(exu_n6490), .Y(exu_n23037));
AND2X1 exu_U2130(.A(exu_n23041), .B(exu_n6491), .Y(ecc_ecc_datain_m[16]));
AND2X1 exu_U2131(.A(exu_n1545), .B(exu_n6492), .Y(exu_n23041));
AND2X1 exu_U2132(.A(ecc_decode_n48), .B(ecc_decode_n18), .Y(ecc_decode_n44));
AND2X1 exu_U2133(.A(exu_n23045), .B(exu_n6493), .Y(ecc_ecc_datain_m[15]));
AND2X1 exu_U2134(.A(exu_n1546), .B(exu_n6494), .Y(exu_n23045));
AND2X1 exu_U2135(.A(exu_n23049), .B(exu_n6495), .Y(ecc_ecc_datain_m[14]));
AND2X1 exu_U2136(.A(exu_n1547), .B(exu_n6496), .Y(exu_n23049));
AND2X1 exu_U2137(.A(ecc_decode_n48), .B(ecc_decode_n21), .Y(ecc_decode_n45));
AND2X1 exu_U2138(.A(exu_n23053), .B(exu_n6497), .Y(ecc_ecc_datain_m[13]));
AND2X1 exu_U2139(.A(exu_n1548), .B(exu_n6498), .Y(exu_n23053));
AND2X1 exu_U2140(.A(exu_n23057), .B(exu_n6499), .Y(ecc_ecc_datain_m[12]));
AND2X1 exu_U2141(.A(exu_n1549), .B(exu_n6500), .Y(exu_n23057));
AND2X1 exu_U2142(.A(ecc_decode_n48), .B(ecc_decode_n22), .Y(ecc_decode_n46));
AND2X1 exu_U2143(.A(exu_n23061), .B(exu_n6501), .Y(ecc_ecc_datain_m[11]));
AND2X1 exu_U2144(.A(exu_n1550), .B(exu_n6502), .Y(exu_n23061));
AND2X1 exu_U2145(.A(ecc_decode_n48), .B(ecc_decode_n24), .Y(ecc_decode_n47));
AND2X1 exu_U2146(.A(exu_n23065), .B(exu_n6503), .Y(ecc_ecc_datain_m[10]));
AND2X1 exu_U2147(.A(exu_n1551), .B(exu_n6504), .Y(exu_n23065));
AND2X1 exu_U2148(.A(exu_n22817), .B(exu_n6379), .Y(ecc_ecc_datain_m[9]));
AND2X1 exu_U2149(.A(exu_n1489), .B(exu_n6380), .Y(exu_n22817));
AND2X1 exu_U2150(.A(exu_n22821), .B(exu_n6381), .Y(ecc_ecc_datain_m[8]));
AND2X1 exu_U2151(.A(exu_n1490), .B(exu_n6382), .Y(exu_n22821));
AND2X1 exu_U2152(.A(exu_n22825), .B(exu_n6383), .Y(ecc_ecc_datain_m[7]));
AND2X1 exu_U2153(.A(exu_n1491), .B(exu_n6384), .Y(exu_n22825));
AND2X1 exu_U2154(.A(exu_n22829), .B(exu_n6385), .Y(ecc_ecc_datain_m[6]));
AND2X1 exu_U2155(.A(exu_n1492), .B(exu_n6386), .Y(exu_n22829));
AND2X1 exu_U2156(.A(exu_n22849), .B(exu_n6395), .Y(ecc_ecc_datain_m[5]));
AND2X1 exu_U2157(.A(exu_n1497), .B(exu_n6396), .Y(exu_n22849));
AND2X1 exu_U2158(.A(exu_n22893), .B(exu_n6417), .Y(ecc_ecc_datain_m[4]));
AND2X1 exu_U2159(.A(exu_n1508), .B(exu_n6418), .Y(exu_n22893));
OR2X1 exu_U2160(.A(exu_n15516), .B(exu_n14775), .Y(ecc_error_data_m[4]));
AND2X1 exu_U2161(.A(exu_n22937), .B(exu_n6439), .Y(ecc_ecc_datain_m[3]));
AND2X1 exu_U2162(.A(exu_n1519), .B(exu_n6440), .Y(exu_n22937));
AND2X1 exu_U2163(.A(exu_tlu_wsr_data_m[2]), .B(exu_n16615), .Y(ecl_byp_3lsb_m[2]));
AND2X1 exu_U2164(.A(exu_n22981), .B(exu_n6461), .Y(ecc_ecc_datain_m[2]));
AND2X1 exu_U2165(.A(exu_n1530), .B(exu_n6462), .Y(exu_n22981));
AND2X1 exu_U2166(.A(ecc_decode_n34), .B(ecc_decode_n18), .Y(ecc_decode_n15));
AND2X1 exu_U2167(.A(exu_tlu_wsr_data_m[1]), .B(exu_n16615), .Y(ecl_byp_3lsb_m[1]));
AND2X1 exu_U2168(.A(exu_n23025), .B(exu_n6483), .Y(ecc_ecc_datain_m[1]));
AND2X1 exu_U2169(.A(exu_n1541), .B(exu_n6484), .Y(exu_n23025));
AND2X1 exu_U2170(.A(ecc_decode_n21), .B(ecc_decode_n34), .Y(ecc_decode_n16));
INVX1 exu_U2171(.A(ecl_read_tlusr_m), .Y(exu_n16582));
AND2X1 exu_U2172(.A(exu_tlu_wsr_data_m[0]), .B(exu_n16615), .Y(ecl_byp_3lsb_m[0]));
AND2X1 exu_U2173(.A(ecc_decode_n22), .B(ecc_decode_n34), .Y(ecc_decode_n17));
AND2X1 exu_U2174(.A(exu_n23069), .B(exu_n6505), .Y(ecc_ecc_datain_m[0]));
AND2X1 exu_U2175(.A(exu_n1552), .B(exu_n6506), .Y(exu_n23069));
INVX1 exu_U2176(.A(exu_n16195), .Y(exu_n16202));
INVX1 exu_U2177(.A(exu_n16194), .Y(exu_n16200));
AND2X1 exu_U2178(.A(ecl_byp_rcc_mux1_sel_w2), .B(ecl_byplog_rs1_n32), .Y(ecl_byplog_rs1_n30));
AND2X1 exu_U2179(.A(exu_n22065), .B(exu_n6066), .Y(bypass_rs2_data_w2[63]));
AND2X1 exu_U2180(.A(exu_n1238), .B(exu_n6067), .Y(exu_n22065));
AND2X1 exu_U2181(.A(exu_n22069), .B(exu_n6068), .Y(bypass_rs2_data_w2[62]));
AND2X1 exu_U2182(.A(exu_n1239), .B(exu_n6069), .Y(exu_n22069));
AND2X1 exu_U2183(.A(exu_n22073), .B(exu_n6070), .Y(bypass_rs2_data_w2[61]));
AND2X1 exu_U2184(.A(exu_n1240), .B(exu_n6071), .Y(exu_n22073));
AND2X1 exu_U2185(.A(exu_n22077), .B(exu_n6072), .Y(bypass_rs2_data_w2[60]));
AND2X1 exu_U2186(.A(exu_n1241), .B(exu_n6073), .Y(exu_n22077));
AND2X1 exu_U2187(.A(exu_n22085), .B(exu_n6076), .Y(bypass_rs2_data_w2[59]));
AND2X1 exu_U2188(.A(exu_n1243), .B(exu_n6077), .Y(exu_n22085));
AND2X1 exu_U2189(.A(exu_n22089), .B(exu_n6078), .Y(bypass_rs2_data_w2[58]));
AND2X1 exu_U2190(.A(exu_n1244), .B(exu_n6079), .Y(exu_n22089));
AND2X1 exu_U2191(.A(exu_n22093), .B(exu_n6080), .Y(bypass_rs2_data_w2[57]));
AND2X1 exu_U2192(.A(exu_n1245), .B(exu_n6081), .Y(exu_n22093));
AND2X1 exu_U2193(.A(exu_n22097), .B(exu_n6082), .Y(bypass_rs2_data_w2[56]));
AND2X1 exu_U2194(.A(exu_n1246), .B(exu_n6083), .Y(exu_n22097));
AND2X1 exu_U2195(.A(exu_n22101), .B(exu_n6084), .Y(bypass_rs2_data_w2[55]));
AND2X1 exu_U2196(.A(exu_n1247), .B(exu_n6085), .Y(exu_n22101));
AND2X1 exu_U2197(.A(exu_n22105), .B(exu_n6086), .Y(bypass_rs2_data_w2[54]));
AND2X1 exu_U2198(.A(exu_n1248), .B(exu_n6087), .Y(exu_n22105));
AND2X1 exu_U2199(.A(exu_n22109), .B(exu_n6088), .Y(bypass_rs2_data_w2[53]));
AND2X1 exu_U2200(.A(exu_n1249), .B(exu_n6089), .Y(exu_n22109));
AND2X1 exu_U2201(.A(exu_n22113), .B(exu_n6090), .Y(bypass_rs2_data_w2[52]));
AND2X1 exu_U2202(.A(exu_n1250), .B(exu_n6091), .Y(exu_n22113));
AND2X1 exu_U2203(.A(exu_n22117), .B(exu_n6092), .Y(bypass_rs2_data_w2[51]));
AND2X1 exu_U2204(.A(exu_n1251), .B(exu_n6093), .Y(exu_n22117));
AND2X1 exu_U2205(.A(exu_n22121), .B(exu_n6094), .Y(bypass_rs2_data_w2[50]));
AND2X1 exu_U2206(.A(exu_n1252), .B(exu_n6095), .Y(exu_n22121));
AND2X1 exu_U2207(.A(exu_n22129), .B(exu_n6098), .Y(bypass_rs2_data_w2[49]));
AND2X1 exu_U2208(.A(exu_n1254), .B(exu_n6099), .Y(exu_n22129));
AND2X1 exu_U2209(.A(exu_n22133), .B(exu_n6100), .Y(bypass_rs2_data_w2[48]));
AND2X1 exu_U2210(.A(exu_n1255), .B(exu_n6101), .Y(exu_n22133));
AND2X1 exu_U2211(.A(exu_n22137), .B(exu_n6102), .Y(bypass_rs2_data_w2[47]));
AND2X1 exu_U2212(.A(exu_n1256), .B(exu_n6103), .Y(exu_n22137));
AND2X1 exu_U2213(.A(exu_n22141), .B(exu_n6104), .Y(bypass_rs2_data_w2[46]));
AND2X1 exu_U2214(.A(exu_n1257), .B(exu_n6105), .Y(exu_n22141));
AND2X1 exu_U2215(.A(exu_n1258), .B(exu_n6107), .Y(exu_n22145));
AND2X1 exu_U2216(.A(exu_n1259), .B(exu_n6109), .Y(exu_n22149));
AND2X1 exu_U2217(.A(exu_n1260), .B(exu_n6111), .Y(exu_n22153));
AND2X1 exu_U2218(.A(exu_n1261), .B(exu_n6113), .Y(exu_n22157));
AND2X1 exu_U2219(.A(exu_n1262), .B(exu_n6115), .Y(exu_n22161));
AND2X1 exu_U2220(.A(exu_n1263), .B(exu_n6117), .Y(exu_n22165));
AND2X1 exu_U2221(.A(exu_n1265), .B(exu_n6121), .Y(exu_n22173));
AND2X1 exu_U2222(.A(exu_n1266), .B(exu_n6123), .Y(exu_n22177));
AND2X1 exu_U2223(.A(exu_n1267), .B(exu_n6125), .Y(exu_n22181));
AND2X1 exu_U2224(.A(exu_n1268), .B(exu_n6127), .Y(exu_n22185));
AND2X1 exu_U2225(.A(exu_n1269), .B(exu_n6129), .Y(exu_n22189));
AND2X1 exu_U2226(.A(exu_n1270), .B(exu_n6131), .Y(exu_n22193));
AND2X1 exu_U2227(.A(exu_n1271), .B(exu_n6133), .Y(exu_n22197));
AND2X1 exu_U2228(.A(exu_n1272), .B(exu_n6135), .Y(exu_n22201));
AND2X1 exu_U2229(.A(exu_n1273), .B(exu_n6137), .Y(exu_n22205));
AND2X1 exu_U2230(.A(exu_n22209), .B(exu_n6138), .Y(bypass_rs2_data_w2[30]));
AND2X1 exu_U2231(.A(exu_n1274), .B(exu_n6139), .Y(exu_n22209));
AND2X1 exu_U2232(.A(exu_n22217), .B(exu_n6142), .Y(bypass_rs2_data_w2[29]));
AND2X1 exu_U2233(.A(exu_n1276), .B(exu_n6143), .Y(exu_n22217));
AND2X1 exu_U2234(.A(exu_n22221), .B(exu_n6144), .Y(bypass_rs2_data_w2[28]));
AND2X1 exu_U2235(.A(exu_n1277), .B(exu_n6145), .Y(exu_n22221));
AND2X1 exu_U2236(.A(exu_n22225), .B(exu_n6146), .Y(bypass_rs2_data_w2[27]));
AND2X1 exu_U2237(.A(exu_n1278), .B(exu_n6147), .Y(exu_n22225));
AND2X1 exu_U2238(.A(exu_n22229), .B(exu_n6148), .Y(bypass_rs2_data_w2[26]));
AND2X1 exu_U2239(.A(exu_n1279), .B(exu_n6149), .Y(exu_n22229));
AND2X1 exu_U2240(.A(exu_n22233), .B(exu_n6150), .Y(bypass_rs2_data_w2[25]));
AND2X1 exu_U2241(.A(exu_n1280), .B(exu_n6151), .Y(exu_n22233));
AND2X1 exu_U2242(.A(exu_n22237), .B(exu_n6152), .Y(bypass_rs2_data_w2[24]));
AND2X1 exu_U2243(.A(exu_n1281), .B(exu_n6153), .Y(exu_n22237));
AND2X1 exu_U2244(.A(exu_n22241), .B(exu_n6154), .Y(bypass_rs2_data_w2[23]));
AND2X1 exu_U2245(.A(exu_n1282), .B(exu_n6155), .Y(exu_n22241));
AND2X1 exu_U2246(.A(exu_n22245), .B(exu_n6156), .Y(bypass_rs2_data_w2[22]));
AND2X1 exu_U2247(.A(exu_n1283), .B(exu_n6157), .Y(exu_n22245));
AND2X1 exu_U2248(.A(exu_n22249), .B(exu_n6158), .Y(bypass_rs2_data_w2[21]));
AND2X1 exu_U2249(.A(exu_n1284), .B(exu_n6159), .Y(exu_n22249));
AND2X1 exu_U2250(.A(exu_n22253), .B(exu_n6160), .Y(bypass_rs2_data_w2[20]));
AND2X1 exu_U2251(.A(exu_n1285), .B(exu_n6161), .Y(exu_n22253));
AND2X1 exu_U2252(.A(exu_n22261), .B(exu_n6164), .Y(bypass_rs2_data_w2[19]));
AND2X1 exu_U2253(.A(exu_n1287), .B(exu_n6165), .Y(exu_n22261));
AND2X1 exu_U2254(.A(exu_n22265), .B(exu_n6166), .Y(bypass_rs2_data_w2[18]));
AND2X1 exu_U2255(.A(exu_n1288), .B(exu_n6167), .Y(exu_n22265));
AND2X1 exu_U2256(.A(exu_n22269), .B(exu_n6168), .Y(bypass_rs2_data_w2[17]));
AND2X1 exu_U2257(.A(exu_n1289), .B(exu_n6169), .Y(exu_n22269));
AND2X1 exu_U2258(.A(exu_n22273), .B(exu_n6170), .Y(bypass_rs2_data_w2[16]));
AND2X1 exu_U2259(.A(exu_n1290), .B(exu_n6171), .Y(exu_n22273));
AND2X1 exu_U2260(.A(exu_n22277), .B(exu_n6172), .Y(bypass_rs2_data_w2[15]));
AND2X1 exu_U2261(.A(exu_n1291), .B(exu_n6173), .Y(exu_n22277));
AND2X1 exu_U2262(.A(exu_n22281), .B(exu_n6174), .Y(bypass_rs2_data_w2[14]));
AND2X1 exu_U2263(.A(exu_n1292), .B(exu_n6175), .Y(exu_n22281));
AND2X1 exu_U2264(.A(exu_n22285), .B(exu_n6176), .Y(bypass_rs2_data_w2[13]));
AND2X1 exu_U2265(.A(exu_n1293), .B(exu_n6177), .Y(exu_n22285));
AND2X1 exu_U2266(.A(exu_n22289), .B(exu_n6178), .Y(bypass_rs2_data_w2[12]));
AND2X1 exu_U2267(.A(exu_n1294), .B(exu_n6179), .Y(exu_n22289));
AND2X1 exu_U2268(.A(exu_n22293), .B(exu_n6180), .Y(bypass_rs2_data_w2[11]));
AND2X1 exu_U2269(.A(exu_n1295), .B(exu_n6181), .Y(exu_n22293));
AND2X1 exu_U2270(.A(exu_n22297), .B(exu_n6182), .Y(bypass_rs2_data_w2[10]));
AND2X1 exu_U2271(.A(exu_n1296), .B(exu_n6183), .Y(exu_n22297));
AND2X1 exu_U2272(.A(exu_n1234), .B(exu_n6059), .Y(exu_n22049));
AND2X1 exu_U2273(.A(exu_n22053), .B(exu_n6060), .Y(bypass_rs2_data_w2[8]));
AND2X1 exu_U2274(.A(exu_n1235), .B(exu_n6061), .Y(exu_n22053));
AND2X1 exu_U2275(.A(exu_n22057), .B(exu_n6062), .Y(bypass_rs2_data_w2[7]));
AND2X1 exu_U2276(.A(exu_n1236), .B(exu_n6063), .Y(exu_n22057));
AND2X1 exu_U2277(.A(exu_n22061), .B(exu_n6064), .Y(bypass_rs2_data_w2[6]));
AND2X1 exu_U2278(.A(exu_n1237), .B(exu_n6065), .Y(exu_n22061));
AND2X1 exu_U2279(.A(exu_n22081), .B(exu_n6074), .Y(bypass_rs2_data_w2[5]));
AND2X1 exu_U2280(.A(exu_n1242), .B(exu_n6075), .Y(exu_n22081));
AND2X1 exu_U2281(.A(exu_n22125), .B(exu_n6096), .Y(bypass_rs2_data_w2[4]));
AND2X1 exu_U2282(.A(exu_n1253), .B(exu_n6097), .Y(exu_n22125));
AND2X1 exu_U2283(.A(exu_n22169), .B(exu_n6118), .Y(bypass_rs2_data_w2[3]));
AND2X1 exu_U2284(.A(exu_n1264), .B(exu_n6119), .Y(exu_n22169));
AND2X1 exu_U2285(.A(exu_n22213), .B(exu_n6140), .Y(bypass_rs2_data_w2[2]));
AND2X1 exu_U2286(.A(exu_n1275), .B(exu_n6141), .Y(exu_n22213));
AND2X1 exu_U2287(.A(exu_n22257), .B(exu_n6162), .Y(bypass_rs2_data_w2[1]));
AND2X1 exu_U2288(.A(exu_n1286), .B(exu_n6163), .Y(exu_n22257));
OR2X1 exu_U2289(.A(exu_n12087), .B(exu_n13503), .Y(ecl_byplog_rs2_N2));
AND2X1 exu_U2290(.A(ecl_byplog_rs2_n24), .B(exu_n9319), .Y(ecl_byplog_rs2_n26));
AND2X1 exu_U2291(.A(ecl_byplog_rs2_n32), .B(ecl_byplog_rs2_n15), .Y(ecl_byplog_rs2_n24));
AND2X1 exu_U2292(.A(exu_n217), .B(exu_n5142), .Y(ecl_byplog_rs2_match_w));
AND2X1 exu_U2293(.A(exu_n15557), .B(ecl_byplog_rs2_n24), .Y(ecl_byplog_rs2_n37));
AND2X1 exu_U2294(.A(exu_n22301), .B(exu_n6184), .Y(bypass_rs2_data_w2[0]));
AND2X1 exu_U2295(.A(exu_n1297), .B(exu_n6185), .Y(exu_n22301));
OR2X1 exu_U2296(.A(exu_n12089), .B(exu_n13505), .Y(ecl_byplog_rs3_N2));
OR2X1 exu_U2297(.A(exu_n12142), .B(exu_n14760), .Y(exu_n19186));
AND2X1 exu_U2298(.A(exu_n157), .B(exu_n16389), .Y(exu_n19213));
AND2X1 exu_U2299(.A(exu_n4072), .B(exu_n9063), .Y(ecl_byplog_rs1_match_w));
AND2X1 exu_U2300(.A(exu_n15557), .B(ecl_byplog_rs1_n35), .Y(ecl_byplog_rs1_n42));
AND2X1 exu_U2301(.A(ecl_byplog_rs1_n35), .B(exu_n9323), .Y(ecl_byplog_rs1_n38));
OR2X1 exu_U2302(.A(ecl_ifu_exu_rs1_d[4]), .B(ecl_ifu_exu_rs1_d[3]), .Y(ecl_byplog_rs1_n41));
AND2X1 exu_U2303(.A(exu_n15), .B(exu_n16389), .Y(ecl_byplog_rs1_n49));
AND2X1 exu_U2304(.A(exu_n854), .B(exu_n5615), .Y(exu_n20681));
AND2X1 exu_U2305(.A(exu_n856), .B(exu_n5617), .Y(exu_n20687));
AND2X1 exu_U2306(.A(exu_n858), .B(exu_n5619), .Y(exu_n20693));
AND2X1 exu_U2307(.A(exu_n860), .B(exu_n5621), .Y(exu_n20699));
AND2X1 exu_U2308(.A(exu_n862), .B(exu_n5623), .Y(exu_n20705));
AND2X1 exu_U2309(.A(exu_n868), .B(exu_n5629), .Y(exu_n20723));
AND2X1 exu_U2310(.A(exu_n890), .B(exu_n5651), .Y(exu_n20789));
AND2X1 exu_U2311(.A(exu_n912), .B(exu_n5673), .Y(exu_n20855));
INVX1 exu_U2312(.A(div_curr_q[30]), .Y(exu_n16434));
INVX1 exu_U2313(.A(div_curr_q[29]), .Y(exu_n16433));
INVX1 exu_U2314(.A(div_curr_q[28]), .Y(exu_n16432));
INVX1 exu_U2315(.A(div_curr_q[27]), .Y(exu_n16431));
INVX1 exu_U2316(.A(div_curr_q[26]), .Y(exu_n16430));
INVX1 exu_U2317(.A(div_curr_q[25]), .Y(exu_n16429));
INVX1 exu_U2318(.A(div_curr_q[24]), .Y(exu_n16428));
INVX1 exu_U2319(.A(div_curr_q[23]), .Y(exu_n16427));
INVX1 exu_U2320(.A(div_curr_q[22]), .Y(exu_n16426));
INVX1 exu_U2321(.A(div_curr_q[21]), .Y(exu_n16425));
INVX1 exu_U2322(.A(div_curr_q[20]), .Y(exu_n16424));
INVX1 exu_U2323(.A(div_curr_q[19]), .Y(exu_n16423));
INVX1 exu_U2324(.A(div_curr_q[18]), .Y(exu_n16422));
INVX1 exu_U2325(.A(div_curr_q[17]), .Y(exu_n16421));
INVX1 exu_U2326(.A(div_curr_q[16]), .Y(exu_n16420));
INVX1 exu_U2327(.A(div_curr_q[15]), .Y(exu_n16419));
INVX1 exu_U2328(.A(div_curr_q[14]), .Y(exu_n16418));
INVX1 exu_U2329(.A(div_curr_q[13]), .Y(exu_n16417));
INVX1 exu_U2330(.A(div_curr_q[12]), .Y(exu_n16416));
INVX1 exu_U2331(.A(div_curr_q[11]), .Y(exu_n16415));
INVX1 exu_U2332(.A(div_curr_q[10]), .Y(exu_n16414));
INVX1 exu_U2333(.A(div_curr_q[9]), .Y(exu_n16413));
INVX1 exu_U2334(.A(div_curr_q[8]), .Y(exu_n16412));
INVX1 exu_U2335(.A(div_curr_q[7]), .Y(exu_n16411));
INVX1 exu_U2336(.A(div_curr_q[6]), .Y(exu_n16410));
INVX1 exu_U2337(.A(div_curr_q[5]), .Y(exu_n16409));
INVX1 exu_U2338(.A(div_curr_q[4]), .Y(exu_n16408));
INVX1 exu_U2339(.A(div_curr_q[3]), .Y(exu_n16407));
INVX1 exu_U2340(.A(div_curr_q[2]), .Y(exu_n16406));
INVX1 exu_U2341(.A(div_curr_q[1]), .Y(exu_n16405));
INVX1 exu_U2342(.A(div_curr_q[0]), .Y(exu_n16404));
AND2X1 exu_U2343(.A(exu_n16558), .B(ecl_divcntl_upper32_equal_d1), .Y(ecl_divcntl_n79));
AND2X1 exu_U2344(.A(exu_n2567), .B(exu_n7595), .Y(exu_n26354));
OR2X1 exu_U2345(.A(exu_n12088), .B(exu_n13504), .Y(ecl_byplog_rs3h_N2));
AND2X1 exu_U2346(.A(exu_n19238), .B(exu_n19222), .Y(exu_n19231));
AND2X1 exu_U2347(.A(exu_n221), .B(exu_n5146), .Y(ecl_byplog_rs3h_match_w));
AND2X1 exu_U2348(.A(exu_n15557), .B(exu_n19231), .Y(exu_n19243));
AND2X1 exu_U2349(.A(exu_n19231), .B(exu_n5537), .Y(exu_n19233));
OR2X1 exu_U2350(.A(exu_n12145), .B(exu_n14760), .Y(exu_n19222));
AND2X1 exu_U2351(.A(exu_n151), .B(exu_n16389), .Y(exu_n19249));
AND2X1 exu_U2352(.A(exu_n4111), .B(exu_n9105), .Y(ecl_ccr_mux_ccr_out_n43));
AND2X1 exu_U2353(.A(exu_n4110), .B(exu_n9104), .Y(ecl_ccr_mux_ccr_out_n44));
AND2X1 exu_U2354(.A(exu_n4109), .B(exu_n9103), .Y(ecl_ccr_mux_ccr_out_n37));
AND2X1 exu_U2355(.A(exu_n4108), .B(exu_n9102), .Y(ecl_ccr_mux_ccr_out_n38));
AND2X1 exu_U2356(.A(exu_n4107), .B(exu_n9101), .Y(ecl_ccr_mux_ccr_out_n31));
AND2X1 exu_U2357(.A(exu_n4106), .B(exu_n9100), .Y(ecl_ccr_mux_ccr_out_n32));
AND2X1 exu_U2358(.A(exu_n4105), .B(exu_n9099), .Y(ecl_ccr_mux_ccr_out_n25));
AND2X1 exu_U2359(.A(exu_n4104), .B(exu_n9098), .Y(ecl_ccr_mux_ccr_out_n26));
AND2X1 exu_U2360(.A(exu_n4103), .B(exu_n9097), .Y(ecl_ccr_mux_ccr_out_n19));
AND2X1 exu_U2361(.A(exu_n4102), .B(exu_n9096), .Y(ecl_ccr_mux_ccr_out_n20));
AND2X1 exu_U2362(.A(exu_n4101), .B(exu_n9095), .Y(ecl_ccr_mux_ccr_out_n13));
AND2X1 exu_U2363(.A(exu_n4100), .B(exu_n9094), .Y(ecl_ccr_mux_ccr_out_n14));
AND2X1 exu_U2364(.A(exu_n4099), .B(exu_n9093), .Y(ecl_ccr_mux_ccr_out_n7));
AND2X1 exu_U2365(.A(exu_n4098), .B(exu_n9092), .Y(ecl_ccr_mux_ccr_out_n8));
AND2X1 exu_U2366(.A(exu_n4097), .B(exu_n9091), .Y(ecl_ccr_mux_ccr_out_n1));
AND2X1 exu_U2367(.A(exu_n4096), .B(exu_n9090), .Y(ecl_ccr_mux_ccr_out_n2));
AND2X1 exu_U2368(.A(exu_n4551), .B(exu_n9342), .Y(ecl_ccr_use_cc_w));
OR2X1 exu_U2369(.A(ecl_eccctl_rs1_ce_m), .B(ecl_eccctl_rs2_ce_m), .Y(ecl_eccctl_n17));
AND2X1 exu_U2370(.A(exu_n16592), .B(exu_n16593), .Y(ecl_eccctl_n35));
INVX1 exu_U2371(.A(ecl_eccctl_rs2_ue_m), .Y(exu_n16593));
INVX1 exu_U2372(.A(ecl_eccctl_rs1_ue_m), .Y(exu_n16594));
AND2X1 exu_U2373(.A(exu_n3990), .B(exu_n9005), .Y(exu_n31670));
AND2X1 exu_U2374(.A(exu_n3989), .B(exu_n9004), .Y(exu_n31671));
AND2X1 exu_U2375(.A(exu_n3986), .B(exu_n9002), .Y(exu_n31665));
AND2X1 exu_U2376(.A(exu_n3971), .B(exu_n8987), .Y(exu_n31621));
AND2X1 exu_U2377(.A(exu_n3974), .B(exu_n8989), .Y(exu_n31627));
AND2X1 exu_U2378(.A(exu_n3976), .B(exu_n8992), .Y(exu_n31635));
AND2X1 exu_U2379(.A(exu_n3979), .B(exu_n8994), .Y(exu_n31641));
AND2X1 exu_U2380(.A(exu_n3981), .B(exu_n8997), .Y(exu_n31651));
AND2X1 exu_U2381(.A(exu_n3984), .B(exu_n8999), .Y(exu_n31657));
INVX1 exu_U2382(.A(tlu_exu_agp_tid[0]), .Y(rml_n35));
INVX1 exu_U2383(.A(ecl_rml_early_flush_w), .Y(exu_n16608));
AND2X1 exu_U2384(.A(exu_n4012), .B(exu_n9028), .Y(rml_cwp_cwp_output_mux_n38));
AND2X1 exu_U2385(.A(exu_n4010), .B(exu_n9026), .Y(rml_cwp_cwp_output_mux_n32));
INVX1 exu_U2386(.A(ecl_wb_byplog_wen_g2), .Y(exu_n16600));
AND2X1 exu_U2387(.A(rml_n106), .B(rml_rml_kill_w), .Y(rml_canrestore_wen_w));
OR2X1 exu_U2388(.A(exu_n13448), .B(rml_rml_canrestore_wen_w), .Y(rml_n106));
AND2X1 exu_U2389(.A(rml_n80), .B(rml_rml_kill_w), .Y(rml_otherwin_wen_w));
OR2X1 exu_U2390(.A(exu_n13443), .B(rml_rml_otherwin_wen_w), .Y(rml_n80));
AND2X1 exu_U2391(.A(rml_n99), .B(rml_rml_kill_w), .Y(rml_cleanwin_wen_w));
OR2X1 exu_U2392(.A(exu_n13446), .B(rml_rml_cleanwin_wen_w), .Y(rml_n99));
AND2X1 exu_U2393(.A(exu_n4539), .B(rml_rml_kill_w), .Y(rml_wstate_wen_w));
INVX1 exu_U2394(.A(rml_cwp_swap_req_vec[2]), .Y(exu_n16625));
INVX1 exu_U2395(.A(rml_cwp_swap_req_vec[1]), .Y(exu_n16626));
INVX1 exu_U2396(.A(rml_cwp_cwp_output_queue_pv[2]), .Y(exu_n16618));
INVX1 exu_U2397(.A(rml_cwp_swap_req_vec[0]), .Y(exu_n16511));
INVX1 exu_U2398(.A(rml_cwp_cwp_output_queue_pv[0]), .Y(exu_n16616));
INVX1 exu_U2399(.A(rml_cwp_swap_req_vec[3]), .Y(exu_n16624));
OR2X1 exu_U2400(.A(rml_cwp_swap_slot0_state[1]), .B(rml_cwp_swap_slot0_state_valid[0]), .Y(rml_cwp_swap_req_vec[0]));
AND2X1 exu_U2401(.A(ecl_tid_d[1]), .B(ecl_tid_d[0]), .Y(ecl_thr_d[3]));
AND2X1 exu_U2402(.A(exu_n3626), .B(exu_n8643), .Y(alu_va_e[63]));
AND2X1 exu_U2403(.A(exu_n4902), .B(exu_n16588), .Y(rml_n79));
INVX1 exu_U2404(.A(rml_save_e), .Y(exu_n16606));
INVX1 exu_U2405(.A(rml_restore_e), .Y(exu_n16604));
AND2X1 exu_U2406(.A(exu_n4540), .B(exu_n9337), .Y(ecl_writeback_n134));
INVX1 exu_U2407(.A(rml_ecl_other_e), .Y(exu_n16603));
OR2X1 exu_U2408(.A(ecl_writeback_sraddr_w[3]), .B(ecl_writeback_sraddr_w[5]), .Y(ecl_writeback_n57));
AND2X1 exu_U2409(.A(exu_n4541), .B(ecl_writeback_wrsr_w), .Y(ecl_writeback_n58));
INVX1 exu_U2410(.A(ecl_writeback_sraddr_w[0]), .Y(exu_n16553));
OR2X1 exu_U2411(.A(exu_n13438), .B(exu_n14758), .Y(ecl_byplog_rs1_n29));
OR2X1 exu_U2412(.A(ecl_ifu_exu_rs2_d[4]), .B(ecl_ifu_exu_rs2_d[3]), .Y(ecl_byplog_rs2_n51));
AND2X1 exu_U2413(.A(exu_n19202), .B(exu_n19186), .Y(exu_n19195));
AND2X1 exu_U2414(.A(exu_n219), .B(exu_n5144), .Y(ecl_byplog_rs3_match_w));
AND2X1 exu_U2415(.A(exu_n15557), .B(exu_n19195), .Y(exu_n19207));
AND2X1 exu_U2416(.A(exu_n19195), .B(exu_n5533), .Y(exu_n19197));
OR2X1 exu_U2417(.A(ecl_ifu_exu_rs3_d[4]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n19219));
OR2X1 exu_U2418(.A(ecc_rs1_err_e[2]), .B(ecc_rs1_err_e[1]), .Y(ecc_chk_rs1_n9));
OR2X1 exu_U2419(.A(ecc_rs2_err_e[2]), .B(ecc_rs2_err_e[1]), .Y(exu_n20002));
OR2X1 exu_U2420(.A(ecc_rs3_err_e[2]), .B(ecc_rs3_err_e[1]), .Y(exu_n20138));
AND2X1 exu_U2421(.A(ecl_n69), .B(exu_n15436), .Y(ecl_cancel_rs3_ecc_e));
INVX1 exu_U2422(.A(ecl_divcntl_subnext_mux_in1[0]), .Y(exu_n16437));
OR2X1 exu_U2423(.A(exu_n15638), .B(exu_n15823), .Y(exu_n17040));
AND2X1 exu_U2424(.A(exu_n4919), .B(exu_n9630), .Y(div_n68));
AND2X1 exu_U2425(.A(exu_n4924), .B(exu_n9635), .Y(div_n67));
OR2X1 exu_U2426(.A(exu_n13497), .B(exu_n14814), .Y(div_ecl_detect_zero_low));
AND2X1 exu_U2427(.A(exu_n4914), .B(exu_n9625), .Y(div_n37));
INVX1 exu_U2428(.A(ecl_flush_w1), .Y(exu_n16607));
AND2X1 exu_U2429(.A(exu_n248), .B(exu_n5175), .Y(exu_n17789));
AND2X1 exu_U2430(.A(exu_n250), .B(exu_n5177), .Y(exu_n17795));
AND2X1 exu_U2431(.A(exu_n306), .B(exu_n5233), .Y(exu_n17963));
AND2X1 exu_U2432(.A(exu_n308), .B(exu_n5235), .Y(exu_n17969));
AND2X1 exu_U2433(.A(exu_n310), .B(exu_n5237), .Y(exu_n17975));
AND2X1 exu_U2434(.A(exu_n4884), .B(exu_n9607), .Y(rml_n36));
AND2X1 exu_U2435(.A(exu_n4155), .B(exu_n9133), .Y(rml_cwp_inc_n3));
INVX1 exu_U2436(.A(rml_rml_ecl_cwp_e[0]), .Y(exu_n16569));
AND2X1 exu_U2437(.A(exu_n16504), .B(exu_n16503), .Y(ecl_divcntl_n66));
AND2X1 exu_U2438(.A(rml_tid_d[1]), .B(rml_tid_d[0]), .Y(exu_n15948));
OR2X1 exu_U2439(.A(exu_n15615), .B(exu_n15898), .Y(exu_n16876));
AND2X1 exu_U2440(.A(exu_n4008), .B(exu_n9024), .Y(rml_cwp_cwp_output_mux_n26));
AND2X1 exu_U2441(.A(rml_cwp_wen_nokill_w), .B(rml_rml_kill_w), .Y(rml_cwp_wen_w));
AND2X1 exu_U2442(.A(rml_n102), .B(rml_rml_kill_w), .Y(rml_cansave_wen_w));
OR2X1 exu_U2443(.A(exu_n13447), .B(rml_rml_cansave_wen_w), .Y(rml_n102));
AND2X1 exu_U2444(.A(tlu_exu_agp_tid[1]), .B(rml_n35), .Y(rml_agp_thr[2]));
INVX1 exu_U2445(.A(rml_tid_e[1]), .Y(exu_n16571));
AND2X1 exu_U2446(.A(exu_n3996), .B(exu_n9013), .Y(exu_n31693));
AND2X1 exu_U2447(.A(exu_n3992), .B(exu_n9008), .Y(exu_n31680));
AND2X1 exu_U2448(.A(exu_n3994), .B(exu_n9010), .Y(exu_n31686));
INVX1 exu_U2449(.A(exu_n16195), .Y(exu_n16201));
AND2X1 exu_U2450(.A(exu_n3764), .B(exu_n8843), .Y(div_gencc_in_15));
AND2X1 exu_U2451(.A(exu_n3766), .B(exu_n8845), .Y(div_gencc_in_13));
AND2X1 exu_U2452(.A(exu_n3768), .B(exu_n8847), .Y(div_gencc_in_11));
AND2X1 exu_U2453(.A(exu_n3770), .B(exu_n8849), .Y(div_gencc_in_0));
AND2X1 exu_U2454(.A(exu_n4416), .B(exu_n9264), .Y(div_low32or_n5));
AND2X1 exu_U2455(.A(exu_n3748), .B(exu_n8827), .Y(div_gencc_in_2));
AND2X1 exu_U2456(.A(exu_n3750), .B(exu_n8829), .Y(div_gencc_in_28));
AND2X1 exu_U2457(.A(exu_n3752), .B(exu_n8831), .Y(div_gencc_in_26));
AND2X1 exu_U2458(.A(exu_n3754), .B(exu_n8833), .Y(div_gencc_in_24));
AND2X1 exu_U2459(.A(exu_n3737), .B(exu_n8816), .Y(div_gencc_in_3));
AND2X1 exu_U2460(.A(exu_n4421), .B(exu_n9269), .Y(div_low32or_n19));
AND2X1 exu_U2461(.A(exu_n4006), .B(exu_n9022), .Y(rml_cwp_cwp_output_mux_n20));
AND2X1 exu_U2462(.A(exu_n16396), .B(rml_cwp_swap_thr[2]), .Y(rml_cwp_swap_sel[2]));
INVX1 exu_U2463(.A(mux_drive_disable), .Y(exu_n16396));
OR2X1 exu_U2464(.A(rml_cwp_swap_tid[1]), .B(rml_cwp_swap_thr[1]), .Y(rml_cwp_n38));
OR2X1 exu_U2465(.A(exu_n13332), .B(exu_n14639), .Y(alu_ecl_log_n64_e));
AND2X1 exu_U2466(.A(exu_n3411), .B(exu_n8492), .Y(exu_n28941));
AND2X1 exu_U2467(.A(exu_n4941), .B(exu_n9655), .Y(alu_n109));
AND2X1 exu_U2468(.A(exu_n4940), .B(exu_n9654), .Y(alu_n110));
AND2X1 exu_U2469(.A(exu_n4937), .B(exu_n9652), .Y(alu_n104));
AND2X1 exu_U2470(.A(exu_n4942), .B(exu_n9657), .Y(alu_n118));
AND2X1 exu_U2471(.A(exu_n4945), .B(exu_n9659), .Y(alu_n124));
INVX1 exu_U2472(.A(alu_logic_rs1_data_bf1[63]), .Y(exu_n16552));
AND2X1 exu_U2473(.A(exu_n148), .B(exu_n5115), .Y(exu_n17357));
OR2X1 exu_U2474(.A(exu_n13367), .B(exu_n14674), .Y(alu_ecl_log_n32_e));
AND2X1 exu_U2475(.A(exu_n3481), .B(exu_n8562), .Y(exu_n29151));
AND2X1 exu_U2476(.A(exu_n4931), .B(exu_n9644), .Y(alu_n79));
AND2X1 exu_U2477(.A(exu_n4930), .B(exu_n9643), .Y(alu_n80));
AND2X1 exu_U2478(.A(exu_n4927), .B(exu_n9641), .Y(alu_n74));
AND2X1 exu_U2479(.A(exu_n4936), .B(exu_n9649), .Y(alu_n93));
AND2X1 exu_U2480(.A(exu_n4935), .B(exu_n9648), .Y(alu_n94));
AND2X1 exu_U2481(.A(exu_n4932), .B(exu_n9646), .Y(alu_n88));
AND2X1 exu_U2482(.A(alu_logic_rs1_data_bf1[31]), .B(exu_n16512), .Y(ecl_n144));
OR2X1 exu_U2483(.A(alu_ecl_adderin2_31_e), .B(alu_logic_rs1_data_bf1[31]), .Y(ecl_n143));
INVX1 exu_U2484(.A(ecl_ccr_setcc_w2), .Y(exu_n16584));
INVX1 exu_U2485(.A(ecl_divcntl_gencc_in_msb_l_d1), .Y(exu_n16558));
AND2X1 exu_U2486(.A(ecl_divcntl_sel_div_d1), .B(exu_n15487), .Y(ecl_divcntl_n80));
INVX1 exu_U2487(.A(ecl_divcntl_low32_nonzero_d1), .Y(exu_n16557));
AND2X1 exu_U2488(.A(exu_n4513), .B(ecl_divcntl_sel_div_d1), .Y(ecl_divcntl_n69));
AND2X1 exu_U2489(.A(exu_n15347), .B(ecl_divcntl_sel_div_d1), .Y(ecl_divcntl_n76));
AND2X1 exu_U2490(.A(ecl_divcntl_sel_div_d1), .B(ecl_div_muls), .Y(ecl_divcntl_n84));
OR2X1 exu_U2491(.A(ecl_ccr_n35), .B(exu_n14772), .Y(ecl_ccr_n14));
AND2X1 exu_U2492(.A(ifu_exu_inst_vld_w), .B(exu_n9343), .Y(ecl_ccr_n36));
AND2X1 exu_U2493(.A(rml_tid_d[1]), .B(rml_tid_d[0]), .Y(rml_thr_d[3]));
INVX1 exu_U2494(.A(ifu_tlu_sraddr_d[1]), .Y(exu_n16375));
AND2X1 exu_U2495(.A(rml_tid_d[1]), .B(rml_tid_d[0]), .Y(exu_n15949));
AND2X1 exu_U2496(.A(exu_n4079), .B(exu_n9074), .Y(ecl_writeback_rdpr_mux1_n2));
AND2X1 exu_U2497(.A(exu_n4081), .B(exu_n9076), .Y(ecl_writeback_rdpr_mux1_n8));
OR2X1 exu_U2498(.A(ifu_tlu_sraddr_d[0]), .B(ifu_tlu_sraddr_d[2]), .Y(ecl_writeback_n91));
AND2X1 exu_U2499(.A(exu_n4083), .B(exu_n9078), .Y(ecl_writeback_rdpr_mux1_n14));
AND2X1 exu_U2500(.A(exu_n15744), .B(ecl_writeback_n85), .Y(ecl_writeback_n180));
AND2X1 exu_U2501(.A(exu_n15743), .B(ecl_writeback_n81), .Y(ecl_writeback_n178));
AND2X1 exu_U2502(.A(ecl_div_muls), .B(ecl_mdqctl_n46), .Y(ecl_mdqctl_wb_yreg_shift_g));
AND2X1 exu_U2503(.A(exu_n15741), .B(ecl_writeback_n77), .Y(ecl_writeback_n175));
AND2X1 exu_U2504(.A(exu_n2575), .B(exu_n7603), .Y(exu_n26378));
AND2X1 exu_U2505(.A(exu_n2577), .B(exu_n7604), .Y(exu_n26383));
AND2X1 exu_U2506(.A(exu_n2579), .B(exu_n7606), .Y(exu_n26389));
AND2X1 exu_U2507(.A(exu_n2581), .B(exu_n7608), .Y(exu_n26395));
AND2X1 exu_U2508(.A(exu_n2585), .B(exu_n7612), .Y(exu_n26407));
AND2X1 exu_U2509(.A(exu_n2587), .B(exu_n7614), .Y(exu_n26413));
AND2X1 exu_U2510(.A(exu_n2589), .B(exu_n7616), .Y(exu_n26419));
AND2X1 exu_U2511(.A(exu_n2591), .B(exu_n7618), .Y(exu_n26425));
AND2X1 exu_U2512(.A(exu_n2593), .B(exu_n7620), .Y(exu_n26431));
AND2X1 exu_U2513(.A(exu_n2595), .B(exu_n7622), .Y(exu_n26437));
AND2X1 exu_U2514(.A(exu_n2597), .B(exu_n7624), .Y(exu_n26443));
AND2X1 exu_U2515(.A(exu_n2599), .B(exu_n7626), .Y(exu_n26449));
AND2X1 exu_U2516(.A(exu_n2601), .B(exu_n7628), .Y(exu_n26455));
AND2X1 exu_U2517(.A(exu_n2603), .B(exu_n7630), .Y(exu_n26461));
AND2X1 exu_U2518(.A(exu_n2607), .B(exu_n7634), .Y(exu_n26473));
AND2X1 exu_U2519(.A(exu_n2609), .B(exu_n7636), .Y(exu_n26479));
AND2X1 exu_U2520(.A(exu_n2611), .B(exu_n7638), .Y(exu_n26485));
AND2X1 exu_U2521(.A(exu_n2613), .B(exu_n7640), .Y(exu_n26491));
AND2X1 exu_U2522(.A(exu_n2615), .B(exu_n7642), .Y(exu_n26497));
AND2X1 exu_U2523(.A(exu_n2617), .B(exu_n7644), .Y(exu_n26503));
AND2X1 exu_U2524(.A(exu_n2619), .B(exu_n7646), .Y(exu_n26509));
AND2X1 exu_U2525(.A(exu_n2621), .B(exu_n7648), .Y(exu_n26515));
AND2X1 exu_U2526(.A(exu_n2623), .B(exu_n7650), .Y(exu_n26521));
AND2X1 exu_U2527(.A(exu_n2625), .B(exu_n7652), .Y(exu_n26527));
AND2X1 exu_U2528(.A(exu_n2629), .B(exu_n7656), .Y(exu_n26539));
AND2X1 exu_U2529(.A(exu_n2631), .B(exu_n7658), .Y(exu_n26545));
AND2X1 exu_U2530(.A(exu_n2633), .B(exu_n7660), .Y(exu_n26551));
AND2X1 exu_U2531(.A(exu_n2635), .B(exu_n7662), .Y(exu_n26557));
AND2X1 exu_U2532(.A(exu_n2637), .B(exu_n7664), .Y(exu_n26563));
AND2X1 exu_U2533(.A(exu_n2639), .B(exu_n7666), .Y(exu_n26569));
AND2X1 exu_U2534(.A(exu_n2641), .B(exu_n7668), .Y(exu_n26575));
AND2X1 exu_U2535(.A(exu_n2643), .B(exu_n7670), .Y(exu_n26581));
AND2X1 exu_U2536(.A(exu_n2645), .B(exu_n7672), .Y(exu_n26587));
AND2X1 exu_U2537(.A(exu_n2647), .B(exu_n7673), .Y(exu_n26592));
AND2X1 exu_U2538(.A(exu_n2651), .B(exu_n7677), .Y(exu_n26604));
AND2X1 exu_U2539(.A(exu_n2653), .B(exu_n7679), .Y(exu_n26610));
AND2X1 exu_U2540(.A(exu_n2655), .B(exu_n7681), .Y(exu_n26616));
AND2X1 exu_U2541(.A(exu_n2657), .B(exu_n7683), .Y(exu_n26622));
AND2X1 exu_U2542(.A(exu_n2659), .B(exu_n7685), .Y(exu_n26628));
AND2X1 exu_U2543(.A(exu_n2661), .B(exu_n7687), .Y(exu_n26634));
AND2X1 exu_U2544(.A(exu_n2663), .B(exu_n7689), .Y(exu_n26640));
AND2X1 exu_U2545(.A(exu_n2665), .B(exu_n7691), .Y(exu_n26646));
AND2X1 exu_U2546(.A(exu_n2667), .B(exu_n7693), .Y(exu_n26652));
AND2X1 exu_U2547(.A(exu_n2669), .B(exu_n7695), .Y(exu_n26658));
AND2X1 exu_U2548(.A(exu_n2673), .B(exu_n7699), .Y(exu_n26670));
AND2X1 exu_U2549(.A(exu_n2675), .B(exu_n7701), .Y(exu_n26676));
AND2X1 exu_U2550(.A(exu_n2677), .B(exu_n7703), .Y(exu_n26682));
AND2X1 exu_U2551(.A(exu_n2679), .B(exu_n7705), .Y(exu_n26688));
AND2X1 exu_U2552(.A(exu_n2681), .B(exu_n7707), .Y(exu_n26694));
AND2X1 exu_U2553(.A(exu_n2683), .B(exu_n7709), .Y(exu_n26700));
AND2X1 exu_U2554(.A(exu_n2685), .B(exu_n7711), .Y(exu_n26706));
AND2X1 exu_U2555(.A(exu_n2687), .B(exu_n7713), .Y(exu_n26712));
AND2X1 exu_U2556(.A(exu_n2689), .B(exu_n7715), .Y(exu_n26718));
AND2X1 exu_U2557(.A(exu_n2691), .B(exu_n7717), .Y(exu_n26724));
INVX1 exu_U2558(.A(ecl_tid_e[0]), .Y(exu_n16579));
AND2X1 exu_U2559(.A(exu_n2569), .B(exu_n7597), .Y(exu_n26360));
AND2X1 exu_U2560(.A(exu_n2571), .B(exu_n7599), .Y(exu_n26366));
AND2X1 exu_U2561(.A(exu_n2573), .B(exu_n7601), .Y(exu_n26372));
AND2X1 exu_U2562(.A(exu_n2583), .B(exu_n7610), .Y(exu_n26401));
AND2X1 exu_U2563(.A(exu_n2605), .B(exu_n7632), .Y(exu_n26467));
AND2X1 exu_U2564(.A(exu_n2627), .B(exu_n7654), .Y(exu_n26533));
AND2X1 exu_U2565(.A(exu_n2649), .B(exu_n7675), .Y(exu_n26598));
AND2X1 exu_U2566(.A(exu_n2671), .B(exu_n7697), .Y(exu_n26664));
AND2X1 exu_U2567(.A(exu_n2693), .B(exu_n7719), .Y(exu_n26730));
INVX1 exu_U2568(.A(se), .Y(exu_n29301));
INVX1 exu_U2569(.A(se), .Y(exu_n29366));
AND2X1 exu_U2570(.A(exu_n4688), .B(exu_n9448), .Y(bypass_sr_out_mux_n17));
AND2X1 exu_U2571(.A(exu_n4689), .B(exu_n9450), .Y(bypass_sr_out_mux_n21));
AND2X1 exu_U2572(.A(exu_n4690), .B(exu_n9452), .Y(bypass_sr_out_mux_n25));
AND2X1 exu_U2573(.A(exu_n4691), .B(exu_n9454), .Y(bypass_sr_out_mux_n29));
AND2X1 exu_U2574(.A(exu_n4693), .B(exu_n9458), .Y(bypass_sr_out_mux_n37));
AND2X1 exu_U2575(.A(exu_n4694), .B(exu_n9460), .Y(bypass_sr_out_mux_n41));
AND2X1 exu_U2576(.A(exu_n4695), .B(exu_n9462), .Y(bypass_sr_out_mux_n45));
AND2X1 exu_U2577(.A(exu_n4696), .B(exu_n9464), .Y(bypass_sr_out_mux_n49));
AND2X1 exu_U2578(.A(exu_n4697), .B(exu_n9466), .Y(bypass_sr_out_mux_n53));
AND2X1 exu_U2579(.A(exu_n4698), .B(exu_n9468), .Y(bypass_sr_out_mux_n57));
AND2X1 exu_U2580(.A(exu_n4699), .B(exu_n9470), .Y(bypass_sr_out_mux_n61));
AND2X1 exu_U2581(.A(exu_n4700), .B(exu_n9472), .Y(bypass_sr_out_mux_n65));
AND2X1 exu_U2582(.A(exu_n4701), .B(exu_n9474), .Y(bypass_sr_out_mux_n69));
AND2X1 exu_U2583(.A(exu_n4702), .B(exu_n9476), .Y(bypass_sr_out_mux_n73));
AND2X1 exu_U2584(.A(exu_n4704), .B(exu_n9480), .Y(bypass_sr_out_mux_n81));
AND2X1 exu_U2585(.A(exu_n4705), .B(exu_n9482), .Y(bypass_sr_out_mux_n85));
AND2X1 exu_U2586(.A(exu_n4706), .B(exu_n9484), .Y(bypass_sr_out_mux_n89));
AND2X1 exu_U2587(.A(exu_n4707), .B(exu_n9486), .Y(bypass_sr_out_mux_n93));
AND2X1 exu_U2588(.A(exu_n4708), .B(exu_n9488), .Y(bypass_sr_out_mux_n97));
AND2X1 exu_U2589(.A(exu_n4709), .B(exu_n9490), .Y(bypass_sr_out_mux_n101));
AND2X1 exu_U2590(.A(exu_n4710), .B(exu_n9492), .Y(bypass_sr_out_mux_n105));
AND2X1 exu_U2591(.A(exu_n4711), .B(exu_n9494), .Y(bypass_sr_out_mux_n109));
AND2X1 exu_U2592(.A(exu_n4712), .B(exu_n9496), .Y(bypass_sr_out_mux_n113));
AND2X1 exu_U2593(.A(exu_n4713), .B(exu_n9498), .Y(bypass_sr_out_mux_n117));
AND2X1 exu_U2594(.A(exu_n4715), .B(exu_n9502), .Y(bypass_sr_out_mux_n125));
AND2X1 exu_U2595(.A(exu_n4716), .B(exu_n9504), .Y(bypass_sr_out_mux_n129));
AND2X1 exu_U2596(.A(exu_n4717), .B(exu_n9506), .Y(bypass_sr_out_mux_n133));
AND2X1 exu_U2597(.A(exu_n4718), .B(exu_n9508), .Y(bypass_sr_out_mux_n137));
AND2X1 exu_U2598(.A(exu_n4719), .B(exu_n9510), .Y(bypass_sr_out_mux_n141));
AND2X1 exu_U2599(.A(exu_n4720), .B(exu_n9512), .Y(bypass_sr_out_mux_n145));
AND2X1 exu_U2600(.A(exu_n4721), .B(exu_n9514), .Y(bypass_sr_out_mux_n149));
AND2X1 exu_U2601(.A(exu_n4722), .B(exu_n9516), .Y(bypass_sr_out_mux_n153));
AND2X1 exu_U2602(.A(exu_n4723), .B(exu_n9518), .Y(bypass_sr_out_mux_n157));
AND2X1 exu_U2603(.A(exu_n4724), .B(exu_n9520), .Y(bypass_sr_out_mux_n161));
AND2X1 exu_U2604(.A(exu_n4726), .B(exu_n9524), .Y(bypass_sr_out_mux_n169));
AND2X1 exu_U2605(.A(exu_n4727), .B(exu_n9526), .Y(bypass_sr_out_mux_n173));
AND2X1 exu_U2606(.A(exu_n4728), .B(exu_n9528), .Y(bypass_sr_out_mux_n177));
AND2X1 exu_U2607(.A(exu_n4729), .B(exu_n9530), .Y(bypass_sr_out_mux_n181));
AND2X1 exu_U2608(.A(exu_n4730), .B(exu_n9532), .Y(bypass_sr_out_mux_n185));
AND2X1 exu_U2609(.A(ecc_decode_n44), .B(ecc_decode_n27), .Y(ecc_error_data_m[25]));
AND2X1 exu_U2610(.A(exu_n4731), .B(exu_n9534), .Y(bypass_sr_out_mux_n189));
AND2X1 exu_U2611(.A(ecc_decode_n44), .B(ecc_decode_n29), .Y(ecc_error_data_m[24]));
AND2X1 exu_U2612(.A(exu_n4732), .B(exu_n9536), .Y(bypass_sr_out_mux_n193));
AND2X1 exu_U2613(.A(ecc_decode_n45), .B(ecc_decode_n27), .Y(ecc_error_data_m[23]));
AND2X1 exu_U2614(.A(exu_n4733), .B(exu_n9538), .Y(bypass_sr_out_mux_n197));
AND2X1 exu_U2615(.A(ecc_decode_n45), .B(ecc_decode_n29), .Y(ecc_error_data_m[22]));
AND2X1 exu_U2616(.A(exu_n4734), .B(exu_n9540), .Y(bypass_sr_out_mux_n201));
AND2X1 exu_U2617(.A(ecc_decode_n46), .B(ecc_decode_n27), .Y(ecc_error_data_m[21]));
AND2X1 exu_U2618(.A(exu_n4735), .B(exu_n9542), .Y(bypass_sr_out_mux_n205));
AND2X1 exu_U2619(.A(ecc_decode_n46), .B(ecc_decode_n29), .Y(ecc_error_data_m[20]));
AND2X1 exu_U2620(.A(exu_n4737), .B(exu_n9546), .Y(bypass_sr_out_mux_n213));
AND2X1 exu_U2621(.A(ecc_decode_n47), .B(ecc_decode_n27), .Y(ecc_error_data_m[19]));
AND2X1 exu_U2622(.A(exu_n4738), .B(exu_n9548), .Y(bypass_sr_out_mux_n217));
AND2X1 exu_U2623(.A(ecc_decode_n47), .B(ecc_decode_n29), .Y(ecc_error_data_m[18]));
AND2X1 exu_U2624(.A(exu_n4739), .B(exu_n9550), .Y(bypass_sr_out_mux_n221));
AND2X1 exu_U2625(.A(ecc_decode_n44), .B(ecc_decode_n35), .Y(ecc_error_data_m[17]));
AND2X1 exu_U2626(.A(exu_n4740), .B(exu_n9552), .Y(bypass_sr_out_mux_n225));
AND2X1 exu_U2627(.A(ecc_decode_n44), .B(ecc_decode_n36), .Y(ecc_error_data_m[16]));
AND2X1 exu_U2628(.A(exu_n4741), .B(exu_n9554), .Y(bypass_sr_out_mux_n229));
AND2X1 exu_U2629(.A(ecc_decode_n45), .B(ecc_decode_n35), .Y(ecc_error_data_m[15]));
AND2X1 exu_U2630(.A(exu_n4742), .B(exu_n9556), .Y(bypass_sr_out_mux_n233));
AND2X1 exu_U2631(.A(ecc_decode_n45), .B(ecc_decode_n36), .Y(ecc_error_data_m[14]));
AND2X1 exu_U2632(.A(exu_n4743), .B(exu_n9558), .Y(bypass_sr_out_mux_n237));
AND2X1 exu_U2633(.A(ecc_decode_n46), .B(ecc_decode_n35), .Y(ecc_error_data_m[13]));
AND2X1 exu_U2634(.A(exu_n4744), .B(exu_n9560), .Y(bypass_sr_out_mux_n241));
AND2X1 exu_U2635(.A(ecc_decode_n46), .B(ecc_decode_n36), .Y(ecc_error_data_m[12]));
AND2X1 exu_U2636(.A(exu_n4745), .B(exu_n9562), .Y(bypass_sr_out_mux_n245));
AND2X1 exu_U2637(.A(ecc_decode_n47), .B(ecc_decode_n35), .Y(ecc_error_data_m[11]));
AND2X1 exu_U2638(.A(exu_n4746), .B(exu_n9564), .Y(bypass_sr_out_mux_n249));
AND2X1 exu_U2639(.A(ecc_decode_n27), .B(ecc_decode_n15), .Y(ecc_error_data_m[10]));
AND2X1 exu_U2640(.A(exu_n4684), .B(exu_n9440), .Y(bypass_sr_out_mux_n1));
AND2X1 exu_U2641(.A(ecc_decode_n29), .B(ecc_decode_n15), .Y(ecc_error_data_m[9]));
AND2X1 exu_U2642(.A(exu_n4685), .B(exu_n9442), .Y(bypass_sr_out_mux_n5));
AND2X1 exu_U2643(.A(ecc_decode_n27), .B(ecc_decode_n16), .Y(ecc_error_data_m[8]));
AND2X1 exu_U2644(.A(exu_n4686), .B(exu_n9444), .Y(bypass_sr_out_mux_n9));
AND2X1 exu_U2645(.A(ecc_decode_n16), .B(ecc_decode_n29), .Y(ecc_error_data_m[7]));
AND2X1 exu_U2646(.A(exu_n4687), .B(exu_n9446), .Y(bypass_sr_out_mux_n13));
AND2X1 exu_U2647(.A(ecc_decode_n17), .B(ecc_decode_n27), .Y(ecc_error_data_m[6]));
AND2X1 exu_U2648(.A(exu_n4692), .B(exu_n9456), .Y(bypass_sr_out_mux_n33));
AND2X1 exu_U2649(.A(ecc_decode_n17), .B(ecc_decode_n29), .Y(ecc_error_data_m[5]));
AND2X1 exu_U2650(.A(exu_n4703), .B(exu_n9478), .Y(bypass_sr_out_mux_n77));
AND2X1 exu_U2651(.A(exu_n4714), .B(exu_n9500), .Y(bypass_sr_out_mux_n121));
AND2X1 exu_U2652(.A(ecc_decode_n35), .B(ecc_decode_n15), .Y(ecc_error_data_m[3]));
AND2X1 exu_U2653(.A(exu_n4725), .B(exu_n9522), .Y(bypass_sr_out_mux_n165));
AND2X1 exu_U2654(.A(ecc_decode_n36), .B(ecc_decode_n15), .Y(ecc_error_data_m[2]));
AND2X1 exu_U2655(.A(exu_n4736), .B(exu_n9544), .Y(bypass_sr_out_mux_n209));
AND2X1 exu_U2656(.A(ecc_decode_n35), .B(ecc_decode_n16), .Y(ecc_error_data_m[1]));
AND2X1 exu_U2657(.A(exu_n4747), .B(exu_n9566), .Y(bypass_sr_out_mux_n253));
AND2X1 exu_U2658(.A(ecc_decode_n35), .B(ecc_decode_n17), .Y(ecc_error_data_m[0]));
INVX1 exu_U2659(.A(se), .Y(exu_n29431));
INVX1 exu_U2660(.A(se), .Y(exu_n29496));
AND2X1 exu_U2661(.A(exu_n1691), .B(exu_n6707), .Y(exu_n23610));
AND2X1 exu_U2662(.A(exu_n1691), .B(exu_n6709), .Y(exu_n23615));
AND2X1 exu_U2663(.A(exu_n1694), .B(exu_n6711), .Y(exu_n23620));
AND2X1 exu_U2664(.A(exu_n1696), .B(exu_n6714), .Y(exu_n23624));
AND2X1 exu_U2665(.A(exu_n1699), .B(exu_n6718), .Y(exu_n23635));
AND2X1 exu_U2666(.A(exu_n1700), .B(exu_n6720), .Y(exu_n23640));
AND2X1 exu_U2667(.A(exu_n1701), .B(exu_n6722), .Y(exu_n23645));
AND2X1 exu_U2668(.A(exu_n1702), .B(exu_n6724), .Y(exu_n23650));
AND2X1 exu_U2669(.A(exu_n1703), .B(exu_n6726), .Y(exu_n23655));
AND2X1 exu_U2670(.A(exu_n1704), .B(exu_n6728), .Y(exu_n23660));
AND2X1 exu_U2671(.A(exu_n1705), .B(exu_n6730), .Y(exu_n23665));
AND2X1 exu_U2672(.A(exu_n1706), .B(exu_n6732), .Y(exu_n23670));
AND2X1 exu_U2673(.A(exu_n1707), .B(exu_n6734), .Y(exu_n23675));
AND2X1 exu_U2674(.A(exu_n1708), .B(exu_n6736), .Y(exu_n23680));
AND2X1 exu_U2675(.A(exu_n1711), .B(exu_n6740), .Y(exu_n23691));
AND2X1 exu_U2676(.A(exu_n1712), .B(exu_n6742), .Y(exu_n23696));
AND2X1 exu_U2677(.A(exu_n1714), .B(exu_n6744), .Y(exu_n23701));
AND2X1 exu_U2678(.A(exu_n1715), .B(exu_n6745), .Y(exu_n23708));
AND2X1 exu_U2679(.A(exu_n1717), .B(exu_n6747), .Y(exu_n23714));
AND2X1 exu_U2680(.A(exu_n1719), .B(exu_n6749), .Y(exu_n23720));
AND2X1 exu_U2681(.A(exu_n1721), .B(exu_n6751), .Y(exu_n23726));
AND2X1 exu_U2682(.A(exu_n1723), .B(exu_n6753), .Y(exu_n23732));
AND2X1 exu_U2683(.A(exu_n1725), .B(exu_n6755), .Y(exu_n23738));
AND2X1 exu_U2684(.A(exu_n1727), .B(exu_n6757), .Y(exu_n23744));
AND2X1 exu_U2685(.A(exu_n1731), .B(exu_n6761), .Y(exu_n23756));
AND2X1 exu_U2686(.A(exu_n1733), .B(exu_n6763), .Y(exu_n23762));
AND2X1 exu_U2687(.A(exu_n1735), .B(exu_n6765), .Y(exu_n23768));
AND2X1 exu_U2688(.A(exu_n1737), .B(exu_n6767), .Y(exu_n23774));
AND2X1 exu_U2689(.A(exu_n1739), .B(exu_n6769), .Y(exu_n23780));
AND2X1 exu_U2690(.A(exu_n1741), .B(exu_n6771), .Y(exu_n23786));
AND2X1 exu_U2691(.A(exu_n1743), .B(exu_n6773), .Y(exu_n23792));
AND2X1 exu_U2692(.A(exu_n1745), .B(exu_n6775), .Y(exu_n23798));
AND2X1 exu_U2693(.A(exu_n1747), .B(exu_n6777), .Y(exu_n23804));
AND2X1 exu_U2694(.A(exu_n1749), .B(exu_n6779), .Y(exu_n23810));
AND2X1 exu_U2695(.A(exu_n1753), .B(exu_n6783), .Y(exu_n23822));
AND2X1 exu_U2696(.A(exu_n1755), .B(exu_n6785), .Y(exu_n23828));
AND2X1 exu_U2697(.A(exu_n1757), .B(exu_n6787), .Y(exu_n23834));
AND2X1 exu_U2698(.A(exu_n1759), .B(exu_n6789), .Y(exu_n23840));
AND2X1 exu_U2699(.A(exu_n1761), .B(exu_n6791), .Y(exu_n23846));
AND2X1 exu_U2700(.A(exu_n1763), .B(exu_n6793), .Y(exu_n23852));
AND2X1 exu_U2701(.A(exu_n1765), .B(exu_n6795), .Y(exu_n23858));
AND2X1 exu_U2702(.A(exu_n1767), .B(exu_n6797), .Y(exu_n23864));
AND2X1 exu_U2703(.A(exu_n1769), .B(exu_n6799), .Y(exu_n23870));
AND2X1 exu_U2704(.A(exu_n1771), .B(exu_n6801), .Y(exu_n23876));
AND2X1 exu_U2705(.A(exu_n1775), .B(exu_n6805), .Y(exu_n23888));
AND2X1 exu_U2706(.A(exu_n1777), .B(exu_n6807), .Y(exu_n23894));
AND2X1 exu_U2707(.A(exu_n1779), .B(exu_n6809), .Y(exu_n23900));
AND2X1 exu_U2708(.A(exu_n1781), .B(exu_n6811), .Y(exu_n23906));
AND2X1 exu_U2709(.A(exu_n1783), .B(exu_n6813), .Y(exu_n23912));
AND2X1 exu_U2710(.A(exu_n1785), .B(exu_n6815), .Y(exu_n23918));
AND2X1 exu_U2711(.A(exu_n1787), .B(exu_n6817), .Y(exu_n23924));
AND2X1 exu_U2712(.A(exu_n1789), .B(exu_n6819), .Y(exu_n23930));
AND2X1 exu_U2713(.A(exu_n1791), .B(exu_n6821), .Y(exu_n23936));
AND2X1 exu_U2714(.A(exu_n1793), .B(exu_n6823), .Y(exu_n23942));
AND2X1 exu_U2715(.A(exu_n1681), .B(exu_n6699), .Y(exu_n23586));
AND2X1 exu_U2716(.A(exu_n1682), .B(exu_n6700), .Y(exu_n23585));
AND2X1 exu_U2717(.A(exu_n1683), .B(exu_n6701), .Y(exu_n23592));
AND2X1 exu_U2718(.A(exu_n1685), .B(exu_n6703), .Y(exu_n23598));
AND2X1 exu_U2719(.A(exu_n1687), .B(exu_n6705), .Y(exu_n23604));
AND2X1 exu_U2720(.A(exu_n1697), .B(exu_n6715), .Y(exu_n23630));
AND2X1 exu_U2721(.A(exu_n1709), .B(exu_n6737), .Y(exu_n23686));
AND2X1 exu_U2722(.A(exu_n1729), .B(exu_n6759), .Y(exu_n23750));
AND2X1 exu_U2723(.A(exu_n1751), .B(exu_n6781), .Y(exu_n23816));
AND2X1 exu_U2724(.A(exu_n1773), .B(exu_n6803), .Y(exu_n23882));
INVX1 exu_U2725(.A(ifu_exu_dbrinst_d), .Y(exu_n16395));
AND2X1 exu_U2726(.A(exu_n1795), .B(exu_n6825), .Y(exu_n23948));
INVX1 exu_U2727(.A(se), .Y(exu_n29561));
AND2X1 exu_U2728(.A(exu_n2127), .B(exu_n7155), .Y(exu_n25002));
AND2X1 exu_U2729(.A(exu_n2127), .B(exu_n7157), .Y(exu_n25007));
AND2X1 exu_U2730(.A(exu_n2130), .B(exu_n7159), .Y(exu_n25012));
AND2X1 exu_U2731(.A(exu_n2133), .B(exu_n7161), .Y(exu_n25017));
AND2X1 exu_U2732(.A(exu_n2138), .B(exu_n7165), .Y(exu_n25028));
AND2X1 exu_U2733(.A(exu_n2141), .B(exu_n7167), .Y(exu_n25033));
AND2X1 exu_U2734(.A(exu_n2144), .B(exu_n7169), .Y(exu_n25038));
AND2X1 exu_U2735(.A(exu_n2147), .B(exu_n7171), .Y(exu_n25043));
AND2X1 exu_U2736(.A(exu_n2150), .B(exu_n7173), .Y(exu_n25048));
AND2X1 exu_U2737(.A(exu_n2153), .B(exu_n7175), .Y(exu_n25053));
AND2X1 exu_U2738(.A(exu_n2156), .B(exu_n7177), .Y(exu_n25058));
AND2X1 exu_U2739(.A(exu_n2159), .B(exu_n7179), .Y(exu_n25063));
AND2X1 exu_U2740(.A(exu_n2162), .B(exu_n7181), .Y(exu_n25068));
AND2X1 exu_U2741(.A(exu_n2165), .B(exu_n7183), .Y(exu_n25073));
AND2X1 exu_U2742(.A(exu_n2170), .B(exu_n7187), .Y(exu_n25084));
AND2X1 exu_U2743(.A(exu_n2173), .B(exu_n7189), .Y(exu_n25089));
AND2X1 exu_U2744(.A(exu_n2176), .B(exu_n7191), .Y(exu_n25094));
AND2X1 exu_U2745(.A(exu_n2179), .B(exu_n7193), .Y(exu_n25099));
AND2X1 exu_U2746(.A(exu_n22145), .B(exu_n6106), .Y(bypass_rs2_data_w2[45]));
AND2X1 exu_U2747(.A(exu_n2181), .B(exu_n7196), .Y(exu_n25103));
AND2X1 exu_U2748(.A(exu_n22149), .B(exu_n6108), .Y(bypass_rs2_data_w2[44]));
AND2X1 exu_U2749(.A(exu_n2182), .B(exu_n7198), .Y(exu_n25108));
AND2X1 exu_U2750(.A(exu_n22153), .B(exu_n6110), .Y(bypass_rs2_data_w2[43]));
AND2X1 exu_U2751(.A(exu_n2183), .B(exu_n7200), .Y(exu_n25113));
AND2X1 exu_U2752(.A(exu_n22157), .B(exu_n6112), .Y(bypass_rs2_data_w2[42]));
AND2X1 exu_U2753(.A(exu_n2184), .B(exu_n7202), .Y(exu_n25118));
AND2X1 exu_U2754(.A(exu_n22161), .B(exu_n6114), .Y(bypass_rs2_data_w2[41]));
AND2X1 exu_U2755(.A(exu_n2185), .B(exu_n7204), .Y(exu_n25123));
AND2X1 exu_U2756(.A(exu_n22165), .B(exu_n6116), .Y(bypass_rs2_data_w2[40]));
AND2X1 exu_U2757(.A(exu_n2186), .B(exu_n7206), .Y(exu_n25128));
AND2X1 exu_U2758(.A(exu_n22173), .B(exu_n6120), .Y(bypass_rs2_data_w2[39]));
AND2X1 exu_U2759(.A(exu_n2189), .B(exu_n7210), .Y(exu_n25139));
AND2X1 exu_U2760(.A(exu_n22177), .B(exu_n6122), .Y(bypass_rs2_data_w2[38]));
AND2X1 exu_U2761(.A(exu_n2190), .B(exu_n7212), .Y(exu_n25144));
AND2X1 exu_U2762(.A(exu_n22181), .B(exu_n6124), .Y(bypass_rs2_data_w2[37]));
AND2X1 exu_U2763(.A(exu_n2191), .B(exu_n7214), .Y(exu_n25149));
AND2X1 exu_U2764(.A(exu_n22185), .B(exu_n6126), .Y(bypass_rs2_data_w2[36]));
AND2X1 exu_U2765(.A(exu_n2192), .B(exu_n7216), .Y(exu_n25154));
AND2X1 exu_U2766(.A(exu_n22189), .B(exu_n6128), .Y(bypass_rs2_data_w2[35]));
AND2X1 exu_U2767(.A(exu_n2193), .B(exu_n7218), .Y(exu_n25159));
AND2X1 exu_U2768(.A(exu_n22193), .B(exu_n6130), .Y(bypass_rs2_data_w2[34]));
AND2X1 exu_U2769(.A(exu_n2194), .B(exu_n7220), .Y(exu_n25164));
AND2X1 exu_U2770(.A(exu_n22197), .B(exu_n6132), .Y(bypass_rs2_data_w2[33]));
AND2X1 exu_U2771(.A(exu_n2195), .B(exu_n7222), .Y(exu_n25169));
AND2X1 exu_U2772(.A(exu_n22201), .B(exu_n6134), .Y(bypass_rs2_data_w2[32]));
AND2X1 exu_U2773(.A(exu_n2196), .B(exu_n7224), .Y(exu_n25174));
AND2X1 exu_U2774(.A(exu_n22205), .B(exu_n6136), .Y(bypass_rs2_data_w2[31]));
AND2X1 exu_U2775(.A(exu_n2198), .B(exu_n7226), .Y(exu_n25179));
AND2X1 exu_U2776(.A(exu_n2199), .B(exu_n7227), .Y(exu_n25186));
AND2X1 exu_U2777(.A(exu_n2203), .B(exu_n7231), .Y(exu_n25198));
AND2X1 exu_U2778(.A(exu_n2205), .B(exu_n7233), .Y(exu_n25204));
AND2X1 exu_U2779(.A(exu_n2207), .B(exu_n7235), .Y(exu_n25210));
AND2X1 exu_U2780(.A(exu_n2209), .B(exu_n7237), .Y(exu_n25216));
AND2X1 exu_U2781(.A(exu_n2211), .B(exu_n7239), .Y(exu_n25222));
AND2X1 exu_U2782(.A(exu_n2213), .B(exu_n7241), .Y(exu_n25228));
AND2X1 exu_U2783(.A(exu_n2215), .B(exu_n7243), .Y(exu_n25234));
AND2X1 exu_U2784(.A(exu_n2217), .B(exu_n7245), .Y(exu_n25240));
AND2X1 exu_U2785(.A(exu_n2219), .B(exu_n7247), .Y(exu_n25246));
AND2X1 exu_U2786(.A(exu_n2221), .B(exu_n7249), .Y(exu_n25252));
AND2X1 exu_U2787(.A(exu_n2225), .B(exu_n7253), .Y(exu_n25264));
AND2X1 exu_U2788(.A(exu_n2227), .B(exu_n7255), .Y(exu_n25270));
AND2X1 exu_U2789(.A(exu_n2229), .B(exu_n7257), .Y(exu_n25276));
AND2X1 exu_U2790(.A(exu_n2231), .B(exu_n7259), .Y(exu_n25282));
AND2X1 exu_U2791(.A(exu_n2233), .B(exu_n7261), .Y(exu_n25288));
AND2X1 exu_U2792(.A(exu_n2235), .B(exu_n7263), .Y(exu_n25294));
AND2X1 exu_U2793(.A(exu_n2237), .B(exu_n7265), .Y(exu_n25300));
AND2X1 exu_U2794(.A(exu_n2239), .B(exu_n7267), .Y(exu_n25306));
AND2X1 exu_U2795(.A(exu_n2241), .B(exu_n7269), .Y(exu_n25312));
AND2X1 exu_U2796(.A(exu_n2243), .B(exu_n7271), .Y(exu_n25318));
AND2X1 exu_U2797(.A(exu_n2117), .B(exu_n7147), .Y(exu_n24978));
AND2X1 exu_U2798(.A(exu_n2118), .B(exu_n7148), .Y(exu_n24977));
AND2X1 exu_U2799(.A(exu_n2119), .B(exu_n7149), .Y(exu_n24984));
AND2X1 exu_U2800(.A(exu_n2121), .B(exu_n7151), .Y(exu_n24990));
AND2X1 exu_U2801(.A(exu_n2123), .B(exu_n7153), .Y(exu_n24996));
AND2X1 exu_U2802(.A(exu_n2135), .B(exu_n7163), .Y(exu_n25022));
AND2X1 exu_U2803(.A(exu_n2167), .B(exu_n7185), .Y(exu_n25078));
AND2X1 exu_U2804(.A(exu_n2187), .B(exu_n7207), .Y(exu_n25134));
AND2X1 exu_U2805(.A(exu_n2201), .B(exu_n7229), .Y(exu_n25192));
AND2X1 exu_U2806(.A(exu_n2223), .B(exu_n7251), .Y(exu_n25258));
OR2X1 exu_U2807(.A(exu_n13435), .B(exu_n14758), .Y(ecl_byplog_rs2_n21));
AND2X1 exu_U2808(.A(ecl_byplog_rs2_n23), .B(ecl_byplog_rs2_n24), .Y(ecl_byplog_rs2_n19));
AND2X1 exu_U2809(.A(exu_n15435), .B(exu_n15423), .Y(ecl_byplog_rs2_n23));
OR2X1 exu_U2810(.A(exu_n13437), .B(exu_n14760), .Y(ecl_byplog_rs2_n15));
AND2X1 exu_U2811(.A(exu_n21), .B(exu_n16389), .Y(ecl_byplog_rs2_n44));
AND2X1 exu_U2812(.A(exu_n2245), .B(exu_n7273), .Y(exu_n25324));
INVX1 exu_U2813(.A(se), .Y(exu_n29626));
AND2X1 exu_U2814(.A(exu_n1306), .B(exu_n6191), .Y(exu_n22321));
AND2X1 exu_U2815(.A(exu_n2379), .B(exu_n7407), .Y(exu_n25729));
AND2X1 exu_U2816(.A(exu_n1308), .B(exu_n6192), .Y(exu_n22325));
AND2X1 exu_U2817(.A(exu_n2380), .B(exu_n7408), .Y(exu_n25733));
AND2X1 exu_U2818(.A(exu_n1310), .B(exu_n6193), .Y(exu_n22329));
AND2X1 exu_U2819(.A(exu_n2381), .B(exu_n7409), .Y(exu_n25737));
AND2X1 exu_U2820(.A(exu_n1312), .B(exu_n6194), .Y(exu_n22333));
AND2X1 exu_U2821(.A(exu_n2382), .B(exu_n7410), .Y(exu_n25741));
AND2X1 exu_U2822(.A(exu_n1316), .B(exu_n6196), .Y(exu_n22341));
AND2X1 exu_U2823(.A(exu_n2384), .B(exu_n7412), .Y(exu_n25749));
AND2X1 exu_U2824(.A(exu_n1318), .B(exu_n6197), .Y(exu_n22345));
AND2X1 exu_U2825(.A(exu_n2385), .B(exu_n7413), .Y(exu_n25753));
AND2X1 exu_U2826(.A(exu_n1320), .B(exu_n6198), .Y(exu_n22349));
AND2X1 exu_U2827(.A(exu_n2386), .B(exu_n7414), .Y(exu_n25757));
AND2X1 exu_U2828(.A(exu_n1322), .B(exu_n6199), .Y(exu_n22353));
AND2X1 exu_U2829(.A(exu_n2387), .B(exu_n7415), .Y(exu_n25761));
AND2X1 exu_U2830(.A(exu_n1324), .B(exu_n6200), .Y(exu_n22357));
AND2X1 exu_U2831(.A(exu_n2388), .B(exu_n7416), .Y(exu_n25765));
AND2X1 exu_U2832(.A(exu_n1326), .B(exu_n6201), .Y(exu_n22361));
AND2X1 exu_U2833(.A(exu_n2389), .B(exu_n7417), .Y(exu_n25769));
AND2X1 exu_U2834(.A(exu_n1328), .B(exu_n6202), .Y(exu_n22365));
AND2X1 exu_U2835(.A(exu_n2390), .B(exu_n7418), .Y(exu_n25773));
AND2X1 exu_U2836(.A(exu_n1330), .B(exu_n6203), .Y(exu_n22369));
AND2X1 exu_U2837(.A(exu_n2391), .B(exu_n7419), .Y(exu_n25777));
AND2X1 exu_U2838(.A(exu_n1332), .B(exu_n6204), .Y(exu_n22373));
AND2X1 exu_U2839(.A(exu_n2392), .B(exu_n7420), .Y(exu_n25781));
AND2X1 exu_U2840(.A(exu_n1334), .B(exu_n6205), .Y(exu_n22377));
AND2X1 exu_U2841(.A(exu_n2393), .B(exu_n7421), .Y(exu_n25785));
AND2X1 exu_U2842(.A(exu_n1338), .B(exu_n6207), .Y(exu_n22385));
AND2X1 exu_U2843(.A(exu_n2395), .B(exu_n7423), .Y(exu_n25793));
AND2X1 exu_U2844(.A(exu_n1340), .B(exu_n6208), .Y(exu_n22389));
AND2X1 exu_U2845(.A(exu_n2396), .B(exu_n7424), .Y(exu_n25797));
AND2X1 exu_U2846(.A(exu_n1342), .B(exu_n6209), .Y(exu_n22393));
AND2X1 exu_U2847(.A(exu_n2397), .B(exu_n7425), .Y(exu_n25801));
AND2X1 exu_U2848(.A(exu_n1344), .B(exu_n6210), .Y(exu_n22397));
AND2X1 exu_U2849(.A(exu_n2398), .B(exu_n7426), .Y(exu_n25805));
AND2X1 exu_U2850(.A(exu_n1346), .B(exu_n6211), .Y(exu_n22401));
AND2X1 exu_U2851(.A(exu_n2399), .B(exu_n7427), .Y(exu_n25809));
AND2X1 exu_U2852(.A(exu_n1348), .B(exu_n6212), .Y(exu_n22405));
AND2X1 exu_U2853(.A(exu_n2400), .B(exu_n7428), .Y(exu_n25813));
AND2X1 exu_U2854(.A(exu_n1350), .B(exu_n6213), .Y(exu_n22409));
AND2X1 exu_U2855(.A(exu_n2401), .B(exu_n7429), .Y(exu_n25817));
AND2X1 exu_U2856(.A(exu_n1352), .B(exu_n6214), .Y(exu_n22413));
AND2X1 exu_U2857(.A(exu_n2402), .B(exu_n7430), .Y(exu_n25821));
AND2X1 exu_U2858(.A(exu_n1354), .B(exu_n6215), .Y(exu_n22417));
AND2X1 exu_U2859(.A(exu_n2403), .B(exu_n7431), .Y(exu_n25825));
AND2X1 exu_U2860(.A(exu_n1356), .B(exu_n6216), .Y(exu_n22421));
AND2X1 exu_U2861(.A(exu_n2404), .B(exu_n7432), .Y(exu_n25829));
AND2X1 exu_U2862(.A(exu_n1360), .B(exu_n6218), .Y(exu_n22429));
AND2X1 exu_U2863(.A(exu_n2406), .B(exu_n7434), .Y(exu_n25837));
AND2X1 exu_U2864(.A(exu_n1362), .B(exu_n6219), .Y(exu_n22433));
AND2X1 exu_U2865(.A(exu_n2407), .B(exu_n7435), .Y(exu_n25841));
AND2X1 exu_U2866(.A(exu_n1364), .B(exu_n6220), .Y(exu_n22437));
AND2X1 exu_U2867(.A(exu_n2408), .B(exu_n7436), .Y(exu_n25845));
AND2X1 exu_U2868(.A(exu_n1366), .B(exu_n6221), .Y(exu_n22441));
AND2X1 exu_U2869(.A(exu_n2409), .B(exu_n7437), .Y(exu_n25849));
AND2X1 exu_U2870(.A(exu_n1368), .B(exu_n6222), .Y(exu_n22445));
AND2X1 exu_U2871(.A(exu_n2410), .B(exu_n7438), .Y(exu_n25853));
AND2X1 exu_U2872(.A(exu_n1370), .B(exu_n6223), .Y(exu_n22449));
AND2X1 exu_U2873(.A(exu_n2411), .B(exu_n7439), .Y(exu_n25857));
AND2X1 exu_U2874(.A(exu_n1372), .B(exu_n6224), .Y(exu_n22453));
AND2X1 exu_U2875(.A(exu_n2412), .B(exu_n7440), .Y(exu_n25861));
AND2X1 exu_U2876(.A(exu_n1374), .B(exu_n6225), .Y(exu_n22457));
AND2X1 exu_U2877(.A(exu_n2413), .B(exu_n7441), .Y(exu_n25865));
AND2X1 exu_U2878(.A(exu_n1376), .B(exu_n6226), .Y(exu_n22461));
AND2X1 exu_U2879(.A(exu_n2414), .B(exu_n7442), .Y(exu_n25869));
AND2X1 exu_U2880(.A(exu_n1378), .B(exu_n6227), .Y(exu_n22465));
AND2X1 exu_U2881(.A(exu_n2415), .B(exu_n7443), .Y(exu_n25873));
AND2X1 exu_U2882(.A(exu_n1382), .B(exu_n6229), .Y(exu_n22473));
AND2X1 exu_U2883(.A(exu_n2417), .B(exu_n7445), .Y(exu_n25881));
AND2X1 exu_U2884(.A(exu_n1384), .B(exu_n6230), .Y(exu_n22477));
AND2X1 exu_U2885(.A(exu_n2418), .B(exu_n7446), .Y(exu_n25885));
AND2X1 exu_U2886(.A(exu_n1386), .B(exu_n6231), .Y(exu_n22481));
AND2X1 exu_U2887(.A(exu_n2419), .B(exu_n7447), .Y(exu_n25889));
AND2X1 exu_U2888(.A(exu_n1388), .B(exu_n6232), .Y(exu_n22485));
AND2X1 exu_U2889(.A(exu_n2420), .B(exu_n7448), .Y(exu_n25893));
AND2X1 exu_U2890(.A(exu_n1390), .B(exu_n6233), .Y(exu_n22489));
AND2X1 exu_U2891(.A(exu_n2421), .B(exu_n7449), .Y(exu_n25897));
AND2X1 exu_U2892(.A(exu_n1392), .B(exu_n6234), .Y(exu_n22493));
AND2X1 exu_U2893(.A(exu_n2422), .B(exu_n7450), .Y(exu_n25901));
AND2X1 exu_U2894(.A(exu_n1394), .B(exu_n6235), .Y(exu_n22497));
AND2X1 exu_U2895(.A(exu_n2423), .B(exu_n7451), .Y(exu_n25905));
AND2X1 exu_U2896(.A(exu_n1396), .B(exu_n6236), .Y(exu_n22501));
AND2X1 exu_U2897(.A(exu_n2424), .B(exu_n7452), .Y(exu_n25909));
AND2X1 exu_U2898(.A(exu_n1398), .B(exu_n6237), .Y(exu_n22505));
AND2X1 exu_U2899(.A(exu_n2425), .B(exu_n7453), .Y(exu_n25913));
AND2X1 exu_U2900(.A(exu_n1400), .B(exu_n6238), .Y(exu_n22509));
AND2X1 exu_U2901(.A(exu_n2426), .B(exu_n7454), .Y(exu_n25917));
AND2X1 exu_U2902(.A(exu_n1404), .B(exu_n6240), .Y(exu_n22517));
AND2X1 exu_U2903(.A(exu_n2428), .B(exu_n7456), .Y(exu_n25925));
AND2X1 exu_U2904(.A(exu_n1406), .B(exu_n6241), .Y(exu_n22521));
AND2X1 exu_U2905(.A(exu_n2429), .B(exu_n7457), .Y(exu_n25929));
AND2X1 exu_U2906(.A(exu_n1408), .B(exu_n6242), .Y(exu_n22525));
AND2X1 exu_U2907(.A(exu_n2430), .B(exu_n7458), .Y(exu_n25933));
AND2X1 exu_U2908(.A(exu_n1410), .B(exu_n6243), .Y(exu_n22529));
AND2X1 exu_U2909(.A(exu_n2431), .B(exu_n7459), .Y(exu_n25937));
AND2X1 exu_U2910(.A(exu_n1412), .B(exu_n6244), .Y(exu_n22533));
AND2X1 exu_U2911(.A(exu_n2432), .B(exu_n7460), .Y(exu_n25941));
AND2X1 exu_U2912(.A(exu_n1414), .B(exu_n6245), .Y(exu_n22537));
AND2X1 exu_U2913(.A(exu_n2433), .B(exu_n7461), .Y(exu_n25945));
AND2X1 exu_U2914(.A(exu_n1416), .B(exu_n6246), .Y(exu_n22541));
AND2X1 exu_U2915(.A(exu_n2434), .B(exu_n7462), .Y(exu_n25949));
AND2X1 exu_U2916(.A(exu_n1418), .B(exu_n6247), .Y(exu_n22545));
AND2X1 exu_U2917(.A(exu_n2435), .B(exu_n7463), .Y(exu_n25953));
AND2X1 exu_U2918(.A(exu_n1420), .B(exu_n6248), .Y(exu_n22549));
AND2X1 exu_U2919(.A(exu_n2436), .B(exu_n7464), .Y(exu_n25957));
AND2X1 exu_U2920(.A(exu_n1422), .B(exu_n6249), .Y(exu_n22553));
AND2X1 exu_U2921(.A(exu_n2437), .B(exu_n7465), .Y(exu_n25961));
AND2X1 exu_U2922(.A(exu_n1298), .B(exu_n6187), .Y(exu_n22305));
AND2X1 exu_U2923(.A(exu_n2375), .B(exu_n7403), .Y(exu_n25713));
AND2X1 exu_U2924(.A(exu_n1300), .B(exu_n6188), .Y(exu_n22309));
AND2X1 exu_U2925(.A(exu_n2376), .B(exu_n7404), .Y(exu_n25717));
AND2X1 exu_U2926(.A(exu_n1302), .B(exu_n6189), .Y(exu_n22313));
AND2X1 exu_U2927(.A(exu_n2377), .B(exu_n7405), .Y(exu_n25721));
AND2X1 exu_U2928(.A(exu_n1304), .B(exu_n6190), .Y(exu_n22317));
AND2X1 exu_U2929(.A(exu_n2378), .B(exu_n7406), .Y(exu_n25725));
AND2X1 exu_U2930(.A(exu_n1314), .B(exu_n6195), .Y(exu_n22337));
AND2X1 exu_U2931(.A(exu_n2383), .B(exu_n7411), .Y(exu_n25745));
AND2X1 exu_U2932(.A(exu_n1336), .B(exu_n6206), .Y(exu_n22381));
AND2X1 exu_U2933(.A(exu_n2394), .B(exu_n7422), .Y(exu_n25789));
AND2X1 exu_U2934(.A(exu_n1358), .B(exu_n6217), .Y(exu_n22425));
AND2X1 exu_U2935(.A(exu_n2405), .B(exu_n7433), .Y(exu_n25833));
AND2X1 exu_U2936(.A(exu_n1380), .B(exu_n6228), .Y(exu_n22469));
AND2X1 exu_U2937(.A(exu_n2416), .B(exu_n7444), .Y(exu_n25877));
AND2X1 exu_U2938(.A(exu_n1402), .B(exu_n6239), .Y(exu_n22513));
AND2X1 exu_U2939(.A(exu_n2427), .B(exu_n7455), .Y(exu_n25921));
OR2X1 exu_U2940(.A(exu_n12140), .B(exu_n14758), .Y(exu_n19192));
AND2X1 exu_U2941(.A(exu_n1424), .B(exu_n6250), .Y(exu_n22557));
AND2X1 exu_U2942(.A(exu_n2438), .B(exu_n7466), .Y(exu_n25965));
INVX1 exu_U2943(.A(se), .Y(exu_n29691));
AND2X1 exu_U2944(.A(exu_n21809), .B(exu_n5939), .Y(bypass_rs1_data_w2[63]));
AND2X1 exu_U2945(.A(exu_n1174), .B(exu_n5940), .Y(exu_n21809));
AND2X1 exu_U2946(.A(exu_n1929), .B(exu_n6959), .Y(exu_n24353));
AND2X1 exu_U2947(.A(exu_n21813), .B(exu_n5941), .Y(bypass_rs1_data_w2[62]));
AND2X1 exu_U2948(.A(exu_n1175), .B(exu_n5942), .Y(exu_n21813));
AND2X1 exu_U2949(.A(exu_n1930), .B(exu_n6960), .Y(exu_n24357));
AND2X1 exu_U2950(.A(exu_n21817), .B(exu_n5943), .Y(bypass_rs1_data_w2[61]));
AND2X1 exu_U2951(.A(exu_n1176), .B(exu_n5944), .Y(exu_n21817));
AND2X1 exu_U2952(.A(exu_n1931), .B(exu_n6961), .Y(exu_n24361));
AND2X1 exu_U2953(.A(exu_n21821), .B(exu_n5945), .Y(bypass_rs1_data_w2[60]));
AND2X1 exu_U2954(.A(exu_n1177), .B(exu_n5946), .Y(exu_n21821));
AND2X1 exu_U2955(.A(exu_n1932), .B(exu_n6962), .Y(exu_n24365));
AND2X1 exu_U2956(.A(exu_n21829), .B(exu_n5949), .Y(bypass_rs1_data_w2[59]));
AND2X1 exu_U2957(.A(exu_n1179), .B(exu_n5950), .Y(exu_n21829));
AND2X1 exu_U2958(.A(exu_n1934), .B(exu_n6964), .Y(exu_n24373));
AND2X1 exu_U2959(.A(exu_n21833), .B(exu_n5951), .Y(bypass_rs1_data_w2[58]));
AND2X1 exu_U2960(.A(exu_n1180), .B(exu_n5952), .Y(exu_n21833));
AND2X1 exu_U2961(.A(exu_n1935), .B(exu_n6965), .Y(exu_n24377));
AND2X1 exu_U2962(.A(exu_n21837), .B(exu_n5953), .Y(bypass_rs1_data_w2[57]));
AND2X1 exu_U2963(.A(exu_n1181), .B(exu_n5954), .Y(exu_n21837));
AND2X1 exu_U2964(.A(exu_n1936), .B(exu_n6966), .Y(exu_n24381));
AND2X1 exu_U2965(.A(exu_n21841), .B(exu_n5955), .Y(bypass_rs1_data_w2[56]));
AND2X1 exu_U2966(.A(exu_n1182), .B(exu_n5956), .Y(exu_n21841));
AND2X1 exu_U2967(.A(exu_n1937), .B(exu_n6967), .Y(exu_n24385));
AND2X1 exu_U2968(.A(exu_n21845), .B(exu_n5957), .Y(bypass_rs1_data_w2[55]));
AND2X1 exu_U2969(.A(exu_n1183), .B(exu_n5958), .Y(exu_n21845));
AND2X1 exu_U2970(.A(exu_n1938), .B(exu_n6968), .Y(exu_n24389));
AND2X1 exu_U2971(.A(exu_n21849), .B(exu_n5959), .Y(bypass_rs1_data_w2[54]));
AND2X1 exu_U2972(.A(exu_n1184), .B(exu_n5960), .Y(exu_n21849));
AND2X1 exu_U2973(.A(exu_n1939), .B(exu_n6969), .Y(exu_n24393));
AND2X1 exu_U2974(.A(exu_n21853), .B(exu_n5961), .Y(bypass_rs1_data_w2[53]));
AND2X1 exu_U2975(.A(exu_n1185), .B(exu_n5962), .Y(exu_n21853));
AND2X1 exu_U2976(.A(exu_n1940), .B(exu_n6970), .Y(exu_n24397));
AND2X1 exu_U2977(.A(exu_n21857), .B(exu_n5963), .Y(bypass_rs1_data_w2[52]));
AND2X1 exu_U2978(.A(exu_n1186), .B(exu_n5964), .Y(exu_n21857));
AND2X1 exu_U2979(.A(exu_n1941), .B(exu_n6971), .Y(exu_n24401));
AND2X1 exu_U2980(.A(exu_n21861), .B(exu_n5965), .Y(bypass_rs1_data_w2[51]));
AND2X1 exu_U2981(.A(exu_n1187), .B(exu_n5966), .Y(exu_n21861));
AND2X1 exu_U2982(.A(exu_n1942), .B(exu_n6972), .Y(exu_n24405));
AND2X1 exu_U2983(.A(exu_n21865), .B(exu_n5967), .Y(bypass_rs1_data_w2[50]));
AND2X1 exu_U2984(.A(exu_n1188), .B(exu_n5968), .Y(exu_n21865));
AND2X1 exu_U2985(.A(exu_n1943), .B(exu_n6973), .Y(exu_n24409));
AND2X1 exu_U2986(.A(exu_n21873), .B(exu_n5971), .Y(bypass_rs1_data_w2[49]));
AND2X1 exu_U2987(.A(exu_n1190), .B(exu_n5972), .Y(exu_n21873));
AND2X1 exu_U2988(.A(exu_n1945), .B(exu_n6975), .Y(exu_n24417));
AND2X1 exu_U2989(.A(exu_n21877), .B(exu_n5973), .Y(bypass_rs1_data_w2[48]));
AND2X1 exu_U2990(.A(exu_n1191), .B(exu_n5974), .Y(exu_n21877));
AND2X1 exu_U2991(.A(exu_n1946), .B(exu_n6976), .Y(exu_n24421));
AND2X1 exu_U2992(.A(exu_n21881), .B(exu_n5975), .Y(bypass_rs1_data_w2[47]));
AND2X1 exu_U2993(.A(exu_n1192), .B(exu_n5976), .Y(exu_n21881));
AND2X1 exu_U2994(.A(exu_n1947), .B(exu_n6977), .Y(exu_n24425));
AND2X1 exu_U2995(.A(exu_n21885), .B(exu_n5977), .Y(bypass_rs1_data_w2[46]));
AND2X1 exu_U2996(.A(exu_n1193), .B(exu_n5978), .Y(exu_n21885));
AND2X1 exu_U2997(.A(exu_n1948), .B(exu_n6978), .Y(exu_n24429));
AND2X1 exu_U2998(.A(exu_n21889), .B(exu_n5979), .Y(bypass_rs1_data_w2[45]));
AND2X1 exu_U2999(.A(exu_n1194), .B(exu_n5980), .Y(exu_n21889));
AND2X1 exu_U3000(.A(exu_n1949), .B(exu_n6979), .Y(exu_n24433));
AND2X1 exu_U3001(.A(exu_n21893), .B(exu_n5981), .Y(bypass_rs1_data_w2[44]));
AND2X1 exu_U3002(.A(exu_n1195), .B(exu_n5982), .Y(exu_n21893));
AND2X1 exu_U3003(.A(exu_n1950), .B(exu_n6980), .Y(exu_n24437));
AND2X1 exu_U3004(.A(exu_n21897), .B(exu_n5983), .Y(bypass_rs1_data_w2[43]));
AND2X1 exu_U3005(.A(exu_n1196), .B(exu_n5984), .Y(exu_n21897));
AND2X1 exu_U3006(.A(exu_n1951), .B(exu_n6981), .Y(exu_n24441));
AND2X1 exu_U3007(.A(exu_n21901), .B(exu_n5985), .Y(bypass_rs1_data_w2[42]));
AND2X1 exu_U3008(.A(exu_n1197), .B(exu_n5986), .Y(exu_n21901));
AND2X1 exu_U3009(.A(exu_n1952), .B(exu_n6982), .Y(exu_n24445));
AND2X1 exu_U3010(.A(exu_n21905), .B(exu_n5987), .Y(bypass_rs1_data_w2[41]));
AND2X1 exu_U3011(.A(exu_n1198), .B(exu_n5988), .Y(exu_n21905));
AND2X1 exu_U3012(.A(exu_n1953), .B(exu_n6983), .Y(exu_n24449));
AND2X1 exu_U3013(.A(exu_n21909), .B(exu_n5989), .Y(bypass_rs1_data_w2[40]));
AND2X1 exu_U3014(.A(exu_n1199), .B(exu_n5990), .Y(exu_n21909));
AND2X1 exu_U3015(.A(exu_n1954), .B(exu_n6984), .Y(exu_n24453));
AND2X1 exu_U3016(.A(exu_n21917), .B(exu_n5993), .Y(bypass_rs1_data_w2[39]));
AND2X1 exu_U3017(.A(exu_n1201), .B(exu_n5994), .Y(exu_n21917));
AND2X1 exu_U3018(.A(exu_n1956), .B(exu_n6986), .Y(exu_n24461));
AND2X1 exu_U3019(.A(exu_n21921), .B(exu_n5995), .Y(bypass_rs1_data_w2[38]));
AND2X1 exu_U3020(.A(exu_n1202), .B(exu_n5996), .Y(exu_n21921));
AND2X1 exu_U3021(.A(exu_n1957), .B(exu_n6987), .Y(exu_n24465));
AND2X1 exu_U3022(.A(exu_n21925), .B(exu_n5997), .Y(bypass_rs1_data_w2[37]));
AND2X1 exu_U3023(.A(exu_n1203), .B(exu_n5998), .Y(exu_n21925));
AND2X1 exu_U3024(.A(exu_n1958), .B(exu_n6988), .Y(exu_n24469));
AND2X1 exu_U3025(.A(exu_n21929), .B(exu_n5999), .Y(bypass_rs1_data_w2[36]));
AND2X1 exu_U3026(.A(exu_n1204), .B(exu_n6000), .Y(exu_n21929));
AND2X1 exu_U3027(.A(exu_n1959), .B(exu_n6989), .Y(exu_n24473));
AND2X1 exu_U3028(.A(exu_n21933), .B(exu_n6001), .Y(bypass_rs1_data_w2[35]));
AND2X1 exu_U3029(.A(exu_n1205), .B(exu_n6002), .Y(exu_n21933));
AND2X1 exu_U3030(.A(exu_n1960), .B(exu_n6990), .Y(exu_n24477));
AND2X1 exu_U3031(.A(exu_n21937), .B(exu_n6003), .Y(bypass_rs1_data_w2[34]));
AND2X1 exu_U3032(.A(exu_n1206), .B(exu_n6004), .Y(exu_n21937));
AND2X1 exu_U3033(.A(exu_n1961), .B(exu_n6991), .Y(exu_n24481));
AND2X1 exu_U3034(.A(exu_n21941), .B(exu_n6005), .Y(bypass_rs1_data_w2[33]));
AND2X1 exu_U3035(.A(exu_n1207), .B(exu_n6006), .Y(exu_n21941));
AND2X1 exu_U3036(.A(exu_n1962), .B(exu_n6992), .Y(exu_n24485));
AND2X1 exu_U3037(.A(exu_n21945), .B(exu_n6007), .Y(bypass_rs1_data_w2[32]));
AND2X1 exu_U3038(.A(exu_n1208), .B(exu_n6008), .Y(exu_n21945));
AND2X1 exu_U3039(.A(exu_n1963), .B(exu_n6993), .Y(exu_n24489));
AND2X1 exu_U3040(.A(exu_n21949), .B(exu_n6009), .Y(bypass_rs1_data_w2[31]));
AND2X1 exu_U3041(.A(exu_n1209), .B(exu_n6010), .Y(exu_n21949));
AND2X1 exu_U3042(.A(exu_n1964), .B(exu_n6994), .Y(exu_n24493));
AND2X1 exu_U3043(.A(exu_n21953), .B(exu_n6011), .Y(bypass_rs1_data_w2[30]));
AND2X1 exu_U3044(.A(exu_n1210), .B(exu_n6012), .Y(exu_n21953));
AND2X1 exu_U3045(.A(exu_n1965), .B(exu_n6995), .Y(exu_n24497));
AND2X1 exu_U3046(.A(exu_n21961), .B(exu_n6015), .Y(bypass_rs1_data_w2[29]));
AND2X1 exu_U3047(.A(exu_n1212), .B(exu_n6016), .Y(exu_n21961));
AND2X1 exu_U3048(.A(exu_n1967), .B(exu_n6997), .Y(exu_n24505));
AND2X1 exu_U3049(.A(exu_n21965), .B(exu_n6017), .Y(bypass_rs1_data_w2[28]));
AND2X1 exu_U3050(.A(exu_n1213), .B(exu_n6018), .Y(exu_n21965));
AND2X1 exu_U3051(.A(exu_n1968), .B(exu_n6998), .Y(exu_n24509));
AND2X1 exu_U3052(.A(exu_n21969), .B(exu_n6019), .Y(bypass_rs1_data_w2[27]));
AND2X1 exu_U3053(.A(exu_n1214), .B(exu_n6020), .Y(exu_n21969));
AND2X1 exu_U3054(.A(exu_n1969), .B(exu_n6999), .Y(exu_n24513));
AND2X1 exu_U3055(.A(exu_n21973), .B(exu_n6021), .Y(bypass_rs1_data_w2[26]));
AND2X1 exu_U3056(.A(exu_n1215), .B(exu_n6022), .Y(exu_n21973));
AND2X1 exu_U3057(.A(exu_n1970), .B(exu_n7000), .Y(exu_n24517));
AND2X1 exu_U3058(.A(exu_n21977), .B(exu_n6023), .Y(bypass_rs1_data_w2[25]));
AND2X1 exu_U3059(.A(exu_n1216), .B(exu_n6024), .Y(exu_n21977));
AND2X1 exu_U3060(.A(exu_n1971), .B(exu_n7001), .Y(exu_n24521));
AND2X1 exu_U3061(.A(exu_n21981), .B(exu_n6025), .Y(bypass_rs1_data_w2[24]));
AND2X1 exu_U3062(.A(exu_n1217), .B(exu_n6026), .Y(exu_n21981));
AND2X1 exu_U3063(.A(exu_n1972), .B(exu_n7002), .Y(exu_n24525));
AND2X1 exu_U3064(.A(exu_n21985), .B(exu_n6027), .Y(bypass_rs1_data_w2[23]));
AND2X1 exu_U3065(.A(exu_n1218), .B(exu_n6028), .Y(exu_n21985));
AND2X1 exu_U3066(.A(exu_n1973), .B(exu_n7003), .Y(exu_n24529));
AND2X1 exu_U3067(.A(exu_n21989), .B(exu_n6029), .Y(bypass_rs1_data_w2[22]));
AND2X1 exu_U3068(.A(exu_n1219), .B(exu_n6030), .Y(exu_n21989));
AND2X1 exu_U3069(.A(exu_n1974), .B(exu_n7004), .Y(exu_n24533));
AND2X1 exu_U3070(.A(exu_n21993), .B(exu_n6031), .Y(bypass_rs1_data_w2[21]));
AND2X1 exu_U3071(.A(exu_n1220), .B(exu_n6032), .Y(exu_n21993));
AND2X1 exu_U3072(.A(exu_n1975), .B(exu_n7005), .Y(exu_n24537));
AND2X1 exu_U3073(.A(exu_n21997), .B(exu_n6033), .Y(bypass_rs1_data_w2[20]));
AND2X1 exu_U3074(.A(exu_n1221), .B(exu_n6034), .Y(exu_n21997));
AND2X1 exu_U3075(.A(exu_n1976), .B(exu_n7006), .Y(exu_n24541));
AND2X1 exu_U3076(.A(exu_n22005), .B(exu_n6037), .Y(bypass_rs1_data_w2[19]));
AND2X1 exu_U3077(.A(exu_n1223), .B(exu_n6038), .Y(exu_n22005));
AND2X1 exu_U3078(.A(exu_n1978), .B(exu_n7008), .Y(exu_n24549));
AND2X1 exu_U3079(.A(exu_n22009), .B(exu_n6039), .Y(bypass_rs1_data_w2[18]));
AND2X1 exu_U3080(.A(exu_n1224), .B(exu_n6040), .Y(exu_n22009));
AND2X1 exu_U3081(.A(exu_n1979), .B(exu_n7009), .Y(exu_n24553));
AND2X1 exu_U3082(.A(exu_n22013), .B(exu_n6041), .Y(bypass_rs1_data_w2[17]));
AND2X1 exu_U3083(.A(exu_n1225), .B(exu_n6042), .Y(exu_n22013));
AND2X1 exu_U3084(.A(exu_n1980), .B(exu_n7010), .Y(exu_n24557));
AND2X1 exu_U3085(.A(exu_n22017), .B(exu_n6043), .Y(bypass_rs1_data_w2[16]));
AND2X1 exu_U3086(.A(exu_n1226), .B(exu_n6044), .Y(exu_n22017));
AND2X1 exu_U3087(.A(exu_n1981), .B(exu_n7011), .Y(exu_n24561));
AND2X1 exu_U3088(.A(exu_n22021), .B(exu_n6045), .Y(bypass_rs1_data_w2[15]));
AND2X1 exu_U3089(.A(exu_n1227), .B(exu_n6046), .Y(exu_n22021));
AND2X1 exu_U3090(.A(exu_n1982), .B(exu_n7012), .Y(exu_n24565));
AND2X1 exu_U3091(.A(exu_n22025), .B(exu_n6047), .Y(bypass_rs1_data_w2[14]));
AND2X1 exu_U3092(.A(exu_n1228), .B(exu_n6048), .Y(exu_n22025));
AND2X1 exu_U3093(.A(exu_n1983), .B(exu_n7013), .Y(exu_n24569));
AND2X1 exu_U3094(.A(exu_n22029), .B(exu_n6049), .Y(bypass_rs1_data_w2[13]));
AND2X1 exu_U3095(.A(exu_n1229), .B(exu_n6050), .Y(exu_n22029));
AND2X1 exu_U3096(.A(exu_n1984), .B(exu_n7014), .Y(exu_n24573));
AND2X1 exu_U3097(.A(exu_n22033), .B(exu_n6051), .Y(bypass_rs1_data_w2[12]));
AND2X1 exu_U3098(.A(exu_n1230), .B(exu_n6052), .Y(exu_n22033));
AND2X1 exu_U3099(.A(exu_n1985), .B(exu_n7015), .Y(exu_n24577));
AND2X1 exu_U3100(.A(exu_n22037), .B(exu_n6053), .Y(bypass_rs1_data_w2[11]));
AND2X1 exu_U3101(.A(exu_n1231), .B(exu_n6054), .Y(exu_n22037));
AND2X1 exu_U3102(.A(exu_n1986), .B(exu_n7016), .Y(exu_n24581));
AND2X1 exu_U3103(.A(exu_n22041), .B(exu_n6055), .Y(bypass_rs1_data_w2[10]));
AND2X1 exu_U3104(.A(exu_n1232), .B(exu_n6056), .Y(exu_n22041));
AND2X1 exu_U3105(.A(exu_n1987), .B(exu_n7017), .Y(exu_n24585));
AND2X1 exu_U3106(.A(exu_n21793), .B(exu_n5931), .Y(bypass_rs1_data_w2[9]));
AND2X1 exu_U3107(.A(exu_n1170), .B(exu_n5932), .Y(exu_n21793));
AND2X1 exu_U3108(.A(exu_n1925), .B(exu_n6955), .Y(exu_n24337));
AND2X1 exu_U3109(.A(exu_n21797), .B(exu_n5933), .Y(bypass_rs1_data_w2[8]));
AND2X1 exu_U3110(.A(exu_n1171), .B(exu_n5934), .Y(exu_n21797));
AND2X1 exu_U3111(.A(exu_n1926), .B(exu_n6956), .Y(exu_n24341));
AND2X1 exu_U3112(.A(exu_n21801), .B(exu_n5935), .Y(bypass_rs1_data_w2[7]));
AND2X1 exu_U3113(.A(exu_n1172), .B(exu_n5936), .Y(exu_n21801));
AND2X1 exu_U3114(.A(exu_n1927), .B(exu_n6957), .Y(exu_n24345));
AND2X1 exu_U3115(.A(exu_n21805), .B(exu_n5937), .Y(bypass_rs1_data_w2[6]));
AND2X1 exu_U3116(.A(exu_n1173), .B(exu_n5938), .Y(exu_n21805));
AND2X1 exu_U3117(.A(exu_n1928), .B(exu_n6958), .Y(exu_n24349));
AND2X1 exu_U3118(.A(exu_n21825), .B(exu_n5947), .Y(bypass_rs1_data_w2[5]));
AND2X1 exu_U3119(.A(exu_n1178), .B(exu_n5948), .Y(exu_n21825));
AND2X1 exu_U3120(.A(exu_n1933), .B(exu_n6963), .Y(exu_n24369));
AND2X1 exu_U3121(.A(exu_n21869), .B(exu_n5969), .Y(bypass_rs1_data_w2[4]));
AND2X1 exu_U3122(.A(exu_n1189), .B(exu_n5970), .Y(exu_n21869));
AND2X1 exu_U3123(.A(exu_n1944), .B(exu_n6974), .Y(exu_n24413));
AND2X1 exu_U3124(.A(exu_n21913), .B(exu_n5991), .Y(bypass_rs1_data_w2[3]));
AND2X1 exu_U3125(.A(exu_n1200), .B(exu_n5992), .Y(exu_n21913));
AND2X1 exu_U3126(.A(exu_n1955), .B(exu_n6985), .Y(exu_n24457));
AND2X1 exu_U3127(.A(exu_n21957), .B(exu_n6013), .Y(bypass_rs1_data_w2[2]));
AND2X1 exu_U3128(.A(exu_n1211), .B(exu_n6014), .Y(exu_n21957));
AND2X1 exu_U3129(.A(exu_n1966), .B(exu_n6996), .Y(exu_n24501));
AND2X1 exu_U3130(.A(exu_n22001), .B(exu_n6035), .Y(bypass_rs1_data_w2[1]));
AND2X1 exu_U3131(.A(exu_n1222), .B(exu_n6036), .Y(exu_n22001));
AND2X1 exu_U3132(.A(exu_n1977), .B(exu_n7007), .Y(exu_n24545));
OR2X1 exu_U3133(.A(exu_n13439), .B(exu_n14757), .Y(ecl_byplog_rs1_n21));
AND2X1 exu_U3134(.A(exu_n22045), .B(exu_n6057), .Y(bypass_rs1_data_w2[0]));
AND2X1 exu_U3135(.A(exu_n1233), .B(exu_n6058), .Y(exu_n22045));
AND2X1 exu_U3136(.A(exu_n1988), .B(exu_n7018), .Y(exu_n24589));
INVX1 exu_U3137(.A(se), .Y(exu_n29756));
INVX1 exu_U3138(.A(se), .Y(exu_n29821));
INVX1 exu_U3139(.A(se), .Y(exu_n29886));
INVX1 exu_U3140(.A(se), .Y(exu_n29950));
AND2X1 exu_U3141(.A(exu_n16216), .B(ecl_divcntl_div_state_1), .Y(ecl_divcntl_n85));
INVX1 exu_U3142(.A(se), .Y(exu_n30015));
INVX1 exu_U3143(.A(se), .Y(exu_n30080));
AND2X1 exu_U3144(.A(exu_n15740), .B(rml_cwp_full_swap_w), .Y(rml_cwp_n28));
OR2X1 exu_U3145(.A(rml_save_e), .B(rml_restore_e), .Y(rml_cwp_n104));
AND2X1 exu_U3146(.A(exu_n228), .B(exu_n5155), .Y(exu_n17729));
AND2X1 exu_U3147(.A(exu_n230), .B(exu_n5157), .Y(exu_n17735));
AND2X1 exu_U3148(.A(exu_n232), .B(exu_n5159), .Y(exu_n17741));
AND2X1 exu_U3149(.A(ecl_divcntl_cntr[4]), .B(ecl_divcntl_cntr[3]), .Y(ecl_divcntl_n88));
INVX1 exu_U3150(.A(ecl_tid_m[1]), .Y(exu_n16578));
INVX1 exu_U3151(.A(ecl_tid_m[0]), .Y(exu_n16577));
OR2X1 exu_U3152(.A(exu_n15637), .B(exu_n15864), .Y(exu_n17035));
OR2X1 exu_U3153(.A(exu_n15636), .B(exu_n15865), .Y(exu_n17030));
OR2X1 exu_U3154(.A(exu_n15635), .B(exu_n15866), .Y(exu_n17023));
OR2X1 exu_U3155(.A(exu_n15634), .B(exu_n15868), .Y(exu_n17018));
OR2X1 exu_U3156(.A(exu_n15633), .B(exu_n15869), .Y(exu_n17013));
OR2X1 exu_U3157(.A(exu_n15632), .B(exu_n15870), .Y(exu_n17008));
OR2X1 exu_U3158(.A(exu_n15631), .B(exu_n15871), .Y(exu_n17003));
OR2X1 exu_U3159(.A(exu_n15630), .B(exu_n15872), .Y(exu_n16998));
OR2X1 exu_U3160(.A(exu_n15629), .B(exu_n15873), .Y(exu_n16993));
OR2X1 exu_U3161(.A(exu_n15628), .B(exu_n15874), .Y(exu_n16988));
OR2X1 exu_U3162(.A(exu_n15627), .B(exu_n15875), .Y(exu_n16983));
OR2X1 exu_U3163(.A(exu_n15626), .B(exu_n15876), .Y(exu_n16978));
OR2X1 exu_U3164(.A(exu_n15625), .B(exu_n15877), .Y(exu_n16971));
OR2X1 exu_U3165(.A(exu_n15624), .B(exu_n15879), .Y(exu_n16966));
OR2X1 exu_U3166(.A(exu_n15623), .B(exu_n15880), .Y(exu_n16961));
OR2X1 exu_U3167(.A(exu_n15622), .B(exu_n15881), .Y(exu_n16956));
OR2X1 exu_U3168(.A(exu_n15621), .B(exu_n15882), .Y(exu_n16951));
OR2X1 exu_U3169(.A(exu_n15620), .B(exu_n15883), .Y(exu_n16946));
OR2X1 exu_U3170(.A(exu_n15619), .B(exu_n15884), .Y(exu_n16941));
OR2X1 exu_U3171(.A(exu_n15618), .B(exu_n15885), .Y(exu_n16936));
OR2X1 exu_U3172(.A(exu_n15617), .B(exu_n15886), .Y(exu_n16931));
OR2X1 exu_U3173(.A(exu_n15576), .B(exu_n15887), .Y(exu_n16926));
OR2X1 exu_U3174(.A(exu_n15575), .B(exu_n15888), .Y(exu_n16923));
OR2X1 exu_U3175(.A(exu_n15574), .B(exu_n15890), .Y(exu_n16920));
OR2X1 exu_U3176(.A(exu_n15573), .B(exu_n15891), .Y(exu_n16917));
OR2X1 exu_U3177(.A(exu_n15572), .B(exu_n15892), .Y(exu_n16914));
OR2X1 exu_U3178(.A(exu_n15571), .B(exu_n15893), .Y(exu_n16911));
OR2X1 exu_U3179(.A(exu_n15570), .B(exu_n15894), .Y(exu_n16908));
OR2X1 exu_U3180(.A(exu_n15569), .B(exu_n15895), .Y(exu_n16905));
OR2X1 exu_U3181(.A(exu_n15568), .B(exu_n15896), .Y(exu_n16902));
OR2X1 exu_U3182(.A(div_adderin2[32]), .B(exu_n15858), .Y(exu_n16899));
OR2X1 exu_U3183(.A(exu_n15616), .B(exu_n15897), .Y(exu_n16881));
OR2X1 exu_U3184(.A(exu_n15614), .B(exu_n15900), .Y(exu_n16871));
OR2X1 exu_U3185(.A(exu_n15613), .B(exu_n15901), .Y(exu_n16864));
OR2X1 exu_U3186(.A(exu_n15612), .B(exu_n15902), .Y(exu_n16859));
OR2X1 exu_U3187(.A(exu_n15611), .B(exu_n15903), .Y(exu_n16854));
OR2X1 exu_U3188(.A(exu_n15610), .B(exu_n15904), .Y(exu_n16849));
OR2X1 exu_U3189(.A(exu_n15609), .B(exu_n15905), .Y(exu_n16844));
OR2X1 exu_U3190(.A(exu_n15608), .B(exu_n15906), .Y(exu_n16839));
OR2X1 exu_U3191(.A(exu_n15607), .B(exu_n15907), .Y(exu_n16834));
OR2X1 exu_U3192(.A(exu_n15606), .B(exu_n15908), .Y(exu_n16829));
OR2X1 exu_U3193(.A(exu_n15605), .B(exu_n15909), .Y(exu_n16824));
OR2X1 exu_U3194(.A(exu_n15604), .B(exu_n15911), .Y(exu_n16819));
OR2X1 exu_U3195(.A(exu_n15603), .B(exu_n15912), .Y(exu_n16812));
OR2X1 exu_U3196(.A(exu_n15602), .B(exu_n15913), .Y(exu_n16807));
OR2X1 exu_U3197(.A(exu_n15601), .B(exu_n15914), .Y(exu_n16802));
OR2X1 exu_U3198(.A(exu_n15600), .B(exu_n15915), .Y(exu_n16797));
OR2X1 exu_U3199(.A(exu_n15599), .B(exu_n15916), .Y(exu_n16792));
OR2X1 exu_U3200(.A(exu_n15598), .B(exu_n15917), .Y(exu_n16787));
OR2X1 exu_U3201(.A(exu_n15597), .B(exu_n15918), .Y(exu_n16782));
OR2X1 exu_U3202(.A(exu_n15596), .B(exu_n15919), .Y(exu_n16777));
OR2X1 exu_U3203(.A(exu_n15595), .B(exu_n15920), .Y(exu_n16772));
OR2X1 exu_U3204(.A(exu_n15567), .B(exu_n15860), .Y(exu_n16767));
OR2X1 exu_U3205(.A(exu_n15566), .B(exu_n15861), .Y(exu_n16764));
OR2X1 exu_U3206(.A(exu_n15565), .B(exu_n15862), .Y(exu_n16761));
OR2X1 exu_U3207(.A(exu_n15564), .B(exu_n15863), .Y(exu_n16758));
OR2X1 exu_U3208(.A(exu_n15563), .B(exu_n15867), .Y(exu_n16755));
OR2X1 exu_U3209(.A(exu_n15562), .B(exu_n15878), .Y(exu_n16752));
OR2X1 exu_U3210(.A(exu_n15561), .B(exu_n15889), .Y(exu_n16749));
OR2X1 exu_U3211(.A(exu_n15560), .B(exu_n15899), .Y(exu_n16746));
OR2X1 exu_U3212(.A(exu_n15559), .B(exu_n15910), .Y(exu_n16743));
OR2X1 exu_U3213(.A(div_adderin2[0]), .B(exu_n15859), .Y(exu_n16740));
OR2X1 exu_U3214(.A(exu_n12180), .B(exu_n13592), .Y(div_byp_yreg_e[7]));
AND2X1 exu_U3215(.A(exu_n855), .B(exu_n5616), .Y(exu_n20680));
OR2X1 exu_U3216(.A(exu_n12181), .B(exu_n13593), .Y(div_byp_yreg_e[6]));
AND2X1 exu_U3217(.A(exu_n857), .B(exu_n5618), .Y(exu_n20686));
OR2X1 exu_U3218(.A(exu_n12182), .B(exu_n13594), .Y(div_byp_yreg_e[5]));
AND2X1 exu_U3219(.A(exu_n859), .B(exu_n5620), .Y(exu_n20692));
OR2X1 exu_U3220(.A(exu_n12183), .B(exu_n13595), .Y(div_byp_yreg_e[4]));
AND2X1 exu_U3221(.A(exu_n861), .B(exu_n5622), .Y(exu_n20698));
OR2X1 exu_U3222(.A(exu_n12184), .B(exu_n13596), .Y(div_byp_yreg_e[3]));
AND2X1 exu_U3223(.A(exu_n863), .B(exu_n5624), .Y(exu_n20704));
OR2X1 exu_U3224(.A(exu_n12187), .B(exu_n13599), .Y(div_byp_yreg_e[2]));
AND2X1 exu_U3225(.A(exu_n869), .B(exu_n5630), .Y(exu_n20722));
OR2X1 exu_U3226(.A(exu_n12198), .B(exu_n13610), .Y(div_byp_yreg_e[1]));
AND2X1 exu_U3227(.A(exu_n891), .B(exu_n5652), .Y(exu_n20788));
OR2X1 exu_U3228(.A(exu_n12209), .B(exu_n13621), .Y(div_byp_yreg_e[0]));
AND2X1 exu_U3229(.A(exu_n913), .B(exu_n5674), .Y(exu_n20854));
INVX1 exu_U3230(.A(div_curr_q[31]), .Y(exu_n16435));
AND2X1 exu_U3231(.A(div_curr_q[30]), .B(ecl_divcntl_n60), .Y(div_neg32[30]));
AND2X1 exu_U3232(.A(div_curr_q[29]), .B(ecl_divcntl_n60), .Y(div_neg32[29]));
AND2X1 exu_U3233(.A(div_curr_q[28]), .B(ecl_divcntl_n60), .Y(div_neg32[28]));
AND2X1 exu_U3234(.A(div_curr_q[27]), .B(ecl_divcntl_n60), .Y(div_neg32[27]));
AND2X1 exu_U3235(.A(div_curr_q[26]), .B(ecl_divcntl_n60), .Y(div_neg32[26]));
AND2X1 exu_U3236(.A(div_curr_q[25]), .B(ecl_divcntl_n60), .Y(div_neg32[25]));
AND2X1 exu_U3237(.A(div_curr_q[24]), .B(ecl_divcntl_n60), .Y(div_neg32[24]));
AND2X1 exu_U3238(.A(div_curr_q[23]), .B(ecl_divcntl_n60), .Y(div_neg32[23]));
AND2X1 exu_U3239(.A(div_curr_q[22]), .B(ecl_divcntl_n60), .Y(div_neg32[22]));
AND2X1 exu_U3240(.A(div_curr_q[21]), .B(ecl_divcntl_n60), .Y(div_neg32[21]));
AND2X1 exu_U3241(.A(div_curr_q[20]), .B(ecl_divcntl_n60), .Y(div_neg32[20]));
AND2X1 exu_U3242(.A(div_curr_q[19]), .B(ecl_divcntl_n60), .Y(div_neg32[19]));
AND2X1 exu_U3243(.A(div_curr_q[18]), .B(ecl_divcntl_n60), .Y(div_neg32[18]));
AND2X1 exu_U3244(.A(div_curr_q[17]), .B(ecl_divcntl_n60), .Y(div_neg32[17]));
AND2X1 exu_U3245(.A(div_curr_q[16]), .B(ecl_divcntl_n60), .Y(div_neg32[16]));
AND2X1 exu_U3246(.A(div_curr_q[15]), .B(ecl_divcntl_n60), .Y(div_neg32[15]));
AND2X1 exu_U3247(.A(div_curr_q[14]), .B(ecl_divcntl_n60), .Y(div_neg32[14]));
AND2X1 exu_U3248(.A(div_curr_q[13]), .B(ecl_divcntl_n60), .Y(div_neg32[13]));
AND2X1 exu_U3249(.A(div_curr_q[12]), .B(ecl_divcntl_n60), .Y(div_neg32[12]));
AND2X1 exu_U3250(.A(div_curr_q[11]), .B(ecl_divcntl_n60), .Y(div_neg32[11]));
AND2X1 exu_U3251(.A(div_curr_q[10]), .B(ecl_divcntl_n60), .Y(div_neg32[10]));
AND2X1 exu_U3252(.A(ecl_divcntl_n60), .B(div_curr_q[9]), .Y(div_neg32[9]));
AND2X1 exu_U3253(.A(div_curr_q[8]), .B(ecl_divcntl_n60), .Y(div_neg32[8]));
AND2X1 exu_U3254(.A(div_curr_q[7]), .B(ecl_divcntl_n60), .Y(div_neg32[7]));
AND2X1 exu_U3255(.A(div_curr_q[6]), .B(ecl_divcntl_n60), .Y(div_neg32[6]));
AND2X1 exu_U3256(.A(div_curr_q[5]), .B(ecl_divcntl_n60), .Y(div_neg32[5]));
AND2X1 exu_U3257(.A(div_curr_q[4]), .B(ecl_divcntl_n60), .Y(div_neg32[4]));
AND2X1 exu_U3258(.A(div_curr_q[3]), .B(ecl_divcntl_n60), .Y(div_neg32[3]));
AND2X1 exu_U3259(.A(div_curr_q[2]), .B(ecl_divcntl_n60), .Y(div_neg32[2]));
AND2X1 exu_U3260(.A(div_curr_q[1]), .B(ecl_divcntl_n60), .Y(div_neg32[1]));
AND2X1 exu_U3261(.A(div_curr_q[0]), .B(ecl_divcntl_n60), .Y(div_neg32[0]));
INVX1 exu_U3262(.A(ecl_tid_w[0]), .Y(exu_n16576));
AND2X1 exu_U3263(.A(exu_n4635), .B(exu_n9415), .Y(bypass_rs3h_w2_mux_n29));
AND2X1 exu_U3264(.A(exu_n4596), .B(exu_n9382), .Y(bypass_mux_rs3h_data_1_n43));
AND2X1 exu_U3265(.A(exu_n4637), .B(exu_n9416), .Y(bypass_rs3h_w2_mux_n33));
AND2X1 exu_U3266(.A(exu_n4597), .B(exu_n9383), .Y(bypass_mux_rs3h_data_1_n49));
AND2X1 exu_U3267(.A(exu_n4641), .B(exu_n9418), .Y(bypass_rs3h_w2_mux_n41));
AND2X1 exu_U3268(.A(exu_n4599), .B(exu_n9385), .Y(bypass_mux_rs3h_data_1_n61));
AND2X1 exu_U3269(.A(exu_n4643), .B(exu_n9419), .Y(bypass_rs3h_w2_mux_n45));
AND2X1 exu_U3270(.A(exu_n4600), .B(exu_n9386), .Y(bypass_mux_rs3h_data_1_n67));
AND2X1 exu_U3271(.A(exu_n4645), .B(exu_n9420), .Y(bypass_rs3h_w2_mux_n49));
AND2X1 exu_U3272(.A(exu_n4601), .B(exu_n9387), .Y(bypass_mux_rs3h_data_1_n73));
AND2X1 exu_U3273(.A(exu_n4647), .B(exu_n9421), .Y(bypass_rs3h_w2_mux_n53));
AND2X1 exu_U3274(.A(exu_n4602), .B(exu_n9388), .Y(bypass_mux_rs3h_data_1_n79));
AND2X1 exu_U3275(.A(exu_n4649), .B(exu_n9422), .Y(bypass_rs3h_w2_mux_n57));
AND2X1 exu_U3276(.A(exu_n4603), .B(exu_n9389), .Y(bypass_mux_rs3h_data_1_n85));
AND2X1 exu_U3277(.A(exu_n4651), .B(exu_n9423), .Y(bypass_rs3h_w2_mux_n61));
AND2X1 exu_U3278(.A(exu_n4604), .B(exu_n9390), .Y(bypass_mux_rs3h_data_1_n91));
AND2X1 exu_U3279(.A(exu_n4653), .B(exu_n9424), .Y(bypass_rs3h_w2_mux_n65));
AND2X1 exu_U3280(.A(exu_n4605), .B(exu_n9391), .Y(bypass_mux_rs3h_data_1_n97));
AND2X1 exu_U3281(.A(exu_n4655), .B(exu_n9425), .Y(bypass_rs3h_w2_mux_n69));
AND2X1 exu_U3282(.A(exu_n4606), .B(exu_n9392), .Y(bypass_mux_rs3h_data_1_n103));
AND2X1 exu_U3283(.A(exu_n4657), .B(exu_n9426), .Y(bypass_rs3h_w2_mux_n73));
AND2X1 exu_U3284(.A(exu_n4607), .B(exu_n9393), .Y(bypass_mux_rs3h_data_1_n109));
AND2X1 exu_U3285(.A(exu_n4659), .B(exu_n9427), .Y(bypass_rs3h_w2_mux_n77));
AND2X1 exu_U3286(.A(exu_n4608), .B(exu_n9394), .Y(bypass_mux_rs3h_data_1_n115));
AND2X1 exu_U3287(.A(exu_n4663), .B(exu_n9429), .Y(bypass_rs3h_w2_mux_n85));
AND2X1 exu_U3288(.A(exu_n4610), .B(exu_n9396), .Y(bypass_mux_rs3h_data_1_n127));
AND2X1 exu_U3289(.A(exu_n4665), .B(exu_n9430), .Y(bypass_rs3h_w2_mux_n89));
AND2X1 exu_U3290(.A(exu_n4611), .B(exu_n9397), .Y(bypass_mux_rs3h_data_1_n133));
AND2X1 exu_U3291(.A(exu_n4667), .B(exu_n9431), .Y(bypass_rs3h_w2_mux_n93));
AND2X1 exu_U3292(.A(exu_n4612), .B(exu_n9398), .Y(bypass_mux_rs3h_data_1_n139));
AND2X1 exu_U3293(.A(exu_n4669), .B(exu_n9432), .Y(bypass_rs3h_w2_mux_n97));
AND2X1 exu_U3294(.A(exu_n4613), .B(exu_n9399), .Y(bypass_mux_rs3h_data_1_n145));
AND2X1 exu_U3295(.A(exu_n4671), .B(exu_n9433), .Y(bypass_rs3h_w2_mux_n101));
AND2X1 exu_U3296(.A(exu_n4614), .B(exu_n9400), .Y(bypass_mux_rs3h_data_1_n151));
AND2X1 exu_U3297(.A(exu_n4673), .B(exu_n9434), .Y(bypass_rs3h_w2_mux_n105));
AND2X1 exu_U3298(.A(exu_n4615), .B(exu_n9401), .Y(bypass_mux_rs3h_data_1_n157));
AND2X1 exu_U3299(.A(exu_n4675), .B(exu_n9435), .Y(bypass_rs3h_w2_mux_n109));
AND2X1 exu_U3300(.A(exu_n4616), .B(exu_n9402), .Y(bypass_mux_rs3h_data_1_n163));
AND2X1 exu_U3301(.A(exu_n4677), .B(exu_n9436), .Y(bypass_rs3h_w2_mux_n113));
AND2X1 exu_U3302(.A(exu_n4617), .B(exu_n9403), .Y(bypass_mux_rs3h_data_1_n169));
AND2X1 exu_U3303(.A(exu_n4679), .B(exu_n9437), .Y(bypass_rs3h_w2_mux_n117));
AND2X1 exu_U3304(.A(exu_n4618), .B(exu_n9404), .Y(bypass_mux_rs3h_data_1_n175));
AND2X1 exu_U3305(.A(exu_n4681), .B(exu_n9438), .Y(bypass_rs3h_w2_mux_n121));
AND2X1 exu_U3306(.A(exu_n4619), .B(exu_n9405), .Y(bypass_mux_rs3h_data_1_n181));
OR2X1 exu_U3307(.A(exu_n12914), .B(exu_n14198), .Y(alu_byp_rd_data_e[9]));
AND2X1 exu_U3308(.A(exu_n2568), .B(exu_n7596), .Y(exu_n26353));
AND2X1 exu_U3309(.A(exu_n4621), .B(exu_n9408), .Y(bypass_rs3h_w2_mux_n1));
AND2X1 exu_U3310(.A(exu_n4589), .B(exu_n9375), .Y(bypass_mux_rs3h_data_1_n1));
AND2X1 exu_U3311(.A(exu_n4623), .B(exu_n9409), .Y(bypass_rs3h_w2_mux_n5));
AND2X1 exu_U3312(.A(exu_n4590), .B(exu_n9376), .Y(bypass_mux_rs3h_data_1_n7));
AND2X1 exu_U3313(.A(exu_n4625), .B(exu_n9410), .Y(bypass_rs3h_w2_mux_n9));
AND2X1 exu_U3314(.A(exu_n4591), .B(exu_n9377), .Y(bypass_mux_rs3h_data_1_n13));
AND2X1 exu_U3315(.A(exu_n4627), .B(exu_n9411), .Y(bypass_rs3h_w2_mux_n13));
AND2X1 exu_U3316(.A(exu_n4592), .B(exu_n9378), .Y(bypass_mux_rs3h_data_1_n19));
AND2X1 exu_U3317(.A(exu_n4629), .B(exu_n9412), .Y(bypass_rs3h_w2_mux_n17));
AND2X1 exu_U3318(.A(exu_n4593), .B(exu_n9379), .Y(bypass_mux_rs3h_data_1_n25));
AND2X1 exu_U3319(.A(exu_n4631), .B(exu_n9413), .Y(bypass_rs3h_w2_mux_n21));
AND2X1 exu_U3320(.A(exu_n4594), .B(exu_n9380), .Y(bypass_mux_rs3h_data_1_n31));
AND2X1 exu_U3321(.A(exu_n4633), .B(exu_n9414), .Y(bypass_rs3h_w2_mux_n25));
AND2X1 exu_U3322(.A(exu_n4595), .B(exu_n9381), .Y(bypass_mux_rs3h_data_1_n37));
AND2X1 exu_U3323(.A(exu_n4639), .B(exu_n9417), .Y(bypass_rs3h_w2_mux_n37));
AND2X1 exu_U3324(.A(exu_n4598), .B(exu_n9384), .Y(bypass_mux_rs3h_data_1_n55));
AND2X1 exu_U3325(.A(exu_n4661), .B(exu_n9428), .Y(bypass_rs3h_w2_mux_n81));
AND2X1 exu_U3326(.A(exu_n4609), .B(exu_n9395), .Y(bypass_mux_rs3h_data_1_n121));
OR2X1 exu_U3327(.A(exu_n12143), .B(exu_n14758), .Y(exu_n19228));
AND2X1 exu_U3328(.A(exu_n15819), .B(exu_n19228), .Y(exu_n19225));
AND2X1 exu_U3329(.A(exu_n19230), .B(exu_n19231), .Y(exu_n19226));
AND2X1 exu_U3330(.A(exu_n15434), .B(exu_n15422), .Y(exu_n19230));
AND2X1 exu_U3331(.A(exu_n4683), .B(exu_n9439), .Y(bypass_rs3h_w2_mux_n125));
AND2X1 exu_U3332(.A(exu_n4620), .B(exu_n9406), .Y(bypass_mux_rs3h_data_1_n187));
INVX1 exu_U3333(.A(se), .Y(bypass_dfill_data_dff_n1));
INVX1 exu_U3334(.A(ecl_eccctl_rs3_ue_m), .Y(exu_n16592));
OR2X1 exu_U3335(.A(exu_n15639), .B(alu_logic_rs1_data_bf1[10]), .Y(exu_n17090));
OR2X1 exu_U3336(.A(exu_n15640), .B(alu_logic_rs1_data_bf1[11]), .Y(exu_n17095));
OR2X1 exu_U3337(.A(exu_n15641), .B(alu_logic_rs1_data_bf1[12]), .Y(exu_n17100));
OR2X1 exu_U3338(.A(exu_n15642), .B(alu_logic_rs1_data_bf1[13]), .Y(exu_n17105));
OR2X1 exu_U3339(.A(exu_n15643), .B(alu_logic_rs1_data_bf1[14]), .Y(exu_n17110));
OR2X1 exu_U3340(.A(exu_n15644), .B(alu_logic_rs1_data_bf1[15]), .Y(exu_n17115));
OR2X1 exu_U3341(.A(exu_n15645), .B(alu_logic_rs1_data_bf1[16]), .Y(exu_n17120));
OR2X1 exu_U3342(.A(exu_n15646), .B(alu_logic_rs1_data_bf1[17]), .Y(exu_n17125));
OR2X1 exu_U3343(.A(exu_n15647), .B(alu_logic_rs1_data_bf1[18]), .Y(exu_n17130));
OR2X1 exu_U3344(.A(exu_n15648), .B(alu_logic_rs1_data_bf1[19]), .Y(exu_n17137));
OR2X1 exu_U3345(.A(exu_n15649), .B(alu_logic_rs1_data_bf1[20]), .Y(exu_n17142));
OR2X1 exu_U3346(.A(exu_n15650), .B(alu_logic_rs1_data_bf1[21]), .Y(exu_n17147));
OR2X1 exu_U3347(.A(exu_n15651), .B(alu_logic_rs1_data_bf1[22]), .Y(exu_n17152));
OR2X1 exu_U3348(.A(exu_n15652), .B(alu_logic_rs1_data_bf1[23]), .Y(exu_n17157));
OR2X1 exu_U3349(.A(exu_n15653), .B(alu_logic_rs1_data_bf1[24]), .Y(exu_n17162));
OR2X1 exu_U3350(.A(exu_n15654), .B(alu_logic_rs1_data_bf1[25]), .Y(exu_n17167));
OR2X1 exu_U3351(.A(exu_n15655), .B(alu_logic_rs1_data_bf1[26]), .Y(exu_n17172));
OR2X1 exu_U3352(.A(exu_n15656), .B(alu_logic_rs1_data_bf1[27]), .Y(exu_n17177));
OR2X1 exu_U3353(.A(exu_n15657), .B(alu_logic_rs1_data_bf1[28]), .Y(exu_n17182));
OR2X1 exu_U3354(.A(exu_n15658), .B(alu_logic_rs1_data_bf1[29]), .Y(exu_n17189));
OR2X1 exu_U3355(.A(exu_n15659), .B(alu_logic_rs1_data_bf1[30]), .Y(exu_n17194));
OR2X1 exu_U3356(.A(exu_n15660), .B(alu_logic_rs1_data_bf1[31]), .Y(exu_n17199));
OR2X1 exu_U3357(.A(alu_addsub_rs2_data[32]), .B(alu_logic_rs1_data_bf1[32]), .Y(exu_n17217));
OR2X1 exu_U3358(.A(exu_n15586), .B(alu_logic_rs1_data_bf1[33]), .Y(exu_n17220));
OR2X1 exu_U3359(.A(exu_n15587), .B(alu_logic_rs1_data_bf1[34]), .Y(exu_n17223));
OR2X1 exu_U3360(.A(exu_n15588), .B(alu_logic_rs1_data_bf1[35]), .Y(exu_n17226));
OR2X1 exu_U3361(.A(exu_n15589), .B(alu_logic_rs1_data_bf1[36]), .Y(exu_n17229));
OR2X1 exu_U3362(.A(exu_n15590), .B(alu_logic_rs1_data_bf1[37]), .Y(exu_n17232));
OR2X1 exu_U3363(.A(exu_n15591), .B(alu_logic_rs1_data_bf1[38]), .Y(exu_n17235));
OR2X1 exu_U3364(.A(exu_n15592), .B(alu_logic_rs1_data_bf1[39]), .Y(exu_n17238));
OR2X1 exu_U3365(.A(exu_n15593), .B(alu_logic_rs1_data_bf1[40]), .Y(exu_n17241));
OR2X1 exu_U3366(.A(exu_n15594), .B(alu_logic_rs1_data_bf1[41]), .Y(exu_n17244));
OR2X1 exu_U3367(.A(exu_n15661), .B(alu_logic_rs1_data_bf1[42]), .Y(exu_n17249));
OR2X1 exu_U3368(.A(exu_n15662), .B(alu_logic_rs1_data_bf1[43]), .Y(exu_n17254));
OR2X1 exu_U3369(.A(exu_n15663), .B(alu_logic_rs1_data_bf1[44]), .Y(exu_n17259));
OR2X1 exu_U3370(.A(exu_n15664), .B(alu_logic_rs1_data_bf1[45]), .Y(exu_n17264));
OR2X1 exu_U3371(.A(exu_n15665), .B(alu_logic_rs1_data_bf1[46]), .Y(exu_n17269));
OR2X1 exu_U3372(.A(exu_n13427), .B(exu_n14740), .Y(ecl_ccr_ccr_d[0]));
OR2X1 exu_U3373(.A(exu_n13426), .B(exu_n14739), .Y(ecl_ccr_ccr_d[1]));
OR2X1 exu_U3374(.A(exu_n13425), .B(exu_n14738), .Y(ecl_ccr_ccr_d[2]));
OR2X1 exu_U3375(.A(exu_n13424), .B(exu_n14737), .Y(ecl_ccr_ccr_d[3]));
OR2X1 exu_U3376(.A(exu_n13423), .B(exu_n14736), .Y(ecl_ccr_ccr_d[4]));
OR2X1 exu_U3377(.A(exu_n13422), .B(exu_n14735), .Y(ecl_ccr_ccr_d[5]));
OR2X1 exu_U3378(.A(exu_n13421), .B(exu_n14734), .Y(ecl_ccr_ccr_d[6]));
OR2X1 exu_U3379(.A(exu_n13420), .B(exu_n14733), .Y(ecl_ccr_ccr_d[7]));
AND2X1 exu_U3380(.A(ecl_eccctl_n15), .B(exu_n9324), .Y(ecl_ecc_log_rs3_m));
AND2X1 exu_U3381(.A(exu_n16593), .B(exu_n16594), .Y(ecl_eccctl_n15));
AND2X1 exu_U3382(.A(exu_n16594), .B(exu_n9326), .Y(ecl_ecc_log_rs1_m));
AND2X1 exu_U3383(.A(exu_n4524), .B(exu_n16594), .Y(ecl_ecc_log_rs2_m));
AND2X1 exu_U3384(.A(exu_n4537), .B(exu_n9335), .Y(ecl_writeback_n98));
AND2X1 exu_U3385(.A(exu_n4536), .B(exu_n9334), .Y(ecl_writeback_n97));
INVX1 exu_U3386(.A(ecl_writeback_short_longop_done_m), .Y(exu_n16596));
AND2X1 exu_U3387(.A(ecl_flush_w1), .B(ecl_thr_match_mw1), .Y(ecl_ecl_exu_kill_m));
AND2X1 exu_U3388(.A(exu_n3988), .B(exu_n9001), .Y(exu_n31646));
AND2X1 exu_U3389(.A(exu_n3973), .B(exu_n8986), .Y(exu_n31617));
AND2X1 exu_U3390(.A(exu_n3978), .B(exu_n8991), .Y(exu_n31616));
AND2X1 exu_U3391(.A(exu_n3983), .B(exu_n8996), .Y(exu_n31647));
OR2X1 exu_U3392(.A(exu_n15583), .B(alu_logic_rs1_data_bf1[7]), .Y(exu_n17079));
OR2X1 exu_U3393(.A(exu_n15584), .B(alu_logic_rs1_data_bf1[8]), .Y(exu_n17082));
OR2X1 exu_U3394(.A(exu_n15585), .B(alu_logic_rs1_data_bf1[9]), .Y(exu_n17085));
OR2X1 exu_U3395(.A(alu_addsub_rs2_data_0), .B(alu_logic_rs1_data_bf1[0]), .Y(exu_n17058));
OR2X1 exu_U3396(.A(exu_n15577), .B(alu_logic_rs1_data_bf1[1]), .Y(exu_n17061));
OR2X1 exu_U3397(.A(exu_n15578), .B(alu_logic_rs1_data_bf1[2]), .Y(exu_n17064));
OR2X1 exu_U3398(.A(exu_n15579), .B(alu_logic_rs1_data_bf1[3]), .Y(exu_n17067));
OR2X1 exu_U3399(.A(exu_n15580), .B(alu_logic_rs1_data_bf1[4]), .Y(exu_n17070));
OR2X1 exu_U3400(.A(exu_n15581), .B(alu_logic_rs1_data_bf1[5]), .Y(exu_n17073));
OR2X1 exu_U3401(.A(exu_n15582), .B(alu_logic_rs1_data_bf1[6]), .Y(exu_n17076));
AND2X1 exu_U3402(.A(tlu_exu_agp_tid[1]), .B(tlu_exu_agp_tid[0]), .Y(rml_agp_thr[3]));
OR2X1 exu_U3403(.A(ecl_kill_rml_w), .B(ecl_tlu_priv_trap_w), .Y(ecl_rml_kill_w));
AND2X1 exu_U3404(.A(exu_n4020), .B(exu_n9036), .Y(rml_cwp_cwp_output_mux_n62));
AND2X1 exu_U3405(.A(exu_n4021), .B(exu_n9037), .Y(rml_cwp_cwp_output_mux_n61));
OR2X1 exu_U3406(.A(rml_restore_e), .B(rml_cwp_n96), .Y(rml_n48));
OR2X1 exu_U3407(.A(exu_n13403), .B(exu_n14714), .Y(rml_cwp_new_swap_cwp[0]));
AND2X1 exu_U3408(.A(exu_n4013), .B(exu_n9029), .Y(rml_cwp_cwp_output_mux_n37));
OR2X1 exu_U3409(.A(exu_n13402), .B(exu_n14713), .Y(rml_cwp_new_swap_cwp[1]));
AND2X1 exu_U3410(.A(exu_n4011), .B(exu_n9027), .Y(rml_cwp_cwp_output_mux_n31));
AND2X1 exu_U3411(.A(exu_n244), .B(exu_n5171), .Y(exu_n17777));
AND2X1 exu_U3412(.A(exu_n4028), .B(exu_n9044), .Y(rml_cwp_cwp_output_mux_n86));
AND2X1 exu_U3413(.A(exu_n4029), .B(exu_n9045), .Y(rml_cwp_cwp_output_mux_n85));
AND2X1 exu_U3414(.A(exu_n242), .B(exu_n5169), .Y(exu_n17771));
AND2X1 exu_U3415(.A(exu_n4016), .B(exu_n9032), .Y(rml_cwp_cwp_output_mux_n50));
AND2X1 exu_U3416(.A(exu_n4017), .B(exu_n9033), .Y(rml_cwp_cwp_output_mux_n49));
AND2X1 exu_U3417(.A(exu_n240), .B(exu_n5167), .Y(exu_n17765));
AND2X1 exu_U3418(.A(exu_n4014), .B(exu_n9030), .Y(rml_cwp_cwp_output_mux_n44));
AND2X1 exu_U3419(.A(exu_n4015), .B(exu_n9031), .Y(rml_cwp_cwp_output_mux_n43));
AND2X1 exu_U3420(.A(exu_n16196), .B(exu_n15398), .Y(ecl_writeback_ecl_sel_mul_g));
AND2X1 exu_U3421(.A(ecl_div_sel_div), .B(exu_n15398), .Y(ecl_writeback_ecl_sel_div_g));
AND2X1 exu_U3422(.A(ecl_eccctl_ecc_rd_mux_n17), .B(exu_n9072), .Y(ecl_eccctl_wb_rd_m[0]));
AND2X1 exu_U3423(.A(exu_n4078), .B(exu_n9073), .Y(ecl_eccctl_ecc_rd_mux_n17));
AND2X1 exu_U3424(.A(ecl_eccctl_ecc_rd_mux_n13), .B(exu_n9070), .Y(ecl_eccctl_wb_rd_m[1]));
AND2X1 exu_U3425(.A(exu_n4077), .B(exu_n9071), .Y(ecl_eccctl_ecc_rd_mux_n13));
AND2X1 exu_U3426(.A(ecl_eccctl_ecc_rd_mux_n9), .B(exu_n9068), .Y(ecl_eccctl_wb_rd_m[2]));
AND2X1 exu_U3427(.A(exu_n4076), .B(exu_n9069), .Y(ecl_eccctl_ecc_rd_mux_n9));
AND2X1 exu_U3428(.A(ecl_eccctl_ecc_rd_mux_n5), .B(exu_n9066), .Y(ecl_eccctl_wb_rd_m[3]));
AND2X1 exu_U3429(.A(exu_n4075), .B(exu_n9067), .Y(ecl_eccctl_ecc_rd_mux_n5));
AND2X1 exu_U3430(.A(exu_n4074), .B(exu_n9065), .Y(ecl_eccctl_ecc_rd_mux_n1));
AND2X1 exu_U3431(.A(rml_tid_e[1]), .B(exu_n16570), .Y(rml_cwp_thr_e[2]));
AND2X1 exu_U3432(.A(rml_tid_e[1]), .B(rml_tid_e[0]), .Y(rml_cwp_thr_e[3]));
INVX1 exu_U3433(.A(ecl_divcntl_cntr[3]), .Y(exu_n16623));
OR2X1 exu_U3434(.A(ecl_divcntl_cntr[1]), .B(exu_n16438), .Y(ecl_divcntl_cnt6_n31));
INVX1 exu_U3435(.A(ecl_divcntl_cntr[2]), .Y(exu_n16622));
INVX1 exu_U3436(.A(ecl_divcntl_cntr[0]), .Y(exu_n16621));
OR2X1 exu_U3437(.A(rml_cwp_swap_slot3_state[1]), .B(rml_cwp_swap_slot3_state_valid[0]), .Y(rml_cwp_swap_req_vec[3]));
AND2X1 exu_U3438(.A(exu_n16625), .B(exu_n16626), .Y(rml_cwp_cwp_output_queue_n20));
OR2X1 exu_U3439(.A(rml_cwp_swap_slot2_state[1]), .B(rml_cwp_swap_slot2_state_valid[0]), .Y(rml_cwp_swap_req_vec[2]));
AND2X1 exu_U3440(.A(rml_cwp_cwp_output_queue_n26), .B(exu_n9048), .Y(rml_cwp_cwp_output_queue_n25));
OR2X1 exu_U3441(.A(rml_cwp_swap_slot1_state[1]), .B(rml_cwp_swap_slot1_state_valid[0]), .Y(rml_cwp_swap_req_vec[1]));
AND2X1 exu_U3442(.A(exu_n16624), .B(exu_n16511), .Y(rml_cwp_cwp_output_queue_n30));
AND2X1 exu_U3443(.A(exu_n16616), .B(exu_n9050), .Y(rml_cwp_cwp_output_queue_n26));
AND2X1 exu_U3444(.A(exu_n11558), .B(exu_n9052), .Y(rml_cwp_cwp_output_queue_n35));
INVX1 exu_U3445(.A(rml_cwp_swap_tid[1]), .Y(exu_n16620));
INVX1 exu_U3446(.A(rml_cwp_swap_tid[0]), .Y(exu_n16619));
AND2X1 exu_U3447(.A(exu_n4004), .B(exu_n9020), .Y(rml_cwp_cwp_output_mux_n14));
AND2X1 exu_U3448(.A(exu_n4018), .B(exu_n9034), .Y(rml_cwp_cwp_output_mux_n56));
AND2X1 exu_U3449(.A(exu_n4019), .B(exu_n9035), .Y(rml_cwp_cwp_output_mux_n55));
INVX1 exu_U3450(.A(se), .Y(exu_n18474));
INVX1 exu_U3451(.A(exu_n18474), .Y(exu_n16000));
INVX1 exu_U3452(.A(exu_n18474), .Y(exu_n16001));
INVX1 exu_U3453(.A(exu_n18474), .Y(exu_n16002));
INVX1 exu_U3454(.A(exu_n15821), .Y(exu_n16556));
AND2X1 exu_U3455(.A(exu_n4578), .B(exu_n9358), .Y(ecl_yreg0_mux_n2));
AND2X1 exu_U3456(.A(ecl_n84), .B(exu_n9662), .Y(ecl_n83));
AND2X1 exu_U3457(.A(exu_n4964), .B(exu_n9663), .Y(ecl_n84));
AND2X1 exu_U3458(.A(ecl_n88), .B(exu_n9664), .Y(ecl_n82));
AND2X1 exu_U3459(.A(exu_n4965), .B(exu_n9666), .Y(ecl_n88));
INVX1 exu_U3460(.A(rml_ecl_clean_window_e), .Y(exu_n16392));
AND2X1 exu_U3461(.A(ifu_exu_flushw_e), .B(exu_n9619), .Y(rml_n52));
OR2X1 exu_U3462(.A(exu_n13444), .B(exu_n14766), .Y(ecl_writeback_n135));
AND2X1 exu_U3463(.A(exu_n4901), .B(exu_n9617), .Y(rml_n103));
INVX1 exu_U3464(.A(ifu_exu_restored_e), .Y(exu_n16385));
INVX1 exu_U3465(.A(ifu_exu_saved_e), .Y(exu_n16383));
AND2X1 exu_U3466(.A(exu_n4544), .B(exu_n15768), .Y(ecl_writeback_n153));
AND2X1 exu_U3467(.A(ecl_writeback_n55), .B(exu_n9329), .Y(ecl_writeback_n44));
AND2X1 exu_U3468(.A(exu_n16553), .B(ecl_writeback_n58), .Y(ecl_writeback_n55));
OR2X1 exu_U3469(.A(ecl_writeback_return_e), .B(ecl_wb_e), .Y(ecl_writeback_n68));
INVX1 exu_U3470(.A(ecl_restore_e), .Y(exu_n16611));
AND2X1 exu_U3471(.A(exu_n4885), .B(exu_n9609), .Y(rml_ecl_rmlop_done_e));
OR2X1 exu_U3472(.A(exu_n15767), .B(ecl_byplog_rs1_n28), .Y(ecl_byplog_rs1_n19));
OR2X1 exu_U3473(.A(exu_n15345), .B(exu_n15769), .Y(ecl_byplog_rs1_n28));
AND2X1 exu_U3474(.A(exu_n15820), .B(ecl_byplog_rs2_n21), .Y(ecl_byplog_rs2_n18));
AND2X1 exu_U3475(.A(exu_n15818), .B(exu_n19192), .Y(exu_n19189));
AND2X1 exu_U3476(.A(exu_n19194), .B(exu_n19195), .Y(exu_n19190));
AND2X1 exu_U3477(.A(exu_n15433), .B(exu_n15421), .Y(exu_n19194));
AND2X1 exu_U3478(.A(exu_n4543), .B(ecl_wb_byplog_wen_g2), .Y(ecl_writeback_n51));
OR2X1 exu_U3479(.A(ecl_writeback_restore_w), .B(ecl_writeback_restore_ready), .Y(ecl_writeback_n54));
AND2X1 exu_U3480(.A(exu_n4588), .B(exu_n9374), .Y(ecc_chk_rs1_n6));
AND2X1 exu_U3481(.A(ecl_eccctl_n30), .B(ecl_rs1_vld_e), .Y(ecl_ecc_rs1_use_rf_e));
AND2X1 exu_U3482(.A(ecl_eccctl_rs1_sel_rf_e), .B(ifu_exu_inst_vld_e), .Y(ecl_eccctl_n30));
AND2X1 exu_U3483(.A(exu_n783), .B(exu_n5545), .Y(exu_n19999));
AND2X1 exu_U3484(.A(ecl_eccctl_n29), .B(ecl_rs2_vld_e), .Y(ecl_ecc_rs2_use_rf_e));
AND2X1 exu_U3485(.A(ecl_eccctl_rs2_sel_rf_e), .B(ifu_exu_inst_vld_e), .Y(ecl_eccctl_n29));
AND2X1 exu_U3486(.A(exu_n785), .B(exu_n5546), .Y(exu_n20135));
INVX1 exu_U3487(.A(ecc_chk_rs3_parity), .Y(exu_n16513));
AND2X1 exu_U3488(.A(ecl_eccctl_n28), .B(ecl_rs3_vld_e), .Y(ecl_ecc_rs3_use_rf_e));
AND2X1 exu_U3489(.A(ecl_eccctl_rs3_sel_rf_e), .B(ifu_exu_inst_vld_e), .Y(ecl_eccctl_n28));
INVX1 exu_U3490(.A(ecl_cancel_rs3_ecc_e), .Y(exu_n16394));
OR2X1 exu_U3491(.A(exu_n13433), .B(exu_n14752), .Y(ecl_divcntl_firstlast_sub));
AND2X1 exu_U3492(.A(exu_n16583), .B(ecl_divcntl_muls_rs1_data_31_w), .Y(ecl_divcntl_n43));
INVX1 exu_U3493(.A(ecl_divcntl_div_adder_out_31_w), .Y(exu_n16583));
OR2X1 exu_U3494(.A(exu_n13498), .B(exu_n14815), .Y(div_ecl_detect_zero_high));
INVX1 exu_U3495(.A(ifu_exu_inst_vld_w), .Y(exu_n16390));
AND2X1 exu_U3496(.A(exu_n15458), .B(exu_n9306), .Y(ecl_mdqctl_n20));
AND2X1 exu_U3497(.A(exu_n247), .B(exu_n5174), .Y(exu_n17782));
AND2X1 exu_U3498(.A(exu_n246), .B(exu_n5173), .Y(exu_n17783));
OR2X1 exu_U3499(.A(exu_n12100), .B(exu_n13516), .Y(rml_cwp_trap_old_cwp_m[1]));
AND2X1 exu_U3500(.A(exu_n249), .B(exu_n5176), .Y(exu_n17788));
OR2X1 exu_U3501(.A(exu_n12101), .B(exu_n13517), .Y(rml_cwp_trap_old_cwp_m[0]));
AND2X1 exu_U3502(.A(exu_n251), .B(exu_n5178), .Y(exu_n17794));
OR2X1 exu_U3503(.A(exu_n12129), .B(exu_n13545), .Y(rml_ecl_wstate_d[2]));
AND2X1 exu_U3504(.A(exu_n307), .B(exu_n5234), .Y(exu_n17962));
OR2X1 exu_U3505(.A(exu_n12130), .B(exu_n13546), .Y(rml_ecl_wstate_d[1]));
AND2X1 exu_U3506(.A(exu_n309), .B(exu_n5236), .Y(exu_n17968));
INVX1 exu_U3507(.A(rml_rml_ecl_other_d), .Y(exu_n16572));
OR2X1 exu_U3508(.A(exu_n12131), .B(exu_n13547), .Y(rml_ecl_wstate_d[0]));
AND2X1 exu_U3509(.A(exu_n311), .B(exu_n5238), .Y(exu_n17974));
AND2X1 exu_U3510(.A(exu_n452), .B(exu_n5300), .Y(exu_n18423));
INVX1 exu_U3511(.A(rml_cansave_wen_e), .Y(exu_n16382));
INVX1 exu_U3512(.A(rml_rml_ecl_cansave_e[0]), .Y(exu_n16589));
AND2X1 exu_U3513(.A(exu_n453), .B(exu_n5301), .Y(exu_n18428));
INVX1 exu_U3514(.A(rml_canrestore_wen_e), .Y(exu_n16384));
INVX1 exu_U3515(.A(rml_rml_ecl_canrestore_e[0]), .Y(exu_n16588));
INVX1 exu_U3516(.A(rml_rml_ecl_otherwin_e[0]), .Y(exu_n16587));
INVX1 exu_U3517(.A(rml_rml_ecl_cleanwin_e[2]), .Y(exu_n16586));
AND2X1 exu_U3518(.A(exu_n276), .B(exu_n5203), .Y(exu_n17873));
AND2X1 exu_U3519(.A(exu_n278), .B(exu_n5205), .Y(exu_n17879));
AND2X1 exu_U3520(.A(exu_n280), .B(exu_n5207), .Y(exu_n17885));
AND2X1 exu_U3521(.A(exu_n282), .B(exu_n5209), .Y(exu_n17891));
AND2X1 exu_U3522(.A(exu_n284), .B(exu_n5211), .Y(exu_n17897));
AND2X1 exu_U3523(.A(exu_n286), .B(exu_n5213), .Y(exu_n17903));
AND2X1 exu_U3524(.A(exu_n288), .B(exu_n5215), .Y(exu_n17909));
AND2X1 exu_U3525(.A(exu_n290), .B(exu_n5217), .Y(exu_n17915));
AND2X1 exu_U3526(.A(exu_n292), .B(exu_n5219), .Y(exu_n17921));
AND2X1 exu_U3527(.A(exu_n294), .B(exu_n5221), .Y(exu_n17927));
AND2X1 exu_U3528(.A(exu_n296), .B(exu_n5223), .Y(exu_n17933));
AND2X1 exu_U3529(.A(exu_n298), .B(exu_n5225), .Y(exu_n17939));
AND2X1 exu_U3530(.A(exu_n16505), .B(exu_n9313), .Y(ecl_divcntl_wb_req_g));
AND2X1 exu_U3531(.A(exu_n234), .B(exu_n5161), .Y(exu_n17747));
AND2X1 exu_U3532(.A(exu_n236), .B(exu_n5163), .Y(exu_n17753));
AND2X1 exu_U3533(.A(exu_n238), .B(exu_n5165), .Y(exu_n17759));
AND2X1 exu_U3534(.A(exu_n3810), .B(exu_n8889), .Y(div_adderin1[31]));
AND2X1 exu_U3535(.A(exu_n52), .B(exu_n5019), .Y(exu_n16880));
AND2X1 exu_U3536(.A(exu_n15475), .B(exu_n15960), .Y(rml_cwp_n94));
OR2X1 exu_U3537(.A(exu_n15216), .B(exu_n14746), .Y(rml_cwp_cwp_wen_tlu_w[0]));
AND2X1 exu_U3538(.A(exu_n15216), .B(exu_n9122), .Y(rml_cwp_cwp_next0_mux_sel0));
AND2X1 exu_U3539(.A(exu_n256), .B(exu_n5183), .Y(exu_n17813));
AND2X1 exu_U3540(.A(exu_n15474), .B(exu_n15958), .Y(rml_cwp_n93));
OR2X1 exu_U3541(.A(exu_n15215), .B(exu_n14745), .Y(rml_cwp_cwp_wen_tlu_w[1]));
AND2X1 exu_U3542(.A(exu_n15215), .B(exu_n9123), .Y(rml_cwp_cwp_next1_mux_sel0));
AND2X1 exu_U3543(.A(exu_n262), .B(exu_n5189), .Y(exu_n17831));
AND2X1 exu_U3544(.A(exu_n15473), .B(ecl_rml_thr_w[2]), .Y(rml_cwp_n92));
OR2X1 exu_U3545(.A(exu_n15214), .B(exu_n14744), .Y(rml_cwp_cwp_wen_tlu_w[2]));
AND2X1 exu_U3546(.A(exu_n15214), .B(exu_n9124), .Y(rml_cwp_cwp_next2_mux_sel0));
AND2X1 exu_U3547(.A(exu_n268), .B(exu_n5195), .Y(exu_n17849));
OR2X1 exu_U3548(.A(exu_n13401), .B(exu_n14712), .Y(rml_cwp_new_swap_cwp[2]));
AND2X1 exu_U3549(.A(exu_n4009), .B(exu_n9025), .Y(rml_cwp_cwp_output_mux_n25));
AND2X1 exu_U3550(.A(exu_n15472), .B(ecl_rml_thr_w[3]), .Y(rml_cwp_n91));
OR2X1 exu_U3551(.A(exu_n15213), .B(exu_n14743), .Y(rml_cwp_cwp_wen_tlu_w[3]));
AND2X1 exu_U3552(.A(exu_n15213), .B(exu_n9125), .Y(rml_cwp_cwp_next3_mux_sel0));
AND2X1 exu_U3553(.A(exu_n274), .B(exu_n5201), .Y(exu_n17867));
OR2X1 exu_U3554(.A(tlu_exu_agp[1]), .B(exu_n16556), .Y(rml_new_agp[1]));
OR2X1 exu_U3555(.A(tlu_exu_agp[0]), .B(exu_n16556), .Y(rml_new_agp[0]));
AND2X1 exu_U3556(.A(exu_n4890), .B(exu_n15355), .Y(rml_n70));
AND2X1 exu_U3557(.A(exu_n3999), .B(exu_n9015), .Y(exu_n31699));
AND2X1 exu_U3558(.A(exu_n3998), .B(exu_n9014), .Y(exu_n31700));
AND2X1 exu_U3559(.A(exu_n3995), .B(exu_n9012), .Y(exu_n31694));
AND2X1 exu_U3560(.A(exu_n3991), .B(exu_n9007), .Y(exu_n31681));
AND2X1 exu_U3561(.A(exu_n1), .B(exu_n9009), .Y(exu_n31687));
AND2X1 exu_U3562(.A(exu_n4419), .B(exu_n9266), .Y(div_low32or_n11));
AND2X1 exu_U3563(.A(exu_n4418), .B(exu_n9265), .Y(div_low32or_n12));
AND2X1 exu_U3564(.A(exu_n4415), .B(exu_n9263), .Y(div_low32or_n6));
AND2X1 exu_U3565(.A(exu_n4424), .B(exu_n9271), .Y(div_low32or_n25));
AND2X1 exu_U3566(.A(exu_n4423), .B(exu_n9270), .Y(div_low32or_n26));
AND2X1 exu_U3567(.A(exu_n4420), .B(exu_n9268), .Y(div_low32or_n20));
OR2X1 exu_U3568(.A(exu_n13400), .B(exu_n14711), .Y(rml_cwp_swap_data[6]));
AND2X1 exu_U3569(.A(exu_n4007), .B(exu_n9023), .Y(rml_cwp_cwp_output_mux_n19));
AND2X1 exu_U3570(.A(exu_n16396), .B(rml_cwp_swap_thr[3]), .Y(rml_cwp_swap_sel[3]));
AND2X1 exu_U3571(.A(exu_n16396), .B(rml_cwp_swap_thr[1]), .Y(rml_cwp_swap_sel[1]));
AND2X1 exu_U3572(.A(exu_n4939), .B(exu_n9651), .Y(alu_n100));
AND2X1 exu_U3573(.A(exu_n4944), .B(exu_n9656), .Y(alu_n99));
OR2X1 exu_U3574(.A(exu_n15682), .B(alu_logic_rs1_data_bf1[63]), .Y(exu_n17358));
AND2X1 exu_U3575(.A(exu_n4929), .B(exu_n9640), .Y(alu_n70));
AND2X1 exu_U3576(.A(exu_n4934), .B(exu_n9645), .Y(alu_n69));
AND2X1 exu_U3577(.A(alu_ecl_adderin2_31_e), .B(ecl_n144), .Y(ecl_n141));
INVX1 exu_U3578(.A(tlu_exu_cwpccr_update_m), .Y(exu_n16319));
AND2X1 exu_U3579(.A(exu_n15960), .B(ecl_ccr_n20), .Y(ecl_ccr_wen_thr0_w));
AND2X1 exu_U3580(.A(exu_n15926), .B(exu_n15469), .Y(ecl_ccr_n20));
AND2X1 exu_U3581(.A(exu_n4558), .B(exu_n15469), .Y(ecl_ccr_mux_ccrin0_sel2));
AND2X1 exu_U3582(.A(exu_n15958), .B(ecl_ccr_n18), .Y(ecl_ccr_wen_thr1_w));
AND2X1 exu_U3583(.A(exu_n15926), .B(exu_n15468), .Y(ecl_ccr_n18));
AND2X1 exu_U3584(.A(exu_n4556), .B(exu_n15468), .Y(ecl_ccr_mux_ccrin1_sel2));
AND2X1 exu_U3585(.A(ecl_rml_thr_w[2]), .B(ecl_ccr_n16), .Y(ecl_ccr_wen_thr2_w));
AND2X1 exu_U3586(.A(exu_n15926), .B(exu_n15467), .Y(ecl_ccr_n16));
AND2X1 exu_U3587(.A(exu_n4554), .B(exu_n15467), .Y(ecl_ccr_mux_ccrin2_sel2));
AND2X1 exu_U3588(.A(exu_n385), .B(exu_n5296), .Y(ecl_ccr_exu_ifu_cc_w[7]));
AND2X1 exu_U3589(.A(exu_n15198), .B(ecl_divcntl_n68), .Y(ecl_divcntl_ccr_cc_w2[7]));
AND2X1 exu_U3590(.A(exu_n15684), .B(exu_n16558), .Y(ecl_divcntl_n68));
AND2X1 exu_U3591(.A(exu_n16557), .B(ecl_divcntl_n70), .Y(ecl_divcntl_ccr_cc_w2[6]));
AND2X1 exu_U3592(.A(exu_n384), .B(exu_n5295), .Y(ecl_ccr_exu_ifu_cc_w[6]));
AND2X1 exu_U3593(.A(exu_n383), .B(exu_n5294), .Y(ecl_ccr_exu_ifu_cc_w[5]));
AND2X1 exu_U3594(.A(exu_n382), .B(exu_n5293), .Y(ecl_ccr_exu_ifu_cc_w[4]));
AND2X1 exu_U3595(.A(ecl_divcntl_n72), .B(exu_n9314), .Y(ecl_divcntl_ccr_cc_w2[3]));
AND2X1 exu_U3596(.A(exu_n381), .B(exu_n5292), .Y(ecl_ccr_exu_ifu_cc_w[3]));
OR2X1 exu_U3597(.A(exu_n15388), .B(exu_n14753), .Y(ecl_divcntl_ccr_cc_w2[2]));
AND2X1 exu_U3598(.A(exu_n380), .B(exu_n5291), .Y(ecl_ccr_exu_ifu_cc_w[2]));
AND2X1 exu_U3599(.A(exu_n4515), .B(exu_n15684), .Y(ecl_divcntl_n74));
AND2X1 exu_U3600(.A(exu_n379), .B(exu_n5290), .Y(ecl_ccr_exu_ifu_cc_w[1]));
AND2X1 exu_U3601(.A(ecl_ccr_thr_w2[0]), .B(ecl_ccr_setcc_w2), .Y(ecl_ccr_n28));
AND2X1 exu_U3602(.A(ecl_divcntl_muls_c), .B(ecl_divcntl_n84), .Y(ecl_divcntl_ccr_cc_w2[0]));
AND2X1 exu_U3603(.A(ecl_rml_thr_w[3]), .B(ecl_ccr_n13), .Y(ecl_ccr_wen_thr3_w));
AND2X1 exu_U3604(.A(exu_n15926), .B(exu_n15466), .Y(ecl_ccr_n13));
AND2X1 exu_U3605(.A(exu_n378), .B(exu_n5289), .Y(ecl_ccr_exu_ifu_cc_w[0]));
AND2X1 exu_U3606(.A(exu_n4552), .B(exu_n15466), .Y(ecl_ccr_mux_ccrin3_sel2));
AND2X1 exu_U3607(.A(exu_n300), .B(exu_n5227), .Y(exu_n17945));
AND2X1 exu_U3608(.A(exu_n302), .B(exu_n5229), .Y(exu_n17951));
INVX1 exu_U3609(.A(ifu_tlu_sraddr_d[2]), .Y(exu_n16374));
AND2X1 exu_U3610(.A(exu_n304), .B(exu_n5231), .Y(exu_n17957));
OR2X1 exu_U3611(.A(exu_n13412), .B(exu_n14725), .Y(ecl_writeback_rdpr_mux1_out[2]));
AND2X1 exu_U3612(.A(exu_n4080), .B(exu_n9075), .Y(ecl_writeback_rdpr_mux1_n1));
OR2X1 exu_U3613(.A(exu_n13413), .B(exu_n14726), .Y(ecl_writeback_rdpr_mux1_out[1]));
AND2X1 exu_U3614(.A(exu_n4082), .B(exu_n9077), .Y(ecl_writeback_rdpr_mux1_n7));
AND2X1 exu_U3615(.A(exu_n4531), .B(ifu_tlu_sraddr_d[3]), .Y(ecl_writeback_rdpr_mux2_sel3));
AND2X1 exu_U3616(.A(ecl_writeback_n91), .B(exu_n15354), .Y(ecl_writeback_n89));
OR2X1 exu_U3617(.A(exu_n13414), .B(exu_n14727), .Y(ecl_writeback_rdpr_mux1_out[0]));
AND2X1 exu_U3618(.A(exu_n4084), .B(exu_n9079), .Y(ecl_writeback_rdpr_mux1_n13));
OR2X1 exu_U3619(.A(exu_n15390), .B(exu_n14762), .Y(ecl_writeback_sel_cwp_d));
INVX1 exu_U3620(.A(exu_n21628), .Y(exu_n16009));
INVX1 exu_U3621(.A(se), .Y(exu_n21628));
INVX1 exu_U3622(.A(exu_n21661), .Y(exu_n16013));
INVX1 exu_U3623(.A(se), .Y(exu_n21661));
INVX1 exu_U3624(.A(ecl_mdqctl_wb_divthr_g[0]), .Y(exu_n16506));
INVX1 exu_U3625(.A(exu_n21694), .Y(exu_n16017));
INVX1 exu_U3626(.A(se), .Y(exu_n21694));
INVX1 exu_U3627(.A(ecl_mdqctl_wb_divthr_g[1]), .Y(exu_n16507));
INVX1 exu_U3628(.A(exu_n21727), .Y(exu_n16021));
INVX1 exu_U3629(.A(se), .Y(exu_n21727));
AND2X1 exu_U3630(.A(ecl_mdqctl_wb_divthr_g[1]), .B(ecl_mdqctl_wb_divthr_g[0]), .Y(ecl_writeback_n192));
INVX1 exu_U3631(.A(exu_n21760), .Y(exu_n16025));
INVX1 exu_U3632(.A(se), .Y(exu_n21760));
OR2X1 exu_U3633(.A(exu_n12918), .B(exu_n14202), .Y(alu_byp_rd_data_e[63]));
AND2X1 exu_U3634(.A(exu_n2576), .B(exu_n9673), .Y(exu_n26377));
OR2X1 exu_U3635(.A(exu_n12919), .B(exu_n14203), .Y(alu_byp_rd_data_e[62]));
AND2X1 exu_U3636(.A(exu_n2578), .B(exu_n7605), .Y(exu_n26382));
OR2X1 exu_U3637(.A(exu_n12920), .B(exu_n14204), .Y(alu_byp_rd_data_e[61]));
AND2X1 exu_U3638(.A(exu_n2580), .B(exu_n7607), .Y(exu_n26388));
OR2X1 exu_U3639(.A(exu_n12921), .B(exu_n14205), .Y(alu_byp_rd_data_e[60]));
AND2X1 exu_U3640(.A(exu_n2582), .B(exu_n7609), .Y(exu_n26394));
OR2X1 exu_U3641(.A(exu_n12923), .B(exu_n14207), .Y(alu_byp_rd_data_e[59]));
AND2X1 exu_U3642(.A(exu_n2586), .B(exu_n7613), .Y(exu_n26406));
OR2X1 exu_U3643(.A(exu_n12924), .B(exu_n14208), .Y(alu_byp_rd_data_e[58]));
AND2X1 exu_U3644(.A(exu_n2588), .B(exu_n7615), .Y(exu_n26412));
OR2X1 exu_U3645(.A(exu_n12925), .B(exu_n14209), .Y(alu_byp_rd_data_e[57]));
AND2X1 exu_U3646(.A(exu_n2590), .B(exu_n7617), .Y(exu_n26418));
OR2X1 exu_U3647(.A(exu_n12926), .B(exu_n14210), .Y(alu_byp_rd_data_e[56]));
AND2X1 exu_U3648(.A(exu_n2592), .B(exu_n7619), .Y(exu_n26424));
OR2X1 exu_U3649(.A(exu_n12927), .B(exu_n14211), .Y(alu_byp_rd_data_e[55]));
AND2X1 exu_U3650(.A(exu_n2594), .B(exu_n7621), .Y(exu_n26430));
OR2X1 exu_U3651(.A(exu_n12928), .B(exu_n14212), .Y(alu_byp_rd_data_e[54]));
AND2X1 exu_U3652(.A(exu_n2596), .B(exu_n7623), .Y(exu_n26436));
OR2X1 exu_U3653(.A(exu_n12929), .B(exu_n14213), .Y(alu_byp_rd_data_e[53]));
AND2X1 exu_U3654(.A(exu_n2598), .B(exu_n7625), .Y(exu_n26442));
OR2X1 exu_U3655(.A(exu_n12930), .B(exu_n14214), .Y(alu_byp_rd_data_e[52]));
AND2X1 exu_U3656(.A(exu_n2600), .B(exu_n7627), .Y(exu_n26448));
OR2X1 exu_U3657(.A(exu_n12931), .B(exu_n14215), .Y(alu_byp_rd_data_e[51]));
AND2X1 exu_U3658(.A(exu_n2602), .B(exu_n7629), .Y(exu_n26454));
OR2X1 exu_U3659(.A(exu_n12932), .B(exu_n14216), .Y(alu_byp_rd_data_e[50]));
AND2X1 exu_U3660(.A(exu_n2604), .B(exu_n7631), .Y(exu_n26460));
OR2X1 exu_U3661(.A(exu_n12934), .B(exu_n14218), .Y(alu_byp_rd_data_e[49]));
AND2X1 exu_U3662(.A(exu_n2608), .B(exu_n7635), .Y(exu_n26472));
OR2X1 exu_U3663(.A(exu_n12935), .B(exu_n14219), .Y(alu_byp_rd_data_e[48]));
AND2X1 exu_U3664(.A(exu_n2610), .B(exu_n7637), .Y(exu_n26478));
OR2X1 exu_U3665(.A(exu_n12936), .B(exu_n14220), .Y(alu_byp_rd_data_e[47]));
AND2X1 exu_U3666(.A(exu_n2612), .B(exu_n7639), .Y(exu_n26484));
OR2X1 exu_U3667(.A(exu_n12937), .B(exu_n14221), .Y(alu_byp_rd_data_e[46]));
AND2X1 exu_U3668(.A(exu_n2614), .B(exu_n7641), .Y(exu_n26490));
OR2X1 exu_U3669(.A(exu_n12938), .B(exu_n14222), .Y(alu_byp_rd_data_e[45]));
AND2X1 exu_U3670(.A(exu_n2616), .B(exu_n7643), .Y(exu_n26496));
OR2X1 exu_U3671(.A(exu_n12939), .B(exu_n14223), .Y(alu_byp_rd_data_e[44]));
AND2X1 exu_U3672(.A(exu_n2618), .B(exu_n7645), .Y(exu_n26502));
OR2X1 exu_U3673(.A(exu_n12940), .B(exu_n14224), .Y(alu_byp_rd_data_e[43]));
AND2X1 exu_U3674(.A(exu_n2620), .B(exu_n7647), .Y(exu_n26508));
OR2X1 exu_U3675(.A(exu_n12941), .B(exu_n14225), .Y(alu_byp_rd_data_e[42]));
AND2X1 exu_U3676(.A(exu_n2622), .B(exu_n7649), .Y(exu_n26514));
OR2X1 exu_U3677(.A(exu_n12942), .B(exu_n14226), .Y(alu_byp_rd_data_e[41]));
AND2X1 exu_U3678(.A(exu_n2624), .B(exu_n7651), .Y(exu_n26520));
OR2X1 exu_U3679(.A(exu_n12943), .B(exu_n14227), .Y(alu_byp_rd_data_e[40]));
AND2X1 exu_U3680(.A(exu_n2626), .B(exu_n7653), .Y(exu_n26526));
OR2X1 exu_U3681(.A(exu_n12945), .B(exu_n14229), .Y(alu_byp_rd_data_e[39]));
AND2X1 exu_U3682(.A(exu_n2630), .B(exu_n7657), .Y(exu_n26538));
OR2X1 exu_U3683(.A(exu_n12946), .B(exu_n14230), .Y(alu_byp_rd_data_e[38]));
AND2X1 exu_U3684(.A(exu_n2632), .B(exu_n7659), .Y(exu_n26544));
OR2X1 exu_U3685(.A(exu_n12947), .B(exu_n14231), .Y(alu_byp_rd_data_e[37]));
AND2X1 exu_U3686(.A(exu_n2634), .B(exu_n7661), .Y(exu_n26550));
OR2X1 exu_U3687(.A(exu_n12948), .B(exu_n14232), .Y(alu_byp_rd_data_e[36]));
AND2X1 exu_U3688(.A(exu_n2636), .B(exu_n7663), .Y(exu_n26556));
OR2X1 exu_U3689(.A(exu_n12949), .B(exu_n14233), .Y(alu_byp_rd_data_e[35]));
AND2X1 exu_U3690(.A(exu_n2638), .B(exu_n7665), .Y(exu_n26562));
OR2X1 exu_U3691(.A(exu_n12950), .B(exu_n14234), .Y(alu_byp_rd_data_e[34]));
AND2X1 exu_U3692(.A(exu_n2640), .B(exu_n7667), .Y(exu_n26568));
OR2X1 exu_U3693(.A(exu_n12951), .B(exu_n14235), .Y(alu_byp_rd_data_e[33]));
AND2X1 exu_U3694(.A(exu_n2642), .B(exu_n7669), .Y(exu_n26574));
OR2X1 exu_U3695(.A(exu_n12952), .B(exu_n14236), .Y(alu_byp_rd_data_e[32]));
AND2X1 exu_U3696(.A(exu_n2644), .B(exu_n7671), .Y(exu_n26580));
AND2X1 exu_U3697(.A(exu_n864), .B(exu_n5625), .Y(exu_n20711));
OR2X1 exu_U3698(.A(exu_n12953), .B(exu_n14237), .Y(alu_byp_rd_data_e[31]));
AND2X1 exu_U3699(.A(exu_n2646), .B(exu_n9674), .Y(exu_n26586));
AND2X1 exu_U3700(.A(exu_n866), .B(exu_n5627), .Y(exu_n20717));
OR2X1 exu_U3701(.A(exu_n12954), .B(exu_n14238), .Y(alu_byp_rd_data_e[30]));
AND2X1 exu_U3702(.A(exu_n2648), .B(exu_n7674), .Y(exu_n26591));
AND2X1 exu_U3703(.A(exu_n870), .B(exu_n5631), .Y(exu_n20729));
OR2X1 exu_U3704(.A(exu_n12956), .B(exu_n14240), .Y(alu_byp_rd_data_e[29]));
AND2X1 exu_U3705(.A(exu_n2652), .B(exu_n7678), .Y(exu_n26603));
AND2X1 exu_U3706(.A(exu_n872), .B(exu_n5633), .Y(exu_n20735));
OR2X1 exu_U3707(.A(exu_n12957), .B(exu_n14241), .Y(alu_byp_rd_data_e[28]));
AND2X1 exu_U3708(.A(exu_n2654), .B(exu_n7680), .Y(exu_n26609));
AND2X1 exu_U3709(.A(exu_n874), .B(exu_n5635), .Y(exu_n20741));
OR2X1 exu_U3710(.A(exu_n12958), .B(exu_n14242), .Y(alu_byp_rd_data_e[27]));
AND2X1 exu_U3711(.A(exu_n2656), .B(exu_n7682), .Y(exu_n26615));
AND2X1 exu_U3712(.A(exu_n876), .B(exu_n5637), .Y(exu_n20747));
OR2X1 exu_U3713(.A(exu_n12959), .B(exu_n14243), .Y(alu_byp_rd_data_e[26]));
AND2X1 exu_U3714(.A(exu_n2658), .B(exu_n7684), .Y(exu_n26621));
AND2X1 exu_U3715(.A(exu_n878), .B(exu_n5639), .Y(exu_n20753));
OR2X1 exu_U3716(.A(exu_n12960), .B(exu_n14244), .Y(alu_byp_rd_data_e[25]));
AND2X1 exu_U3717(.A(exu_n2660), .B(exu_n7686), .Y(exu_n26627));
AND2X1 exu_U3718(.A(exu_n880), .B(exu_n5641), .Y(exu_n20759));
OR2X1 exu_U3719(.A(exu_n12961), .B(exu_n14245), .Y(alu_byp_rd_data_e[24]));
AND2X1 exu_U3720(.A(exu_n2662), .B(exu_n7688), .Y(exu_n26633));
AND2X1 exu_U3721(.A(exu_n882), .B(exu_n5643), .Y(exu_n20765));
OR2X1 exu_U3722(.A(exu_n12962), .B(exu_n14246), .Y(alu_byp_rd_data_e[23]));
AND2X1 exu_U3723(.A(exu_n2664), .B(exu_n7690), .Y(exu_n26639));
AND2X1 exu_U3724(.A(exu_n884), .B(exu_n5645), .Y(exu_n20771));
OR2X1 exu_U3725(.A(exu_n12963), .B(exu_n14247), .Y(alu_byp_rd_data_e[22]));
AND2X1 exu_U3726(.A(exu_n2666), .B(exu_n7692), .Y(exu_n26645));
AND2X1 exu_U3727(.A(exu_n886), .B(exu_n5647), .Y(exu_n20777));
OR2X1 exu_U3728(.A(exu_n12964), .B(exu_n14248), .Y(alu_byp_rd_data_e[21]));
AND2X1 exu_U3729(.A(exu_n2668), .B(exu_n7694), .Y(exu_n26651));
AND2X1 exu_U3730(.A(exu_n888), .B(exu_n5649), .Y(exu_n20783));
OR2X1 exu_U3731(.A(exu_n12965), .B(exu_n14249), .Y(alu_byp_rd_data_e[20]));
AND2X1 exu_U3732(.A(exu_n2670), .B(exu_n7696), .Y(exu_n26657));
AND2X1 exu_U3733(.A(exu_n892), .B(exu_n5653), .Y(exu_n20795));
OR2X1 exu_U3734(.A(exu_n12967), .B(exu_n14251), .Y(alu_byp_rd_data_e[19]));
AND2X1 exu_U3735(.A(exu_n2674), .B(exu_n7700), .Y(exu_n26669));
AND2X1 exu_U3736(.A(exu_n894), .B(exu_n5655), .Y(exu_n20801));
OR2X1 exu_U3737(.A(exu_n12968), .B(exu_n14252), .Y(alu_byp_rd_data_e[18]));
AND2X1 exu_U3738(.A(exu_n2676), .B(exu_n7702), .Y(exu_n26675));
AND2X1 exu_U3739(.A(exu_n896), .B(exu_n5657), .Y(exu_n20807));
OR2X1 exu_U3740(.A(exu_n12969), .B(exu_n14253), .Y(alu_byp_rd_data_e[17]));
AND2X1 exu_U3741(.A(exu_n2678), .B(exu_n7704), .Y(exu_n26681));
AND2X1 exu_U3742(.A(exu_n898), .B(exu_n5659), .Y(exu_n20813));
OR2X1 exu_U3743(.A(exu_n12970), .B(exu_n14254), .Y(alu_byp_rd_data_e[16]));
AND2X1 exu_U3744(.A(exu_n2680), .B(exu_n7706), .Y(exu_n26687));
AND2X1 exu_U3745(.A(exu_n900), .B(exu_n5661), .Y(exu_n20819));
OR2X1 exu_U3746(.A(exu_n12971), .B(exu_n14255), .Y(alu_byp_rd_data_e[15]));
AND2X1 exu_U3747(.A(exu_n2682), .B(exu_n7708), .Y(exu_n26693));
AND2X1 exu_U3748(.A(exu_n902), .B(exu_n5663), .Y(exu_n20825));
OR2X1 exu_U3749(.A(exu_n12972), .B(exu_n14256), .Y(alu_byp_rd_data_e[14]));
AND2X1 exu_U3750(.A(exu_n2684), .B(exu_n7710), .Y(exu_n26699));
AND2X1 exu_U3751(.A(exu_n904), .B(exu_n5665), .Y(exu_n20831));
OR2X1 exu_U3752(.A(exu_n12973), .B(exu_n14257), .Y(alu_byp_rd_data_e[13]));
AND2X1 exu_U3753(.A(exu_n2686), .B(exu_n7712), .Y(exu_n26705));
AND2X1 exu_U3754(.A(exu_n906), .B(exu_n5667), .Y(exu_n20837));
OR2X1 exu_U3755(.A(exu_n12974), .B(exu_n14258), .Y(alu_byp_rd_data_e[12]));
AND2X1 exu_U3756(.A(exu_n2688), .B(exu_n7714), .Y(exu_n26711));
AND2X1 exu_U3757(.A(exu_n908), .B(exu_n5669), .Y(exu_n20843));
OR2X1 exu_U3758(.A(exu_n12975), .B(exu_n14259), .Y(alu_byp_rd_data_e[11]));
AND2X1 exu_U3759(.A(exu_n2690), .B(exu_n7716), .Y(exu_n26717));
AND2X1 exu_U3760(.A(exu_n910), .B(exu_n5671), .Y(exu_n20849));
OR2X1 exu_U3761(.A(exu_n12976), .B(exu_n14260), .Y(alu_byp_rd_data_e[10]));
AND2X1 exu_U3762(.A(exu_n2692), .B(exu_n7718), .Y(exu_n26723));
AND2X1 exu_U3763(.A(exu_n850), .B(exu_n5611), .Y(exu_n20669));
AND2X1 exu_U3764(.A(exu_n852), .B(exu_n5613), .Y(exu_n20675));
OR2X1 exu_U3765(.A(exu_n12915), .B(exu_n14199), .Y(alu_byp_rd_data_e[8]));
AND2X1 exu_U3766(.A(exu_n2570), .B(exu_n7598), .Y(exu_n26359));
OR2X1 exu_U3767(.A(exu_n12916), .B(exu_n14200), .Y(alu_byp_rd_data_e[7]));
AND2X1 exu_U3768(.A(exu_n2572), .B(exu_n7600), .Y(exu_n26365));
OR2X1 exu_U3769(.A(exu_n12917), .B(exu_n14201), .Y(alu_byp_rd_data_e[6]));
AND2X1 exu_U3770(.A(exu_n2574), .B(exu_n7602), .Y(exu_n26371));
OR2X1 exu_U3771(.A(exu_n12922), .B(exu_n14206), .Y(alu_byp_rd_data_e[5]));
AND2X1 exu_U3772(.A(exu_n2584), .B(exu_n7611), .Y(exu_n26400));
OR2X1 exu_U3773(.A(exu_n12933), .B(exu_n14217), .Y(alu_byp_rd_data_e[4]));
AND2X1 exu_U3774(.A(exu_n2606), .B(exu_n7633), .Y(exu_n26466));
OR2X1 exu_U3775(.A(exu_n12944), .B(exu_n14228), .Y(alu_byp_rd_data_e[3]));
AND2X1 exu_U3776(.A(exu_n2628), .B(exu_n7655), .Y(exu_n26532));
OR2X1 exu_U3777(.A(exu_n12955), .B(exu_n14239), .Y(alu_byp_rd_data_e[2]));
AND2X1 exu_U3778(.A(exu_n2650), .B(exu_n7676), .Y(exu_n26597));
OR2X1 exu_U3779(.A(exu_n12966), .B(exu_n14250), .Y(alu_byp_rd_data_e[1]));
AND2X1 exu_U3780(.A(exu_n2672), .B(exu_n7698), .Y(exu_n26663));
INVX1 exu_U3781(.A(exu_n29301), .Y(exu_n16031));
OR2X1 exu_U3782(.A(exu_n12977), .B(exu_n14261), .Y(alu_byp_rd_data_e[0]));
AND2X1 exu_U3783(.A(exu_n2694), .B(exu_n7720), .Y(exu_n26729));
AND2X1 exu_U3784(.A(exu_n15420), .B(ecl_read_yreg_e), .Y(ecl_byp_sel_eclpr_e));
INVX1 exu_U3785(.A(exu_n29301), .Y(exu_n16032));
INVX1 exu_U3786(.A(exu_n29366), .Y(exu_n16038));
INVX1 exu_U3787(.A(exu_n29366), .Y(exu_n16039));
AND2X1 exu_U3788(.A(bypass_sr_out_mux_n17), .B(exu_n9447), .Y(bypass_full_rd_data_m[63]));
AND2X1 exu_U3789(.A(exu_n1561), .B(exu_n6579), .Y(exu_n23226));
AND2X1 exu_U3790(.A(bypass_sr_out_mux_n21), .B(exu_n9449), .Y(bypass_full_rd_data_m[62]));
AND2X1 exu_U3791(.A(exu_n1563), .B(exu_n6581), .Y(exu_n23232));
AND2X1 exu_U3792(.A(bypass_sr_out_mux_n25), .B(exu_n9451), .Y(bypass_full_rd_data_m[61]));
AND2X1 exu_U3793(.A(exu_n1565), .B(exu_n6583), .Y(exu_n23238));
AND2X1 exu_U3794(.A(bypass_sr_out_mux_n29), .B(exu_n9453), .Y(bypass_full_rd_data_m[60]));
AND2X1 exu_U3795(.A(exu_n1567), .B(exu_n6585), .Y(exu_n23244));
AND2X1 exu_U3796(.A(bypass_sr_out_mux_n37), .B(exu_n9457), .Y(bypass_full_rd_data_m[59]));
AND2X1 exu_U3797(.A(exu_n1571), .B(exu_n6589), .Y(exu_n23256));
AND2X1 exu_U3798(.A(bypass_sr_out_mux_n41), .B(exu_n9459), .Y(bypass_full_rd_data_m[58]));
AND2X1 exu_U3799(.A(exu_n1573), .B(exu_n6591), .Y(exu_n23262));
AND2X1 exu_U3800(.A(bypass_sr_out_mux_n45), .B(exu_n9461), .Y(bypass_full_rd_data_m[57]));
AND2X1 exu_U3801(.A(exu_n1575), .B(exu_n6593), .Y(exu_n23268));
AND2X1 exu_U3802(.A(bypass_sr_out_mux_n49), .B(exu_n9463), .Y(bypass_full_rd_data_m[56]));
AND2X1 exu_U3803(.A(exu_n1577), .B(exu_n6595), .Y(exu_n23274));
AND2X1 exu_U3804(.A(bypass_sr_out_mux_n53), .B(exu_n9465), .Y(bypass_full_rd_data_m[55]));
AND2X1 exu_U3805(.A(exu_n1579), .B(exu_n6597), .Y(exu_n23280));
AND2X1 exu_U3806(.A(bypass_sr_out_mux_n57), .B(exu_n9467), .Y(bypass_full_rd_data_m[54]));
AND2X1 exu_U3807(.A(exu_n1581), .B(exu_n6599), .Y(exu_n23286));
AND2X1 exu_U3808(.A(bypass_sr_out_mux_n61), .B(exu_n9469), .Y(bypass_full_rd_data_m[53]));
AND2X1 exu_U3809(.A(exu_n1583), .B(exu_n6601), .Y(exu_n23292));
AND2X1 exu_U3810(.A(bypass_sr_out_mux_n65), .B(exu_n9471), .Y(bypass_full_rd_data_m[52]));
AND2X1 exu_U3811(.A(exu_n1585), .B(exu_n6603), .Y(exu_n23298));
AND2X1 exu_U3812(.A(bypass_sr_out_mux_n69), .B(exu_n9473), .Y(bypass_full_rd_data_m[51]));
AND2X1 exu_U3813(.A(exu_n1587), .B(exu_n6605), .Y(exu_n23304));
AND2X1 exu_U3814(.A(bypass_sr_out_mux_n73), .B(exu_n9475), .Y(bypass_full_rd_data_m[50]));
AND2X1 exu_U3815(.A(exu_n1589), .B(exu_n6607), .Y(exu_n23310));
AND2X1 exu_U3816(.A(bypass_sr_out_mux_n81), .B(exu_n9479), .Y(bypass_full_rd_data_m[49]));
AND2X1 exu_U3817(.A(exu_n1593), .B(exu_n6611), .Y(exu_n23322));
AND2X1 exu_U3818(.A(bypass_sr_out_mux_n85), .B(exu_n9481), .Y(bypass_full_rd_data_m[48]));
AND2X1 exu_U3819(.A(exu_n1595), .B(exu_n6613), .Y(exu_n23328));
AND2X1 exu_U3820(.A(bypass_sr_out_mux_n89), .B(exu_n9483), .Y(bypass_full_rd_data_m[47]));
AND2X1 exu_U3821(.A(exu_n1597), .B(exu_n6615), .Y(exu_n23334));
AND2X1 exu_U3822(.A(bypass_sr_out_mux_n93), .B(exu_n9485), .Y(bypass_full_rd_data_m[46]));
AND2X1 exu_U3823(.A(exu_n1599), .B(exu_n6617), .Y(exu_n23340));
AND2X1 exu_U3824(.A(bypass_sr_out_mux_n97), .B(exu_n9487), .Y(bypass_full_rd_data_m[45]));
AND2X1 exu_U3825(.A(exu_n1601), .B(exu_n6619), .Y(exu_n23346));
AND2X1 exu_U3826(.A(bypass_sr_out_mux_n101), .B(exu_n9489), .Y(bypass_full_rd_data_m[44]));
AND2X1 exu_U3827(.A(exu_n1603), .B(exu_n6621), .Y(exu_n23352));
AND2X1 exu_U3828(.A(bypass_sr_out_mux_n105), .B(exu_n9491), .Y(bypass_full_rd_data_m[43]));
AND2X1 exu_U3829(.A(exu_n1605), .B(exu_n6623), .Y(exu_n23358));
AND2X1 exu_U3830(.A(bypass_sr_out_mux_n109), .B(exu_n9493), .Y(bypass_full_rd_data_m[42]));
AND2X1 exu_U3831(.A(exu_n1607), .B(exu_n6625), .Y(exu_n23364));
AND2X1 exu_U3832(.A(bypass_sr_out_mux_n113), .B(exu_n9495), .Y(bypass_full_rd_data_m[41]));
AND2X1 exu_U3833(.A(exu_n1609), .B(exu_n6627), .Y(exu_n23370));
AND2X1 exu_U3834(.A(bypass_sr_out_mux_n117), .B(exu_n9497), .Y(bypass_full_rd_data_m[40]));
AND2X1 exu_U3835(.A(exu_n1611), .B(exu_n6629), .Y(exu_n23376));
AND2X1 exu_U3836(.A(bypass_sr_out_mux_n125), .B(exu_n9501), .Y(bypass_full_rd_data_m[39]));
AND2X1 exu_U3837(.A(exu_n1615), .B(exu_n6633), .Y(exu_n23388));
AND2X1 exu_U3838(.A(bypass_sr_out_mux_n129), .B(exu_n9503), .Y(bypass_full_rd_data_m[38]));
AND2X1 exu_U3839(.A(exu_n1617), .B(exu_n6635), .Y(exu_n23394));
AND2X1 exu_U3840(.A(bypass_sr_out_mux_n133), .B(exu_n9505), .Y(bypass_full_rd_data_m[37]));
AND2X1 exu_U3841(.A(exu_n1619), .B(exu_n6637), .Y(exu_n23400));
AND2X1 exu_U3842(.A(bypass_sr_out_mux_n137), .B(exu_n9507), .Y(bypass_full_rd_data_m[36]));
AND2X1 exu_U3843(.A(exu_n1621), .B(exu_n6639), .Y(exu_n23406));
AND2X1 exu_U3844(.A(bypass_sr_out_mux_n141), .B(exu_n9509), .Y(bypass_full_rd_data_m[35]));
AND2X1 exu_U3845(.A(exu_n1623), .B(exu_n6641), .Y(exu_n23412));
AND2X1 exu_U3846(.A(bypass_sr_out_mux_n145), .B(exu_n9511), .Y(bypass_full_rd_data_m[34]));
AND2X1 exu_U3847(.A(exu_n1625), .B(exu_n6643), .Y(exu_n23418));
AND2X1 exu_U3848(.A(bypass_sr_out_mux_n149), .B(exu_n9513), .Y(bypass_full_rd_data_m[33]));
AND2X1 exu_U3849(.A(exu_n1627), .B(exu_n6645), .Y(exu_n23424));
AND2X1 exu_U3850(.A(bypass_sr_out_mux_n153), .B(exu_n9515), .Y(bypass_full_rd_data_m[32]));
AND2X1 exu_U3851(.A(exu_n1629), .B(exu_n6647), .Y(exu_n23430));
AND2X1 exu_U3852(.A(bypass_sr_out_mux_n157), .B(exu_n9517), .Y(bypass_full_rd_data_m[31]));
AND2X1 exu_U3853(.A(exu_n1631), .B(exu_n6649), .Y(exu_n23436));
AND2X1 exu_U3854(.A(bypass_sr_out_mux_n161), .B(exu_n9519), .Y(bypass_full_rd_data_m[30]));
AND2X1 exu_U3855(.A(exu_n1633), .B(exu_n6651), .Y(exu_n23442));
AND2X1 exu_U3856(.A(bypass_sr_out_mux_n169), .B(exu_n9523), .Y(bypass_full_rd_data_m[29]));
AND2X1 exu_U3857(.A(exu_n1637), .B(exu_n6655), .Y(exu_n23454));
AND2X1 exu_U3858(.A(bypass_sr_out_mux_n173), .B(exu_n9525), .Y(bypass_full_rd_data_m[28]));
AND2X1 exu_U3859(.A(exu_n1639), .B(exu_n6657), .Y(exu_n23460));
AND2X1 exu_U3860(.A(bypass_sr_out_mux_n177), .B(exu_n9527), .Y(bypass_full_rd_data_m[27]));
AND2X1 exu_U3861(.A(exu_n1641), .B(exu_n6659), .Y(exu_n23466));
AND2X1 exu_U3862(.A(bypass_sr_out_mux_n181), .B(exu_n9529), .Y(bypass_full_rd_data_m[26]));
AND2X1 exu_U3863(.A(exu_n1643), .B(exu_n6661), .Y(exu_n23472));
AND2X1 exu_U3864(.A(bypass_sr_out_mux_n185), .B(exu_n9531), .Y(bypass_full_rd_data_m[25]));
AND2X1 exu_U3865(.A(exu_n1645), .B(exu_n6663), .Y(exu_n23478));
AND2X1 exu_U3866(.A(bypass_sr_out_mux_n189), .B(exu_n9533), .Y(bypass_full_rd_data_m[24]));
AND2X1 exu_U3867(.A(exu_n1647), .B(exu_n6665), .Y(exu_n23484));
AND2X1 exu_U3868(.A(bypass_sr_out_mux_n193), .B(exu_n9535), .Y(bypass_full_rd_data_m[23]));
AND2X1 exu_U3869(.A(exu_n1649), .B(exu_n6667), .Y(exu_n23490));
AND2X1 exu_U3870(.A(bypass_sr_out_mux_n197), .B(exu_n9537), .Y(bypass_full_rd_data_m[22]));
AND2X1 exu_U3871(.A(exu_n1651), .B(exu_n6669), .Y(exu_n23496));
AND2X1 exu_U3872(.A(bypass_sr_out_mux_n201), .B(exu_n9539), .Y(bypass_full_rd_data_m[21]));
AND2X1 exu_U3873(.A(exu_n1653), .B(exu_n6671), .Y(exu_n23502));
AND2X1 exu_U3874(.A(bypass_sr_out_mux_n205), .B(exu_n9541), .Y(bypass_full_rd_data_m[20]));
AND2X1 exu_U3875(.A(exu_n1655), .B(exu_n6673), .Y(exu_n23508));
AND2X1 exu_U3876(.A(bypass_sr_out_mux_n213), .B(exu_n9545), .Y(bypass_full_rd_data_m[19]));
AND2X1 exu_U3877(.A(exu_n1659), .B(exu_n6677), .Y(exu_n23520));
AND2X1 exu_U3878(.A(bypass_sr_out_mux_n217), .B(exu_n9547), .Y(bypass_full_rd_data_m[18]));
AND2X1 exu_U3879(.A(exu_n1661), .B(exu_n6679), .Y(exu_n23526));
AND2X1 exu_U3880(.A(bypass_sr_out_mux_n221), .B(exu_n9549), .Y(bypass_full_rd_data_m[17]));
AND2X1 exu_U3881(.A(exu_n1663), .B(exu_n6681), .Y(exu_n23532));
AND2X1 exu_U3882(.A(bypass_sr_out_mux_n225), .B(exu_n9551), .Y(bypass_full_rd_data_m[16]));
AND2X1 exu_U3883(.A(exu_n1665), .B(exu_n6683), .Y(exu_n23538));
AND2X1 exu_U3884(.A(bypass_sr_out_mux_n229), .B(exu_n9553), .Y(bypass_full_rd_data_m[15]));
AND2X1 exu_U3885(.A(exu_n1667), .B(exu_n6685), .Y(exu_n23544));
AND2X1 exu_U3886(.A(bypass_sr_out_mux_n233), .B(exu_n9555), .Y(bypass_full_rd_data_m[14]));
AND2X1 exu_U3887(.A(exu_n1669), .B(exu_n6687), .Y(exu_n23550));
AND2X1 exu_U3888(.A(bypass_sr_out_mux_n237), .B(exu_n9557), .Y(bypass_full_rd_data_m[13]));
AND2X1 exu_U3889(.A(exu_n1671), .B(exu_n6689), .Y(exu_n23556));
AND2X1 exu_U3890(.A(bypass_sr_out_mux_n241), .B(exu_n9559), .Y(bypass_full_rd_data_m[12]));
AND2X1 exu_U3891(.A(exu_n1673), .B(exu_n6691), .Y(exu_n23562));
AND2X1 exu_U3892(.A(bypass_sr_out_mux_n245), .B(exu_n9561), .Y(bypass_full_rd_data_m[11]));
AND2X1 exu_U3893(.A(exu_n1675), .B(exu_n6693), .Y(exu_n23568));
AND2X1 exu_U3894(.A(bypass_sr_out_mux_n249), .B(exu_n9563), .Y(bypass_full_rd_data_m[10]));
AND2X1 exu_U3895(.A(exu_n1677), .B(exu_n6695), .Y(exu_n23574));
AND2X1 exu_U3896(.A(exu_n1553), .B(exu_n6571), .Y(exu_n23202));
AND2X1 exu_U3897(.A(bypass_sr_out_mux_n5), .B(exu_n9441), .Y(bypass_full_rd_data_m[8]));
AND2X1 exu_U3898(.A(exu_n1555), .B(exu_n6573), .Y(exu_n23208));
AND2X1 exu_U3899(.A(bypass_sr_out_mux_n9), .B(exu_n9443), .Y(bypass_full_rd_data_m[7]));
AND2X1 exu_U3900(.A(exu_n1557), .B(exu_n6575), .Y(exu_n23214));
AND2X1 exu_U3901(.A(bypass_sr_out_mux_n13), .B(exu_n9445), .Y(bypass_full_rd_data_m[6]));
AND2X1 exu_U3902(.A(exu_n1559), .B(exu_n6577), .Y(exu_n23220));
AND2X1 exu_U3903(.A(bypass_sr_out_mux_n33), .B(exu_n9455), .Y(bypass_full_rd_data_m[5]));
AND2X1 exu_U3904(.A(exu_n1569), .B(exu_n6587), .Y(exu_n23250));
AND2X1 exu_U3905(.A(bypass_sr_out_mux_n77), .B(exu_n9477), .Y(bypass_full_rd_data_m[4]));
AND2X1 exu_U3906(.A(exu_n1591), .B(exu_n6609), .Y(exu_n23316));
AND2X1 exu_U3907(.A(bypass_sr_out_mux_n121), .B(exu_n9499), .Y(bypass_full_rd_data_m[3]));
AND2X1 exu_U3908(.A(exu_n1613), .B(exu_n6631), .Y(exu_n23382));
AND2X1 exu_U3909(.A(bypass_sr_out_mux_n165), .B(exu_n9521), .Y(bypass_full_rd_data_m[2]));
AND2X1 exu_U3910(.A(exu_n1635), .B(exu_n6653), .Y(exu_n23448));
AND2X1 exu_U3911(.A(bypass_sr_out_mux_n209), .B(exu_n9543), .Y(bypass_full_rd_data_m[1]));
AND2X1 exu_U3912(.A(exu_n1657), .B(exu_n6675), .Y(exu_n23514));
INVX1 exu_U3913(.A(exu_n29431), .Y(exu_n16045));
AND2X1 exu_U3914(.A(bypass_sr_out_mux_n253), .B(exu_n9565), .Y(bypass_full_rd_data_m[0]));
AND2X1 exu_U3915(.A(exu_n1679), .B(exu_n6697), .Y(exu_n23580));
INVX1 exu_U3916(.A(exu_n29431), .Y(exu_n16046));
AND2X1 exu_U3917(.A(exu_n11369), .B(exu_n8790), .Y(div_byp_muldivout_g[63]));
AND2X1 exu_U3918(.A(exu_n11371), .B(exu_n8791), .Y(div_byp_muldivout_g[62]));
AND2X1 exu_U3919(.A(exu_n11373), .B(exu_n8792), .Y(div_byp_muldivout_g[61]));
AND2X1 exu_U3920(.A(exu_n11375), .B(exu_n8793), .Y(div_byp_muldivout_g[60]));
AND2X1 exu_U3921(.A(exu_n11379), .B(exu_n8795), .Y(div_byp_muldivout_g[59]));
AND2X1 exu_U3922(.A(exu_n11381), .B(exu_n8796), .Y(div_byp_muldivout_g[58]));
AND2X1 exu_U3923(.A(exu_n11383), .B(exu_n8797), .Y(div_byp_muldivout_g[57]));
AND2X1 exu_U3924(.A(exu_n11385), .B(exu_n8798), .Y(div_byp_muldivout_g[56]));
AND2X1 exu_U3925(.A(exu_n11387), .B(exu_n8799), .Y(div_byp_muldivout_g[55]));
AND2X1 exu_U3926(.A(exu_n11389), .B(exu_n8800), .Y(div_byp_muldivout_g[54]));
AND2X1 exu_U3927(.A(exu_n11391), .B(exu_n8801), .Y(div_byp_muldivout_g[53]));
AND2X1 exu_U3928(.A(exu_n11393), .B(exu_n8802), .Y(div_byp_muldivout_g[52]));
AND2X1 exu_U3929(.A(exu_n11395), .B(exu_n8803), .Y(div_byp_muldivout_g[51]));
AND2X1 exu_U3930(.A(exu_n11397), .B(exu_n8804), .Y(div_byp_muldivout_g[50]));
AND2X1 exu_U3931(.A(exu_n11401), .B(exu_n8806), .Y(div_byp_muldivout_g[49]));
AND2X1 exu_U3932(.A(exu_n11403), .B(exu_n8807), .Y(div_byp_muldivout_g[48]));
AND2X1 exu_U3933(.A(exu_n11405), .B(exu_n8808), .Y(div_byp_muldivout_g[47]));
AND2X1 exu_U3934(.A(exu_n11407), .B(exu_n8809), .Y(div_byp_muldivout_g[46]));
AND2X1 exu_U3935(.A(exu_n11409), .B(exu_n8810), .Y(div_byp_muldivout_g[45]));
AND2X1 exu_U3936(.A(exu_n11411), .B(exu_n8811), .Y(div_byp_muldivout_g[44]));
AND2X1 exu_U3937(.A(exu_n11413), .B(exu_n8812), .Y(div_byp_muldivout_g[43]));
AND2X1 exu_U3938(.A(exu_n11415), .B(exu_n8813), .Y(div_byp_muldivout_g[42]));
AND2X1 exu_U3939(.A(exu_n11417), .B(exu_n8814), .Y(div_byp_muldivout_g[41]));
AND2X1 exu_U3940(.A(exu_n11419), .B(exu_n8815), .Y(div_byp_muldivout_g[40]));
AND2X1 exu_U3941(.A(exu_n11423), .B(exu_n8817), .Y(div_byp_muldivout_g[39]));
AND2X1 exu_U3942(.A(exu_n11425), .B(exu_n8818), .Y(div_byp_muldivout_g[38]));
AND2X1 exu_U3943(.A(exu_n11427), .B(exu_n8819), .Y(div_byp_muldivout_g[37]));
AND2X1 exu_U3944(.A(exu_n11429), .B(exu_n8820), .Y(div_byp_muldivout_g[36]));
AND2X1 exu_U3945(.A(exu_n11431), .B(exu_n8821), .Y(div_byp_muldivout_g[35]));
AND2X1 exu_U3946(.A(exu_n11433), .B(exu_n8822), .Y(div_byp_muldivout_g[34]));
AND2X1 exu_U3947(.A(exu_n11435), .B(exu_n8823), .Y(div_byp_muldivout_g[33]));
AND2X1 exu_U3948(.A(exu_n11437), .B(exu_n8824), .Y(div_byp_muldivout_g[32]));
AND2X1 exu_U3949(.A(exu_n11439), .B(exu_n8825), .Y(div_byp_muldivout_g[31]));
AND2X1 exu_U3950(.A(exu_n11441), .B(exu_n8826), .Y(div_byp_muldivout_g[30]));
AND2X1 exu_U3951(.A(exu_n11445), .B(exu_n8828), .Y(div_byp_muldivout_g[29]));
AND2X1 exu_U3952(.A(exu_n11447), .B(exu_n8829), .Y(div_byp_muldivout_g[28]));
AND2X1 exu_U3953(.A(exu_n11449), .B(exu_n8830), .Y(div_byp_muldivout_g[27]));
AND2X1 exu_U3954(.A(exu_n11451), .B(exu_n8831), .Y(div_byp_muldivout_g[26]));
AND2X1 exu_U3955(.A(exu_n11453), .B(exu_n8832), .Y(div_byp_muldivout_g[25]));
AND2X1 exu_U3956(.A(exu_n11455), .B(exu_n8833), .Y(div_byp_muldivout_g[24]));
AND2X1 exu_U3957(.A(exu_n11457), .B(exu_n8834), .Y(div_byp_muldivout_g[23]));
AND2X1 exu_U3958(.A(exu_n11459), .B(exu_n8835), .Y(div_byp_muldivout_g[22]));
AND2X1 exu_U3959(.A(exu_n11461), .B(exu_n8836), .Y(div_byp_muldivout_g[21]));
AND2X1 exu_U3960(.A(exu_n11463), .B(exu_n8837), .Y(div_byp_muldivout_g[20]));
AND2X1 exu_U3961(.A(exu_n11467), .B(exu_n8839), .Y(div_byp_muldivout_g[19]));
AND2X1 exu_U3962(.A(exu_n11469), .B(exu_n8840), .Y(div_byp_muldivout_g[18]));
AND2X1 exu_U3963(.A(exu_n11471), .B(exu_n8841), .Y(div_byp_muldivout_g[17]));
AND2X1 exu_U3964(.A(exu_n11473), .B(exu_n8842), .Y(div_byp_muldivout_g[16]));
AND2X1 exu_U3965(.A(exu_n11475), .B(exu_n8843), .Y(div_byp_muldivout_g[15]));
AND2X1 exu_U3966(.A(exu_n11477), .B(exu_n8844), .Y(div_byp_muldivout_g[14]));
AND2X1 exu_U3967(.A(exu_n11479), .B(exu_n8845), .Y(div_byp_muldivout_g[13]));
AND2X1 exu_U3968(.A(exu_n11481), .B(exu_n8846), .Y(div_byp_muldivout_g[12]));
AND2X1 exu_U3969(.A(exu_n11483), .B(exu_n8847), .Y(div_byp_muldivout_g[11]));
AND2X1 exu_U3970(.A(exu_n11485), .B(exu_n8848), .Y(div_byp_muldivout_g[10]));
AND2X1 exu_U3971(.A(exu_n11363), .B(exu_n8787), .Y(div_byp_muldivout_g[8]));
AND2X1 exu_U3972(.A(exu_n11365), .B(exu_n8788), .Y(div_byp_muldivout_g[7]));
AND2X1 exu_U3973(.A(exu_n11367), .B(exu_n8789), .Y(div_byp_muldivout_g[6]));
AND2X1 exu_U3974(.A(exu_n11377), .B(exu_n8794), .Y(div_byp_muldivout_g[5]));
AND2X1 exu_U3975(.A(exu_n11399), .B(exu_n8805), .Y(div_byp_muldivout_g[4]));
AND2X1 exu_U3976(.A(exu_n11421), .B(exu_n8816), .Y(div_byp_muldivout_g[3]));
AND2X1 exu_U3977(.A(exu_n11443), .B(exu_n8827), .Y(div_byp_muldivout_g[2]));
AND2X1 exu_U3978(.A(exu_n11465), .B(exu_n8838), .Y(div_byp_muldivout_g[1]));
INVX1 exu_U3979(.A(exu_n29496), .Y(exu_n16052));
AND2X1 exu_U3980(.A(exu_n11487), .B(exu_n8849), .Y(div_byp_muldivout_g[0]));
INVX1 exu_U3981(.A(exu_n29496), .Y(exu_n16053));
OR2X1 exu_U3982(.A(exu_n12406), .B(exu_n13818), .Y(bypass_rs1_data_btwn_mux[63]));
AND2X1 exu_U3983(.A(exu_n1689), .B(exu_n6708), .Y(exu_n23609));
OR2X1 exu_U3984(.A(exu_n12407), .B(exu_n13819), .Y(bypass_rs1_data_btwn_mux[62]));
AND2X1 exu_U3985(.A(exu_n1692), .B(exu_n6710), .Y(exu_n23614));
OR2X1 exu_U3986(.A(exu_n12408), .B(exu_n13820), .Y(bypass_rs1_data_btwn_mux[61]));
AND2X1 exu_U3987(.A(exu_n1695), .B(exu_n6712), .Y(exu_n23619));
OR2X1 exu_U3988(.A(exu_n12409), .B(exu_n13821), .Y(bypass_rs1_data_btwn_mux[60]));
AND2X1 exu_U3989(.A(exu_n1713), .B(exu_n6713), .Y(exu_n23625));
OR2X1 exu_U3990(.A(exu_n12411), .B(exu_n13823), .Y(bypass_rs1_data_btwn_mux[59]));
AND2X1 exu_U3991(.A(exu_n1713), .B(exu_n6717), .Y(exu_n23636));
OR2X1 exu_U3992(.A(exu_n12412), .B(exu_n13824), .Y(bypass_rs1_data_btwn_mux[58]));
AND2X1 exu_U3993(.A(exu_n1713), .B(exu_n6719), .Y(exu_n23641));
OR2X1 exu_U3994(.A(exu_n12413), .B(exu_n13825), .Y(bypass_rs1_data_btwn_mux[57]));
AND2X1 exu_U3995(.A(exu_n1713), .B(exu_n6721), .Y(exu_n23646));
OR2X1 exu_U3996(.A(exu_n12414), .B(exu_n13826), .Y(bypass_rs1_data_btwn_mux[56]));
AND2X1 exu_U3997(.A(exu_n1713), .B(exu_n6723), .Y(exu_n23651));
OR2X1 exu_U3998(.A(exu_n12415), .B(exu_n13827), .Y(bypass_rs1_data_btwn_mux[55]));
AND2X1 exu_U3999(.A(exu_n1713), .B(exu_n6725), .Y(exu_n23656));
OR2X1 exu_U4000(.A(exu_n12416), .B(exu_n13828), .Y(bypass_rs1_data_btwn_mux[54]));
AND2X1 exu_U4001(.A(exu_n1713), .B(exu_n6727), .Y(exu_n23661));
OR2X1 exu_U4002(.A(exu_n12417), .B(exu_n13829), .Y(bypass_rs1_data_btwn_mux[53]));
AND2X1 exu_U4003(.A(exu_n1713), .B(exu_n6729), .Y(exu_n23666));
OR2X1 exu_U4004(.A(exu_n12418), .B(exu_n13830), .Y(bypass_rs1_data_btwn_mux[52]));
AND2X1 exu_U4005(.A(exu_n1713), .B(exu_n6731), .Y(exu_n23671));
OR2X1 exu_U4006(.A(exu_n12419), .B(exu_n13831), .Y(bypass_rs1_data_btwn_mux[51]));
AND2X1 exu_U4007(.A(exu_n1713), .B(exu_n6733), .Y(exu_n23676));
OR2X1 exu_U4008(.A(exu_n12420), .B(exu_n13832), .Y(bypass_rs1_data_btwn_mux[50]));
AND2X1 exu_U4009(.A(exu_n1713), .B(exu_n6735), .Y(exu_n23681));
OR2X1 exu_U4010(.A(exu_n12422), .B(exu_n13834), .Y(bypass_rs1_data_btwn_mux[49]));
AND2X1 exu_U4011(.A(exu_n1713), .B(exu_n6739), .Y(exu_n23692));
OR2X1 exu_U4012(.A(exu_n12423), .B(exu_n13835), .Y(bypass_rs1_data_btwn_mux[48]));
AND2X1 exu_U4013(.A(exu_n1713), .B(exu_n6741), .Y(exu_n23697));
OR2X1 exu_U4014(.A(exu_n12424), .B(exu_n13836), .Y(bypass_rs1_data_btwn_mux[47]));
AND2X1 exu_U4015(.A(exu_n1713), .B(exu_n6743), .Y(exu_n23702));
OR2X1 exu_U4016(.A(exu_n12425), .B(exu_n13837), .Y(bypass_rs1_data_btwn_mux[46]));
AND2X1 exu_U4017(.A(exu_n1716), .B(exu_n6746), .Y(exu_n23707));
OR2X1 exu_U4018(.A(exu_n12426), .B(exu_n13838), .Y(bypass_rs1_data_btwn_mux[45]));
AND2X1 exu_U4019(.A(exu_n1718), .B(exu_n6748), .Y(exu_n23713));
OR2X1 exu_U4020(.A(exu_n12427), .B(exu_n13839), .Y(bypass_rs1_data_btwn_mux[44]));
AND2X1 exu_U4021(.A(exu_n1720), .B(exu_n6750), .Y(exu_n23719));
OR2X1 exu_U4022(.A(exu_n12428), .B(exu_n13840), .Y(bypass_rs1_data_btwn_mux[43]));
AND2X1 exu_U4023(.A(exu_n1722), .B(exu_n6752), .Y(exu_n23725));
OR2X1 exu_U4024(.A(exu_n12429), .B(exu_n13841), .Y(bypass_rs1_data_btwn_mux[42]));
AND2X1 exu_U4025(.A(exu_n1724), .B(exu_n6754), .Y(exu_n23731));
OR2X1 exu_U4026(.A(exu_n12430), .B(exu_n13842), .Y(bypass_rs1_data_btwn_mux[41]));
AND2X1 exu_U4027(.A(exu_n1726), .B(exu_n6756), .Y(exu_n23737));
OR2X1 exu_U4028(.A(exu_n12431), .B(exu_n13843), .Y(bypass_rs1_data_btwn_mux[40]));
AND2X1 exu_U4029(.A(exu_n1728), .B(exu_n6758), .Y(exu_n23743));
OR2X1 exu_U4030(.A(exu_n12433), .B(exu_n13845), .Y(bypass_rs1_data_btwn_mux[39]));
AND2X1 exu_U4031(.A(exu_n1732), .B(exu_n6762), .Y(exu_n23755));
OR2X1 exu_U4032(.A(exu_n12434), .B(exu_n13846), .Y(bypass_rs1_data_btwn_mux[38]));
AND2X1 exu_U4033(.A(exu_n1734), .B(exu_n6764), .Y(exu_n23761));
OR2X1 exu_U4034(.A(exu_n12435), .B(exu_n13847), .Y(bypass_rs1_data_btwn_mux[37]));
AND2X1 exu_U4035(.A(exu_n1736), .B(exu_n6766), .Y(exu_n23767));
OR2X1 exu_U4036(.A(exu_n12436), .B(exu_n13848), .Y(bypass_rs1_data_btwn_mux[36]));
AND2X1 exu_U4037(.A(exu_n1738), .B(exu_n6768), .Y(exu_n23773));
OR2X1 exu_U4038(.A(exu_n12437), .B(exu_n13849), .Y(bypass_rs1_data_btwn_mux[35]));
AND2X1 exu_U4039(.A(exu_n1740), .B(exu_n6770), .Y(exu_n23779));
OR2X1 exu_U4040(.A(exu_n12438), .B(exu_n13850), .Y(bypass_rs1_data_btwn_mux[34]));
AND2X1 exu_U4041(.A(exu_n1742), .B(exu_n6772), .Y(exu_n23785));
OR2X1 exu_U4042(.A(exu_n12439), .B(exu_n13851), .Y(bypass_rs1_data_btwn_mux[33]));
AND2X1 exu_U4043(.A(exu_n1744), .B(exu_n6774), .Y(exu_n23791));
OR2X1 exu_U4044(.A(exu_n12440), .B(exu_n13852), .Y(bypass_rs1_data_btwn_mux[32]));
AND2X1 exu_U4045(.A(exu_n1746), .B(exu_n6776), .Y(exu_n23797));
OR2X1 exu_U4046(.A(exu_n12441), .B(exu_n13853), .Y(bypass_rs1_data_btwn_mux[31]));
AND2X1 exu_U4047(.A(exu_n1748), .B(exu_n6778), .Y(exu_n23803));
OR2X1 exu_U4048(.A(exu_n12442), .B(exu_n13854), .Y(bypass_rs1_data_btwn_mux[30]));
AND2X1 exu_U4049(.A(exu_n1750), .B(exu_n6780), .Y(exu_n23809));
OR2X1 exu_U4050(.A(exu_n12444), .B(exu_n13856), .Y(bypass_rs1_data_btwn_mux[29]));
AND2X1 exu_U4051(.A(exu_n1754), .B(exu_n6784), .Y(exu_n23821));
OR2X1 exu_U4052(.A(exu_n12445), .B(exu_n13857), .Y(bypass_rs1_data_btwn_mux[28]));
AND2X1 exu_U4053(.A(exu_n1756), .B(exu_n6786), .Y(exu_n23827));
OR2X1 exu_U4054(.A(exu_n12446), .B(exu_n13858), .Y(bypass_rs1_data_btwn_mux[27]));
AND2X1 exu_U4055(.A(exu_n1758), .B(exu_n6788), .Y(exu_n23833));
OR2X1 exu_U4056(.A(exu_n12447), .B(exu_n13859), .Y(bypass_rs1_data_btwn_mux[26]));
AND2X1 exu_U4057(.A(exu_n1760), .B(exu_n6790), .Y(exu_n23839));
OR2X1 exu_U4058(.A(exu_n12448), .B(exu_n13860), .Y(bypass_rs1_data_btwn_mux[25]));
AND2X1 exu_U4059(.A(exu_n1762), .B(exu_n6792), .Y(exu_n23845));
OR2X1 exu_U4060(.A(exu_n12449), .B(exu_n13861), .Y(bypass_rs1_data_btwn_mux[24]));
AND2X1 exu_U4061(.A(exu_n1764), .B(exu_n6794), .Y(exu_n23851));
OR2X1 exu_U4062(.A(exu_n12450), .B(exu_n13862), .Y(bypass_rs1_data_btwn_mux[23]));
AND2X1 exu_U4063(.A(exu_n1766), .B(exu_n6796), .Y(exu_n23857));
OR2X1 exu_U4064(.A(exu_n12451), .B(exu_n13863), .Y(bypass_rs1_data_btwn_mux[22]));
AND2X1 exu_U4065(.A(exu_n1768), .B(exu_n6798), .Y(exu_n23863));
OR2X1 exu_U4066(.A(exu_n12452), .B(exu_n13864), .Y(bypass_rs1_data_btwn_mux[21]));
AND2X1 exu_U4067(.A(exu_n1770), .B(exu_n6800), .Y(exu_n23869));
OR2X1 exu_U4068(.A(exu_n12453), .B(exu_n13865), .Y(bypass_rs1_data_btwn_mux[20]));
AND2X1 exu_U4069(.A(exu_n1772), .B(exu_n6802), .Y(exu_n23875));
OR2X1 exu_U4070(.A(exu_n12455), .B(exu_n13867), .Y(bypass_rs1_data_btwn_mux[19]));
AND2X1 exu_U4071(.A(exu_n1776), .B(exu_n6806), .Y(exu_n23887));
OR2X1 exu_U4072(.A(exu_n12456), .B(exu_n13868), .Y(bypass_rs1_data_btwn_mux[18]));
AND2X1 exu_U4073(.A(exu_n1778), .B(exu_n6808), .Y(exu_n23893));
OR2X1 exu_U4074(.A(exu_n12457), .B(exu_n13869), .Y(bypass_rs1_data_btwn_mux[17]));
AND2X1 exu_U4075(.A(exu_n1780), .B(exu_n6810), .Y(exu_n23899));
OR2X1 exu_U4076(.A(exu_n12458), .B(exu_n13870), .Y(bypass_rs1_data_btwn_mux[16]));
AND2X1 exu_U4077(.A(exu_n1782), .B(exu_n6812), .Y(exu_n23905));
OR2X1 exu_U4078(.A(exu_n12459), .B(exu_n13871), .Y(bypass_rs1_data_btwn_mux[15]));
AND2X1 exu_U4079(.A(exu_n1784), .B(exu_n6814), .Y(exu_n23911));
OR2X1 exu_U4080(.A(exu_n12460), .B(exu_n13872), .Y(bypass_rs1_data_btwn_mux[14]));
AND2X1 exu_U4081(.A(exu_n1786), .B(exu_n6816), .Y(exu_n23917));
OR2X1 exu_U4082(.A(exu_n12461), .B(exu_n13873), .Y(bypass_rs1_data_btwn_mux[13]));
AND2X1 exu_U4083(.A(exu_n1788), .B(exu_n6818), .Y(exu_n23923));
OR2X1 exu_U4084(.A(exu_n12462), .B(exu_n13874), .Y(bypass_rs1_data_btwn_mux[12]));
AND2X1 exu_U4085(.A(exu_n1790), .B(exu_n6820), .Y(exu_n23929));
OR2X1 exu_U4086(.A(exu_n12463), .B(exu_n13875), .Y(bypass_rs1_data_btwn_mux[11]));
AND2X1 exu_U4087(.A(exu_n1792), .B(exu_n6822), .Y(exu_n23935));
OR2X1 exu_U4088(.A(exu_n12464), .B(exu_n13876), .Y(bypass_rs1_data_btwn_mux[10]));
AND2X1 exu_U4089(.A(exu_n1794), .B(exu_n6824), .Y(exu_n23941));
OR2X1 exu_U4090(.A(exu_n12402), .B(exu_n13814), .Y(bypass_rs1_data_btwn_mux[9]));
OR2X1 exu_U4091(.A(exu_n12403), .B(exu_n13815), .Y(bypass_rs1_data_btwn_mux[8]));
AND2X1 exu_U4092(.A(exu_n1684), .B(exu_n6702), .Y(exu_n23591));
OR2X1 exu_U4093(.A(exu_n12404), .B(exu_n13816), .Y(bypass_rs1_data_btwn_mux[7]));
AND2X1 exu_U4094(.A(exu_n1686), .B(exu_n6704), .Y(exu_n23597));
OR2X1 exu_U4095(.A(exu_n12405), .B(exu_n13817), .Y(bypass_rs1_data_btwn_mux[6]));
AND2X1 exu_U4096(.A(exu_n1688), .B(exu_n6706), .Y(exu_n23603));
OR2X1 exu_U4097(.A(exu_n12410), .B(exu_n13822), .Y(bypass_rs1_data_btwn_mux[5]));
AND2X1 exu_U4098(.A(exu_n1698), .B(exu_n6716), .Y(exu_n23629));
OR2X1 exu_U4099(.A(exu_n12421), .B(exu_n13833), .Y(bypass_rs1_data_btwn_mux[4]));
AND2X1 exu_U4100(.A(exu_n1710), .B(exu_n6738), .Y(exu_n23685));
OR2X1 exu_U4101(.A(exu_n12432), .B(exu_n13844), .Y(bypass_rs1_data_btwn_mux[3]));
AND2X1 exu_U4102(.A(exu_n1730), .B(exu_n6760), .Y(exu_n23749));
OR2X1 exu_U4103(.A(exu_n12443), .B(exu_n13855), .Y(bypass_rs1_data_btwn_mux[2]));
AND2X1 exu_U4104(.A(exu_n1752), .B(exu_n6782), .Y(exu_n23815));
OR2X1 exu_U4105(.A(exu_n12454), .B(exu_n13866), .Y(bypass_rs1_data_btwn_mux[1]));
AND2X1 exu_U4106(.A(exu_n1774), .B(exu_n6804), .Y(exu_n23881));
INVX1 exu_U4107(.A(exu_n29561), .Y(exu_n16059));
OR2X1 exu_U4108(.A(exu_n16395), .B(sehold), .Y(ecl_byplog_rs1_n14));
OR2X1 exu_U4109(.A(exu_n12465), .B(exu_n13877), .Y(bypass_rs1_data_btwn_mux[0]));
AND2X1 exu_U4110(.A(exu_n1796), .B(exu_n6826), .Y(exu_n23947));
INVX1 exu_U4111(.A(exu_n29561), .Y(exu_n16060));
OR2X1 exu_U4112(.A(exu_n12662), .B(exu_n14010), .Y(bypass_rs2_data_btwn_mux[63]));
AND2X1 exu_U4113(.A(exu_n2125), .B(exu_n7156), .Y(exu_n25001));
INVX1 exu_U4114(.A(irf_byp_rs2_data_d_l[63]), .Y(bypass_mux_rs2_data_2_in1[63]));
OR2X1 exu_U4115(.A(exu_n12663), .B(exu_n14011), .Y(bypass_rs2_data_btwn_mux[62]));
AND2X1 exu_U4116(.A(exu_n2128), .B(exu_n7158), .Y(exu_n25006));
INVX1 exu_U4117(.A(irf_byp_rs2_data_d_l[62]), .Y(bypass_mux_rs2_data_2_in1[62]));
OR2X1 exu_U4118(.A(exu_n12664), .B(exu_n14012), .Y(bypass_rs2_data_btwn_mux[61]));
AND2X1 exu_U4119(.A(exu_n2131), .B(exu_n7160), .Y(exu_n25011));
INVX1 exu_U4120(.A(irf_byp_rs2_data_d_l[61]), .Y(bypass_mux_rs2_data_2_in1[61]));
OR2X1 exu_U4121(.A(exu_n12665), .B(exu_n14013), .Y(bypass_rs2_data_btwn_mux[60]));
AND2X1 exu_U4122(.A(exu_n2134), .B(exu_n7162), .Y(exu_n25016));
INVX1 exu_U4123(.A(irf_byp_rs2_data_d_l[60]), .Y(bypass_mux_rs2_data_2_in1[60]));
OR2X1 exu_U4124(.A(exu_n12667), .B(exu_n14015), .Y(bypass_rs2_data_btwn_mux[59]));
AND2X1 exu_U4125(.A(exu_n2139), .B(exu_n7166), .Y(exu_n25027));
INVX1 exu_U4126(.A(irf_byp_rs2_data_d_l[59]), .Y(bypass_mux_rs2_data_2_in1[59]));
OR2X1 exu_U4127(.A(exu_n12668), .B(exu_n14016), .Y(bypass_rs2_data_btwn_mux[58]));
AND2X1 exu_U4128(.A(exu_n2142), .B(exu_n7168), .Y(exu_n25032));
INVX1 exu_U4129(.A(irf_byp_rs2_data_d_l[58]), .Y(bypass_mux_rs2_data_2_in1[58]));
OR2X1 exu_U4130(.A(exu_n12669), .B(exu_n14017), .Y(bypass_rs2_data_btwn_mux[57]));
AND2X1 exu_U4131(.A(exu_n2145), .B(exu_n7170), .Y(exu_n25037));
INVX1 exu_U4132(.A(irf_byp_rs2_data_d_l[57]), .Y(bypass_mux_rs2_data_2_in1[57]));
OR2X1 exu_U4133(.A(exu_n12670), .B(exu_n14018), .Y(bypass_rs2_data_btwn_mux[56]));
AND2X1 exu_U4134(.A(exu_n2148), .B(exu_n7172), .Y(exu_n25042));
INVX1 exu_U4135(.A(irf_byp_rs2_data_d_l[56]), .Y(bypass_mux_rs2_data_2_in1[56]));
OR2X1 exu_U4136(.A(exu_n12671), .B(exu_n14019), .Y(bypass_rs2_data_btwn_mux[55]));
AND2X1 exu_U4137(.A(exu_n2151), .B(exu_n7174), .Y(exu_n25047));
INVX1 exu_U4138(.A(irf_byp_rs2_data_d_l[55]), .Y(bypass_mux_rs2_data_2_in1[55]));
OR2X1 exu_U4139(.A(exu_n12672), .B(exu_n14020), .Y(bypass_rs2_data_btwn_mux[54]));
AND2X1 exu_U4140(.A(exu_n2154), .B(exu_n7176), .Y(exu_n25052));
INVX1 exu_U4141(.A(irf_byp_rs2_data_d_l[54]), .Y(bypass_mux_rs2_data_2_in1[54]));
OR2X1 exu_U4142(.A(exu_n12673), .B(exu_n14021), .Y(bypass_rs2_data_btwn_mux[53]));
AND2X1 exu_U4143(.A(exu_n2157), .B(exu_n7178), .Y(exu_n25057));
INVX1 exu_U4144(.A(irf_byp_rs2_data_d_l[53]), .Y(bypass_mux_rs2_data_2_in1[53]));
OR2X1 exu_U4145(.A(exu_n12674), .B(exu_n14022), .Y(bypass_rs2_data_btwn_mux[52]));
AND2X1 exu_U4146(.A(exu_n2160), .B(exu_n7180), .Y(exu_n25062));
INVX1 exu_U4147(.A(irf_byp_rs2_data_d_l[52]), .Y(bypass_mux_rs2_data_2_in1[52]));
OR2X1 exu_U4148(.A(exu_n12675), .B(exu_n14023), .Y(bypass_rs2_data_btwn_mux[51]));
AND2X1 exu_U4149(.A(exu_n2163), .B(exu_n7182), .Y(exu_n25067));
INVX1 exu_U4150(.A(irf_byp_rs2_data_d_l[51]), .Y(bypass_mux_rs2_data_2_in1[51]));
OR2X1 exu_U4151(.A(exu_n12676), .B(exu_n14024), .Y(bypass_rs2_data_btwn_mux[50]));
AND2X1 exu_U4152(.A(exu_n2166), .B(exu_n7184), .Y(exu_n25072));
INVX1 exu_U4153(.A(irf_byp_rs2_data_d_l[50]), .Y(bypass_mux_rs2_data_2_in1[50]));
OR2X1 exu_U4154(.A(exu_n12678), .B(exu_n14026), .Y(bypass_rs2_data_btwn_mux[49]));
AND2X1 exu_U4155(.A(exu_n2171), .B(exu_n7188), .Y(exu_n25083));
INVX1 exu_U4156(.A(irf_byp_rs2_data_d_l[49]), .Y(bypass_mux_rs2_data_2_in1[49]));
OR2X1 exu_U4157(.A(exu_n12679), .B(exu_n14027), .Y(bypass_rs2_data_btwn_mux[48]));
AND2X1 exu_U4158(.A(exu_n2174), .B(exu_n7190), .Y(exu_n25088));
INVX1 exu_U4159(.A(irf_byp_rs2_data_d_l[48]), .Y(bypass_mux_rs2_data_2_in1[48]));
OR2X1 exu_U4160(.A(exu_n12680), .B(exu_n14028), .Y(bypass_rs2_data_btwn_mux[47]));
AND2X1 exu_U4161(.A(exu_n2177), .B(exu_n7192), .Y(exu_n25093));
INVX1 exu_U4162(.A(irf_byp_rs2_data_d_l[47]), .Y(bypass_mux_rs2_data_2_in1[47]));
OR2X1 exu_U4163(.A(exu_n12681), .B(exu_n14029), .Y(bypass_rs2_data_btwn_mux[46]));
AND2X1 exu_U4164(.A(exu_n2180), .B(exu_n7194), .Y(exu_n25098));
INVX1 exu_U4165(.A(irf_byp_rs2_data_d_l[46]), .Y(bypass_mux_rs2_data_2_in1[46]));
OR2X1 exu_U4166(.A(exu_n12682), .B(exu_n14030), .Y(bypass_rs2_data_btwn_mux[45]));
AND2X1 exu_U4167(.A(exu_n2197), .B(exu_n7195), .Y(exu_n25104));
INVX1 exu_U4168(.A(irf_byp_rs2_data_d_l[45]), .Y(bypass_mux_rs2_data_2_in1[45]));
OR2X1 exu_U4169(.A(exu_n12683), .B(exu_n14031), .Y(bypass_rs2_data_btwn_mux[44]));
AND2X1 exu_U4170(.A(exu_n2197), .B(exu_n7197), .Y(exu_n25109));
INVX1 exu_U4171(.A(irf_byp_rs2_data_d_l[44]), .Y(bypass_mux_rs2_data_2_in1[44]));
OR2X1 exu_U4172(.A(exu_n12684), .B(exu_n14032), .Y(bypass_rs2_data_btwn_mux[43]));
AND2X1 exu_U4173(.A(exu_n2197), .B(exu_n7199), .Y(exu_n25114));
INVX1 exu_U4174(.A(irf_byp_rs2_data_d_l[43]), .Y(bypass_mux_rs2_data_2_in1[43]));
OR2X1 exu_U4175(.A(exu_n12685), .B(exu_n14033), .Y(bypass_rs2_data_btwn_mux[42]));
AND2X1 exu_U4176(.A(exu_n2197), .B(exu_n7201), .Y(exu_n25119));
INVX1 exu_U4177(.A(irf_byp_rs2_data_d_l[42]), .Y(bypass_mux_rs2_data_2_in1[42]));
OR2X1 exu_U4178(.A(exu_n12686), .B(exu_n14034), .Y(bypass_rs2_data_btwn_mux[41]));
AND2X1 exu_U4179(.A(exu_n2197), .B(exu_n7203), .Y(exu_n25124));
INVX1 exu_U4180(.A(irf_byp_rs2_data_d_l[41]), .Y(bypass_mux_rs2_data_2_in1[41]));
OR2X1 exu_U4181(.A(exu_n12687), .B(exu_n14035), .Y(bypass_rs2_data_btwn_mux[40]));
AND2X1 exu_U4182(.A(exu_n2197), .B(exu_n7205), .Y(exu_n25129));
INVX1 exu_U4183(.A(irf_byp_rs2_data_d_l[40]), .Y(bypass_mux_rs2_data_2_in1[40]));
OR2X1 exu_U4184(.A(exu_n12689), .B(exu_n14037), .Y(bypass_rs2_data_btwn_mux[39]));
AND2X1 exu_U4185(.A(exu_n2197), .B(exu_n7209), .Y(exu_n25140));
INVX1 exu_U4186(.A(irf_byp_rs2_data_d_l[39]), .Y(bypass_mux_rs2_data_2_in1[39]));
OR2X1 exu_U4187(.A(exu_n12690), .B(exu_n14038), .Y(bypass_rs2_data_btwn_mux[38]));
AND2X1 exu_U4188(.A(exu_n2197), .B(exu_n7211), .Y(exu_n25145));
INVX1 exu_U4189(.A(irf_byp_rs2_data_d_l[38]), .Y(bypass_mux_rs2_data_2_in1[38]));
OR2X1 exu_U4190(.A(exu_n12691), .B(exu_n14039), .Y(bypass_rs2_data_btwn_mux[37]));
AND2X1 exu_U4191(.A(exu_n2197), .B(exu_n7213), .Y(exu_n25150));
INVX1 exu_U4192(.A(irf_byp_rs2_data_d_l[37]), .Y(bypass_mux_rs2_data_2_in1[37]));
OR2X1 exu_U4193(.A(exu_n12692), .B(exu_n14040), .Y(bypass_rs2_data_btwn_mux[36]));
AND2X1 exu_U4194(.A(exu_n2197), .B(exu_n7215), .Y(exu_n25155));
INVX1 exu_U4195(.A(irf_byp_rs2_data_d_l[36]), .Y(bypass_mux_rs2_data_2_in1[36]));
OR2X1 exu_U4196(.A(exu_n12693), .B(exu_n14041), .Y(bypass_rs2_data_btwn_mux[35]));
AND2X1 exu_U4197(.A(exu_n2197), .B(exu_n7217), .Y(exu_n25160));
INVX1 exu_U4198(.A(irf_byp_rs2_data_d_l[35]), .Y(bypass_mux_rs2_data_2_in1[35]));
OR2X1 exu_U4199(.A(exu_n12694), .B(exu_n14042), .Y(bypass_rs2_data_btwn_mux[34]));
AND2X1 exu_U4200(.A(exu_n2197), .B(exu_n7219), .Y(exu_n25165));
INVX1 exu_U4201(.A(irf_byp_rs2_data_d_l[34]), .Y(bypass_mux_rs2_data_2_in1[34]));
OR2X1 exu_U4202(.A(exu_n12695), .B(exu_n14043), .Y(bypass_rs2_data_btwn_mux[33]));
AND2X1 exu_U4203(.A(exu_n2197), .B(exu_n7221), .Y(exu_n25170));
INVX1 exu_U4204(.A(irf_byp_rs2_data_d_l[33]), .Y(bypass_mux_rs2_data_2_in1[33]));
OR2X1 exu_U4205(.A(exu_n12696), .B(exu_n14044), .Y(bypass_rs2_data_btwn_mux[32]));
AND2X1 exu_U4206(.A(exu_n2197), .B(exu_n7223), .Y(exu_n25175));
INVX1 exu_U4207(.A(irf_byp_rs2_data_d_l[32]), .Y(bypass_mux_rs2_data_2_in1[32]));
OR2X1 exu_U4208(.A(exu_n12697), .B(exu_n14045), .Y(bypass_rs2_data_btwn_mux[31]));
AND2X1 exu_U4209(.A(exu_n2197), .B(exu_n7225), .Y(exu_n25180));
INVX1 exu_U4210(.A(irf_byp_rs2_data_d_l[31]), .Y(bypass_mux_rs2_data_2_in1[31]));
OR2X1 exu_U4211(.A(exu_n12698), .B(exu_n14046), .Y(bypass_rs2_data_btwn_mux[30]));
AND2X1 exu_U4212(.A(exu_n2200), .B(exu_n7228), .Y(exu_n25185));
INVX1 exu_U4213(.A(irf_byp_rs2_data_d_l[30]), .Y(bypass_mux_rs2_data_2_in1[30]));
OR2X1 exu_U4214(.A(exu_n12700), .B(exu_n14048), .Y(bypass_rs2_data_btwn_mux[29]));
AND2X1 exu_U4215(.A(exu_n2204), .B(exu_n7232), .Y(exu_n25197));
INVX1 exu_U4216(.A(irf_byp_rs2_data_d_l[29]), .Y(bypass_mux_rs2_data_2_in1[29]));
OR2X1 exu_U4217(.A(exu_n12701), .B(exu_n14049), .Y(bypass_rs2_data_btwn_mux[28]));
AND2X1 exu_U4218(.A(exu_n2206), .B(exu_n7234), .Y(exu_n25203));
INVX1 exu_U4219(.A(irf_byp_rs2_data_d_l[28]), .Y(bypass_mux_rs2_data_2_in1[28]));
OR2X1 exu_U4220(.A(exu_n12702), .B(exu_n14050), .Y(bypass_rs2_data_btwn_mux[27]));
AND2X1 exu_U4221(.A(exu_n2208), .B(exu_n7236), .Y(exu_n25209));
INVX1 exu_U4222(.A(irf_byp_rs2_data_d_l[27]), .Y(bypass_mux_rs2_data_2_in1[27]));
OR2X1 exu_U4223(.A(exu_n12703), .B(exu_n14051), .Y(bypass_rs2_data_btwn_mux[26]));
AND2X1 exu_U4224(.A(exu_n2210), .B(exu_n7238), .Y(exu_n25215));
INVX1 exu_U4225(.A(irf_byp_rs2_data_d_l[26]), .Y(bypass_mux_rs2_data_2_in1[26]));
OR2X1 exu_U4226(.A(exu_n12704), .B(exu_n14052), .Y(bypass_rs2_data_btwn_mux[25]));
AND2X1 exu_U4227(.A(exu_n2212), .B(exu_n7240), .Y(exu_n25221));
INVX1 exu_U4228(.A(irf_byp_rs2_data_d_l[25]), .Y(bypass_mux_rs2_data_2_in1[25]));
OR2X1 exu_U4229(.A(exu_n12705), .B(exu_n14053), .Y(bypass_rs2_data_btwn_mux[24]));
AND2X1 exu_U4230(.A(exu_n2214), .B(exu_n7242), .Y(exu_n25227));
INVX1 exu_U4231(.A(irf_byp_rs2_data_d_l[24]), .Y(bypass_mux_rs2_data_2_in1[24]));
OR2X1 exu_U4232(.A(exu_n12706), .B(exu_n14054), .Y(bypass_rs2_data_btwn_mux[23]));
AND2X1 exu_U4233(.A(exu_n2216), .B(exu_n7244), .Y(exu_n25233));
INVX1 exu_U4234(.A(irf_byp_rs2_data_d_l[23]), .Y(bypass_mux_rs2_data_2_in1[23]));
OR2X1 exu_U4235(.A(exu_n12707), .B(exu_n14055), .Y(bypass_rs2_data_btwn_mux[22]));
AND2X1 exu_U4236(.A(exu_n2218), .B(exu_n7246), .Y(exu_n25239));
INVX1 exu_U4237(.A(irf_byp_rs2_data_d_l[22]), .Y(bypass_mux_rs2_data_2_in1[22]));
OR2X1 exu_U4238(.A(exu_n12708), .B(exu_n14056), .Y(bypass_rs2_data_btwn_mux[21]));
AND2X1 exu_U4239(.A(exu_n2220), .B(exu_n7248), .Y(exu_n25245));
INVX1 exu_U4240(.A(irf_byp_rs2_data_d_l[21]), .Y(bypass_mux_rs2_data_2_in1[21]));
OR2X1 exu_U4241(.A(exu_n12709), .B(exu_n14057), .Y(bypass_rs2_data_btwn_mux[20]));
AND2X1 exu_U4242(.A(exu_n2222), .B(exu_n7250), .Y(exu_n25251));
INVX1 exu_U4243(.A(irf_byp_rs2_data_d_l[20]), .Y(bypass_mux_rs2_data_2_in1[20]));
OR2X1 exu_U4244(.A(exu_n12711), .B(exu_n14059), .Y(bypass_rs2_data_btwn_mux[19]));
AND2X1 exu_U4245(.A(exu_n2226), .B(exu_n7254), .Y(exu_n25263));
INVX1 exu_U4246(.A(irf_byp_rs2_data_d_l[19]), .Y(bypass_mux_rs2_data_2_in1[19]));
OR2X1 exu_U4247(.A(exu_n12712), .B(exu_n14060), .Y(bypass_rs2_data_btwn_mux[18]));
AND2X1 exu_U4248(.A(exu_n2228), .B(exu_n7256), .Y(exu_n25269));
INVX1 exu_U4249(.A(irf_byp_rs2_data_d_l[18]), .Y(bypass_mux_rs2_data_2_in1[18]));
OR2X1 exu_U4250(.A(exu_n12713), .B(exu_n14061), .Y(bypass_rs2_data_btwn_mux[17]));
AND2X1 exu_U4251(.A(exu_n2230), .B(exu_n7258), .Y(exu_n25275));
INVX1 exu_U4252(.A(irf_byp_rs2_data_d_l[17]), .Y(bypass_mux_rs2_data_2_in1[17]));
OR2X1 exu_U4253(.A(exu_n12714), .B(exu_n14062), .Y(bypass_rs2_data_btwn_mux[16]));
AND2X1 exu_U4254(.A(exu_n2232), .B(exu_n7260), .Y(exu_n25281));
INVX1 exu_U4255(.A(irf_byp_rs2_data_d_l[16]), .Y(bypass_mux_rs2_data_2_in1[16]));
OR2X1 exu_U4256(.A(exu_n12715), .B(exu_n14063), .Y(bypass_rs2_data_btwn_mux[15]));
AND2X1 exu_U4257(.A(exu_n2234), .B(exu_n7262), .Y(exu_n25287));
INVX1 exu_U4258(.A(irf_byp_rs2_data_d_l[15]), .Y(bypass_mux_rs2_data_2_in1[15]));
OR2X1 exu_U4259(.A(exu_n12716), .B(exu_n14064), .Y(bypass_rs2_data_btwn_mux[14]));
AND2X1 exu_U4260(.A(exu_n2236), .B(exu_n7264), .Y(exu_n25293));
INVX1 exu_U4261(.A(irf_byp_rs2_data_d_l[14]), .Y(bypass_mux_rs2_data_2_in1[14]));
OR2X1 exu_U4262(.A(exu_n12717), .B(exu_n14065), .Y(bypass_rs2_data_btwn_mux[13]));
AND2X1 exu_U4263(.A(exu_n2238), .B(exu_n7266), .Y(exu_n25299));
INVX1 exu_U4264(.A(irf_byp_rs2_data_d_l[13]), .Y(bypass_mux_rs2_data_2_in1[13]));
OR2X1 exu_U4265(.A(exu_n12718), .B(exu_n14066), .Y(bypass_rs2_data_btwn_mux[12]));
AND2X1 exu_U4266(.A(exu_n2240), .B(exu_n7268), .Y(exu_n25305));
INVX1 exu_U4267(.A(irf_byp_rs2_data_d_l[12]), .Y(bypass_mux_rs2_data_2_in1[12]));
OR2X1 exu_U4268(.A(exu_n12719), .B(exu_n14067), .Y(bypass_rs2_data_btwn_mux[11]));
AND2X1 exu_U4269(.A(exu_n2242), .B(exu_n7270), .Y(exu_n25311));
INVX1 exu_U4270(.A(irf_byp_rs2_data_d_l[11]), .Y(bypass_mux_rs2_data_2_in1[11]));
OR2X1 exu_U4271(.A(exu_n12720), .B(exu_n14068), .Y(bypass_rs2_data_btwn_mux[10]));
AND2X1 exu_U4272(.A(exu_n2244), .B(exu_n7272), .Y(exu_n25317));
INVX1 exu_U4273(.A(irf_byp_rs2_data_d_l[10]), .Y(bypass_mux_rs2_data_2_in1[10]));
INVX1 exu_U4274(.A(irf_byp_rs2_data_d_l[9]), .Y(bypass_mux_rs2_data_2_in1[9]));
OR2X1 exu_U4275(.A(exu_n12658), .B(exu_n14006), .Y(bypass_rs2_data_btwn_mux[9]));
OR2X1 exu_U4276(.A(exu_n12659), .B(exu_n14007), .Y(bypass_rs2_data_btwn_mux[8]));
AND2X1 exu_U4277(.A(exu_n2120), .B(exu_n7150), .Y(exu_n24983));
INVX1 exu_U4278(.A(irf_byp_rs2_data_d_l[8]), .Y(bypass_mux_rs2_data_2_in1[8]));
OR2X1 exu_U4279(.A(exu_n12660), .B(exu_n14008), .Y(bypass_rs2_data_btwn_mux[7]));
AND2X1 exu_U4280(.A(exu_n2122), .B(exu_n7152), .Y(exu_n24989));
INVX1 exu_U4281(.A(irf_byp_rs2_data_d_l[7]), .Y(bypass_mux_rs2_data_2_in1[7]));
OR2X1 exu_U4282(.A(exu_n12661), .B(exu_n14009), .Y(bypass_rs2_data_btwn_mux[6]));
AND2X1 exu_U4283(.A(exu_n2124), .B(exu_n7154), .Y(exu_n24995));
INVX1 exu_U4284(.A(irf_byp_rs2_data_d_l[6]), .Y(bypass_mux_rs2_data_2_in1[6]));
OR2X1 exu_U4285(.A(exu_n12666), .B(exu_n14014), .Y(bypass_rs2_data_btwn_mux[5]));
AND2X1 exu_U4286(.A(exu_n2136), .B(exu_n7164), .Y(exu_n25021));
INVX1 exu_U4287(.A(irf_byp_rs2_data_d_l[5]), .Y(bypass_mux_rs2_data_2_in1[5]));
OR2X1 exu_U4288(.A(exu_n12677), .B(exu_n14025), .Y(bypass_rs2_data_btwn_mux[4]));
AND2X1 exu_U4289(.A(exu_n2168), .B(exu_n7186), .Y(exu_n25077));
INVX1 exu_U4290(.A(irf_byp_rs2_data_d_l[4]), .Y(bypass_mux_rs2_data_2_in1[4]));
OR2X1 exu_U4291(.A(exu_n12688), .B(exu_n14036), .Y(bypass_rs2_data_btwn_mux[3]));
AND2X1 exu_U4292(.A(exu_n2188), .B(exu_n7208), .Y(exu_n25133));
INVX1 exu_U4293(.A(irf_byp_rs2_data_d_l[3]), .Y(bypass_mux_rs2_data_2_in1[3]));
OR2X1 exu_U4294(.A(exu_n12699), .B(exu_n14047), .Y(bypass_rs2_data_btwn_mux[2]));
AND2X1 exu_U4295(.A(exu_n2202), .B(exu_n7230), .Y(exu_n25191));
INVX1 exu_U4296(.A(irf_byp_rs2_data_d_l[2]), .Y(bypass_mux_rs2_data_2_in1[2]));
OR2X1 exu_U4297(.A(exu_n12710), .B(exu_n14058), .Y(bypass_rs2_data_btwn_mux[1]));
AND2X1 exu_U4298(.A(exu_n2224), .B(exu_n7252), .Y(exu_n25257));
INVX1 exu_U4299(.A(irf_byp_rs2_data_d_l[1]), .Y(bypass_mux_rs2_data_2_in1[1]));
INVX1 exu_U4300(.A(exu_n29626), .Y(exu_n16066));
OR2X1 exu_U4301(.A(exu_n12721), .B(exu_n14069), .Y(bypass_rs2_data_btwn_mux[0]));
AND2X1 exu_U4302(.A(exu_n2246), .B(exu_n7274), .Y(exu_n25323));
INVX1 exu_U4303(.A(irf_byp_rs2_data_d_l[0]), .Y(bypass_mux_rs2_data_2_in1[0]));
INVX1 exu_U4304(.A(exu_n29626), .Y(exu_n16067));
INVX1 exu_U4305(.A(irf_byp_rs3_data_d_l[63]), .Y(bypass_mux_rs3_data_2_in1[63]));
OR2X1 exu_U4306(.A(exu_n12790), .B(exu_n25730), .Y(bypass_rs3_data_btwn_mux[63]));
INVX1 exu_U4307(.A(irf_byp_rs3_data_d_l[62]), .Y(bypass_mux_rs3_data_2_in1[62]));
OR2X1 exu_U4308(.A(exu_n12791), .B(exu_n25734), .Y(bypass_rs3_data_btwn_mux[62]));
INVX1 exu_U4309(.A(irf_byp_rs3_data_d_l[61]), .Y(bypass_mux_rs3_data_2_in1[61]));
OR2X1 exu_U4310(.A(exu_n12792), .B(exu_n25738), .Y(bypass_rs3_data_btwn_mux[61]));
INVX1 exu_U4311(.A(irf_byp_rs3_data_d_l[60]), .Y(bypass_mux_rs3_data_2_in1[60]));
OR2X1 exu_U4312(.A(exu_n12793), .B(exu_n25742), .Y(bypass_rs3_data_btwn_mux[60]));
INVX1 exu_U4313(.A(irf_byp_rs3_data_d_l[59]), .Y(bypass_mux_rs3_data_2_in1[59]));
OR2X1 exu_U4314(.A(exu_n12795), .B(exu_n25750), .Y(bypass_rs3_data_btwn_mux[59]));
INVX1 exu_U4315(.A(irf_byp_rs3_data_d_l[58]), .Y(bypass_mux_rs3_data_2_in1[58]));
OR2X1 exu_U4316(.A(exu_n12796), .B(exu_n25754), .Y(bypass_rs3_data_btwn_mux[58]));
INVX1 exu_U4317(.A(irf_byp_rs3_data_d_l[57]), .Y(bypass_mux_rs3_data_2_in1[57]));
OR2X1 exu_U4318(.A(exu_n12797), .B(exu_n25758), .Y(bypass_rs3_data_btwn_mux[57]));
INVX1 exu_U4319(.A(irf_byp_rs3_data_d_l[56]), .Y(bypass_mux_rs3_data_2_in1[56]));
OR2X1 exu_U4320(.A(exu_n12798), .B(exu_n25762), .Y(bypass_rs3_data_btwn_mux[56]));
INVX1 exu_U4321(.A(irf_byp_rs3_data_d_l[55]), .Y(bypass_mux_rs3_data_2_in1[55]));
OR2X1 exu_U4322(.A(exu_n12799), .B(exu_n25766), .Y(bypass_rs3_data_btwn_mux[55]));
INVX1 exu_U4323(.A(irf_byp_rs3_data_d_l[54]), .Y(bypass_mux_rs3_data_2_in1[54]));
OR2X1 exu_U4324(.A(exu_n12800), .B(exu_n25770), .Y(bypass_rs3_data_btwn_mux[54]));
INVX1 exu_U4325(.A(irf_byp_rs3_data_d_l[53]), .Y(bypass_mux_rs3_data_2_in1[53]));
OR2X1 exu_U4326(.A(exu_n12801), .B(exu_n25774), .Y(bypass_rs3_data_btwn_mux[53]));
INVX1 exu_U4327(.A(irf_byp_rs3_data_d_l[52]), .Y(bypass_mux_rs3_data_2_in1[52]));
OR2X1 exu_U4328(.A(exu_n12802), .B(exu_n25778), .Y(bypass_rs3_data_btwn_mux[52]));
INVX1 exu_U4329(.A(irf_byp_rs3_data_d_l[51]), .Y(bypass_mux_rs3_data_2_in1[51]));
OR2X1 exu_U4330(.A(exu_n12803), .B(exu_n25782), .Y(bypass_rs3_data_btwn_mux[51]));
INVX1 exu_U4331(.A(irf_byp_rs3_data_d_l[50]), .Y(bypass_mux_rs3_data_2_in1[50]));
OR2X1 exu_U4332(.A(exu_n12804), .B(exu_n25786), .Y(bypass_rs3_data_btwn_mux[50]));
INVX1 exu_U4333(.A(irf_byp_rs3_data_d_l[49]), .Y(bypass_mux_rs3_data_2_in1[49]));
OR2X1 exu_U4334(.A(exu_n12806), .B(exu_n25794), .Y(bypass_rs3_data_btwn_mux[49]));
INVX1 exu_U4335(.A(irf_byp_rs3_data_d_l[48]), .Y(bypass_mux_rs3_data_2_in1[48]));
OR2X1 exu_U4336(.A(exu_n12807), .B(exu_n25798), .Y(bypass_rs3_data_btwn_mux[48]));
INVX1 exu_U4337(.A(irf_byp_rs3_data_d_l[47]), .Y(bypass_mux_rs3_data_2_in1[47]));
OR2X1 exu_U4338(.A(exu_n12808), .B(exu_n25802), .Y(bypass_rs3_data_btwn_mux[47]));
INVX1 exu_U4339(.A(irf_byp_rs3_data_d_l[46]), .Y(bypass_mux_rs3_data_2_in1[46]));
OR2X1 exu_U4340(.A(exu_n12809), .B(exu_n25806), .Y(bypass_rs3_data_btwn_mux[46]));
INVX1 exu_U4341(.A(irf_byp_rs3_data_d_l[45]), .Y(bypass_mux_rs3_data_2_in1[45]));
OR2X1 exu_U4342(.A(exu_n12810), .B(exu_n25810), .Y(bypass_rs3_data_btwn_mux[45]));
INVX1 exu_U4343(.A(irf_byp_rs3_data_d_l[44]), .Y(bypass_mux_rs3_data_2_in1[44]));
OR2X1 exu_U4344(.A(exu_n12811), .B(exu_n25814), .Y(bypass_rs3_data_btwn_mux[44]));
INVX1 exu_U4345(.A(irf_byp_rs3_data_d_l[43]), .Y(bypass_mux_rs3_data_2_in1[43]));
OR2X1 exu_U4346(.A(exu_n12812), .B(exu_n25818), .Y(bypass_rs3_data_btwn_mux[43]));
INVX1 exu_U4347(.A(irf_byp_rs3_data_d_l[42]), .Y(bypass_mux_rs3_data_2_in1[42]));
OR2X1 exu_U4348(.A(exu_n12813), .B(exu_n25822), .Y(bypass_rs3_data_btwn_mux[42]));
INVX1 exu_U4349(.A(irf_byp_rs3_data_d_l[41]), .Y(bypass_mux_rs3_data_2_in1[41]));
OR2X1 exu_U4350(.A(exu_n12814), .B(exu_n25826), .Y(bypass_rs3_data_btwn_mux[41]));
INVX1 exu_U4351(.A(irf_byp_rs3_data_d_l[40]), .Y(bypass_mux_rs3_data_2_in1[40]));
OR2X1 exu_U4352(.A(exu_n12815), .B(exu_n25830), .Y(bypass_rs3_data_btwn_mux[40]));
INVX1 exu_U4353(.A(irf_byp_rs3_data_d_l[39]), .Y(bypass_mux_rs3_data_2_in1[39]));
OR2X1 exu_U4354(.A(exu_n12817), .B(exu_n25838), .Y(bypass_rs3_data_btwn_mux[39]));
INVX1 exu_U4355(.A(irf_byp_rs3_data_d_l[38]), .Y(bypass_mux_rs3_data_2_in1[38]));
OR2X1 exu_U4356(.A(exu_n12818), .B(exu_n25842), .Y(bypass_rs3_data_btwn_mux[38]));
INVX1 exu_U4357(.A(irf_byp_rs3_data_d_l[37]), .Y(bypass_mux_rs3_data_2_in1[37]));
OR2X1 exu_U4358(.A(exu_n12819), .B(exu_n25846), .Y(bypass_rs3_data_btwn_mux[37]));
INVX1 exu_U4359(.A(irf_byp_rs3_data_d_l[36]), .Y(bypass_mux_rs3_data_2_in1[36]));
OR2X1 exu_U4360(.A(exu_n12820), .B(exu_n25850), .Y(bypass_rs3_data_btwn_mux[36]));
INVX1 exu_U4361(.A(irf_byp_rs3_data_d_l[35]), .Y(bypass_mux_rs3_data_2_in1[35]));
OR2X1 exu_U4362(.A(exu_n12821), .B(exu_n25854), .Y(bypass_rs3_data_btwn_mux[35]));
INVX1 exu_U4363(.A(irf_byp_rs3_data_d_l[34]), .Y(bypass_mux_rs3_data_2_in1[34]));
OR2X1 exu_U4364(.A(exu_n12822), .B(exu_n25858), .Y(bypass_rs3_data_btwn_mux[34]));
INVX1 exu_U4365(.A(irf_byp_rs3_data_d_l[33]), .Y(bypass_mux_rs3_data_2_in1[33]));
OR2X1 exu_U4366(.A(exu_n12823), .B(exu_n25862), .Y(bypass_rs3_data_btwn_mux[33]));
INVX1 exu_U4367(.A(irf_byp_rs3_data_d_l[32]), .Y(bypass_mux_rs3_data_2_in1[32]));
OR2X1 exu_U4368(.A(exu_n12824), .B(exu_n25866), .Y(bypass_rs3_data_btwn_mux[32]));
INVX1 exu_U4369(.A(irf_byp_rs3_data_d_l[31]), .Y(bypass_mux_rs3_data_2_in1[31]));
OR2X1 exu_U4370(.A(exu_n12825), .B(exu_n25870), .Y(bypass_rs3_data_btwn_mux[31]));
INVX1 exu_U4371(.A(irf_byp_rs3_data_d_l[30]), .Y(bypass_mux_rs3_data_2_in1[30]));
OR2X1 exu_U4372(.A(exu_n12826), .B(exu_n25874), .Y(bypass_rs3_data_btwn_mux[30]));
INVX1 exu_U4373(.A(irf_byp_rs3_data_d_l[29]), .Y(bypass_mux_rs3_data_2_in1[29]));
OR2X1 exu_U4374(.A(exu_n12828), .B(exu_n25882), .Y(bypass_rs3_data_btwn_mux[29]));
INVX1 exu_U4375(.A(irf_byp_rs3_data_d_l[28]), .Y(bypass_mux_rs3_data_2_in1[28]));
OR2X1 exu_U4376(.A(exu_n12829), .B(exu_n25886), .Y(bypass_rs3_data_btwn_mux[28]));
INVX1 exu_U4377(.A(irf_byp_rs3_data_d_l[27]), .Y(bypass_mux_rs3_data_2_in1[27]));
OR2X1 exu_U4378(.A(exu_n12830), .B(exu_n25890), .Y(bypass_rs3_data_btwn_mux[27]));
INVX1 exu_U4379(.A(irf_byp_rs3_data_d_l[26]), .Y(bypass_mux_rs3_data_2_in1[26]));
OR2X1 exu_U4380(.A(exu_n12831), .B(exu_n25894), .Y(bypass_rs3_data_btwn_mux[26]));
INVX1 exu_U4381(.A(irf_byp_rs3_data_d_l[25]), .Y(bypass_mux_rs3_data_2_in1[25]));
OR2X1 exu_U4382(.A(exu_n12832), .B(exu_n25898), .Y(bypass_rs3_data_btwn_mux[25]));
INVX1 exu_U4383(.A(irf_byp_rs3_data_d_l[24]), .Y(bypass_mux_rs3_data_2_in1[24]));
OR2X1 exu_U4384(.A(exu_n12833), .B(exu_n25902), .Y(bypass_rs3_data_btwn_mux[24]));
INVX1 exu_U4385(.A(irf_byp_rs3_data_d_l[23]), .Y(bypass_mux_rs3_data_2_in1[23]));
OR2X1 exu_U4386(.A(exu_n12834), .B(exu_n25906), .Y(bypass_rs3_data_btwn_mux[23]));
INVX1 exu_U4387(.A(irf_byp_rs3_data_d_l[22]), .Y(bypass_mux_rs3_data_2_in1[22]));
OR2X1 exu_U4388(.A(exu_n12835), .B(exu_n25910), .Y(bypass_rs3_data_btwn_mux[22]));
INVX1 exu_U4389(.A(irf_byp_rs3_data_d_l[21]), .Y(bypass_mux_rs3_data_2_in1[21]));
OR2X1 exu_U4390(.A(exu_n12836), .B(exu_n25914), .Y(bypass_rs3_data_btwn_mux[21]));
INVX1 exu_U4391(.A(irf_byp_rs3_data_d_l[20]), .Y(bypass_mux_rs3_data_2_in1[20]));
OR2X1 exu_U4392(.A(exu_n12837), .B(exu_n25918), .Y(bypass_rs3_data_btwn_mux[20]));
INVX1 exu_U4393(.A(irf_byp_rs3_data_d_l[19]), .Y(bypass_mux_rs3_data_2_in1[19]));
OR2X1 exu_U4394(.A(exu_n12839), .B(exu_n25926), .Y(bypass_rs3_data_btwn_mux[19]));
INVX1 exu_U4395(.A(irf_byp_rs3_data_d_l[18]), .Y(bypass_mux_rs3_data_2_in1[18]));
OR2X1 exu_U4396(.A(exu_n12840), .B(exu_n25930), .Y(bypass_rs3_data_btwn_mux[18]));
INVX1 exu_U4397(.A(irf_byp_rs3_data_d_l[17]), .Y(bypass_mux_rs3_data_2_in1[17]));
OR2X1 exu_U4398(.A(exu_n12841), .B(exu_n25934), .Y(bypass_rs3_data_btwn_mux[17]));
INVX1 exu_U4399(.A(irf_byp_rs3_data_d_l[16]), .Y(bypass_mux_rs3_data_2_in1[16]));
OR2X1 exu_U4400(.A(exu_n12842), .B(exu_n25938), .Y(bypass_rs3_data_btwn_mux[16]));
INVX1 exu_U4401(.A(irf_byp_rs3_data_d_l[15]), .Y(bypass_mux_rs3_data_2_in1[15]));
OR2X1 exu_U4402(.A(exu_n12843), .B(exu_n25942), .Y(bypass_rs3_data_btwn_mux[15]));
INVX1 exu_U4403(.A(irf_byp_rs3_data_d_l[14]), .Y(bypass_mux_rs3_data_2_in1[14]));
OR2X1 exu_U4404(.A(exu_n12844), .B(exu_n25946), .Y(bypass_rs3_data_btwn_mux[14]));
INVX1 exu_U4405(.A(irf_byp_rs3_data_d_l[13]), .Y(bypass_mux_rs3_data_2_in1[13]));
OR2X1 exu_U4406(.A(exu_n12845), .B(exu_n25950), .Y(bypass_rs3_data_btwn_mux[13]));
INVX1 exu_U4407(.A(irf_byp_rs3_data_d_l[12]), .Y(bypass_mux_rs3_data_2_in1[12]));
OR2X1 exu_U4408(.A(exu_n12846), .B(exu_n25954), .Y(bypass_rs3_data_btwn_mux[12]));
INVX1 exu_U4409(.A(irf_byp_rs3_data_d_l[11]), .Y(bypass_mux_rs3_data_2_in1[11]));
OR2X1 exu_U4410(.A(exu_n12847), .B(exu_n25958), .Y(bypass_rs3_data_btwn_mux[11]));
INVX1 exu_U4411(.A(irf_byp_rs3_data_d_l[10]), .Y(bypass_mux_rs3_data_2_in1[10]));
OR2X1 exu_U4412(.A(exu_n12848), .B(exu_n25962), .Y(bypass_rs3_data_btwn_mux[10]));
INVX1 exu_U4413(.A(irf_byp_rs3_data_d_l[9]), .Y(bypass_mux_rs3_data_2_in1[9]));
OR2X1 exu_U4414(.A(exu_n12786), .B(exu_n25714), .Y(bypass_rs3_data_btwn_mux[9]));
INVX1 exu_U4415(.A(irf_byp_rs3_data_d_l[8]), .Y(bypass_mux_rs3_data_2_in1[8]));
OR2X1 exu_U4416(.A(exu_n12787), .B(exu_n25718), .Y(bypass_rs3_data_btwn_mux[8]));
INVX1 exu_U4417(.A(irf_byp_rs3_data_d_l[7]), .Y(bypass_mux_rs3_data_2_in1[7]));
OR2X1 exu_U4418(.A(exu_n12788), .B(exu_n25722), .Y(bypass_rs3_data_btwn_mux[7]));
INVX1 exu_U4419(.A(irf_byp_rs3_data_d_l[6]), .Y(bypass_mux_rs3_data_2_in1[6]));
OR2X1 exu_U4420(.A(exu_n12789), .B(exu_n25726), .Y(bypass_rs3_data_btwn_mux[6]));
INVX1 exu_U4421(.A(irf_byp_rs3_data_d_l[5]), .Y(bypass_mux_rs3_data_2_in1[5]));
OR2X1 exu_U4422(.A(exu_n12794), .B(exu_n25746), .Y(bypass_rs3_data_btwn_mux[5]));
INVX1 exu_U4423(.A(irf_byp_rs3_data_d_l[4]), .Y(bypass_mux_rs3_data_2_in1[4]));
OR2X1 exu_U4424(.A(exu_n12805), .B(exu_n25790), .Y(bypass_rs3_data_btwn_mux[4]));
INVX1 exu_U4425(.A(irf_byp_rs3_data_d_l[3]), .Y(bypass_mux_rs3_data_2_in1[3]));
OR2X1 exu_U4426(.A(exu_n12816), .B(exu_n25834), .Y(bypass_rs3_data_btwn_mux[3]));
INVX1 exu_U4427(.A(irf_byp_rs3_data_d_l[2]), .Y(bypass_mux_rs3_data_2_in1[2]));
OR2X1 exu_U4428(.A(exu_n12827), .B(exu_n25878), .Y(bypass_rs3_data_btwn_mux[2]));
INVX1 exu_U4429(.A(irf_byp_rs3_data_d_l[1]), .Y(bypass_mux_rs3_data_2_in1[1]));
OR2X1 exu_U4430(.A(exu_n12838), .B(exu_n25922), .Y(bypass_rs3_data_btwn_mux[1]));
INVX1 exu_U4431(.A(exu_n29691), .Y(exu_n16073));
INVX1 exu_U4432(.A(irf_byp_rs3_data_d_l[0]), .Y(bypass_mux_rs3_data_2_in1[0]));
OR2X1 exu_U4433(.A(exu_n12849), .B(exu_n25966), .Y(bypass_rs3_data_btwn_mux[0]));
INVX1 exu_U4434(.A(exu_n29691), .Y(exu_n16074));
INVX1 exu_U4435(.A(irf_byp_rs1_data_d_l[63]), .Y(bypass_mux_rcc_data_2_in1[63]));
OR2X1 exu_U4436(.A(exu_n12534), .B(exu_n24354), .Y(bypass_rcc_data_btwn_mux[63]));
INVX1 exu_U4437(.A(irf_byp_rs1_data_d_l[62]), .Y(bypass_mux_rcc_data_2_in1[62]));
OR2X1 exu_U4438(.A(exu_n12535), .B(exu_n24358), .Y(bypass_rcc_data_btwn_mux[62]));
INVX1 exu_U4439(.A(irf_byp_rs1_data_d_l[61]), .Y(bypass_mux_rcc_data_2_in1[61]));
OR2X1 exu_U4440(.A(exu_n12536), .B(exu_n24362), .Y(bypass_rcc_data_btwn_mux[61]));
INVX1 exu_U4441(.A(irf_byp_rs1_data_d_l[60]), .Y(bypass_mux_rcc_data_2_in1[60]));
OR2X1 exu_U4442(.A(exu_n12537), .B(exu_n24366), .Y(bypass_rcc_data_btwn_mux[60]));
INVX1 exu_U4443(.A(irf_byp_rs1_data_d_l[59]), .Y(bypass_mux_rcc_data_2_in1[59]));
OR2X1 exu_U4444(.A(exu_n12539), .B(exu_n24374), .Y(bypass_rcc_data_btwn_mux[59]));
INVX1 exu_U4445(.A(irf_byp_rs1_data_d_l[58]), .Y(bypass_mux_rcc_data_2_in1[58]));
OR2X1 exu_U4446(.A(exu_n12540), .B(exu_n24378), .Y(bypass_rcc_data_btwn_mux[58]));
INVX1 exu_U4447(.A(irf_byp_rs1_data_d_l[57]), .Y(bypass_mux_rcc_data_2_in1[57]));
OR2X1 exu_U4448(.A(exu_n12541), .B(exu_n24382), .Y(bypass_rcc_data_btwn_mux[57]));
INVX1 exu_U4449(.A(irf_byp_rs1_data_d_l[56]), .Y(bypass_mux_rcc_data_2_in1[56]));
OR2X1 exu_U4450(.A(exu_n12542), .B(exu_n24386), .Y(bypass_rcc_data_btwn_mux[56]));
INVX1 exu_U4451(.A(irf_byp_rs1_data_d_l[55]), .Y(bypass_mux_rcc_data_2_in1[55]));
OR2X1 exu_U4452(.A(exu_n12543), .B(exu_n24390), .Y(bypass_rcc_data_btwn_mux[55]));
INVX1 exu_U4453(.A(irf_byp_rs1_data_d_l[54]), .Y(bypass_mux_rcc_data_2_in1[54]));
OR2X1 exu_U4454(.A(exu_n12544), .B(exu_n24394), .Y(bypass_rcc_data_btwn_mux[54]));
INVX1 exu_U4455(.A(irf_byp_rs1_data_d_l[53]), .Y(bypass_mux_rcc_data_2_in1[53]));
OR2X1 exu_U4456(.A(exu_n12545), .B(exu_n24398), .Y(bypass_rcc_data_btwn_mux[53]));
INVX1 exu_U4457(.A(irf_byp_rs1_data_d_l[52]), .Y(bypass_mux_rcc_data_2_in1[52]));
OR2X1 exu_U4458(.A(exu_n12546), .B(exu_n24402), .Y(bypass_rcc_data_btwn_mux[52]));
INVX1 exu_U4459(.A(irf_byp_rs1_data_d_l[51]), .Y(bypass_mux_rcc_data_2_in1[51]));
OR2X1 exu_U4460(.A(exu_n12547), .B(exu_n24406), .Y(bypass_rcc_data_btwn_mux[51]));
INVX1 exu_U4461(.A(irf_byp_rs1_data_d_l[50]), .Y(bypass_mux_rcc_data_2_in1[50]));
OR2X1 exu_U4462(.A(exu_n12548), .B(exu_n24410), .Y(bypass_rcc_data_btwn_mux[50]));
INVX1 exu_U4463(.A(irf_byp_rs1_data_d_l[49]), .Y(bypass_mux_rcc_data_2_in1[49]));
OR2X1 exu_U4464(.A(exu_n12550), .B(exu_n24418), .Y(bypass_rcc_data_btwn_mux[49]));
INVX1 exu_U4465(.A(irf_byp_rs1_data_d_l[48]), .Y(bypass_mux_rcc_data_2_in1[48]));
OR2X1 exu_U4466(.A(exu_n12551), .B(exu_n24422), .Y(bypass_rcc_data_btwn_mux[48]));
INVX1 exu_U4467(.A(irf_byp_rs1_data_d_l[47]), .Y(bypass_mux_rcc_data_2_in1[47]));
OR2X1 exu_U4468(.A(exu_n12552), .B(exu_n24426), .Y(bypass_rcc_data_btwn_mux[47]));
INVX1 exu_U4469(.A(irf_byp_rs1_data_d_l[46]), .Y(bypass_mux_rcc_data_2_in1[46]));
OR2X1 exu_U4470(.A(exu_n12553), .B(exu_n24430), .Y(bypass_rcc_data_btwn_mux[46]));
INVX1 exu_U4471(.A(irf_byp_rs1_data_d_l[45]), .Y(bypass_mux_rcc_data_2_in1[45]));
OR2X1 exu_U4472(.A(exu_n12554), .B(exu_n24434), .Y(bypass_rcc_data_btwn_mux[45]));
INVX1 exu_U4473(.A(irf_byp_rs1_data_d_l[44]), .Y(bypass_mux_rcc_data_2_in1[44]));
OR2X1 exu_U4474(.A(exu_n12555), .B(exu_n24438), .Y(bypass_rcc_data_btwn_mux[44]));
INVX1 exu_U4475(.A(irf_byp_rs1_data_d_l[43]), .Y(bypass_mux_rcc_data_2_in1[43]));
OR2X1 exu_U4476(.A(exu_n12556), .B(exu_n24442), .Y(bypass_rcc_data_btwn_mux[43]));
INVX1 exu_U4477(.A(irf_byp_rs1_data_d_l[42]), .Y(bypass_mux_rcc_data_2_in1[42]));
OR2X1 exu_U4478(.A(exu_n12557), .B(exu_n24446), .Y(bypass_rcc_data_btwn_mux[42]));
INVX1 exu_U4479(.A(irf_byp_rs1_data_d_l[41]), .Y(bypass_mux_rcc_data_2_in1[41]));
OR2X1 exu_U4480(.A(exu_n12558), .B(exu_n24450), .Y(bypass_rcc_data_btwn_mux[41]));
INVX1 exu_U4481(.A(irf_byp_rs1_data_d_l[40]), .Y(bypass_mux_rcc_data_2_in1[40]));
OR2X1 exu_U4482(.A(exu_n12559), .B(exu_n24454), .Y(bypass_rcc_data_btwn_mux[40]));
INVX1 exu_U4483(.A(irf_byp_rs1_data_d_l[39]), .Y(bypass_mux_rcc_data_2_in1[39]));
OR2X1 exu_U4484(.A(exu_n12561), .B(exu_n24462), .Y(bypass_rcc_data_btwn_mux[39]));
INVX1 exu_U4485(.A(irf_byp_rs1_data_d_l[38]), .Y(bypass_mux_rcc_data_2_in1[38]));
OR2X1 exu_U4486(.A(exu_n12562), .B(exu_n24466), .Y(bypass_rcc_data_btwn_mux[38]));
INVX1 exu_U4487(.A(irf_byp_rs1_data_d_l[37]), .Y(bypass_mux_rcc_data_2_in1[37]));
OR2X1 exu_U4488(.A(exu_n12563), .B(exu_n24470), .Y(bypass_rcc_data_btwn_mux[37]));
INVX1 exu_U4489(.A(irf_byp_rs1_data_d_l[36]), .Y(bypass_mux_rcc_data_2_in1[36]));
OR2X1 exu_U4490(.A(exu_n12564), .B(exu_n24474), .Y(bypass_rcc_data_btwn_mux[36]));
INVX1 exu_U4491(.A(irf_byp_rs1_data_d_l[35]), .Y(bypass_mux_rcc_data_2_in1[35]));
OR2X1 exu_U4492(.A(exu_n12565), .B(exu_n24478), .Y(bypass_rcc_data_btwn_mux[35]));
INVX1 exu_U4493(.A(irf_byp_rs1_data_d_l[34]), .Y(bypass_mux_rcc_data_2_in1[34]));
OR2X1 exu_U4494(.A(exu_n12566), .B(exu_n24482), .Y(bypass_rcc_data_btwn_mux[34]));
INVX1 exu_U4495(.A(irf_byp_rs1_data_d_l[33]), .Y(bypass_mux_rcc_data_2_in1[33]));
OR2X1 exu_U4496(.A(exu_n12567), .B(exu_n24486), .Y(bypass_rcc_data_btwn_mux[33]));
INVX1 exu_U4497(.A(irf_byp_rs1_data_d_l[32]), .Y(bypass_mux_rcc_data_2_in1[32]));
OR2X1 exu_U4498(.A(exu_n12568), .B(exu_n24490), .Y(bypass_rcc_data_btwn_mux[32]));
INVX1 exu_U4499(.A(irf_byp_rs1_data_d_l[31]), .Y(bypass_mux_rcc_data_2_in1[31]));
OR2X1 exu_U4500(.A(exu_n12569), .B(exu_n24494), .Y(bypass_rcc_data_btwn_mux[31]));
INVX1 exu_U4501(.A(irf_byp_rs1_data_d_l[30]), .Y(bypass_mux_rcc_data_2_in1[30]));
OR2X1 exu_U4502(.A(exu_n12570), .B(exu_n24498), .Y(bypass_rcc_data_btwn_mux[30]));
INVX1 exu_U4503(.A(irf_byp_rs1_data_d_l[29]), .Y(bypass_mux_rcc_data_2_in1[29]));
OR2X1 exu_U4504(.A(exu_n12572), .B(exu_n24506), .Y(bypass_rcc_data_btwn_mux[29]));
INVX1 exu_U4505(.A(irf_byp_rs1_data_d_l[28]), .Y(bypass_mux_rcc_data_2_in1[28]));
OR2X1 exu_U4506(.A(exu_n12573), .B(exu_n24510), .Y(bypass_rcc_data_btwn_mux[28]));
INVX1 exu_U4507(.A(irf_byp_rs1_data_d_l[27]), .Y(bypass_mux_rcc_data_2_in1[27]));
OR2X1 exu_U4508(.A(exu_n12574), .B(exu_n24514), .Y(bypass_rcc_data_btwn_mux[27]));
INVX1 exu_U4509(.A(irf_byp_rs1_data_d_l[26]), .Y(bypass_mux_rcc_data_2_in1[26]));
OR2X1 exu_U4510(.A(exu_n12575), .B(exu_n24518), .Y(bypass_rcc_data_btwn_mux[26]));
INVX1 exu_U4511(.A(irf_byp_rs1_data_d_l[25]), .Y(bypass_mux_rcc_data_2_in1[25]));
OR2X1 exu_U4512(.A(exu_n12576), .B(exu_n24522), .Y(bypass_rcc_data_btwn_mux[25]));
INVX1 exu_U4513(.A(irf_byp_rs1_data_d_l[24]), .Y(bypass_mux_rcc_data_2_in1[24]));
OR2X1 exu_U4514(.A(exu_n12577), .B(exu_n24526), .Y(bypass_rcc_data_btwn_mux[24]));
INVX1 exu_U4515(.A(irf_byp_rs1_data_d_l[23]), .Y(bypass_mux_rcc_data_2_in1[23]));
OR2X1 exu_U4516(.A(exu_n12578), .B(exu_n24530), .Y(bypass_rcc_data_btwn_mux[23]));
INVX1 exu_U4517(.A(irf_byp_rs1_data_d_l[22]), .Y(bypass_mux_rcc_data_2_in1[22]));
OR2X1 exu_U4518(.A(exu_n12579), .B(exu_n24534), .Y(bypass_rcc_data_btwn_mux[22]));
INVX1 exu_U4519(.A(irf_byp_rs1_data_d_l[21]), .Y(bypass_mux_rcc_data_2_in1[21]));
OR2X1 exu_U4520(.A(exu_n12580), .B(exu_n24538), .Y(bypass_rcc_data_btwn_mux[21]));
INVX1 exu_U4521(.A(irf_byp_rs1_data_d_l[20]), .Y(bypass_mux_rcc_data_2_in1[20]));
OR2X1 exu_U4522(.A(exu_n12581), .B(exu_n24542), .Y(bypass_rcc_data_btwn_mux[20]));
INVX1 exu_U4523(.A(irf_byp_rs1_data_d_l[19]), .Y(bypass_mux_rcc_data_2_in1[19]));
OR2X1 exu_U4524(.A(exu_n12583), .B(exu_n24550), .Y(bypass_rcc_data_btwn_mux[19]));
INVX1 exu_U4525(.A(irf_byp_rs1_data_d_l[18]), .Y(bypass_mux_rcc_data_2_in1[18]));
OR2X1 exu_U4526(.A(exu_n12584), .B(exu_n24554), .Y(bypass_rcc_data_btwn_mux[18]));
INVX1 exu_U4527(.A(irf_byp_rs1_data_d_l[17]), .Y(bypass_mux_rcc_data_2_in1[17]));
OR2X1 exu_U4528(.A(exu_n12585), .B(exu_n24558), .Y(bypass_rcc_data_btwn_mux[17]));
INVX1 exu_U4529(.A(irf_byp_rs1_data_d_l[16]), .Y(bypass_mux_rcc_data_2_in1[16]));
OR2X1 exu_U4530(.A(exu_n12586), .B(exu_n24562), .Y(bypass_rcc_data_btwn_mux[16]));
INVX1 exu_U4531(.A(irf_byp_rs1_data_d_l[15]), .Y(bypass_mux_rcc_data_2_in1[15]));
OR2X1 exu_U4532(.A(exu_n12587), .B(exu_n24566), .Y(bypass_rcc_data_btwn_mux[15]));
INVX1 exu_U4533(.A(irf_byp_rs1_data_d_l[14]), .Y(bypass_mux_rcc_data_2_in1[14]));
OR2X1 exu_U4534(.A(exu_n12588), .B(exu_n24570), .Y(bypass_rcc_data_btwn_mux[14]));
INVX1 exu_U4535(.A(irf_byp_rs1_data_d_l[13]), .Y(bypass_mux_rcc_data_2_in1[13]));
OR2X1 exu_U4536(.A(exu_n12589), .B(exu_n24574), .Y(bypass_rcc_data_btwn_mux[13]));
INVX1 exu_U4537(.A(irf_byp_rs1_data_d_l[12]), .Y(bypass_mux_rcc_data_2_in1[12]));
OR2X1 exu_U4538(.A(exu_n12590), .B(exu_n24578), .Y(bypass_rcc_data_btwn_mux[12]));
INVX1 exu_U4539(.A(irf_byp_rs1_data_d_l[11]), .Y(bypass_mux_rcc_data_2_in1[11]));
OR2X1 exu_U4540(.A(exu_n12591), .B(exu_n24582), .Y(bypass_rcc_data_btwn_mux[11]));
INVX1 exu_U4541(.A(irf_byp_rs1_data_d_l[10]), .Y(bypass_mux_rcc_data_2_in1[10]));
OR2X1 exu_U4542(.A(exu_n12592), .B(exu_n24586), .Y(bypass_rcc_data_btwn_mux[10]));
INVX1 exu_U4543(.A(irf_byp_rs1_data_d_l[9]), .Y(bypass_mux_rcc_data_2_in1[9]));
OR2X1 exu_U4544(.A(exu_n12530), .B(exu_n24338), .Y(bypass_rcc_data_btwn_mux[9]));
INVX1 exu_U4545(.A(irf_byp_rs1_data_d_l[8]), .Y(bypass_mux_rcc_data_2_in1[8]));
OR2X1 exu_U4546(.A(exu_n12531), .B(exu_n24342), .Y(bypass_rcc_data_btwn_mux[8]));
INVX1 exu_U4547(.A(irf_byp_rs1_data_d_l[7]), .Y(bypass_mux_rcc_data_2_in1[7]));
OR2X1 exu_U4548(.A(exu_n12532), .B(exu_n24346), .Y(bypass_rcc_data_btwn_mux[7]));
INVX1 exu_U4549(.A(irf_byp_rs1_data_d_l[6]), .Y(bypass_mux_rcc_data_2_in1[6]));
OR2X1 exu_U4550(.A(exu_n12533), .B(exu_n24350), .Y(bypass_rcc_data_btwn_mux[6]));
INVX1 exu_U4551(.A(irf_byp_rs1_data_d_l[5]), .Y(bypass_mux_rcc_data_2_in1[5]));
OR2X1 exu_U4552(.A(exu_n12538), .B(exu_n24370), .Y(bypass_rcc_data_btwn_mux[5]));
INVX1 exu_U4553(.A(irf_byp_rs1_data_d_l[4]), .Y(bypass_mux_rcc_data_2_in1[4]));
OR2X1 exu_U4554(.A(exu_n12549), .B(exu_n24414), .Y(bypass_rcc_data_btwn_mux[4]));
INVX1 exu_U4555(.A(irf_byp_rs1_data_d_l[3]), .Y(bypass_mux_rcc_data_2_in1[3]));
OR2X1 exu_U4556(.A(exu_n12560), .B(exu_n24458), .Y(bypass_rcc_data_btwn_mux[3]));
INVX1 exu_U4557(.A(irf_byp_rs1_data_d_l[2]), .Y(bypass_mux_rcc_data_2_in1[2]));
OR2X1 exu_U4558(.A(exu_n12571), .B(exu_n24502), .Y(bypass_rcc_data_btwn_mux[2]));
INVX1 exu_U4559(.A(irf_byp_rs1_data_d_l[1]), .Y(bypass_mux_rcc_data_2_in1[1]));
OR2X1 exu_U4560(.A(exu_n12582), .B(exu_n24546), .Y(bypass_rcc_data_btwn_mux[1]));
INVX1 exu_U4561(.A(exu_n29756), .Y(exu_n16080));
INVX1 exu_U4562(.A(irf_byp_rs1_data_d_l[0]), .Y(bypass_mux_rcc_data_2_in1[0]));
OR2X1 exu_U4563(.A(exu_n12593), .B(exu_n24590), .Y(bypass_rcc_data_btwn_mux[0]));
INVX1 exu_U4564(.A(exu_n29756), .Y(exu_n16081));
INVX1 exu_U4565(.A(exu_n29821), .Y(exu_n16087));
INVX1 exu_U4566(.A(exu_n29821), .Y(exu_n16088));
INVX1 exu_U4567(.A(exu_n29886), .Y(exu_n16094));
INVX1 exu_U4568(.A(exu_n29886), .Y(exu_n16095));
INVX1 exu_U4569(.A(exu_n29950), .Y(exu_n16101));
INVX1 exu_U4570(.A(exu_n29950), .Y(exu_n16102));
INVX1 exu_U4571(.A(exu_n30015), .Y(exu_n16108));
INVX1 exu_U4572(.A(exu_n30015), .Y(exu_n16109));
INVX1 exu_U4573(.A(exu_n30080), .Y(exu_n16115));
INVX1 exu_U4574(.A(exu_n30080), .Y(exu_n16116));
OR2X1 exu_U4575(.A(exu_n12090), .B(exu_n13506), .Y(rml_cwp_old_cwp_w[2]));
AND2X1 exu_U4576(.A(exu_n229), .B(exu_n5156), .Y(exu_n17728));
OR2X1 exu_U4577(.A(exu_n12091), .B(exu_n13507), .Y(rml_cwp_old_cwp_w[1]));
AND2X1 exu_U4578(.A(exu_n231), .B(exu_n5158), .Y(exu_n17734));
OR2X1 exu_U4579(.A(exu_n12092), .B(exu_n13508), .Y(rml_cwp_old_cwp_w[0]));
AND2X1 exu_U4580(.A(exu_n233), .B(exu_n5160), .Y(exu_n17740));
INVX1 exu_U4581(.A(ifu_exu_muldivop_d[4]), .Y(exu_n16388));
AND2X1 exu_U4582(.A(ecl_mdqctl_n63), .B(ecl_div_sel_div), .Y(ecl_mdqctl_n46));
AND2X1 exu_U4583(.A(exu_n739), .B(exu_n5437), .Y(div_ecl_dividend_msb));
OR2X1 exu_U4584(.A(exu_n16213), .B(se), .Y(ecl_divcntl_inputs_neg_dff_n6));
INVX1 exu_U4585(.A(ecl_divcntl_div_state[5]), .Y(exu_n16505));
OR2X1 exu_U4586(.A(exu_n13434), .B(exu_n14754), .Y(ecl_divcntl_n30));
AND2X1 exu_U4587(.A(rml_next_cwp_m[0]), .B(rml_rml_cwp_wen_m), .Y(rml_n84));
AND2X1 exu_U4588(.A(exu_n84), .B(exu_n5051), .Y(exu_n17039));
AND2X1 exu_U4589(.A(exu_n3775), .B(exu_n8854), .Y(div_adderin1[63]));
AND2X1 exu_U4590(.A(exu_n83), .B(exu_n5050), .Y(exu_n17034));
AND2X1 exu_U4591(.A(exu_n3776), .B(exu_n8855), .Y(div_adderin1[62]));
AND2X1 exu_U4592(.A(exu_n82), .B(exu_n5049), .Y(exu_n17029));
AND2X1 exu_U4593(.A(exu_n3777), .B(exu_n8856), .Y(div_adderin1[61]));
AND2X1 exu_U4594(.A(exu_n81), .B(exu_n5048), .Y(exu_n17022));
AND2X1 exu_U4595(.A(exu_n3778), .B(exu_n8857), .Y(div_adderin1[60]));
AND2X1 exu_U4596(.A(exu_n80), .B(exu_n5047), .Y(exu_n17017));
AND2X1 exu_U4597(.A(exu_n3780), .B(exu_n8859), .Y(div_adderin1[59]));
AND2X1 exu_U4598(.A(exu_n79), .B(exu_n5046), .Y(exu_n17012));
AND2X1 exu_U4599(.A(exu_n3781), .B(exu_n8860), .Y(div_adderin1[58]));
AND2X1 exu_U4600(.A(exu_n78), .B(exu_n5045), .Y(exu_n17007));
AND2X1 exu_U4601(.A(exu_n3782), .B(exu_n8861), .Y(div_adderin1[57]));
AND2X1 exu_U4602(.A(exu_n77), .B(exu_n5044), .Y(exu_n17002));
AND2X1 exu_U4603(.A(exu_n3783), .B(exu_n8862), .Y(div_adderin1[56]));
AND2X1 exu_U4604(.A(exu_n76), .B(exu_n5043), .Y(exu_n16997));
AND2X1 exu_U4605(.A(exu_n3784), .B(exu_n8863), .Y(div_adderin1[55]));
AND2X1 exu_U4606(.A(exu_n75), .B(exu_n5042), .Y(exu_n16992));
AND2X1 exu_U4607(.A(exu_n3785), .B(exu_n8864), .Y(div_adderin1[54]));
AND2X1 exu_U4608(.A(exu_n74), .B(exu_n5041), .Y(exu_n16987));
AND2X1 exu_U4609(.A(exu_n3786), .B(exu_n8865), .Y(div_adderin1[53]));
AND2X1 exu_U4610(.A(exu_n73), .B(exu_n5040), .Y(exu_n16982));
AND2X1 exu_U4611(.A(exu_n3787), .B(exu_n8866), .Y(div_adderin1[52]));
AND2X1 exu_U4612(.A(exu_n72), .B(exu_n5039), .Y(exu_n16977));
AND2X1 exu_U4613(.A(exu_n3788), .B(exu_n8867), .Y(div_adderin1[51]));
AND2X1 exu_U4614(.A(exu_n71), .B(exu_n5038), .Y(exu_n16970));
AND2X1 exu_U4615(.A(exu_n3789), .B(exu_n8868), .Y(div_adderin1[50]));
AND2X1 exu_U4616(.A(exu_n70), .B(exu_n5037), .Y(exu_n16965));
AND2X1 exu_U4617(.A(exu_n3791), .B(exu_n8870), .Y(div_adderin1[49]));
AND2X1 exu_U4618(.A(exu_n69), .B(exu_n5036), .Y(exu_n16960));
AND2X1 exu_U4619(.A(exu_n3792), .B(exu_n8871), .Y(div_adderin1[48]));
AND2X1 exu_U4620(.A(exu_n68), .B(exu_n5035), .Y(exu_n16955));
AND2X1 exu_U4621(.A(exu_n3793), .B(exu_n8872), .Y(div_adderin1[47]));
AND2X1 exu_U4622(.A(exu_n67), .B(exu_n5034), .Y(exu_n16950));
AND2X1 exu_U4623(.A(exu_n3794), .B(exu_n8873), .Y(div_adderin1[46]));
AND2X1 exu_U4624(.A(exu_n66), .B(exu_n5033), .Y(exu_n16945));
AND2X1 exu_U4625(.A(exu_n3795), .B(exu_n8874), .Y(div_adderin1[45]));
AND2X1 exu_U4626(.A(exu_n65), .B(exu_n5032), .Y(exu_n16940));
AND2X1 exu_U4627(.A(exu_n3796), .B(exu_n8875), .Y(div_adderin1[44]));
AND2X1 exu_U4628(.A(exu_n64), .B(exu_n5031), .Y(exu_n16935));
AND2X1 exu_U4629(.A(exu_n3797), .B(exu_n8876), .Y(div_adderin1[43]));
AND2X1 exu_U4630(.A(exu_n63), .B(exu_n5030), .Y(exu_n16930));
AND2X1 exu_U4631(.A(exu_n3798), .B(exu_n8877), .Y(div_adderin1[42]));
AND2X1 exu_U4632(.A(exu_n62), .B(exu_n5029), .Y(exu_n17056));
AND2X1 exu_U4633(.A(exu_n3799), .B(exu_n8878), .Y(div_adderin1[41]));
AND2X1 exu_U4634(.A(exu_n61), .B(exu_n5028), .Y(exu_n17054));
AND2X1 exu_U4635(.A(exu_n3800), .B(exu_n8879), .Y(div_adderin1[40]));
AND2X1 exu_U4636(.A(exu_n60), .B(exu_n5027), .Y(exu_n17052));
AND2X1 exu_U4637(.A(exu_n3802), .B(exu_n8881), .Y(div_adderin1[39]));
AND2X1 exu_U4638(.A(exu_n59), .B(exu_n5026), .Y(exu_n17050));
AND2X1 exu_U4639(.A(exu_n3803), .B(exu_n8882), .Y(div_adderin1[38]));
AND2X1 exu_U4640(.A(exu_n58), .B(exu_n5025), .Y(exu_n17048));
AND2X1 exu_U4641(.A(exu_n3804), .B(exu_n8883), .Y(div_adderin1[37]));
AND2X1 exu_U4642(.A(exu_n57), .B(exu_n5024), .Y(exu_n17046));
AND2X1 exu_U4643(.A(exu_n3805), .B(exu_n8884), .Y(div_adderin1[36]));
AND2X1 exu_U4644(.A(exu_n15814), .B(ecl_ecl_div_signed_div), .Y(ecl_div_dividend_sign));
INVX1 exu_U4645(.A(exu_n16216), .Y(exu_n16214));
AND2X1 exu_U4646(.A(exu_n56), .B(exu_n5023), .Y(exu_n17044));
AND2X1 exu_U4647(.A(exu_n3806), .B(exu_n8885), .Y(div_adderin1[35]));
AND2X1 exu_U4648(.A(exu_n55), .B(exu_n5022), .Y(exu_n17028));
AND2X1 exu_U4649(.A(exu_n3807), .B(exu_n8886), .Y(div_adderin1[34]));
AND2X1 exu_U4650(.A(exu_n54), .B(exu_n5021), .Y(exu_n16976));
AND2X1 exu_U4651(.A(exu_n3808), .B(exu_n8887), .Y(div_adderin1[33]));
AND2X1 exu_U4652(.A(exu_n3809), .B(exu_n8888), .Y(div_adderin1[32]));
AND2X1 exu_U4653(.A(exu_n53), .B(exu_n5020), .Y(div_ecl_cout32));
AND2X1 exu_U4654(.A(exu_n51), .B(exu_n5018), .Y(exu_n16875));
AND2X1 exu_U4655(.A(exu_n3811), .B(exu_n8890), .Y(div_adderin1[30]));
INVX1 exu_U4656(.A(ecl_div_muls_rs1_31_e_l), .Y(exu_n16581));
AND2X1 exu_U4657(.A(exu_n50), .B(exu_n5017), .Y(exu_n16870));
AND2X1 exu_U4658(.A(exu_n3813), .B(exu_n8892), .Y(div_adderin1[29]));
AND2X1 exu_U4659(.A(exu_n49), .B(exu_n5016), .Y(exu_n16863));
AND2X1 exu_U4660(.A(exu_n3814), .B(exu_n8893), .Y(div_adderin1[28]));
AND2X1 exu_U4661(.A(exu_n48), .B(exu_n5015), .Y(exu_n16858));
AND2X1 exu_U4662(.A(exu_n3815), .B(exu_n8894), .Y(div_adderin1[27]));
AND2X1 exu_U4663(.A(exu_n47), .B(exu_n5014), .Y(exu_n16853));
AND2X1 exu_U4664(.A(exu_n3816), .B(exu_n8895), .Y(div_adderin1[26]));
AND2X1 exu_U4665(.A(exu_n46), .B(exu_n5013), .Y(exu_n16848));
AND2X1 exu_U4666(.A(exu_n3817), .B(exu_n8896), .Y(div_adderin1[25]));
AND2X1 exu_U4667(.A(exu_n45), .B(exu_n5012), .Y(exu_n16843));
AND2X1 exu_U4668(.A(exu_n3818), .B(exu_n8897), .Y(div_adderin1[24]));
AND2X1 exu_U4669(.A(exu_n44), .B(exu_n5011), .Y(exu_n16838));
AND2X1 exu_U4670(.A(exu_n3819), .B(exu_n8898), .Y(div_adderin1[23]));
AND2X1 exu_U4671(.A(exu_n43), .B(exu_n5010), .Y(exu_n16833));
AND2X1 exu_U4672(.A(exu_n3820), .B(exu_n8899), .Y(div_adderin1[22]));
AND2X1 exu_U4673(.A(exu_n42), .B(exu_n5009), .Y(exu_n16828));
AND2X1 exu_U4674(.A(exu_n3821), .B(exu_n8900), .Y(div_adderin1[21]));
AND2X1 exu_U4675(.A(exu_n41), .B(exu_n5008), .Y(exu_n16823));
AND2X1 exu_U4676(.A(exu_n3822), .B(exu_n8901), .Y(div_adderin1[20]));
AND2X1 exu_U4677(.A(exu_n40), .B(exu_n5007), .Y(exu_n16818));
AND2X1 exu_U4678(.A(exu_n3824), .B(exu_n8903), .Y(div_adderin1[19]));
AND2X1 exu_U4679(.A(exu_n39), .B(exu_n5006), .Y(exu_n16811));
AND2X1 exu_U4680(.A(exu_n3825), .B(exu_n8904), .Y(div_adderin1[18]));
AND2X1 exu_U4681(.A(exu_n38), .B(exu_n5005), .Y(exu_n16806));
AND2X1 exu_U4682(.A(exu_n3826), .B(exu_n8905), .Y(div_adderin1[17]));
AND2X1 exu_U4683(.A(exu_n37), .B(exu_n5004), .Y(exu_n16801));
AND2X1 exu_U4684(.A(exu_n3827), .B(exu_n8906), .Y(div_adderin1[16]));
AND2X1 exu_U4685(.A(exu_n36), .B(exu_n5003), .Y(exu_n16796));
AND2X1 exu_U4686(.A(exu_n3828), .B(exu_n8907), .Y(div_adderin1[15]));
AND2X1 exu_U4687(.A(exu_n35), .B(exu_n5002), .Y(exu_n16791));
AND2X1 exu_U4688(.A(exu_n3829), .B(exu_n8908), .Y(div_adderin1[14]));
AND2X1 exu_U4689(.A(exu_n34), .B(exu_n5001), .Y(exu_n16786));
AND2X1 exu_U4690(.A(exu_n3830), .B(exu_n8909), .Y(div_adderin1[13]));
AND2X1 exu_U4691(.A(exu_n33), .B(exu_n5000), .Y(exu_n16781));
AND2X1 exu_U4692(.A(exu_n3831), .B(exu_n8910), .Y(div_adderin1[12]));
AND2X1 exu_U4693(.A(exu_n32), .B(exu_n4999), .Y(exu_n16776));
AND2X1 exu_U4694(.A(exu_n3832), .B(exu_n8911), .Y(div_adderin1[11]));
AND2X1 exu_U4695(.A(exu_n31), .B(exu_n4998), .Y(exu_n16771));
AND2X1 exu_U4696(.A(exu_n3833), .B(exu_n8912), .Y(div_adderin1[10]));
AND2X1 exu_U4697(.A(exu_n30), .B(exu_n4997), .Y(exu_n16897));
AND2X1 exu_U4698(.A(exu_n3771), .B(exu_n8850), .Y(div_adderin1[9]));
AND2X1 exu_U4699(.A(exu_n29), .B(exu_n4996), .Y(exu_n16895));
AND2X1 exu_U4700(.A(exu_n3772), .B(exu_n8851), .Y(div_adderin1[8]));
AND2X1 exu_U4701(.A(exu_n28), .B(exu_n4995), .Y(exu_n16893));
AND2X1 exu_U4702(.A(exu_n3773), .B(exu_n8852), .Y(div_adderin1[7]));
AND2X1 exu_U4703(.A(exu_n27), .B(exu_n4994), .Y(exu_n16891));
AND2X1 exu_U4704(.A(exu_n3774), .B(exu_n8853), .Y(div_adderin1[6]));
AND2X1 exu_U4705(.A(exu_n26), .B(exu_n4993), .Y(exu_n16889));
AND2X1 exu_U4706(.A(exu_n3779), .B(exu_n8858), .Y(div_adderin1[5]));
AND2X1 exu_U4707(.A(exu_n25), .B(exu_n4992), .Y(exu_n16887));
AND2X1 exu_U4708(.A(exu_n3790), .B(exu_n8869), .Y(div_adderin1[4]));
AND2X1 exu_U4709(.A(exu_n24), .B(exu_n4991), .Y(exu_n16885));
AND2X1 exu_U4710(.A(exu_n3801), .B(exu_n8880), .Y(div_adderin1[3]));
AND2X1 exu_U4711(.A(exu_n23), .B(exu_n4990), .Y(exu_n16869));
AND2X1 exu_U4712(.A(exu_n3812), .B(exu_n8891), .Y(div_adderin1[2]));
AND2X1 exu_U4713(.A(exu_n22), .B(exu_n4989), .Y(exu_n16817));
AND2X1 exu_U4714(.A(exu_n3823), .B(exu_n8902), .Y(div_adderin1[1]));
AND2X1 exu_U4715(.A(exu_n3834), .B(exu_n8913), .Y(div_adderin1[0]));
AND2X1 exu_U4716(.A(exu_n4511), .B(exu_n9312), .Y(ecl_div_cin));
AND2X1 exu_U4717(.A(exu_n3353), .B(exu_n8434), .Y(exu_n28770));
AND2X1 exu_U4718(.A(exu_n3355), .B(exu_n8436), .Y(exu_n28773));
AND2X1 exu_U4719(.A(exu_n3354), .B(exu_n8435), .Y(exu_n28774));
AND2X1 exu_U4720(.A(exu_n3359), .B(exu_n8440), .Y(exu_n28785));
AND2X1 exu_U4721(.A(exu_n3358), .B(exu_n8439), .Y(exu_n28786));
AND2X1 exu_U4722(.A(exu_n3361), .B(exu_n8442), .Y(exu_n28791));
AND2X1 exu_U4723(.A(exu_n3360), .B(exu_n8441), .Y(exu_n28792));
AND2X1 exu_U4724(.A(exu_n3363), .B(exu_n8444), .Y(exu_n28797));
AND2X1 exu_U4725(.A(exu_n3362), .B(exu_n8443), .Y(exu_n28798));
AND2X1 exu_U4726(.A(exu_n3365), .B(exu_n8446), .Y(exu_n28803));
AND2X1 exu_U4727(.A(exu_n3364), .B(exu_n8445), .Y(exu_n28804));
AND2X1 exu_U4728(.A(exu_n3367), .B(exu_n8448), .Y(exu_n28809));
AND2X1 exu_U4729(.A(exu_n3366), .B(exu_n8447), .Y(exu_n28810));
AND2X1 exu_U4730(.A(exu_n3369), .B(exu_n8450), .Y(exu_n28815));
AND2X1 exu_U4731(.A(exu_n3368), .B(exu_n8449), .Y(exu_n28816));
AND2X1 exu_U4732(.A(exu_n3371), .B(exu_n8452), .Y(exu_n28821));
AND2X1 exu_U4733(.A(exu_n3370), .B(exu_n8451), .Y(exu_n28822));
AND2X1 exu_U4734(.A(exu_n3373), .B(exu_n8454), .Y(exu_n28827));
AND2X1 exu_U4735(.A(exu_n3372), .B(exu_n8453), .Y(exu_n28828));
AND2X1 exu_U4736(.A(exu_n3375), .B(exu_n8456), .Y(exu_n28833));
AND2X1 exu_U4737(.A(exu_n3374), .B(exu_n8455), .Y(exu_n28834));
AND2X1 exu_U4738(.A(exu_n3377), .B(exu_n8458), .Y(exu_n28839));
AND2X1 exu_U4739(.A(exu_n3376), .B(exu_n8457), .Y(exu_n28840));
AND2X1 exu_U4740(.A(exu_n3381), .B(exu_n8462), .Y(exu_n28851));
AND2X1 exu_U4741(.A(exu_n3380), .B(exu_n8461), .Y(exu_n28852));
AND2X1 exu_U4742(.A(exu_n3383), .B(exu_n8464), .Y(exu_n28857));
AND2X1 exu_U4743(.A(exu_n3382), .B(exu_n8463), .Y(exu_n28858));
AND2X1 exu_U4744(.A(exu_n3385), .B(exu_n8466), .Y(exu_n28863));
AND2X1 exu_U4745(.A(exu_n3384), .B(exu_n8465), .Y(exu_n28864));
AND2X1 exu_U4746(.A(exu_n3387), .B(exu_n8468), .Y(exu_n28869));
AND2X1 exu_U4747(.A(exu_n3386), .B(exu_n8467), .Y(exu_n28870));
AND2X1 exu_U4748(.A(exu_n3389), .B(exu_n8470), .Y(exu_n28875));
AND2X1 exu_U4749(.A(exu_n3388), .B(exu_n8469), .Y(exu_n28876));
AND2X1 exu_U4750(.A(exu_n3391), .B(exu_n8472), .Y(exu_n28881));
AND2X1 exu_U4751(.A(exu_n3390), .B(exu_n8471), .Y(exu_n28882));
AND2X1 exu_U4752(.A(exu_n3393), .B(exu_n8474), .Y(exu_n28887));
AND2X1 exu_U4753(.A(exu_n3392), .B(exu_n8473), .Y(exu_n28888));
AND2X1 exu_U4754(.A(exu_n3395), .B(exu_n8476), .Y(exu_n28893));
AND2X1 exu_U4755(.A(exu_n3394), .B(exu_n8475), .Y(exu_n28894));
INVX1 exu_U4756(.A(exu_n16218), .Y(exu_n16207));
AND2X1 exu_U4757(.A(exu_n3397), .B(exu_n8478), .Y(exu_n28899));
AND2X1 exu_U4758(.A(exu_n3396), .B(exu_n8477), .Y(exu_n28900));
AND2X1 exu_U4759(.A(exu_n3399), .B(exu_n8480), .Y(exu_n28905));
AND2X1 exu_U4760(.A(exu_n3398), .B(exu_n8479), .Y(exu_n28906));
AND2X1 exu_U4761(.A(exu_n3340), .B(exu_n8421), .Y(exu_n28696));
AND2X1 exu_U4762(.A(exu_n3339), .B(exu_n8420), .Y(exu_n28697));
AND2X1 exu_U4763(.A(exu_n3342), .B(exu_n8423), .Y(exu_n28702));
AND2X1 exu_U4764(.A(exu_n3341), .B(exu_n8422), .Y(exu_n28703));
INVX1 exu_U4765(.A(exu_n16206), .Y(exu_n16212));
AND2X1 exu_U4766(.A(exu_n3344), .B(exu_n8425), .Y(exu_n28708));
AND2X1 exu_U4767(.A(exu_n3343), .B(exu_n8424), .Y(exu_n28709));
INVX1 exu_U4768(.A(se), .Y(div_d_dff_n1));
AND2X1 exu_U4769(.A(exu_n3346), .B(exu_n8427), .Y(exu_n28714));
AND2X1 exu_U4770(.A(exu_n3345), .B(exu_n8426), .Y(exu_n28715));
INVX1 exu_U4771(.A(exu_n16206), .Y(exu_n16211));
AND2X1 exu_U4772(.A(exu_n3348), .B(exu_n8429), .Y(exu_n28724));
AND2X1 exu_U4773(.A(exu_n3347), .B(exu_n8428), .Y(exu_n28725));
INVX1 exu_U4774(.A(exu_n16217), .Y(exu_n16210));
AND2X1 exu_U4775(.A(exu_n3350), .B(exu_n8431), .Y(exu_n28740));
AND2X1 exu_U4776(.A(exu_n3349), .B(exu_n8430), .Y(exu_n28741));
INVX1 exu_U4777(.A(exu_n16217), .Y(exu_n16209));
INVX1 exu_U4778(.A(div_d_dff_n1), .Y(exu_n16127));
AND2X1 exu_U4779(.A(exu_n3352), .B(exu_n8433), .Y(exu_n28756));
AND2X1 exu_U4780(.A(exu_n3351), .B(exu_n8432), .Y(exu_n28757));
AND2X1 exu_U4781(.A(exu_n3357), .B(exu_n8438), .Y(exu_n28779));
AND2X1 exu_U4782(.A(exu_n3356), .B(exu_n8437), .Y(exu_n28780));
AND2X1 exu_U4783(.A(exu_n3379), .B(exu_n8460), .Y(exu_n28845));
AND2X1 exu_U4784(.A(exu_n3378), .B(exu_n8459), .Y(exu_n28846));
INVX1 exu_U4785(.A(exu_n16218), .Y(exu_n16208));
INVX1 exu_U4786(.A(div_d_dff_n1), .Y(exu_n16128));
AND2X1 exu_U4787(.A(exu_n3401), .B(exu_n8482), .Y(exu_n28911));
AND2X1 exu_U4788(.A(exu_n3400), .B(exu_n8481), .Y(exu_n28912));
INVX1 exu_U4789(.A(div_d_dff_n1), .Y(exu_n16129));
OR2X1 exu_U4790(.A(exu_n15493), .B(ecl_div_ld_inputs), .Y(ecl_n116));
INVX1 exu_U4791(.A(ifu_exu_tcc_e), .Y(exu_n16381));
OR2X1 exu_U4792(.A(ifu_exu_tcc_e), .B(exu_n15393), .Y(ecl_pick_normal_ttype));
AND2X1 exu_U4793(.A(ecl_tid_w[1]), .B(ecl_tid_w[0]), .Y(ecl_rml_thr_w[3]));
BUFX2 exu_U4794(.A(exu_n15404), .Y(exu_n15958));
BUFX2 exu_U4795(.A(exu_n15405), .Y(exu_n15960));
INVX1 exu_U4796(.A(exu_n15458), .Y(exu_n16398));
INVX1 exu_U4797(.A(irf_byp_rs3h_data_d_l[31]), .Y(bypass_mux_rs3h_data_2_in1[31]));
OR2X1 exu_U4798(.A(exu_n13462), .B(bypass_mux_rs3h_data_1_n46), .Y(bypass_rs3h_data_btwn_mux[31]));
INVX1 exu_U4799(.A(irf_byp_rs3h_data_d_l[30]), .Y(bypass_mux_rs3h_data_2_in1[30]));
OR2X1 exu_U4800(.A(exu_n13463), .B(bypass_mux_rs3h_data_1_n52), .Y(bypass_rs3h_data_btwn_mux[30]));
INVX1 exu_U4801(.A(irf_byp_rs3h_data_d_l[29]), .Y(bypass_mux_rs3h_data_2_in1[29]));
OR2X1 exu_U4802(.A(exu_n13465), .B(bypass_mux_rs3h_data_1_n64), .Y(bypass_rs3h_data_btwn_mux[29]));
INVX1 exu_U4803(.A(irf_byp_rs3h_data_d_l[28]), .Y(bypass_mux_rs3h_data_2_in1[28]));
OR2X1 exu_U4804(.A(exu_n13466), .B(bypass_mux_rs3h_data_1_n70), .Y(bypass_rs3h_data_btwn_mux[28]));
INVX1 exu_U4805(.A(irf_byp_rs3h_data_d_l[27]), .Y(bypass_mux_rs3h_data_2_in1[27]));
OR2X1 exu_U4806(.A(exu_n13467), .B(bypass_mux_rs3h_data_1_n76), .Y(bypass_rs3h_data_btwn_mux[27]));
INVX1 exu_U4807(.A(irf_byp_rs3h_data_d_l[26]), .Y(bypass_mux_rs3h_data_2_in1[26]));
OR2X1 exu_U4808(.A(exu_n13468), .B(bypass_mux_rs3h_data_1_n82), .Y(bypass_rs3h_data_btwn_mux[26]));
INVX1 exu_U4809(.A(irf_byp_rs3h_data_d_l[25]), .Y(bypass_mux_rs3h_data_2_in1[25]));
OR2X1 exu_U4810(.A(exu_n13469), .B(bypass_mux_rs3h_data_1_n88), .Y(bypass_rs3h_data_btwn_mux[25]));
INVX1 exu_U4811(.A(irf_byp_rs3h_data_d_l[24]), .Y(bypass_mux_rs3h_data_2_in1[24]));
OR2X1 exu_U4812(.A(exu_n13470), .B(bypass_mux_rs3h_data_1_n94), .Y(bypass_rs3h_data_btwn_mux[24]));
INVX1 exu_U4813(.A(irf_byp_rs3h_data_d_l[23]), .Y(bypass_mux_rs3h_data_2_in1[23]));
OR2X1 exu_U4814(.A(exu_n13471), .B(bypass_mux_rs3h_data_1_n100), .Y(bypass_rs3h_data_btwn_mux[23]));
INVX1 exu_U4815(.A(irf_byp_rs3h_data_d_l[22]), .Y(bypass_mux_rs3h_data_2_in1[22]));
OR2X1 exu_U4816(.A(exu_n13472), .B(bypass_mux_rs3h_data_1_n106), .Y(bypass_rs3h_data_btwn_mux[22]));
INVX1 exu_U4817(.A(irf_byp_rs3h_data_d_l[21]), .Y(bypass_mux_rs3h_data_2_in1[21]));
OR2X1 exu_U4818(.A(exu_n13473), .B(bypass_mux_rs3h_data_1_n112), .Y(bypass_rs3h_data_btwn_mux[21]));
INVX1 exu_U4819(.A(irf_byp_rs3h_data_d_l[20]), .Y(bypass_mux_rs3h_data_2_in1[20]));
OR2X1 exu_U4820(.A(exu_n13474), .B(bypass_mux_rs3h_data_1_n118), .Y(bypass_rs3h_data_btwn_mux[20]));
INVX1 exu_U4821(.A(irf_byp_rs3h_data_d_l[19]), .Y(bypass_mux_rs3h_data_2_in1[19]));
OR2X1 exu_U4822(.A(exu_n13476), .B(bypass_mux_rs3h_data_1_n130), .Y(bypass_rs3h_data_btwn_mux[19]));
INVX1 exu_U4823(.A(irf_byp_rs3h_data_d_l[18]), .Y(bypass_mux_rs3h_data_2_in1[18]));
OR2X1 exu_U4824(.A(exu_n13477), .B(bypass_mux_rs3h_data_1_n136), .Y(bypass_rs3h_data_btwn_mux[18]));
INVX1 exu_U4825(.A(irf_byp_rs3h_data_d_l[17]), .Y(bypass_mux_rs3h_data_2_in1[17]));
OR2X1 exu_U4826(.A(exu_n13478), .B(bypass_mux_rs3h_data_1_n142), .Y(bypass_rs3h_data_btwn_mux[17]));
INVX1 exu_U4827(.A(irf_byp_rs3h_data_d_l[16]), .Y(bypass_mux_rs3h_data_2_in1[16]));
OR2X1 exu_U4828(.A(exu_n13479), .B(bypass_mux_rs3h_data_1_n148), .Y(bypass_rs3h_data_btwn_mux[16]));
INVX1 exu_U4829(.A(irf_byp_rs3h_data_d_l[15]), .Y(bypass_mux_rs3h_data_2_in1[15]));
OR2X1 exu_U4830(.A(exu_n13480), .B(bypass_mux_rs3h_data_1_n154), .Y(bypass_rs3h_data_btwn_mux[15]));
INVX1 exu_U4831(.A(irf_byp_rs3h_data_d_l[14]), .Y(bypass_mux_rs3h_data_2_in1[14]));
OR2X1 exu_U4832(.A(exu_n13481), .B(bypass_mux_rs3h_data_1_n160), .Y(bypass_rs3h_data_btwn_mux[14]));
INVX1 exu_U4833(.A(irf_byp_rs3h_data_d_l[13]), .Y(bypass_mux_rs3h_data_2_in1[13]));
OR2X1 exu_U4834(.A(exu_n13482), .B(bypass_mux_rs3h_data_1_n166), .Y(bypass_rs3h_data_btwn_mux[13]));
INVX1 exu_U4835(.A(irf_byp_rs3h_data_d_l[12]), .Y(bypass_mux_rs3h_data_2_in1[12]));
OR2X1 exu_U4836(.A(exu_n13483), .B(bypass_mux_rs3h_data_1_n172), .Y(bypass_rs3h_data_btwn_mux[12]));
INVX1 exu_U4837(.A(irf_byp_rs3h_data_d_l[11]), .Y(bypass_mux_rs3h_data_2_in1[11]));
OR2X1 exu_U4838(.A(exu_n13484), .B(bypass_mux_rs3h_data_1_n178), .Y(bypass_rs3h_data_btwn_mux[11]));
INVX1 exu_U4839(.A(irf_byp_rs3h_data_d_l[10]), .Y(bypass_mux_rs3h_data_2_in1[10]));
OR2X1 exu_U4840(.A(exu_n13485), .B(bypass_mux_rs3h_data_1_n184), .Y(bypass_rs3h_data_btwn_mux[10]));
INVX1 exu_U4841(.A(irf_byp_rs3h_data_d_l[9]), .Y(bypass_mux_rs3h_data_2_in1[9]));
OR2X1 exu_U4842(.A(exu_n13455), .B(bypass_mux_rs3h_data_1_n4), .Y(bypass_rs3h_data_btwn_mux[9]));
INVX1 exu_U4843(.A(irf_byp_rs3h_data_d_l[8]), .Y(bypass_mux_rs3h_data_2_in1[8]));
OR2X1 exu_U4844(.A(exu_n13456), .B(bypass_mux_rs3h_data_1_n10), .Y(bypass_rs3h_data_btwn_mux[8]));
INVX1 exu_U4845(.A(irf_byp_rs3h_data_d_l[7]), .Y(bypass_mux_rs3h_data_2_in1[7]));
OR2X1 exu_U4846(.A(exu_n13457), .B(bypass_mux_rs3h_data_1_n16), .Y(bypass_rs3h_data_btwn_mux[7]));
INVX1 exu_U4847(.A(irf_byp_rs3h_data_d_l[6]), .Y(bypass_mux_rs3h_data_2_in1[6]));
OR2X1 exu_U4848(.A(exu_n13458), .B(bypass_mux_rs3h_data_1_n22), .Y(bypass_rs3h_data_btwn_mux[6]));
INVX1 exu_U4849(.A(irf_byp_rs3h_data_d_l[5]), .Y(bypass_mux_rs3h_data_2_in1[5]));
OR2X1 exu_U4850(.A(exu_n13459), .B(bypass_mux_rs3h_data_1_n28), .Y(bypass_rs3h_data_btwn_mux[5]));
INVX1 exu_U4851(.A(irf_byp_rs3h_data_d_l[4]), .Y(bypass_mux_rs3h_data_2_in1[4]));
OR2X1 exu_U4852(.A(exu_n13460), .B(bypass_mux_rs3h_data_1_n34), .Y(bypass_rs3h_data_btwn_mux[4]));
INVX1 exu_U4853(.A(irf_byp_rs3h_data_d_l[3]), .Y(bypass_mux_rs3h_data_2_in1[3]));
OR2X1 exu_U4854(.A(exu_n13461), .B(bypass_mux_rs3h_data_1_n40), .Y(bypass_rs3h_data_btwn_mux[3]));
INVX1 exu_U4855(.A(irf_byp_rs3h_data_d_l[2]), .Y(bypass_mux_rs3h_data_2_in1[2]));
OR2X1 exu_U4856(.A(exu_n13464), .B(bypass_mux_rs3h_data_1_n58), .Y(bypass_rs3h_data_btwn_mux[2]));
INVX1 exu_U4857(.A(irf_byp_rs3h_data_d_l[1]), .Y(bypass_mux_rs3h_data_2_in1[1]));
OR2X1 exu_U4858(.A(exu_n13475), .B(bypass_mux_rs3h_data_1_n124), .Y(bypass_rs3h_data_btwn_mux[1]));
INVX1 exu_U4859(.A(irf_byp_rs3h_data_d_l[0]), .Y(bypass_mux_rs3h_data_2_in1[0]));
OR2X1 exu_U4860(.A(exu_n13486), .B(bypass_mux_rs3h_data_1_n190), .Y(bypass_rs3h_data_btwn_mux[0]));
INVX1 exu_U4861(.A(bypass_rs3h_data_dff_n1), .Y(exu_n16134));
INVX1 exu_U4862(.A(se), .Y(bypass_rs3h_data_dff_n1));
INVX1 exu_U4863(.A(bypass_dfill_data_dff_n1), .Y(exu_n16140));
INVX1 exu_U4864(.A(bypass_dfill_data_dff_n1), .Y(exu_n16141));
AND2X1 exu_U4865(.A(exu_n96), .B(exu_n5063), .Y(exu_n17094));
AND2X1 exu_U4866(.A(exu_n97), .B(exu_n5064), .Y(exu_n17099));
AND2X1 exu_U4867(.A(exu_n98), .B(exu_n5065), .Y(exu_n17104));
AND2X1 exu_U4868(.A(exu_n99), .B(exu_n5066), .Y(exu_n17109));
AND2X1 exu_U4869(.A(exu_n100), .B(exu_n5067), .Y(exu_n17114));
AND2X1 exu_U4870(.A(exu_n101), .B(exu_n5068), .Y(exu_n17119));
AND2X1 exu_U4871(.A(exu_n102), .B(exu_n5069), .Y(exu_n17124));
AND2X1 exu_U4872(.A(exu_n103), .B(exu_n5070), .Y(exu_n17129));
AND2X1 exu_U4873(.A(exu_n104), .B(exu_n5071), .Y(exu_n17136));
AND2X1 exu_U4874(.A(exu_n105), .B(exu_n5072), .Y(exu_n17141));
AND2X1 exu_U4875(.A(exu_n106), .B(exu_n5073), .Y(exu_n17146));
AND2X1 exu_U4876(.A(exu_n107), .B(exu_n5074), .Y(exu_n17151));
AND2X1 exu_U4877(.A(exu_n108), .B(exu_n5075), .Y(exu_n17156));
AND2X1 exu_U4878(.A(exu_n109), .B(exu_n5076), .Y(exu_n17161));
AND2X1 exu_U4879(.A(exu_n110), .B(exu_n5077), .Y(exu_n17166));
AND2X1 exu_U4880(.A(exu_n111), .B(exu_n5078), .Y(exu_n17171));
AND2X1 exu_U4881(.A(exu_n112), .B(exu_n5079), .Y(exu_n17176));
AND2X1 exu_U4882(.A(exu_n113), .B(exu_n5080), .Y(exu_n17181));
AND2X1 exu_U4883(.A(exu_n114), .B(exu_n5081), .Y(exu_n17188));
AND2X1 exu_U4884(.A(exu_n115), .B(exu_n5082), .Y(exu_n17193));
AND2X1 exu_U4885(.A(exu_n116), .B(exu_n5083), .Y(exu_n17198));
AND2X1 exu_U4886(.A(exu_n117), .B(exu_n5084), .Y(alu_ecl_cout32_e));
AND2X1 exu_U4887(.A(exu_n118), .B(exu_n5085), .Y(exu_n17294));
AND2X1 exu_U4888(.A(exu_n119), .B(exu_n5086), .Y(exu_n17346));
AND2X1 exu_U4889(.A(exu_n120), .B(exu_n5087), .Y(exu_n17362));
AND2X1 exu_U4890(.A(exu_n121), .B(exu_n5088), .Y(exu_n17364));
AND2X1 exu_U4891(.A(exu_n122), .B(exu_n5089), .Y(exu_n17366));
AND2X1 exu_U4892(.A(exu_n123), .B(exu_n5090), .Y(exu_n17368));
AND2X1 exu_U4893(.A(exu_n124), .B(exu_n5091), .Y(exu_n17370));
AND2X1 exu_U4894(.A(exu_n125), .B(exu_n5092), .Y(exu_n17372));
AND2X1 exu_U4895(.A(exu_n126), .B(exu_n5093), .Y(exu_n17374));
AND2X1 exu_U4896(.A(exu_n127), .B(exu_n5094), .Y(exu_n17248));
AND2X1 exu_U4897(.A(exu_n128), .B(exu_n5095), .Y(exu_n17253));
AND2X1 exu_U4898(.A(exu_n129), .B(exu_n5096), .Y(exu_n17258));
AND2X1 exu_U4899(.A(exu_n130), .B(exu_n5097), .Y(exu_n17263));
AND2X1 exu_U4900(.A(exu_n131), .B(exu_n5098), .Y(exu_n17268));
AND2X1 exu_U4901(.A(exu_n132), .B(exu_n5099), .Y(exu_n17273));
AND2X1 exu_U4902(.A(exu_n18149), .B(exu_n5287), .Y(ecl_ccr_partial_cc_d[0]));
AND2X1 exu_U4903(.A(exu_n377), .B(exu_n5288), .Y(exu_n18149));
AND2X1 exu_U4904(.A(exu_n18145), .B(exu_n5285), .Y(ecl_ccr_partial_cc_d[1]));
AND2X1 exu_U4905(.A(exu_n376), .B(exu_n5286), .Y(exu_n18145));
AND2X1 exu_U4906(.A(exu_n18141), .B(exu_n5283), .Y(ecl_ccr_partial_cc_d[2]));
AND2X1 exu_U4907(.A(exu_n375), .B(exu_n5284), .Y(exu_n18141));
AND2X1 exu_U4908(.A(exu_n18137), .B(exu_n5281), .Y(ecl_ccr_partial_cc_d[3]));
AND2X1 exu_U4909(.A(exu_n374), .B(exu_n5282), .Y(exu_n18137));
AND2X1 exu_U4910(.A(exu_n18133), .B(exu_n5279), .Y(ecl_ccr_partial_cc_d[4]));
AND2X1 exu_U4911(.A(exu_n373), .B(exu_n5280), .Y(exu_n18133));
AND2X1 exu_U4912(.A(exu_n18129), .B(exu_n5277), .Y(ecl_ccr_partial_cc_d[5]));
AND2X1 exu_U4913(.A(exu_n372), .B(exu_n5278), .Y(exu_n18129));
AND2X1 exu_U4914(.A(exu_n18125), .B(exu_n5275), .Y(ecl_ccr_partial_cc_d[6]));
AND2X1 exu_U4915(.A(exu_n371), .B(exu_n5276), .Y(exu_n18125));
AND2X1 exu_U4916(.A(exu_n18121), .B(exu_n5273), .Y(ecl_ccr_partial_cc_d[7]));
AND2X1 exu_U4917(.A(exu_n370), .B(exu_n5274), .Y(exu_n18121));
OR2X1 exu_U4918(.A(exu_n15742), .B(exu_n15768), .Y(ecl_writeback_n121));
AND2X1 exu_U4919(.A(ecl_writeback_n110), .B(ecl_writeback_restore_tid[0]), .Y(ecl_writeback_n101));
OR2X1 exu_U4920(.A(exu_n13395), .B(exu_n14706), .Y(alu_regzcmp_high_nonzero));
OR2X1 exu_U4921(.A(exu_n13394), .B(exu_n14705), .Y(alu_regzcmp_low_nonzero));
OR2X1 exu_U4922(.A(rml_rml_ecl_cansave_e[2]), .B(rml_rml_ecl_cansave_e[1]), .Y(rml_n121));
AND2X1 exu_U4923(.A(exu_n93), .B(exu_n5060), .Y(exu_n17213));
AND2X1 exu_U4924(.A(exu_n94), .B(exu_n5061), .Y(exu_n17215));
AND2X1 exu_U4925(.A(exu_n95), .B(exu_n5062), .Y(exu_n17089));
INVX1 exu_U4926(.A(exu_n16162), .Y(exu_n16168));
AND2X1 exu_U4927(.A(exu_n86), .B(exu_n5053), .Y(exu_n17135));
AND2X1 exu_U4928(.A(exu_n87), .B(exu_n5054), .Y(exu_n17187));
AND2X1 exu_U4929(.A(exu_n88), .B(exu_n5055), .Y(exu_n17203));
AND2X1 exu_U4930(.A(exu_n89), .B(exu_n5056), .Y(exu_n17205));
AND2X1 exu_U4931(.A(exu_n90), .B(exu_n5057), .Y(exu_n17207));
AND2X1 exu_U4932(.A(exu_n91), .B(exu_n5058), .Y(exu_n17209));
AND2X1 exu_U4933(.A(exu_n92), .B(exu_n5059), .Y(exu_n17211));
INVX1 exu_U4934(.A(ecl_early_ttype_m[7]), .Y(exu_n16403));
INVX1 exu_U4935(.A(exu_tlu_ue_trap_m), .Y(exu_n16595));
AND2X1 exu_U4936(.A(ecl_mdqctl_div_zero_unqual_m), .B(ecl_mdqctl_isdiv_m), .Y(ecl_div_zero_m));
AND2X1 exu_U4937(.A(exu_n4138), .B(exu_n9114), .Y(rml_mux_agp_out1_n8));
AND2X1 exu_U4938(.A(exu_n4136), .B(exu_n9112), .Y(rml_mux_agp_out1_n2));
AND2X1 exu_U4939(.A(rml_cwp_swap_state[0]), .B(rml_cwp_N99), .Y(rml_swap_locals_ins));
OR2X1 exu_U4940(.A(exu_n13407), .B(exu_n14718), .Y(rml_cwp_swap_state[0]));
OR2X1 exu_U4941(.A(rml_n55), .B(exu_n14808), .Y(rml_n49));
OR2X1 exu_U4942(.A(rml_save_e), .B(rml_swap_locals_ins), .Y(rml_n55));
OR2X1 exu_U4943(.A(exu_n12098), .B(exu_n13514), .Y(rml_rml_ecl_cwp_e[0]));
AND2X1 exu_U4944(.A(exu_n245), .B(exu_n5172), .Y(exu_n17776));
OR2X1 exu_U4945(.A(exu_n13411), .B(exu_n14722), .Y(rml_cwp_old_swap_cwp[0]));
OR2X1 exu_U4946(.A(exu_n12097), .B(exu_n13513), .Y(rml_rml_ecl_cwp_e[1]));
AND2X1 exu_U4947(.A(exu_n243), .B(exu_n5170), .Y(exu_n17770));
OR2X1 exu_U4948(.A(exu_n13405), .B(exu_n14716), .Y(rml_cwp_old_swap_cwp[1]));
OR2X1 exu_U4949(.A(exu_n12096), .B(exu_n13512), .Y(rml_rml_ecl_cwp_e[2]));
AND2X1 exu_U4950(.A(exu_n241), .B(exu_n5168), .Y(exu_n17764));
OR2X1 exu_U4951(.A(exu_n13404), .B(exu_n14715), .Y(rml_cwp_old_swap_cwp[2]));
AND2X1 exu_U4952(.A(exu_n3965), .B(exu_n8980), .Y(exu_n31464));
AND2X1 exu_U4953(.A(exu_n3963), .B(exu_n8978), .Y(exu_n31458));
AND2X1 exu_U4954(.A(exu_n11688), .B(exu_n9341), .Y(ecl_writeback_n172));
AND2X1 exu_U4955(.A(exu_n11685), .B(exu_n9340), .Y(ecl_writeback_n166));
AND2X1 exu_U4956(.A(exu_n4094), .B(exu_n9088), .Y(ecl_writeback_rd_g_mux_n26));
AND2X1 exu_U4957(.A(exu_n4092), .B(exu_n9086), .Y(ecl_writeback_rd_g_mux_n20));
AND2X1 exu_U4958(.A(exu_n4090), .B(exu_n9084), .Y(ecl_writeback_rd_g_mux_n14));
AND2X1 exu_U4959(.A(exu_n4088), .B(exu_n9082), .Y(ecl_writeback_rd_g_mux_n8));
AND2X1 exu_U4960(.A(exu_n4086), .B(exu_n9080), .Y(ecl_writeback_rd_g_mux_n2));
AND2X1 exu_U4961(.A(exu_n320), .B(exu_n5247), .Y(exu_n18006));
AND2X1 exu_U4962(.A(exu_n318), .B(exu_n5245), .Y(exu_n18000));
AND2X1 exu_U4963(.A(exu_n316), .B(exu_n5243), .Y(exu_n17994));
AND2X1 exu_U4964(.A(exu_n314), .B(exu_n5241), .Y(exu_n17988));
AND2X1 exu_U4965(.A(exu_n312), .B(exu_n5239), .Y(exu_n17982));
AND2X1 exu_U4966(.A(ecl_writeback_wb_w), .B(ecl_writeback_n149), .Y(ecl_writeback_n148));
AND2X1 exu_U4967(.A(rml_cwp_swap_slot1_state[1]), .B(exu_n9119), .Y(rml_cwp_swap_slot1_state_valid[1]));
AND2X1 exu_U4968(.A(rml_cwp_n43), .B(exu_n15342), .Y(rml_cwp_swap_keep_state[1]));
AND2X1 exu_U4969(.A(exu_n15554), .B(rml_cwp_cwpccr_update_w), .Y(rml_cwp_n75));
AND2X1 exu_U4970(.A(rml_cwp_swap_slot2_state[1]), .B(exu_n9118), .Y(rml_cwp_swap_slot2_state_valid[1]));
AND2X1 exu_U4971(.A(rml_cwp_n41), .B(exu_n15341), .Y(rml_cwp_swap_keep_state[2]));
AND2X1 exu_U4972(.A(exu_n15555), .B(rml_cwp_cwpccr_update_w), .Y(rml_cwp_n76));
AND2X1 exu_U4973(.A(rml_cwp_swap_slot3_state[1]), .B(exu_n9117), .Y(rml_cwp_swap_slot3_state_valid[1]));
AND2X1 exu_U4974(.A(rml_cwp_n39), .B(exu_n15340), .Y(rml_cwp_swap_keep_state[3]));
AND2X1 exu_U4975(.A(exu_n15556), .B(rml_cwp_cwpccr_update_w), .Y(rml_cwp_n77));
INVX1 exu_U4976(.A(ecl_divcntl_div_state_1), .Y(exu_n16438));
AND2X1 exu_U4977(.A(ecl_divcntl_cnt6_n11), .B(exu_n9060), .Y(ecl_divcntl_cnt6_n10));
AND2X1 exu_U4978(.A(ecl_divcntl_cntr[4]), .B(ecl_divcntl_cntr[3]), .Y(ecl_divcntl_cnt6_n11));
OR2X1 exu_U4979(.A(exu_n16622), .B(ecl_divcntl_cntr[4]), .Y(ecl_divcntl_cnt6_n16));
AND2X1 exu_U4980(.A(ecl_divcntl_cntr[4]), .B(exu_n9061), .Y(ecl_divcntl_cnt6_n14));
INVX1 exu_U4981(.A(se), .Y(exu_n17619));
INVX1 exu_U4982(.A(se), .Y(exu_n18198));
INVX1 exu_U4983(.A(se), .Y(exu_n18202));
INVX1 exu_U4984(.A(se), .Y(exu_n18206));
INVX1 exu_U4985(.A(se), .Y(exu_n18210));
INVX1 exu_U4986(.A(se), .Y(exu_n18242));
INVX1 exu_U4987(.A(se), .Y(exu_n18246));
INVX1 exu_U4988(.A(se), .Y(exu_n18250));
INVX1 exu_U4989(.A(se), .Y(exu_n18254));
INVX1 exu_U4990(.A(se), .Y(exu_n18286));
INVX1 exu_U4991(.A(se), .Y(exu_n18290));
INVX1 exu_U4992(.A(se), .Y(exu_n18294));
INVX1 exu_U4993(.A(se), .Y(exu_n18298));
AND2X1 exu_U4994(.A(rml_hi_wstate_reg_data_thr3[1]), .B(exu_n15194), .Y(exu_n18345));
AND2X1 exu_U4995(.A(rml_hi_wstate_reg_data_thr3[2]), .B(exu_n15194), .Y(exu_n18343));
INVX1 exu_U4996(.A(se), .Y(exu_n18330));
AND2X1 exu_U4997(.A(rml_hi_wstate_reg_data_thr2[1]), .B(exu_n15195), .Y(exu_n18351));
AND2X1 exu_U4998(.A(rml_hi_wstate_reg_data_thr2[2]), .B(exu_n15195), .Y(exu_n18349));
INVX1 exu_U4999(.A(se), .Y(exu_n18334));
AND2X1 exu_U5000(.A(rml_hi_wstate_reg_data_thr1[1]), .B(exu_n15196), .Y(exu_n18357));
AND2X1 exu_U5001(.A(rml_hi_wstate_reg_data_thr1[2]), .B(exu_n15196), .Y(exu_n18355));
INVX1 exu_U5002(.A(se), .Y(exu_n18338));
AND2X1 exu_U5003(.A(rml_hi_wstate_reg_data_thr0[1]), .B(exu_n15197), .Y(exu_n18363));
AND2X1 exu_U5004(.A(rml_hi_wstate_reg_data_thr0[2]), .B(exu_n15197), .Y(exu_n18361));
INVX1 exu_U5005(.A(se), .Y(exu_n18342));
INVX1 exu_U5006(.A(se), .Y(exu_n18370));
INVX1 exu_U5007(.A(se), .Y(exu_n18374));
INVX1 exu_U5008(.A(se), .Y(exu_n18378));
INVX1 exu_U5009(.A(se), .Y(exu_n18382));
AND2X1 exu_U5010(.A(rml_cwp_swap_req_vec[3]), .B(exu_n9046), .Y(rml_cwp_next_swap_thr[3]));
AND2X1 exu_U5011(.A(rml_cwp_swap_req_vec[2]), .B(exu_n9047), .Y(rml_cwp_next_swap_thr[2]));
INVX1 exu_U5012(.A(rml_cwp_cwp_output_queue_pv[1]), .Y(exu_n16617));
AND2X1 exu_U5013(.A(rml_cwp_swap_req_vec[1]), .B(exu_n9049), .Y(rml_cwp_next_swap_thr[1]));
AND2X1 exu_U5014(.A(exu_n4034), .B(exu_n9051), .Y(rml_cwp_next_swap_thr[0]));
INVX1 exu_U5015(.A(se), .Y(exu_n18407));
AND2X1 exu_U5016(.A(exu_n4147), .B(rml_cwp_n96), .Y(rml_cwp_n47));
INVX1 exu_U5017(.A(se), .Y(exu_n18412));
OR2X1 exu_U5018(.A(exu_n13399), .B(exu_n14710), .Y(rml_cwp_swap_data[7]));
AND2X1 exu_U5019(.A(exu_n4005), .B(exu_n9021), .Y(rml_cwp_cwp_output_mux_n13));
OR2X1 exu_U5020(.A(exu_n13406), .B(exu_n14717), .Y(rml_cwp_swap_state[1]));
AND2X1 exu_U5021(.A(exu_n4022), .B(exu_n9038), .Y(rml_cwp_cwp_output_mux_n68));
AND2X1 exu_U5022(.A(exu_n4023), .B(exu_n9039), .Y(rml_cwp_cwp_output_mux_n67));
AND2X1 exu_U5023(.A(exu_n736), .B(exu_n5414), .Y(exu_n19002));
AND2X1 exu_U5024(.A(exu_n736), .B(exu_n5415), .Y(exu_n19005));
AND2X1 exu_U5025(.A(exu_n736), .B(exu_n5416), .Y(exu_n19008));
AND2X1 exu_U5026(.A(exu_n736), .B(exu_n5417), .Y(exu_n19011));
AND2X1 exu_U5027(.A(exu_n736), .B(exu_n5419), .Y(exu_n19018));
AND2X1 exu_U5028(.A(exu_n736), .B(exu_n5420), .Y(exu_n19021));
AND2X1 exu_U5029(.A(exu_n736), .B(exu_n5421), .Y(exu_n19024));
AND2X1 exu_U5030(.A(exu_n736), .B(exu_n5422), .Y(exu_n19027));
AND2X1 exu_U5031(.A(exu_n736), .B(exu_n5423), .Y(exu_n19030));
AND2X1 exu_U5032(.A(exu_n736), .B(exu_n5424), .Y(exu_n19033));
AND2X1 exu_U5033(.A(exu_n736), .B(exu_n5425), .Y(exu_n19036));
AND2X1 exu_U5034(.A(exu_n736), .B(exu_n5426), .Y(exu_n19039));
AND2X1 exu_U5035(.A(exu_n736), .B(exu_n5427), .Y(exu_n19042));
AND2X1 exu_U5036(.A(exu_n736), .B(exu_n5428), .Y(exu_n19045));
AND2X1 exu_U5037(.A(exu_n631), .B(exu_n5363), .Y(exu_n18824));
AND2X1 exu_U5038(.A(exu_n631), .B(exu_n5364), .Y(exu_n18827));
AND2X1 exu_U5039(.A(exu_n631), .B(exu_n5365), .Y(exu_n18830));
AND2X1 exu_U5040(.A(exu_n631), .B(exu_n5366), .Y(exu_n18833));
AND2X1 exu_U5041(.A(exu_n631), .B(exu_n5367), .Y(exu_n18836));
AND2X1 exu_U5042(.A(exu_n631), .B(exu_n5369), .Y(exu_n18843));
AND2X1 exu_U5043(.A(exu_n631), .B(exu_n5370), .Y(exu_n18846));
AND2X1 exu_U5044(.A(exu_n631), .B(exu_n5371), .Y(exu_n18849));
AND2X1 exu_U5045(.A(exu_n631), .B(exu_n5372), .Y(exu_n18852));
AND2X1 exu_U5046(.A(exu_n631), .B(exu_n5373), .Y(exu_n18855));
AND2X1 exu_U5047(.A(exu_n631), .B(exu_n5374), .Y(exu_n18858));
AND2X1 exu_U5048(.A(exu_n631), .B(exu_n5375), .Y(exu_n18861));
AND2X1 exu_U5049(.A(exu_n631), .B(exu_n5376), .Y(exu_n18864));
INVX1 exu_U5050(.A(exu_n16002), .Y(exu_n15992));
INVX1 exu_U5051(.A(exu_n16002), .Y(exu_n15991));
INVX1 exu_U5052(.A(exu_n16003), .Y(exu_n15990));
INVX1 exu_U5053(.A(exu_n18474), .Y(exu_n16003));
INVX1 exu_U5054(.A(exu_n16000), .Y(exu_n15999));
INVX1 exu_U5055(.A(exu_n16000), .Y(exu_n15998));
INVX1 exu_U5056(.A(exu_n16000), .Y(exu_n15997));
INVX1 exu_U5057(.A(exu_n16001), .Y(exu_n15996));
INVX1 exu_U5058(.A(exu_n16001), .Y(exu_n15995));
INVX1 exu_U5059(.A(exu_n16001), .Y(exu_n15994));
INVX1 exu_U5060(.A(exu_n16002), .Y(exu_n15993));
INVX1 exu_U5061(.A(ecl_muls_e), .Y(exu_n16614));
OR2X1 exu_U5062(.A(exu_n13453), .B(exu_n14773), .Y(ecl_div_ecl_yreg_0_d));
AND2X1 exu_U5063(.A(exu_n4579), .B(exu_n9359), .Y(ecl_yreg0_mux_n1));
AND2X1 exu_U5064(.A(exu_n4486), .B(exu_n9305), .Y(alu_chk_mem_addr_n1));
AND2X1 exu_U5065(.A(exu_n4485), .B(exu_n9304), .Y(alu_chk_mem_addr_n2));
INVX1 exu_U5066(.A(ecl_ifu_exu_range_check_jlret_e), .Y(exu_n16609));
OR2X1 exu_U5067(.A(exu_n13500), .B(exu_n14818), .Y(ecl_n62));
AND2X1 exu_U5068(.A(exu_n4966), .B(exu_n16595), .Y(ecl_n81));
AND2X1 exu_U5069(.A(exu_n16392), .B(exu_n15239), .Y(ecl_n112));
AND2X1 exu_U5070(.A(ecl_ifu_exu_range_check_jlret_e), .B(ecl_n113), .Y(ecl_misalign_addr_e));
OR2X1 exu_U5071(.A(exu_ifu_brpc_e[0]), .B(exu_ifu_brpc_e[1]), .Y(ecl_n113));
AND2X1 exu_U5072(.A(exu_n4900), .B(exu_n9618), .Y(rml_ecl_clean_window_e));
OR2X1 exu_U5073(.A(exu_n15940), .B(exu_n15030), .Y(rml_rml_ecl_kill_e));
OR2X1 exu_U5074(.A(rml_ecl_otherwin_d[0]), .B(rml_n95), .Y(rml_rml_ecl_other_d));
OR2X1 exu_U5075(.A(rml_ecl_otherwin_d[2]), .B(rml_ecl_otherwin_d[1]), .Y(rml_n95));
AND2X1 exu_U5076(.A(ecl_rml_cwp_wen_e), .B(exu_n15685), .Y(rml_n50));
INVX1 exu_U5077(.A(rml_save_m), .Y(exu_n16605));
AND2X1 exu_U5078(.A(ecl_rml_cwp_wen_e), .B(exu_n9615), .Y(rml_n97));
OR2X1 exu_U5079(.A(exu_n15360), .B(exu_n14812), .Y(rml_cansave_wen_e));
AND2X1 exu_U5080(.A(exu_n4897), .B(exu_n16383), .Y(rml_n104));
OR2X1 exu_U5081(.A(exu_n15360), .B(exu_n14813), .Y(rml_canrestore_wen_e));
AND2X1 exu_U5082(.A(exu_n4899), .B(exu_n16385), .Y(rml_n109));
AND2X1 exu_U5083(.A(rml_rml_ecl_cleanwin_e[2]), .B(rml_rml_ecl_cleanwin_e[0]), .Y(rml_n101));
INVX1 exu_U5084(.A(ecl_ccr_setcc_e), .Y(exu_n16602));
AND2X1 exu_U5085(.A(ecl_writeback_n153), .B(exu_n9338), .Y(ecl_writeback_n152));
AND2X1 exu_U5086(.A(exu_n11675), .B(exu_n9328), .Y(ecl_writeback_n47));
INVX1 exu_U5087(.A(exu_ffu_wsr_inst_e), .Y(exu_n16598));
AND2X1 exu_U5088(.A(exu_n4527), .B(ifu_exu_inst_vld_e), .Y(ecl_writeback_n59));
INVX1 exu_U5089(.A(ecl_writeback_restore_ready), .Y(exu_n16597));
INVX1 exu_U5090(.A(ecl_rml_kill_e), .Y(exu_n16389));
OR2X1 exu_U5091(.A(exu_n13442), .B(exu_n14809), .Y(ecl_writeback_n66));
AND2X1 exu_U5092(.A(ecc_chk_rs3_parity), .B(ecl_ecc_rs3_use_rf_e), .Y(ecc_ecl_rs3_ce));
AND2X1 exu_U5093(.A(exu_n4522), .B(exu_n15353), .Y(ecl_eccctl_n18));
AND2X1 exu_U5094(.A(ecl_wb_eccctl_spec_wen_next), .B(ifu_exu_inj_irferr), .Y(ecl_eccctl_inj_irferr_m));
OR2X1 exu_U5095(.A(ecl_writeback_n52), .B(ecl_writeback_n53), .Y(ecl_wb_eccctl_spec_wen_next));
OR2X1 exu_U5096(.A(ecl_writeback_valid_m), .B(exu_n15236), .Y(ecl_writeback_n52));
OR2X1 exu_U5097(.A(ecl_writeback_n54), .B(ecl_writeback_n51), .Y(ecl_writeback_n53));
AND2X1 exu_U5098(.A(ecl_ecc_rs1_use_rf_e), .B(ecc_chk_rs1_n2), .Y(ecc_ecl_rs1_ue));
AND2X1 exu_U5099(.A(exu_n4587), .B(exu_n16397), .Y(ecc_chk_rs1_n2));
INVX1 exu_U5100(.A(ecc_chk_rs1_parity), .Y(exu_n16397));
AND2X1 exu_U5101(.A(ecc_chk_rs1_parity), .B(ecl_ecc_rs1_use_rf_e), .Y(ecc_ecl_rs1_ce));
AND2X1 exu_U5102(.A(ecl_ecc_rs2_use_rf_e), .B(exu_n19996), .Y(ecc_ecl_rs2_ue));
AND2X1 exu_U5103(.A(exu_n782), .B(exu_n16515), .Y(exu_n19996));
INVX1 exu_U5104(.A(ecc_chk_rs2_parity), .Y(exu_n16515));
AND2X1 exu_U5105(.A(ecc_chk_rs2_parity), .B(ecl_ecc_rs2_use_rf_e), .Y(ecc_ecl_rs2_ce));
AND2X1 exu_U5106(.A(ecl_ecc_rs3_use_rf_e), .B(exu_n20132), .Y(ecc_ecl_rs3_ue));
AND2X1 exu_U5107(.A(exu_n784), .B(exu_n16513), .Y(exu_n20132));
AND2X1 exu_U5108(.A(exu_n15491), .B(exu_n5297), .Y(ecl_divcntl_qnext_cout_mux_n2));
AND2X1 exu_U5109(.A(exu_n10778), .B(exu_n5298), .Y(ecl_divcntl_q_next_nocout[1]));
AND2X1 exu_U5110(.A(exu_n10781), .B(exu_n9773), .Y(ecl_divcntl_sub_next_nocout[1]));
AND2X1 exu_U5111(.A(exu_n15491), .B(exu_n5299), .Y(exu_n17617));
OR2X1 exu_U5112(.A(ecl_divcntl_n54), .B(ecl_divcntl_zero_rem_q), .Y(ecl_divcntl_n53));
AND2X1 exu_U5113(.A(exu_n4509), .B(exu_n16206), .Y(ecl_divcntl_n52));
INVX1 exu_U5114(.A(ecl_ecl_div_signed_div), .Y(exu_n16508));
OR2X1 exu_U5115(.A(ifu_exu_muldivop_d[3]), .B(ifu_exu_muls_d), .Y(ecl_mdqctl_new_div_vld));
AND2X1 exu_U5116(.A(ecl_mdqctl_n55), .B(exu_n9307), .Y(ecl_mdqctl_n51));
AND2X1 exu_U5117(.A(exu_n4501), .B(exu_n16387), .Y(ecl_mdqctl_n55));
INVX1 exu_U5118(.A(mul_exu_ack), .Y(exu_n16371));
AND2X1 exu_U5119(.A(ecl_mdqctl_n20), .B(exu_n15985), .Y(ecl_mdqctl_n22));
OR2X1 exu_U5120(.A(exu_n16186), .B(ecl_mdqctl_divcntl_muldone), .Y(ecl_mdqctl_n13));
OR2X1 exu_U5121(.A(exu_n12099), .B(exu_n13515), .Y(rml_cwp_trap_old_cwp_m[2]));
INVX1 exu_U5122(.A(se), .Y(exu_n19670));
INVX1 exu_U5123(.A(se), .Y(exu_n19674));
AND2X1 exu_U5124(.A(rml_next_cwp_mux_n1), .B(exu_n9127), .Y(rml_next_cwp_e[2]));
AND2X1 exu_U5125(.A(exu_n4152), .B(exu_n9128), .Y(rml_next_cwp_mux_n1));
AND2X1 exu_U5126(.A(rml_next_cwp_mux_n5), .B(exu_n9129), .Y(rml_next_cwp_e[1]));
AND2X1 exu_U5127(.A(exu_n4153), .B(exu_n9130), .Y(rml_next_cwp_mux_n5));
AND2X1 exu_U5128(.A(rml_next_cwp_mux_n9), .B(exu_n9131), .Y(rml_next_cwp_e[0]));
AND2X1 exu_U5129(.A(exu_n4154), .B(exu_n9132), .Y(rml_next_cwp_mux_n9));
INVX1 exu_U5130(.A(se), .Y(exu_n19678));
INVX1 exu_U5131(.A(se), .Y(exu_n19682));
INVX1 exu_U5132(.A(se), .Y(exu_n19686));
INVX1 exu_U5133(.A(se), .Y(exu_n19690));
INVX1 exu_U5134(.A(se), .Y(exu_n19694));
INVX1 exu_U5135(.A(se), .Y(exu_n19698));
AND2X1 exu_U5136(.A(rml_rml_ecl_otherwin_e[2]), .B(rml_n44), .Y(rml_rml_next_otherwin_e[2]));
OR2X1 exu_U5137(.A(rml_rml_ecl_otherwin_e[1]), .B(rml_rml_ecl_otherwin_e[0]), .Y(rml_n44));
INVX1 exu_U5138(.A(se), .Y(exu_n19702));
INVX1 exu_U5139(.A(se), .Y(exu_n19706));
AND2X1 exu_U5140(.A(exu_n16586), .B(exu_n9608), .Y(rml_rml_next_cleanwin_e[2]));
INVX1 exu_U5141(.A(rml_rml_ecl_cleanwin_e[0]), .Y(exu_n16585));
INVX1 exu_U5142(.A(se), .Y(exu_n19710));
INVX1 exu_U5143(.A(se), .Y(exu_n19714));
OR2X1 exu_U5144(.A(exu_n12114), .B(exu_n13530), .Y(rml_ecl_cansave_d[2]));
AND2X1 exu_U5145(.A(exu_n277), .B(exu_n5204), .Y(exu_n17872));
OR2X1 exu_U5146(.A(exu_n12115), .B(exu_n13531), .Y(rml_ecl_cansave_d[1]));
AND2X1 exu_U5147(.A(exu_n279), .B(exu_n5206), .Y(exu_n17878));
OR2X1 exu_U5148(.A(exu_n12116), .B(exu_n13532), .Y(rml_ecl_cansave_d[0]));
AND2X1 exu_U5149(.A(exu_n281), .B(exu_n5208), .Y(exu_n17884));
INVX1 exu_U5150(.A(se), .Y(exu_n19718));
OR2X1 exu_U5151(.A(exu_n12117), .B(exu_n13533), .Y(rml_ecl_canrestore_d[2]));
AND2X1 exu_U5152(.A(exu_n283), .B(exu_n5210), .Y(exu_n17890));
OR2X1 exu_U5153(.A(exu_n12118), .B(exu_n13534), .Y(rml_ecl_canrestore_d[1]));
AND2X1 exu_U5154(.A(exu_n285), .B(exu_n5212), .Y(exu_n17896));
OR2X1 exu_U5155(.A(exu_n12119), .B(exu_n13535), .Y(rml_ecl_canrestore_d[0]));
AND2X1 exu_U5156(.A(exu_n287), .B(exu_n5214), .Y(exu_n17902));
INVX1 exu_U5157(.A(se), .Y(exu_n19722));
OR2X1 exu_U5158(.A(exu_n12120), .B(exu_n13536), .Y(rml_ecl_otherwin_d[2]));
AND2X1 exu_U5159(.A(exu_n289), .B(exu_n5216), .Y(exu_n17908));
OR2X1 exu_U5160(.A(exu_n12121), .B(exu_n13537), .Y(rml_ecl_otherwin_d[1]));
AND2X1 exu_U5161(.A(exu_n291), .B(exu_n5218), .Y(exu_n17914));
OR2X1 exu_U5162(.A(exu_n12122), .B(exu_n13538), .Y(rml_ecl_otherwin_d[0]));
AND2X1 exu_U5163(.A(exu_n293), .B(exu_n5220), .Y(exu_n17920));
INVX1 exu_U5164(.A(se), .Y(exu_n19726));
OR2X1 exu_U5165(.A(exu_n12123), .B(exu_n13539), .Y(rml_ecl_cleanwin_d[2]));
AND2X1 exu_U5166(.A(exu_n295), .B(exu_n5222), .Y(exu_n17926));
OR2X1 exu_U5167(.A(exu_n12124), .B(exu_n13540), .Y(rml_ecl_cleanwin_d[1]));
AND2X1 exu_U5168(.A(exu_n297), .B(exu_n5224), .Y(exu_n17932));
OR2X1 exu_U5169(.A(exu_n12125), .B(exu_n13541), .Y(rml_ecl_cleanwin_d[0]));
AND2X1 exu_U5170(.A(exu_n299), .B(exu_n5226), .Y(exu_n17938));
INVX1 exu_U5171(.A(se), .Y(exu_n19730));
OR2X1 exu_U5172(.A(ecl_mdqctl_div_data_7), .B(ecl_div_muls), .Y(ecl_mdqctl_wb_divsetcc_g));
OR2X1 exu_U5173(.A(exu_n12093), .B(exu_n13509), .Y(rml_ecl_cwp_d[2]));
AND2X1 exu_U5174(.A(exu_n235), .B(exu_n5162), .Y(exu_n17746));
OR2X1 exu_U5175(.A(exu_n12094), .B(exu_n13510), .Y(rml_ecl_cwp_d[1]));
AND2X1 exu_U5176(.A(exu_n237), .B(exu_n5164), .Y(exu_n17752));
OR2X1 exu_U5177(.A(exu_n12095), .B(exu_n13511), .Y(rml_ecl_cwp_d[0]));
AND2X1 exu_U5178(.A(exu_n239), .B(exu_n5166), .Y(exu_n17758));
INVX1 exu_U5179(.A(se), .Y(exu_n19738));
INVX1 exu_U5180(.A(se), .Y(exu_n19742));
INVX1 exu_U5181(.A(se), .Y(exu_n19746));
AND2X1 exu_U5182(.A(exu_n252), .B(exu_n5179), .Y(exu_n17801));
AND2X1 exu_U5183(.A(exu_n253), .B(exu_n5180), .Y(exu_n17800));
AND2X1 exu_U5184(.A(exu_n254), .B(exu_n5181), .Y(exu_n17807));
AND2X1 exu_U5185(.A(exu_n255), .B(exu_n5182), .Y(exu_n17806));
OR2X1 exu_U5186(.A(exu_n12104), .B(exu_n13520), .Y(rml_oddwin_w[0]));
AND2X1 exu_U5187(.A(exu_n257), .B(exu_n5184), .Y(exu_n17812));
INVX1 exu_U5188(.A(se), .Y(exu_n19750));
AND2X1 exu_U5189(.A(exu_n258), .B(exu_n5185), .Y(exu_n17819));
AND2X1 exu_U5190(.A(exu_n259), .B(exu_n5186), .Y(exu_n17818));
AND2X1 exu_U5191(.A(exu_n260), .B(exu_n5187), .Y(exu_n17825));
AND2X1 exu_U5192(.A(exu_n261), .B(exu_n5188), .Y(exu_n17824));
OR2X1 exu_U5193(.A(exu_n12107), .B(exu_n13523), .Y(rml_oddwin_w[1]));
AND2X1 exu_U5194(.A(exu_n263), .B(exu_n5190), .Y(exu_n17830));
INVX1 exu_U5195(.A(se), .Y(exu_n19754));
AND2X1 exu_U5196(.A(exu_n264), .B(exu_n5191), .Y(exu_n17837));
AND2X1 exu_U5197(.A(exu_n265), .B(exu_n5192), .Y(exu_n17836));
AND2X1 exu_U5198(.A(exu_n266), .B(exu_n5193), .Y(exu_n17843));
AND2X1 exu_U5199(.A(exu_n267), .B(exu_n5194), .Y(exu_n17842));
OR2X1 exu_U5200(.A(exu_n12110), .B(exu_n13526), .Y(rml_oddwin_w[2]));
AND2X1 exu_U5201(.A(exu_n269), .B(exu_n5196), .Y(exu_n17848));
INVX1 exu_U5202(.A(se), .Y(exu_n19758));
AND2X1 exu_U5203(.A(exu_n270), .B(exu_n5197), .Y(exu_n17855));
AND2X1 exu_U5204(.A(exu_n271), .B(exu_n5198), .Y(exu_n17854));
AND2X1 exu_U5205(.A(exu_n272), .B(exu_n5199), .Y(exu_n17861));
AND2X1 exu_U5206(.A(exu_n273), .B(exu_n5200), .Y(exu_n17860));
OR2X1 exu_U5207(.A(exu_n12113), .B(exu_n13529), .Y(rml_oddwin_w[3]));
AND2X1 exu_U5208(.A(exu_n275), .B(exu_n5202), .Y(exu_n17866));
INVX1 exu_U5209(.A(se), .Y(exu_n19762));
INVX1 exu_U5210(.A(se), .Y(exu_n19766));
INVX1 exu_U5211(.A(se), .Y(exu_n19770));
INVX1 exu_U5212(.A(se), .Y(exu_n19774));
INVX1 exu_U5213(.A(se), .Y(exu_n19778));
INVX1 exu_U5214(.A(se), .Y(exu_n19782));
INVX1 exu_U5215(.A(se), .Y(exu_n19785));
INVX1 exu_U5216(.A(se), .Y(exu_n19791));
INVX1 exu_U5217(.A(se), .Y(exu_n19794));
INVX1 exu_U5218(.A(se), .Y(ecl_writeback_restore_tid_dff_n2));
INVX1 exu_U5219(.A(se), .Y(exu_n19797));
INVX1 exu_U5220(.A(se), .Y(exu_n19800));
INVX1 exu_U5221(.A(se), .Y(exu_n19788));
INVX1 exu_U5222(.A(se), .Y(exu_n19803));
INVX1 exu_U5223(.A(se), .Y(exu_n19806));
INVX1 exu_U5224(.A(se), .Y(exu_n19809));
INVX1 exu_U5225(.A(se), .Y(exu_n19812));
INVX1 exu_U5226(.A(se), .Y(exu_n19815));
INVX1 exu_U5227(.A(se), .Y(exu_n19818));
INVX1 exu_U5228(.A(se), .Y(exu_n19734));
AND2X1 exu_U5229(.A(exu_n4886), .B(exu_n9610), .Y(rml_n63));
AND2X1 exu_U5230(.A(exu_n4887), .B(exu_n9611), .Y(rml_n62));
AND2X1 exu_U5231(.A(exu_n4888), .B(exu_n9612), .Y(rml_n72));
AND2X1 exu_U5232(.A(exu_n4889), .B(exu_n9613), .Y(rml_n71));
INVX1 exu_U5233(.A(se), .Y(exu_n19821));
INVX1 exu_U5234(.A(se), .Y(exu_n19824));
INVX1 exu_U5235(.A(se), .Y(exu_n19830));
INVX1 exu_U5236(.A(se), .Y(exu_n19836));
INVX1 exu_U5237(.A(se), .Y(exu_n19842));
INVX1 exu_U5238(.A(se), .Y(exu_n19848));
INVX1 exu_U5239(.A(se), .Y(exu_n19854));
INVX1 exu_U5240(.A(se), .Y(exu_n19860));
INVX1 exu_U5241(.A(se), .Y(exu_n19866));
INVX1 exu_U5242(.A(se), .Y(exu_n19872));
INVX1 exu_U5243(.A(se), .Y(exu_n19878));
OR2X1 exu_U5244(.A(ecl_save_e), .B(ecl_restore_e), .Y(ecl_n44));
INVX1 exu_U5245(.A(se), .Y(exu_n19884));
INVX1 exu_U5246(.A(se), .Y(exu_n19890));
INVX1 exu_U5247(.A(se), .Y(exu_n19896));
INVX1 exu_U5248(.A(se), .Y(exu_n19902));
AND2X1 exu_U5249(.A(exu_n3997), .B(exu_n9011), .Y(exu_n31676));
AND2X1 exu_U5250(.A(exu_n3993), .B(exu_n9006), .Y(exu_n31677));
AND2X1 exu_U5251(.A(exu_n3746), .B(exu_n8825), .Y(div_ecl_gencc_in_31));
INVX1 exu_U5252(.A(exu_n16198), .Y(exu_n16197));
AND2X1 exu_U5253(.A(exu_n4417), .B(exu_n9262), .Y(div_low32or_n2));
AND2X1 exu_U5254(.A(exu_n4422), .B(exu_n9267), .Y(div_low32or_n1));
INVX1 exu_U5255(.A(se), .Y(exu_n19908));
INVX1 exu_U5256(.A(se), .Y(exu_n19914));
INVX1 exu_U5257(.A(se), .Y(exu_n19950));
INVX1 exu_U5258(.A(se), .Y(exu_n19958));
INVX1 exu_U5259(.A(se), .Y(exu_n19966));
INVX1 exu_U5260(.A(se), .Y(exu_n19974));
INVX1 exu_U5261(.A(se), .Y(exu_n19982));
AND2X1 exu_U5262(.A(exu_n4149), .B(rml_cwp_swap_data[6]), .Y(rml_cwp_spill_next));
OR2X1 exu_U5263(.A(rml_cwp_swap_thr[3]), .B(rml_cwp_swap_thr[2]), .Y(rml_cwp_swap_tid[1]));
OR2X1 exu_U5264(.A(rml_cwp_swap_thr[3]), .B(rml_cwp_swap_thr[1]), .Y(rml_cwp_swap_tid[0]));
INVX1 exu_U5265(.A(se), .Y(exu_n18417));
AND2X1 exu_U5266(.A(exu_n4002), .B(exu_n9018), .Y(rml_cwp_cwp_output_mux_n8));
AND2X1 exu_U5267(.A(exu_n4003), .B(exu_n9019), .Y(rml_cwp_cwp_output_mux_n7));
AND2X1 exu_U5268(.A(exu_n4024), .B(exu_n9040), .Y(rml_cwp_cwp_output_mux_n74));
AND2X1 exu_U5269(.A(exu_n4025), .B(exu_n9041), .Y(rml_cwp_cwp_output_mux_n73));
AND2X1 exu_U5270(.A(exu_n4026), .B(exu_n9042), .Y(rml_cwp_cwp_output_mux_n80));
AND2X1 exu_U5271(.A(exu_n4027), .B(exu_n9043), .Y(rml_cwp_cwp_output_mux_n79));
AND2X1 exu_U5272(.A(exu_n4000), .B(exu_n9016), .Y(rml_cwp_cwp_output_mux_n2));
AND2X1 exu_U5273(.A(exu_n4001), .B(exu_n9017), .Y(rml_cwp_cwp_output_mux_n1));
INVX1 exu_U5274(.A(se), .Y(exu_n19990));
INVX1 exu_U5275(.A(se), .Y(exu_n20268));
INVX1 exu_U5276(.A(se), .Y(exu_n20277));
AND2X1 exu_U5277(.A(exu_n8664), .B(exu_n9673), .Y(ecl_alu_xcc_e[3]));
AND2X1 exu_U5278(.A(exu_n15426), .B(exu_n9650), .Y(ecl_alu_xcc_e[2]));
AND2X1 exu_U5279(.A(exu_n4969), .B(exu_n16155), .Y(ecl_adder_xcc[1]));
AND2X1 exu_U5280(.A(ecl_n135), .B(ecl_sel_sum_e), .Y(ecl_adder_xcc[0]));
AND2X1 exu_U5281(.A(exu_n8699), .B(exu_n9674), .Y(ecl_alu_icc_e[3]));
OR2X1 exu_U5282(.A(exu_n13499), .B(exu_n14816), .Y(alu_ecl_zlow_e));
AND2X1 exu_U5283(.A(exu_n4970), .B(ecl_sel_sum_e), .Y(ecl_adder_icc[1]));
AND2X1 exu_U5284(.A(ecl_n145), .B(exu_n16155), .Y(ecl_adder_icc[0]));
INVX1 exu_U5285(.A(se), .Y(exu_n20286));
INVX1 exu_U5286(.A(se), .Y(exu_n20295));
INVX1 exu_U5287(.A(se), .Y(exu_n20304));
INVX1 exu_U5288(.A(se), .Y(exu_n20313));
INVX1 exu_U5289(.A(se), .Y(exu_n20322));
INVX1 exu_U5290(.A(se), .Y(exu_n20331));
OR2X1 exu_U5291(.A(exu_n12126), .B(exu_n13542), .Y(rml_ecl_wstate_d[5]));
AND2X1 exu_U5292(.A(exu_n301), .B(exu_n5228), .Y(exu_n17944));
OR2X1 exu_U5293(.A(exu_n12127), .B(exu_n13543), .Y(rml_ecl_wstate_d[4]));
AND2X1 exu_U5294(.A(exu_n303), .B(exu_n5230), .Y(exu_n17950));
OR2X1 exu_U5295(.A(exu_n16374), .B(exu_n14761), .Y(ecl_writeback_sel_wstate_d));
OR2X1 exu_U5296(.A(exu_n12128), .B(exu_n13544), .Y(rml_ecl_wstate_d[3]));
AND2X1 exu_U5297(.A(exu_n305), .B(exu_n5232), .Y(exu_n17956));
INVX1 exu_U5298(.A(ifu_tlu_sraddr_d[3]), .Y(exu_n16373));
AND2X1 exu_U5299(.A(exu_n322), .B(exu_n5249), .Y(exu_n18020));
AND2X1 exu_U5300(.A(exu_n323), .B(exu_n5250), .Y(exu_n18019));
AND2X1 exu_U5301(.A(exu_n324), .B(exu_n5251), .Y(exu_n18026));
AND2X1 exu_U5302(.A(exu_n325), .B(exu_n5252), .Y(exu_n18025));
AND2X1 exu_U5303(.A(exu_n326), .B(exu_n5253), .Y(exu_n18032));
AND2X1 exu_U5304(.A(exu_n327), .B(exu_n5254), .Y(exu_n18031));
INVX1 exu_U5305(.A(se), .Y(exu_n20340));
INVX1 exu_U5306(.A(exu_n16009), .Y(exu_n16006));
INVX1 exu_U5307(.A(exu_n16009), .Y(exu_n16008));
INVX1 exu_U5308(.A(exu_n16009), .Y(exu_n16007));
AND2X1 exu_U5309(.A(exu_n928), .B(exu_n5689), .Y(exu_n20903));
AND2X1 exu_U5310(.A(exu_n929), .B(exu_n5690), .Y(exu_n20902));
AND2X1 exu_U5311(.A(exu_n930), .B(exu_n5691), .Y(exu_n20909));
AND2X1 exu_U5312(.A(exu_n931), .B(exu_n5692), .Y(exu_n20908));
AND2X1 exu_U5313(.A(exu_n934), .B(exu_n5695), .Y(exu_n20921));
AND2X1 exu_U5314(.A(exu_n935), .B(exu_n5696), .Y(exu_n20920));
AND2X1 exu_U5315(.A(exu_n936), .B(exu_n5697), .Y(exu_n20927));
AND2X1 exu_U5316(.A(exu_n937), .B(exu_n5698), .Y(exu_n20926));
AND2X1 exu_U5317(.A(exu_n938), .B(exu_n5699), .Y(exu_n20933));
AND2X1 exu_U5318(.A(exu_n939), .B(exu_n5700), .Y(exu_n20932));
AND2X1 exu_U5319(.A(exu_n940), .B(exu_n5701), .Y(exu_n20939));
AND2X1 exu_U5320(.A(exu_n941), .B(exu_n5702), .Y(exu_n20938));
AND2X1 exu_U5321(.A(exu_n942), .B(exu_n5703), .Y(exu_n20945));
AND2X1 exu_U5322(.A(exu_n943), .B(exu_n5704), .Y(exu_n20944));
AND2X1 exu_U5323(.A(exu_n944), .B(exu_n5705), .Y(exu_n20951));
AND2X1 exu_U5324(.A(exu_n945), .B(exu_n5706), .Y(exu_n20950));
AND2X1 exu_U5325(.A(exu_n946), .B(exu_n5707), .Y(exu_n20957));
AND2X1 exu_U5326(.A(exu_n947), .B(exu_n5708), .Y(exu_n20956));
AND2X1 exu_U5327(.A(exu_n948), .B(exu_n5709), .Y(exu_n20963));
AND2X1 exu_U5328(.A(exu_n949), .B(exu_n5710), .Y(exu_n20962));
AND2X1 exu_U5329(.A(exu_n950), .B(exu_n5711), .Y(exu_n20969));
AND2X1 exu_U5330(.A(exu_n951), .B(exu_n5712), .Y(exu_n20968));
AND2X1 exu_U5331(.A(exu_n952), .B(exu_n5713), .Y(exu_n20975));
AND2X1 exu_U5332(.A(exu_n953), .B(exu_n5714), .Y(exu_n20974));
AND2X1 exu_U5333(.A(exu_n956), .B(exu_n5717), .Y(exu_n20987));
AND2X1 exu_U5334(.A(exu_n957), .B(exu_n5718), .Y(exu_n20986));
AND2X1 exu_U5335(.A(exu_n958), .B(exu_n5719), .Y(exu_n20993));
AND2X1 exu_U5336(.A(exu_n959), .B(exu_n5720), .Y(exu_n20992));
AND2X1 exu_U5337(.A(exu_n960), .B(exu_n5721), .Y(exu_n20999));
AND2X1 exu_U5338(.A(exu_n961), .B(exu_n5722), .Y(exu_n20998));
AND2X1 exu_U5339(.A(exu_n962), .B(exu_n5723), .Y(exu_n21005));
AND2X1 exu_U5340(.A(exu_n963), .B(exu_n5724), .Y(exu_n21004));
AND2X1 exu_U5341(.A(exu_n964), .B(exu_n5725), .Y(exu_n21011));
AND2X1 exu_U5342(.A(exu_n965), .B(exu_n5726), .Y(exu_n21010));
AND2X1 exu_U5343(.A(exu_n966), .B(exu_n5727), .Y(exu_n21017));
AND2X1 exu_U5344(.A(exu_n967), .B(exu_n5728), .Y(exu_n21016));
AND2X1 exu_U5345(.A(exu_n968), .B(exu_n5729), .Y(exu_n21023));
AND2X1 exu_U5346(.A(exu_n969), .B(exu_n5730), .Y(exu_n21022));
AND2X1 exu_U5347(.A(exu_n970), .B(exu_n5731), .Y(exu_n21029));
AND2X1 exu_U5348(.A(exu_n971), .B(exu_n5732), .Y(exu_n21028));
AND2X1 exu_U5349(.A(exu_n972), .B(exu_n5733), .Y(exu_n21035));
AND2X1 exu_U5350(.A(exu_n973), .B(exu_n5734), .Y(exu_n21034));
AND2X1 exu_U5351(.A(exu_n974), .B(exu_n5735), .Y(exu_n21041));
AND2X1 exu_U5352(.A(exu_n975), .B(exu_n5736), .Y(exu_n21040));
AND2X1 exu_U5353(.A(exu_n914), .B(exu_n5675), .Y(exu_n20861));
AND2X1 exu_U5354(.A(exu_n915), .B(exu_n5676), .Y(exu_n20860));
AND2X1 exu_U5355(.A(exu_n916), .B(exu_n5677), .Y(exu_n20867));
AND2X1 exu_U5356(.A(exu_n917), .B(exu_n5678), .Y(exu_n20866));
AND2X1 exu_U5357(.A(exu_n918), .B(exu_n5679), .Y(exu_n20873));
AND2X1 exu_U5358(.A(exu_n919), .B(exu_n5680), .Y(exu_n20872));
INVX1 exu_U5359(.A(exu_n16013), .Y(exu_n16010));
AND2X1 exu_U5360(.A(exu_n920), .B(exu_n5681), .Y(exu_n20879));
AND2X1 exu_U5361(.A(exu_n921), .B(exu_n5682), .Y(exu_n20878));
AND2X1 exu_U5362(.A(exu_n922), .B(exu_n5683), .Y(exu_n20885));
AND2X1 exu_U5363(.A(exu_n923), .B(exu_n5684), .Y(exu_n20884));
AND2X1 exu_U5364(.A(exu_n924), .B(exu_n5685), .Y(exu_n20891));
AND2X1 exu_U5365(.A(exu_n925), .B(exu_n5686), .Y(exu_n20890));
AND2X1 exu_U5366(.A(exu_n926), .B(exu_n5687), .Y(exu_n20897));
AND2X1 exu_U5367(.A(exu_n927), .B(exu_n5688), .Y(exu_n20896));
AND2X1 exu_U5368(.A(exu_n932), .B(exu_n5693), .Y(exu_n20915));
AND2X1 exu_U5369(.A(exu_n933), .B(exu_n5694), .Y(exu_n20914));
AND2X1 exu_U5370(.A(exu_n954), .B(exu_n5715), .Y(exu_n20981));
AND2X1 exu_U5371(.A(exu_n955), .B(exu_n5716), .Y(exu_n20980));
INVX1 exu_U5372(.A(exu_n16013), .Y(exu_n16012));
AND2X1 exu_U5373(.A(exu_n976), .B(exu_n5737), .Y(exu_n21047));
AND2X1 exu_U5374(.A(exu_n977), .B(exu_n5738), .Y(exu_n21046));
INVX1 exu_U5375(.A(exu_n16013), .Y(exu_n16011));
AND2X1 exu_U5376(.A(exu_n992), .B(exu_n5753), .Y(exu_n21095));
AND2X1 exu_U5377(.A(exu_n993), .B(exu_n5754), .Y(exu_n21094));
AND2X1 exu_U5378(.A(exu_n994), .B(exu_n5755), .Y(exu_n21101));
AND2X1 exu_U5379(.A(exu_n995), .B(exu_n5756), .Y(exu_n21100));
AND2X1 exu_U5380(.A(exu_n998), .B(exu_n5759), .Y(exu_n21113));
AND2X1 exu_U5381(.A(exu_n999), .B(exu_n5760), .Y(exu_n21112));
AND2X1 exu_U5382(.A(exu_n1000), .B(exu_n5761), .Y(exu_n21119));
AND2X1 exu_U5383(.A(exu_n1001), .B(exu_n5762), .Y(exu_n21118));
AND2X1 exu_U5384(.A(exu_n1002), .B(exu_n5763), .Y(exu_n21125));
AND2X1 exu_U5385(.A(exu_n1003), .B(exu_n5764), .Y(exu_n21124));
AND2X1 exu_U5386(.A(exu_n1004), .B(exu_n5765), .Y(exu_n21131));
AND2X1 exu_U5387(.A(exu_n1005), .B(exu_n5766), .Y(exu_n21130));
AND2X1 exu_U5388(.A(exu_n1006), .B(exu_n5767), .Y(exu_n21137));
AND2X1 exu_U5389(.A(exu_n1007), .B(exu_n5768), .Y(exu_n21136));
AND2X1 exu_U5390(.A(exu_n1008), .B(exu_n5769), .Y(exu_n21143));
AND2X1 exu_U5391(.A(exu_n1009), .B(exu_n5770), .Y(exu_n21142));
AND2X1 exu_U5392(.A(exu_n1010), .B(exu_n5771), .Y(exu_n21149));
AND2X1 exu_U5393(.A(exu_n1011), .B(exu_n5772), .Y(exu_n21148));
AND2X1 exu_U5394(.A(exu_n1012), .B(exu_n5773), .Y(exu_n21155));
AND2X1 exu_U5395(.A(exu_n1013), .B(exu_n5774), .Y(exu_n21154));
AND2X1 exu_U5396(.A(exu_n1014), .B(exu_n5775), .Y(exu_n21161));
AND2X1 exu_U5397(.A(exu_n1015), .B(exu_n5776), .Y(exu_n21160));
AND2X1 exu_U5398(.A(exu_n1016), .B(exu_n5777), .Y(exu_n21167));
AND2X1 exu_U5399(.A(exu_n1017), .B(exu_n5778), .Y(exu_n21166));
AND2X1 exu_U5400(.A(exu_n1020), .B(exu_n5781), .Y(exu_n21179));
AND2X1 exu_U5401(.A(exu_n1021), .B(exu_n5782), .Y(exu_n21178));
AND2X1 exu_U5402(.A(exu_n1022), .B(exu_n5783), .Y(exu_n21185));
AND2X1 exu_U5403(.A(exu_n1023), .B(exu_n5784), .Y(exu_n21184));
AND2X1 exu_U5404(.A(exu_n1024), .B(exu_n5785), .Y(exu_n21191));
AND2X1 exu_U5405(.A(exu_n1025), .B(exu_n5786), .Y(exu_n21190));
AND2X1 exu_U5406(.A(exu_n1026), .B(exu_n5787), .Y(exu_n21197));
AND2X1 exu_U5407(.A(exu_n1027), .B(exu_n5788), .Y(exu_n21196));
AND2X1 exu_U5408(.A(exu_n1028), .B(exu_n5789), .Y(exu_n21203));
AND2X1 exu_U5409(.A(exu_n1029), .B(exu_n5790), .Y(exu_n21202));
AND2X1 exu_U5410(.A(exu_n1030), .B(exu_n5791), .Y(exu_n21209));
AND2X1 exu_U5411(.A(exu_n1031), .B(exu_n5792), .Y(exu_n21208));
AND2X1 exu_U5412(.A(exu_n1032), .B(exu_n5793), .Y(exu_n21215));
AND2X1 exu_U5413(.A(exu_n1033), .B(exu_n5794), .Y(exu_n21214));
AND2X1 exu_U5414(.A(exu_n1034), .B(exu_n5795), .Y(exu_n21221));
AND2X1 exu_U5415(.A(exu_n1035), .B(exu_n5796), .Y(exu_n21220));
AND2X1 exu_U5416(.A(exu_n1036), .B(exu_n5797), .Y(exu_n21227));
AND2X1 exu_U5417(.A(exu_n1037), .B(exu_n5798), .Y(exu_n21226));
AND2X1 exu_U5418(.A(exu_n1038), .B(exu_n5799), .Y(exu_n21233));
AND2X1 exu_U5419(.A(exu_n1039), .B(exu_n5800), .Y(exu_n21232));
AND2X1 exu_U5420(.A(exu_n978), .B(exu_n5739), .Y(exu_n21053));
AND2X1 exu_U5421(.A(exu_n979), .B(exu_n5740), .Y(exu_n21052));
AND2X1 exu_U5422(.A(exu_n980), .B(exu_n5741), .Y(exu_n21059));
AND2X1 exu_U5423(.A(exu_n981), .B(exu_n5742), .Y(exu_n21058));
AND2X1 exu_U5424(.A(exu_n982), .B(exu_n5743), .Y(exu_n21065));
AND2X1 exu_U5425(.A(exu_n983), .B(exu_n5744), .Y(exu_n21064));
INVX1 exu_U5426(.A(exu_n16017), .Y(exu_n16014));
AND2X1 exu_U5427(.A(exu_n984), .B(exu_n5745), .Y(exu_n21071));
AND2X1 exu_U5428(.A(exu_n985), .B(exu_n5746), .Y(exu_n21070));
AND2X1 exu_U5429(.A(exu_n986), .B(exu_n5747), .Y(exu_n21077));
AND2X1 exu_U5430(.A(exu_n987), .B(exu_n5748), .Y(exu_n21076));
AND2X1 exu_U5431(.A(exu_n988), .B(exu_n5749), .Y(exu_n21083));
AND2X1 exu_U5432(.A(exu_n989), .B(exu_n5750), .Y(exu_n21082));
AND2X1 exu_U5433(.A(exu_n990), .B(exu_n5751), .Y(exu_n21089));
AND2X1 exu_U5434(.A(exu_n991), .B(exu_n5752), .Y(exu_n21088));
AND2X1 exu_U5435(.A(exu_n996), .B(exu_n5757), .Y(exu_n21107));
AND2X1 exu_U5436(.A(exu_n997), .B(exu_n5758), .Y(exu_n21106));
AND2X1 exu_U5437(.A(exu_n1018), .B(exu_n5779), .Y(exu_n21173));
AND2X1 exu_U5438(.A(exu_n1019), .B(exu_n5780), .Y(exu_n21172));
INVX1 exu_U5439(.A(exu_n16017), .Y(exu_n16016));
AND2X1 exu_U5440(.A(exu_n1040), .B(exu_n5801), .Y(exu_n21239));
AND2X1 exu_U5441(.A(exu_n1041), .B(exu_n5802), .Y(exu_n21238));
INVX1 exu_U5442(.A(exu_n16017), .Y(exu_n16015));
AND2X1 exu_U5443(.A(exu_n1056), .B(exu_n5817), .Y(exu_n21287));
AND2X1 exu_U5444(.A(exu_n1057), .B(exu_n5818), .Y(exu_n21286));
AND2X1 exu_U5445(.A(exu_n1058), .B(exu_n5819), .Y(exu_n21293));
AND2X1 exu_U5446(.A(exu_n1059), .B(exu_n5820), .Y(exu_n21292));
AND2X1 exu_U5447(.A(exu_n1062), .B(exu_n5823), .Y(exu_n21305));
AND2X1 exu_U5448(.A(exu_n1063), .B(exu_n5824), .Y(exu_n21304));
AND2X1 exu_U5449(.A(exu_n1064), .B(exu_n5825), .Y(exu_n21311));
AND2X1 exu_U5450(.A(exu_n1065), .B(exu_n5826), .Y(exu_n21310));
AND2X1 exu_U5451(.A(exu_n1066), .B(exu_n5827), .Y(exu_n21317));
AND2X1 exu_U5452(.A(exu_n1067), .B(exu_n5828), .Y(exu_n21316));
AND2X1 exu_U5453(.A(exu_n1068), .B(exu_n5829), .Y(exu_n21323));
AND2X1 exu_U5454(.A(exu_n1069), .B(exu_n5830), .Y(exu_n21322));
AND2X1 exu_U5455(.A(exu_n1070), .B(exu_n5831), .Y(exu_n21329));
AND2X1 exu_U5456(.A(exu_n1071), .B(exu_n5832), .Y(exu_n21328));
AND2X1 exu_U5457(.A(exu_n1072), .B(exu_n5833), .Y(exu_n21335));
AND2X1 exu_U5458(.A(exu_n1073), .B(exu_n5834), .Y(exu_n21334));
AND2X1 exu_U5459(.A(exu_n1074), .B(exu_n5835), .Y(exu_n21341));
AND2X1 exu_U5460(.A(exu_n1075), .B(exu_n5836), .Y(exu_n21340));
AND2X1 exu_U5461(.A(exu_n1076), .B(exu_n5837), .Y(exu_n21347));
AND2X1 exu_U5462(.A(exu_n1077), .B(exu_n5838), .Y(exu_n21346));
AND2X1 exu_U5463(.A(exu_n1078), .B(exu_n5839), .Y(exu_n21353));
AND2X1 exu_U5464(.A(exu_n1079), .B(exu_n5840), .Y(exu_n21352));
AND2X1 exu_U5465(.A(exu_n1080), .B(exu_n5841), .Y(exu_n21359));
AND2X1 exu_U5466(.A(exu_n1081), .B(exu_n5842), .Y(exu_n21358));
AND2X1 exu_U5467(.A(exu_n1084), .B(exu_n5845), .Y(exu_n21371));
AND2X1 exu_U5468(.A(exu_n1085), .B(exu_n5846), .Y(exu_n21370));
AND2X1 exu_U5469(.A(exu_n1086), .B(exu_n5847), .Y(exu_n21377));
AND2X1 exu_U5470(.A(exu_n1087), .B(exu_n5848), .Y(exu_n21376));
AND2X1 exu_U5471(.A(exu_n1088), .B(exu_n5849), .Y(exu_n21383));
AND2X1 exu_U5472(.A(exu_n1089), .B(exu_n5850), .Y(exu_n21382));
AND2X1 exu_U5473(.A(exu_n1090), .B(exu_n5851), .Y(exu_n21389));
AND2X1 exu_U5474(.A(exu_n1091), .B(exu_n5852), .Y(exu_n21388));
AND2X1 exu_U5475(.A(exu_n1092), .B(exu_n5853), .Y(exu_n21395));
AND2X1 exu_U5476(.A(exu_n1093), .B(exu_n5854), .Y(exu_n21394));
AND2X1 exu_U5477(.A(exu_n1094), .B(exu_n5855), .Y(exu_n21401));
AND2X1 exu_U5478(.A(exu_n1095), .B(exu_n5856), .Y(exu_n21400));
AND2X1 exu_U5479(.A(exu_n1096), .B(exu_n5857), .Y(exu_n21407));
AND2X1 exu_U5480(.A(exu_n1097), .B(exu_n5858), .Y(exu_n21406));
AND2X1 exu_U5481(.A(exu_n1098), .B(exu_n5859), .Y(exu_n21413));
AND2X1 exu_U5482(.A(exu_n1099), .B(exu_n5860), .Y(exu_n21412));
AND2X1 exu_U5483(.A(exu_n1100), .B(exu_n5861), .Y(exu_n21419));
AND2X1 exu_U5484(.A(exu_n1101), .B(exu_n5862), .Y(exu_n21418));
AND2X1 exu_U5485(.A(exu_n1102), .B(exu_n5863), .Y(exu_n21425));
AND2X1 exu_U5486(.A(exu_n1103), .B(exu_n5864), .Y(exu_n21424));
AND2X1 exu_U5487(.A(exu_n1042), .B(exu_n5803), .Y(exu_n21245));
AND2X1 exu_U5488(.A(exu_n1043), .B(exu_n5804), .Y(exu_n21244));
AND2X1 exu_U5489(.A(exu_n1044), .B(exu_n5805), .Y(exu_n21251));
AND2X1 exu_U5490(.A(exu_n1045), .B(exu_n5806), .Y(exu_n21250));
AND2X1 exu_U5491(.A(exu_n1046), .B(exu_n5807), .Y(exu_n21257));
AND2X1 exu_U5492(.A(exu_n1047), .B(exu_n5808), .Y(exu_n21256));
INVX1 exu_U5493(.A(exu_n16021), .Y(exu_n16018));
AND2X1 exu_U5494(.A(exu_n1048), .B(exu_n5809), .Y(exu_n21263));
AND2X1 exu_U5495(.A(exu_n1049), .B(exu_n5810), .Y(exu_n21262));
AND2X1 exu_U5496(.A(exu_n1050), .B(exu_n5811), .Y(exu_n21269));
AND2X1 exu_U5497(.A(exu_n1051), .B(exu_n5812), .Y(exu_n21268));
AND2X1 exu_U5498(.A(exu_n1052), .B(exu_n5813), .Y(exu_n21275));
AND2X1 exu_U5499(.A(exu_n1053), .B(exu_n5814), .Y(exu_n21274));
AND2X1 exu_U5500(.A(exu_n1054), .B(exu_n5815), .Y(exu_n21281));
AND2X1 exu_U5501(.A(exu_n1055), .B(exu_n5816), .Y(exu_n21280));
AND2X1 exu_U5502(.A(exu_n1060), .B(exu_n5821), .Y(exu_n21299));
AND2X1 exu_U5503(.A(exu_n1061), .B(exu_n5822), .Y(exu_n21298));
AND2X1 exu_U5504(.A(exu_n1082), .B(exu_n5843), .Y(exu_n21365));
AND2X1 exu_U5505(.A(exu_n1083), .B(exu_n5844), .Y(exu_n21364));
INVX1 exu_U5506(.A(exu_n16021), .Y(exu_n16020));
AND2X1 exu_U5507(.A(exu_n1104), .B(exu_n5865), .Y(exu_n21431));
AND2X1 exu_U5508(.A(exu_n1105), .B(exu_n5866), .Y(exu_n21430));
INVX1 exu_U5509(.A(exu_n16021), .Y(exu_n16019));
AND2X1 exu_U5510(.A(exu_n1120), .B(exu_n5881), .Y(exu_n21479));
AND2X1 exu_U5511(.A(exu_n1121), .B(exu_n5882), .Y(exu_n21478));
AND2X1 exu_U5512(.A(exu_n1122), .B(exu_n5883), .Y(exu_n21485));
AND2X1 exu_U5513(.A(exu_n1123), .B(exu_n5884), .Y(exu_n21484));
AND2X1 exu_U5514(.A(exu_n1126), .B(exu_n5887), .Y(exu_n21497));
AND2X1 exu_U5515(.A(exu_n1127), .B(exu_n5888), .Y(exu_n21496));
AND2X1 exu_U5516(.A(exu_n1128), .B(exu_n5889), .Y(exu_n21503));
AND2X1 exu_U5517(.A(exu_n1129), .B(exu_n5890), .Y(exu_n21502));
AND2X1 exu_U5518(.A(exu_n1130), .B(exu_n5891), .Y(exu_n21509));
AND2X1 exu_U5519(.A(exu_n1131), .B(exu_n5892), .Y(exu_n21508));
AND2X1 exu_U5520(.A(exu_n1132), .B(exu_n5893), .Y(exu_n21515));
AND2X1 exu_U5521(.A(exu_n1133), .B(exu_n5894), .Y(exu_n21514));
AND2X1 exu_U5522(.A(exu_n1134), .B(exu_n5895), .Y(exu_n21521));
AND2X1 exu_U5523(.A(exu_n1135), .B(exu_n5896), .Y(exu_n21520));
AND2X1 exu_U5524(.A(exu_n1136), .B(exu_n5897), .Y(exu_n21527));
AND2X1 exu_U5525(.A(exu_n1137), .B(exu_n5898), .Y(exu_n21526));
AND2X1 exu_U5526(.A(exu_n1138), .B(exu_n5899), .Y(exu_n21533));
AND2X1 exu_U5527(.A(exu_n1139), .B(exu_n5900), .Y(exu_n21532));
AND2X1 exu_U5528(.A(exu_n1140), .B(exu_n5901), .Y(exu_n21539));
AND2X1 exu_U5529(.A(exu_n1141), .B(exu_n5902), .Y(exu_n21538));
AND2X1 exu_U5530(.A(exu_n1142), .B(exu_n5903), .Y(exu_n21545));
AND2X1 exu_U5531(.A(exu_n1143), .B(exu_n5904), .Y(exu_n21544));
AND2X1 exu_U5532(.A(exu_n1144), .B(exu_n5905), .Y(exu_n21551));
AND2X1 exu_U5533(.A(exu_n1145), .B(exu_n5906), .Y(exu_n21550));
AND2X1 exu_U5534(.A(exu_n1148), .B(exu_n5909), .Y(exu_n21563));
AND2X1 exu_U5535(.A(exu_n1149), .B(exu_n5910), .Y(exu_n21562));
AND2X1 exu_U5536(.A(exu_n1150), .B(exu_n5911), .Y(exu_n21569));
AND2X1 exu_U5537(.A(exu_n1151), .B(exu_n5912), .Y(exu_n21568));
AND2X1 exu_U5538(.A(exu_n1152), .B(exu_n5913), .Y(exu_n21575));
AND2X1 exu_U5539(.A(exu_n1153), .B(exu_n5914), .Y(exu_n21574));
AND2X1 exu_U5540(.A(exu_n1154), .B(exu_n5915), .Y(exu_n21581));
AND2X1 exu_U5541(.A(exu_n1155), .B(exu_n5916), .Y(exu_n21580));
AND2X1 exu_U5542(.A(exu_n1156), .B(exu_n5917), .Y(exu_n21587));
AND2X1 exu_U5543(.A(exu_n1157), .B(exu_n5918), .Y(exu_n21586));
AND2X1 exu_U5544(.A(exu_n1158), .B(exu_n5919), .Y(exu_n21593));
AND2X1 exu_U5545(.A(exu_n1159), .B(exu_n5920), .Y(exu_n21592));
AND2X1 exu_U5546(.A(exu_n1160), .B(exu_n5921), .Y(exu_n21599));
AND2X1 exu_U5547(.A(exu_n1161), .B(exu_n5922), .Y(exu_n21598));
AND2X1 exu_U5548(.A(exu_n1162), .B(exu_n5923), .Y(exu_n21605));
AND2X1 exu_U5549(.A(exu_n1163), .B(exu_n5924), .Y(exu_n21604));
AND2X1 exu_U5550(.A(exu_n1164), .B(exu_n5925), .Y(exu_n21611));
AND2X1 exu_U5551(.A(exu_n1165), .B(exu_n5926), .Y(exu_n21610));
AND2X1 exu_U5552(.A(exu_n1166), .B(exu_n5927), .Y(exu_n21617));
AND2X1 exu_U5553(.A(exu_n1167), .B(exu_n5928), .Y(exu_n21616));
AND2X1 exu_U5554(.A(exu_n1106), .B(exu_n5867), .Y(exu_n21437));
AND2X1 exu_U5555(.A(exu_n1107), .B(exu_n5868), .Y(exu_n21436));
AND2X1 exu_U5556(.A(exu_n1108), .B(exu_n5869), .Y(exu_n21443));
AND2X1 exu_U5557(.A(exu_n1109), .B(exu_n5870), .Y(exu_n21442));
AND2X1 exu_U5558(.A(exu_n1110), .B(exu_n5871), .Y(exu_n21449));
AND2X1 exu_U5559(.A(exu_n1111), .B(exu_n5872), .Y(exu_n21448));
INVX1 exu_U5560(.A(exu_n16025), .Y(exu_n16022));
AND2X1 exu_U5561(.A(exu_n1112), .B(exu_n5873), .Y(exu_n21455));
AND2X1 exu_U5562(.A(exu_n1113), .B(exu_n5874), .Y(exu_n21454));
AND2X1 exu_U5563(.A(exu_n1114), .B(exu_n5875), .Y(exu_n21461));
AND2X1 exu_U5564(.A(exu_n1115), .B(exu_n5876), .Y(exu_n21460));
AND2X1 exu_U5565(.A(exu_n1116), .B(exu_n5877), .Y(exu_n21467));
AND2X1 exu_U5566(.A(exu_n1117), .B(exu_n5878), .Y(exu_n21466));
AND2X1 exu_U5567(.A(exu_n1118), .B(exu_n5879), .Y(exu_n21473));
AND2X1 exu_U5568(.A(exu_n1119), .B(exu_n5880), .Y(exu_n21472));
AND2X1 exu_U5569(.A(exu_n1124), .B(exu_n5885), .Y(exu_n21491));
AND2X1 exu_U5570(.A(exu_n1125), .B(exu_n5886), .Y(exu_n21490));
AND2X1 exu_U5571(.A(exu_n1146), .B(exu_n5907), .Y(exu_n21557));
AND2X1 exu_U5572(.A(exu_n1147), .B(exu_n5908), .Y(exu_n21556));
INVX1 exu_U5573(.A(exu_n16025), .Y(exu_n16024));
AND2X1 exu_U5574(.A(exu_n1168), .B(exu_n5929), .Y(exu_n21623));
AND2X1 exu_U5575(.A(exu_n1169), .B(exu_n5930), .Y(exu_n21622));
INVX1 exu_U5576(.A(exu_n16025), .Y(exu_n16023));
OR2X1 exu_U5577(.A(exu_n12185), .B(exu_n13597), .Y(div_byp_yreg_e[31]));
AND2X1 exu_U5578(.A(exu_n865), .B(exu_n5626), .Y(exu_n20710));
AND2X1 exu_U5579(.A(exu_n4792), .B(exu_n9579), .Y(bypass_ifu_exu_sr_mux_n236));
OR2X1 exu_U5580(.A(exu_n12186), .B(exu_n13598), .Y(div_byp_yreg_e[30]));
AND2X1 exu_U5581(.A(exu_n867), .B(exu_n5628), .Y(exu_n20716));
AND2X1 exu_U5582(.A(exu_n4793), .B(exu_n9580), .Y(bypass_ifu_exu_sr_mux_n242));
OR2X1 exu_U5583(.A(exu_n12188), .B(exu_n13600), .Y(div_byp_yreg_e[29]));
AND2X1 exu_U5584(.A(exu_n871), .B(exu_n5632), .Y(exu_n20728));
AND2X1 exu_U5585(.A(exu_n4796), .B(exu_n9583), .Y(bypass_ifu_exu_sr_mux_n254));
OR2X1 exu_U5586(.A(exu_n12189), .B(exu_n13601), .Y(div_byp_yreg_e[28]));
AND2X1 exu_U5587(.A(exu_n873), .B(exu_n5634), .Y(exu_n20734));
AND2X1 exu_U5588(.A(exu_n4797), .B(exu_n9584), .Y(bypass_ifu_exu_sr_mux_n260));
OR2X1 exu_U5589(.A(exu_n12190), .B(exu_n13602), .Y(div_byp_yreg_e[27]));
AND2X1 exu_U5590(.A(exu_n875), .B(exu_n5636), .Y(exu_n20740));
AND2X1 exu_U5591(.A(exu_n4798), .B(exu_n9585), .Y(bypass_ifu_exu_sr_mux_n266));
OR2X1 exu_U5592(.A(exu_n12191), .B(exu_n13603), .Y(div_byp_yreg_e[26]));
AND2X1 exu_U5593(.A(exu_n877), .B(exu_n5638), .Y(exu_n20746));
AND2X1 exu_U5594(.A(exu_n4799), .B(exu_n9586), .Y(bypass_ifu_exu_sr_mux_n272));
OR2X1 exu_U5595(.A(exu_n12192), .B(exu_n13604), .Y(div_byp_yreg_e[25]));
AND2X1 exu_U5596(.A(exu_n879), .B(exu_n5640), .Y(exu_n20752));
AND2X1 exu_U5597(.A(exu_n4800), .B(exu_n9587), .Y(bypass_ifu_exu_sr_mux_n278));
OR2X1 exu_U5598(.A(exu_n12193), .B(exu_n13605), .Y(div_byp_yreg_e[24]));
AND2X1 exu_U5599(.A(exu_n881), .B(exu_n5642), .Y(exu_n20758));
AND2X1 exu_U5600(.A(exu_n4801), .B(exu_n9588), .Y(bypass_ifu_exu_sr_mux_n284));
OR2X1 exu_U5601(.A(exu_n12194), .B(exu_n13606), .Y(div_byp_yreg_e[23]));
AND2X1 exu_U5602(.A(exu_n883), .B(exu_n5644), .Y(exu_n20764));
AND2X1 exu_U5603(.A(exu_n4802), .B(exu_n9589), .Y(bypass_ifu_exu_sr_mux_n290));
OR2X1 exu_U5604(.A(exu_n12195), .B(exu_n13607), .Y(div_byp_yreg_e[22]));
AND2X1 exu_U5605(.A(exu_n885), .B(exu_n5646), .Y(exu_n20770));
AND2X1 exu_U5606(.A(exu_n4803), .B(exu_n9590), .Y(bypass_ifu_exu_sr_mux_n296));
OR2X1 exu_U5607(.A(exu_n12196), .B(exu_n13608), .Y(div_byp_yreg_e[21]));
AND2X1 exu_U5608(.A(exu_n887), .B(exu_n5648), .Y(exu_n20776));
AND2X1 exu_U5609(.A(exu_n4804), .B(exu_n9591), .Y(bypass_ifu_exu_sr_mux_n302));
OR2X1 exu_U5610(.A(exu_n12197), .B(exu_n13609), .Y(div_byp_yreg_e[20]));
AND2X1 exu_U5611(.A(exu_n889), .B(exu_n5650), .Y(exu_n20782));
AND2X1 exu_U5612(.A(exu_n4805), .B(exu_n9592), .Y(bypass_ifu_exu_sr_mux_n308));
OR2X1 exu_U5613(.A(exu_n12199), .B(exu_n13611), .Y(div_byp_yreg_e[19]));
AND2X1 exu_U5614(.A(exu_n893), .B(exu_n5654), .Y(exu_n20794));
AND2X1 exu_U5615(.A(exu_n4808), .B(exu_n9595), .Y(bypass_ifu_exu_sr_mux_n320));
OR2X1 exu_U5616(.A(exu_n12200), .B(exu_n13612), .Y(div_byp_yreg_e[18]));
AND2X1 exu_U5617(.A(exu_n895), .B(exu_n5656), .Y(exu_n20800));
AND2X1 exu_U5618(.A(exu_n4809), .B(exu_n9596), .Y(bypass_ifu_exu_sr_mux_n326));
OR2X1 exu_U5619(.A(exu_n12201), .B(exu_n13613), .Y(div_byp_yreg_e[17]));
AND2X1 exu_U5620(.A(exu_n897), .B(exu_n5658), .Y(exu_n20806));
AND2X1 exu_U5621(.A(exu_n4810), .B(exu_n9597), .Y(bypass_ifu_exu_sr_mux_n332));
OR2X1 exu_U5622(.A(exu_n12202), .B(exu_n13614), .Y(div_byp_yreg_e[16]));
AND2X1 exu_U5623(.A(exu_n899), .B(exu_n5660), .Y(exu_n20812));
AND2X1 exu_U5624(.A(exu_n4811), .B(exu_n9598), .Y(bypass_ifu_exu_sr_mux_n338));
OR2X1 exu_U5625(.A(exu_n12203), .B(exu_n13615), .Y(div_byp_yreg_e[15]));
AND2X1 exu_U5626(.A(exu_n901), .B(exu_n5662), .Y(exu_n20818));
AND2X1 exu_U5627(.A(exu_n4812), .B(exu_n9599), .Y(bypass_ifu_exu_sr_mux_n344));
OR2X1 exu_U5628(.A(exu_n12204), .B(exu_n13616), .Y(div_byp_yreg_e[14]));
AND2X1 exu_U5629(.A(exu_n903), .B(exu_n5664), .Y(exu_n20824));
AND2X1 exu_U5630(.A(exu_n4813), .B(exu_n9600), .Y(bypass_ifu_exu_sr_mux_n350));
OR2X1 exu_U5631(.A(exu_n12205), .B(exu_n13617), .Y(div_byp_yreg_e[13]));
AND2X1 exu_U5632(.A(exu_n905), .B(exu_n5666), .Y(exu_n20830));
AND2X1 exu_U5633(.A(exu_n4814), .B(exu_n9601), .Y(bypass_ifu_exu_sr_mux_n356));
OR2X1 exu_U5634(.A(exu_n12206), .B(exu_n13618), .Y(div_byp_yreg_e[12]));
AND2X1 exu_U5635(.A(exu_n907), .B(exu_n5668), .Y(exu_n20836));
AND2X1 exu_U5636(.A(exu_n4815), .B(exu_n9602), .Y(bypass_ifu_exu_sr_mux_n362));
OR2X1 exu_U5637(.A(exu_n12207), .B(exu_n13619), .Y(div_byp_yreg_e[11]));
AND2X1 exu_U5638(.A(exu_n909), .B(exu_n5670), .Y(exu_n20842));
AND2X1 exu_U5639(.A(exu_n4816), .B(exu_n9603), .Y(bypass_ifu_exu_sr_mux_n368));
OR2X1 exu_U5640(.A(exu_n12208), .B(exu_n13620), .Y(div_byp_yreg_e[10]));
AND2X1 exu_U5641(.A(exu_n911), .B(exu_n5672), .Y(exu_n20848));
AND2X1 exu_U5642(.A(exu_n4817), .B(exu_n9604), .Y(bypass_ifu_exu_sr_mux_n374));
OR2X1 exu_U5643(.A(exu_n12178), .B(exu_n13590), .Y(div_byp_yreg_e[9]));
AND2X1 exu_U5644(.A(exu_n851), .B(exu_n5612), .Y(exu_n20668));
AND2X1 exu_U5645(.A(exu_n4748), .B(exu_n9567), .Y(bypass_ifu_exu_sr_mux_n2));
OR2X1 exu_U5646(.A(exu_n12179), .B(exu_n13591), .Y(div_byp_yreg_e[8]));
AND2X1 exu_U5647(.A(exu_n853), .B(exu_n5614), .Y(exu_n20674));
AND2X1 exu_U5648(.A(exu_n4749), .B(exu_n9568), .Y(bypass_ifu_exu_sr_mux_n8));
AND2X1 exu_U5649(.A(exu_n4750), .B(exu_n9569), .Y(bypass_ifu_exu_sr_mux_n14));
AND2X1 exu_U5650(.A(exu_n4751), .B(exu_n9570), .Y(bypass_ifu_exu_sr_mux_n13));
INVX1 exu_U5651(.A(exu_n16032), .Y(exu_n16026));
AND2X1 exu_U5652(.A(exu_n4752), .B(exu_n9571), .Y(bypass_ifu_exu_sr_mux_n20));
AND2X1 exu_U5653(.A(exu_n4753), .B(exu_n9572), .Y(bypass_ifu_exu_sr_mux_n19));
AND2X1 exu_U5654(.A(exu_n4758), .B(exu_n9573), .Y(bypass_ifu_exu_sr_mux_n50));
AND2X1 exu_U5655(.A(exu_n4759), .B(exu_n9574), .Y(bypass_ifu_exu_sr_mux_n49));
AND2X1 exu_U5656(.A(exu_n4770), .B(exu_n9575), .Y(bypass_ifu_exu_sr_mux_n116));
AND2X1 exu_U5657(.A(exu_n4771), .B(exu_n9576), .Y(bypass_ifu_exu_sr_mux_n115));
AND2X1 exu_U5658(.A(exu_n4782), .B(exu_n9577), .Y(bypass_ifu_exu_sr_mux_n182));
AND2X1 exu_U5659(.A(exu_n4783), .B(exu_n9578), .Y(bypass_ifu_exu_sr_mux_n181));
INVX1 exu_U5660(.A(exu_n16031), .Y(exu_n16030));
AND2X1 exu_U5661(.A(exu_n4794), .B(exu_n9581), .Y(bypass_ifu_exu_sr_mux_n248));
AND2X1 exu_U5662(.A(exu_n4795), .B(exu_n9582), .Y(bypass_ifu_exu_sr_mux_n247));
INVX1 exu_U5663(.A(exu_n16031), .Y(exu_n16029));
AND2X1 exu_U5664(.A(exu_n4806), .B(exu_n9593), .Y(bypass_ifu_exu_sr_mux_n314));
AND2X1 exu_U5665(.A(exu_n4807), .B(exu_n9594), .Y(bypass_ifu_exu_sr_mux_n313));
INVX1 exu_U5666(.A(exu_n16031), .Y(exu_n16028));
AND2X1 exu_U5667(.A(exu_n4818), .B(exu_n9605), .Y(bypass_ifu_exu_sr_mux_n380));
AND2X1 exu_U5668(.A(exu_n4819), .B(exu_n9606), .Y(bypass_ifu_exu_sr_mux_n379));
INVX1 exu_U5669(.A(exu_n16032), .Y(exu_n16027));
INVX1 exu_U5670(.A(exu_n16039), .Y(exu_n16033));
INVX1 exu_U5671(.A(exu_n16038), .Y(exu_n16037));
INVX1 exu_U5672(.A(exu_n16038), .Y(exu_n16036));
INVX1 exu_U5673(.A(exu_n16038), .Y(exu_n16035));
INVX1 exu_U5674(.A(exu_n16039), .Y(exu_n16034));
OR2X1 exu_U5675(.A(exu_n12342), .B(exu_n13754), .Y(bypass_byp_irf_rd_data_m[63]));
AND2X1 exu_U5676(.A(exu_n1562), .B(exu_n6580), .Y(exu_n23225));
OR2X1 exu_U5677(.A(exu_n12343), .B(exu_n13755), .Y(bypass_byp_irf_rd_data_m[62]));
AND2X1 exu_U5678(.A(exu_n1564), .B(exu_n6582), .Y(exu_n23231));
OR2X1 exu_U5679(.A(exu_n12344), .B(exu_n13756), .Y(bypass_byp_irf_rd_data_m[61]));
AND2X1 exu_U5680(.A(exu_n1566), .B(exu_n6584), .Y(exu_n23237));
OR2X1 exu_U5681(.A(exu_n12345), .B(exu_n13757), .Y(bypass_byp_irf_rd_data_m[60]));
AND2X1 exu_U5682(.A(exu_n1568), .B(exu_n6586), .Y(exu_n23243));
OR2X1 exu_U5683(.A(exu_n12347), .B(exu_n13759), .Y(bypass_byp_irf_rd_data_m[59]));
AND2X1 exu_U5684(.A(exu_n1572), .B(exu_n6590), .Y(exu_n23255));
OR2X1 exu_U5685(.A(exu_n12348), .B(exu_n13760), .Y(bypass_byp_irf_rd_data_m[58]));
AND2X1 exu_U5686(.A(exu_n1574), .B(exu_n6592), .Y(exu_n23261));
OR2X1 exu_U5687(.A(exu_n12349), .B(exu_n13761), .Y(bypass_byp_irf_rd_data_m[57]));
AND2X1 exu_U5688(.A(exu_n1576), .B(exu_n6594), .Y(exu_n23267));
OR2X1 exu_U5689(.A(exu_n12350), .B(exu_n13762), .Y(bypass_byp_irf_rd_data_m[56]));
AND2X1 exu_U5690(.A(exu_n1578), .B(exu_n6596), .Y(exu_n23273));
OR2X1 exu_U5691(.A(exu_n12351), .B(exu_n13763), .Y(bypass_byp_irf_rd_data_m[55]));
AND2X1 exu_U5692(.A(exu_n1580), .B(exu_n6598), .Y(exu_n23279));
OR2X1 exu_U5693(.A(exu_n12352), .B(exu_n13764), .Y(bypass_byp_irf_rd_data_m[54]));
AND2X1 exu_U5694(.A(exu_n1582), .B(exu_n6600), .Y(exu_n23285));
OR2X1 exu_U5695(.A(exu_n12353), .B(exu_n13765), .Y(bypass_byp_irf_rd_data_m[53]));
AND2X1 exu_U5696(.A(exu_n1584), .B(exu_n6602), .Y(exu_n23291));
OR2X1 exu_U5697(.A(exu_n12354), .B(exu_n13766), .Y(bypass_byp_irf_rd_data_m[52]));
AND2X1 exu_U5698(.A(exu_n1586), .B(exu_n6604), .Y(exu_n23297));
OR2X1 exu_U5699(.A(exu_n12355), .B(exu_n13767), .Y(bypass_byp_irf_rd_data_m[51]));
AND2X1 exu_U5700(.A(exu_n1588), .B(exu_n6606), .Y(exu_n23303));
OR2X1 exu_U5701(.A(exu_n12356), .B(exu_n13768), .Y(bypass_byp_irf_rd_data_m[50]));
AND2X1 exu_U5702(.A(exu_n1590), .B(exu_n6608), .Y(exu_n23309));
OR2X1 exu_U5703(.A(exu_n12358), .B(exu_n13770), .Y(bypass_byp_irf_rd_data_m[49]));
AND2X1 exu_U5704(.A(exu_n1594), .B(exu_n6612), .Y(exu_n23321));
OR2X1 exu_U5705(.A(exu_n12359), .B(exu_n13771), .Y(bypass_byp_irf_rd_data_m[48]));
AND2X1 exu_U5706(.A(exu_n1596), .B(exu_n6614), .Y(exu_n23327));
OR2X1 exu_U5707(.A(exu_n12360), .B(exu_n13772), .Y(bypass_byp_irf_rd_data_m[47]));
AND2X1 exu_U5708(.A(exu_n1598), .B(exu_n6616), .Y(exu_n23333));
OR2X1 exu_U5709(.A(exu_n12361), .B(exu_n13773), .Y(bypass_byp_irf_rd_data_m[46]));
AND2X1 exu_U5710(.A(exu_n1600), .B(exu_n6618), .Y(exu_n23339));
OR2X1 exu_U5711(.A(exu_n12362), .B(exu_n13774), .Y(bypass_byp_irf_rd_data_m[45]));
AND2X1 exu_U5712(.A(exu_n1602), .B(exu_n6620), .Y(exu_n23345));
OR2X1 exu_U5713(.A(exu_n12363), .B(exu_n13775), .Y(bypass_byp_irf_rd_data_m[44]));
AND2X1 exu_U5714(.A(exu_n1604), .B(exu_n6622), .Y(exu_n23351));
OR2X1 exu_U5715(.A(exu_n12364), .B(exu_n13776), .Y(bypass_byp_irf_rd_data_m[43]));
AND2X1 exu_U5716(.A(exu_n1606), .B(exu_n6624), .Y(exu_n23357));
OR2X1 exu_U5717(.A(exu_n12365), .B(exu_n13777), .Y(bypass_byp_irf_rd_data_m[42]));
AND2X1 exu_U5718(.A(exu_n1608), .B(exu_n6626), .Y(exu_n23363));
OR2X1 exu_U5719(.A(exu_n12366), .B(exu_n13778), .Y(bypass_byp_irf_rd_data_m[41]));
AND2X1 exu_U5720(.A(exu_n1610), .B(exu_n6628), .Y(exu_n23369));
OR2X1 exu_U5721(.A(exu_n12367), .B(exu_n13779), .Y(bypass_byp_irf_rd_data_m[40]));
AND2X1 exu_U5722(.A(exu_n1612), .B(exu_n6630), .Y(exu_n23375));
OR2X1 exu_U5723(.A(exu_n12369), .B(exu_n13781), .Y(bypass_byp_irf_rd_data_m[39]));
AND2X1 exu_U5724(.A(exu_n1616), .B(exu_n6634), .Y(exu_n23387));
OR2X1 exu_U5725(.A(exu_n12370), .B(exu_n13782), .Y(bypass_byp_irf_rd_data_m[38]));
AND2X1 exu_U5726(.A(exu_n1618), .B(exu_n6636), .Y(exu_n23393));
OR2X1 exu_U5727(.A(exu_n12371), .B(exu_n13783), .Y(bypass_byp_irf_rd_data_m[37]));
AND2X1 exu_U5728(.A(exu_n1620), .B(exu_n6638), .Y(exu_n23399));
OR2X1 exu_U5729(.A(exu_n12372), .B(exu_n13784), .Y(bypass_byp_irf_rd_data_m[36]));
AND2X1 exu_U5730(.A(exu_n1622), .B(exu_n6640), .Y(exu_n23405));
OR2X1 exu_U5731(.A(exu_n12373), .B(exu_n13785), .Y(bypass_byp_irf_rd_data_m[35]));
AND2X1 exu_U5732(.A(exu_n1624), .B(exu_n6642), .Y(exu_n23411));
OR2X1 exu_U5733(.A(exu_n12374), .B(exu_n13786), .Y(bypass_byp_irf_rd_data_m[34]));
AND2X1 exu_U5734(.A(exu_n1626), .B(exu_n6644), .Y(exu_n23417));
OR2X1 exu_U5735(.A(exu_n12375), .B(exu_n13787), .Y(bypass_byp_irf_rd_data_m[33]));
AND2X1 exu_U5736(.A(exu_n1628), .B(exu_n6646), .Y(exu_n23423));
OR2X1 exu_U5737(.A(exu_n12376), .B(exu_n13788), .Y(bypass_byp_irf_rd_data_m[32]));
AND2X1 exu_U5738(.A(exu_n1630), .B(exu_n6648), .Y(exu_n23429));
OR2X1 exu_U5739(.A(exu_n12377), .B(exu_n13789), .Y(bypass_byp_irf_rd_data_m[31]));
AND2X1 exu_U5740(.A(exu_n1632), .B(exu_n6650), .Y(exu_n23435));
OR2X1 exu_U5741(.A(exu_n12378), .B(exu_n13790), .Y(bypass_byp_irf_rd_data_m[30]));
AND2X1 exu_U5742(.A(exu_n1634), .B(exu_n6652), .Y(exu_n23441));
OR2X1 exu_U5743(.A(exu_n12380), .B(exu_n13792), .Y(bypass_byp_irf_rd_data_m[29]));
AND2X1 exu_U5744(.A(exu_n1638), .B(exu_n6656), .Y(exu_n23453));
OR2X1 exu_U5745(.A(exu_n12381), .B(exu_n13793), .Y(bypass_byp_irf_rd_data_m[28]));
AND2X1 exu_U5746(.A(exu_n1640), .B(exu_n6658), .Y(exu_n23459));
OR2X1 exu_U5747(.A(exu_n12382), .B(exu_n13794), .Y(bypass_byp_irf_rd_data_m[27]));
AND2X1 exu_U5748(.A(exu_n1642), .B(exu_n6660), .Y(exu_n23465));
OR2X1 exu_U5749(.A(exu_n12383), .B(exu_n13795), .Y(bypass_byp_irf_rd_data_m[26]));
AND2X1 exu_U5750(.A(exu_n1644), .B(exu_n6662), .Y(exu_n23471));
OR2X1 exu_U5751(.A(exu_n12384), .B(exu_n13796), .Y(bypass_byp_irf_rd_data_m[25]));
AND2X1 exu_U5752(.A(exu_n1646), .B(exu_n6664), .Y(exu_n23477));
OR2X1 exu_U5753(.A(exu_n12385), .B(exu_n13797), .Y(bypass_byp_irf_rd_data_m[24]));
AND2X1 exu_U5754(.A(exu_n1648), .B(exu_n6666), .Y(exu_n23483));
OR2X1 exu_U5755(.A(exu_n12386), .B(exu_n13798), .Y(bypass_byp_irf_rd_data_m[23]));
AND2X1 exu_U5756(.A(exu_n1650), .B(exu_n6668), .Y(exu_n23489));
OR2X1 exu_U5757(.A(exu_n12387), .B(exu_n13799), .Y(bypass_byp_irf_rd_data_m[22]));
AND2X1 exu_U5758(.A(exu_n1652), .B(exu_n6670), .Y(exu_n23495));
OR2X1 exu_U5759(.A(exu_n12388), .B(exu_n13800), .Y(bypass_byp_irf_rd_data_m[21]));
AND2X1 exu_U5760(.A(exu_n1654), .B(exu_n6672), .Y(exu_n23501));
OR2X1 exu_U5761(.A(exu_n12389), .B(exu_n13801), .Y(bypass_byp_irf_rd_data_m[20]));
AND2X1 exu_U5762(.A(exu_n1656), .B(exu_n6674), .Y(exu_n23507));
OR2X1 exu_U5763(.A(exu_n12391), .B(exu_n13803), .Y(bypass_byp_irf_rd_data_m[19]));
AND2X1 exu_U5764(.A(exu_n1660), .B(exu_n6678), .Y(exu_n23519));
OR2X1 exu_U5765(.A(exu_n12392), .B(exu_n13804), .Y(bypass_byp_irf_rd_data_m[18]));
AND2X1 exu_U5766(.A(exu_n1662), .B(exu_n6680), .Y(exu_n23525));
OR2X1 exu_U5767(.A(exu_n12393), .B(exu_n13805), .Y(bypass_byp_irf_rd_data_m[17]));
AND2X1 exu_U5768(.A(exu_n1664), .B(exu_n6682), .Y(exu_n23531));
OR2X1 exu_U5769(.A(exu_n12394), .B(exu_n13806), .Y(bypass_byp_irf_rd_data_m[16]));
AND2X1 exu_U5770(.A(exu_n1666), .B(exu_n6684), .Y(exu_n23537));
OR2X1 exu_U5771(.A(exu_n12395), .B(exu_n13807), .Y(bypass_byp_irf_rd_data_m[15]));
AND2X1 exu_U5772(.A(exu_n1668), .B(exu_n6686), .Y(exu_n23543));
OR2X1 exu_U5773(.A(exu_n12396), .B(exu_n13808), .Y(bypass_byp_irf_rd_data_m[14]));
AND2X1 exu_U5774(.A(exu_n1670), .B(exu_n6688), .Y(exu_n23549));
OR2X1 exu_U5775(.A(exu_n12397), .B(exu_n13809), .Y(bypass_byp_irf_rd_data_m[13]));
AND2X1 exu_U5776(.A(exu_n1672), .B(exu_n6690), .Y(exu_n23555));
OR2X1 exu_U5777(.A(exu_n12398), .B(exu_n13810), .Y(bypass_byp_irf_rd_data_m[12]));
AND2X1 exu_U5778(.A(exu_n1674), .B(exu_n6692), .Y(exu_n23561));
OR2X1 exu_U5779(.A(exu_n12399), .B(exu_n13811), .Y(bypass_byp_irf_rd_data_m[11]));
AND2X1 exu_U5780(.A(exu_n1676), .B(exu_n6694), .Y(exu_n23567));
OR2X1 exu_U5781(.A(exu_n12400), .B(exu_n13812), .Y(bypass_byp_irf_rd_data_m[10]));
AND2X1 exu_U5782(.A(exu_n1678), .B(exu_n6696), .Y(exu_n23573));
OR2X1 exu_U5783(.A(exu_n12338), .B(exu_n13750), .Y(bypass_byp_irf_rd_data_m[9]));
AND2X1 exu_U5784(.A(exu_n1554), .B(exu_n6572), .Y(exu_n23201));
OR2X1 exu_U5785(.A(exu_n12339), .B(exu_n13751), .Y(bypass_byp_irf_rd_data_m[8]));
AND2X1 exu_U5786(.A(exu_n1556), .B(exu_n6574), .Y(exu_n23207));
OR2X1 exu_U5787(.A(exu_n12340), .B(exu_n13752), .Y(bypass_byp_irf_rd_data_m[7]));
AND2X1 exu_U5788(.A(exu_n1558), .B(exu_n6576), .Y(exu_n23213));
INVX1 exu_U5789(.A(exu_n16046), .Y(exu_n16040));
OR2X1 exu_U5790(.A(exu_n12341), .B(exu_n13753), .Y(bypass_byp_irf_rd_data_m[6]));
AND2X1 exu_U5791(.A(exu_n1560), .B(exu_n6578), .Y(exu_n23219));
OR2X1 exu_U5792(.A(exu_n12346), .B(exu_n13758), .Y(bypass_byp_irf_rd_data_m[5]));
AND2X1 exu_U5793(.A(exu_n1570), .B(exu_n6588), .Y(exu_n23249));
OR2X1 exu_U5794(.A(exu_n12357), .B(exu_n13769), .Y(bypass_byp_irf_rd_data_m[4]));
AND2X1 exu_U5795(.A(exu_n1592), .B(exu_n6610), .Y(exu_n23315));
OR2X1 exu_U5796(.A(exu_n12368), .B(exu_n13780), .Y(bypass_byp_irf_rd_data_m[3]));
AND2X1 exu_U5797(.A(exu_n1614), .B(exu_n6632), .Y(exu_n23381));
INVX1 exu_U5798(.A(exu_n16045), .Y(exu_n16044));
OR2X1 exu_U5799(.A(exu_n12379), .B(exu_n13791), .Y(bypass_byp_irf_rd_data_m[2]));
AND2X1 exu_U5800(.A(exu_n1636), .B(exu_n6654), .Y(exu_n23447));
INVX1 exu_U5801(.A(exu_n16045), .Y(exu_n16043));
OR2X1 exu_U5802(.A(exu_n12390), .B(exu_n13802), .Y(bypass_byp_irf_rd_data_m[1]));
AND2X1 exu_U5803(.A(exu_n1658), .B(exu_n6676), .Y(exu_n23513));
INVX1 exu_U5804(.A(exu_n16045), .Y(exu_n16042));
OR2X1 exu_U5805(.A(exu_n12401), .B(exu_n13813), .Y(bypass_byp_irf_rd_data_m[0]));
AND2X1 exu_U5806(.A(exu_n1680), .B(exu_n6698), .Y(exu_n23579));
INVX1 exu_U5807(.A(exu_n16046), .Y(exu_n16041));
AND2X1 exu_U5808(.A(exu_n22577), .B(exu_n6259), .Y(bypass_rd_data_g[63]));
AND2X1 exu_U5809(.A(exu_n1429), .B(exu_n6260), .Y(exu_n22577));
AND2X1 exu_U5810(.A(exu_n22581), .B(exu_n6261), .Y(bypass_rd_data_g[62]));
AND2X1 exu_U5811(.A(exu_n1430), .B(exu_n6262), .Y(exu_n22581));
AND2X1 exu_U5812(.A(exu_n22585), .B(exu_n6263), .Y(bypass_rd_data_g[61]));
AND2X1 exu_U5813(.A(exu_n1431), .B(exu_n6264), .Y(exu_n22585));
AND2X1 exu_U5814(.A(exu_n22589), .B(exu_n6265), .Y(bypass_rd_data_g[60]));
AND2X1 exu_U5815(.A(exu_n1432), .B(exu_n6266), .Y(exu_n22589));
AND2X1 exu_U5816(.A(exu_n22597), .B(exu_n6269), .Y(bypass_rd_data_g[59]));
AND2X1 exu_U5817(.A(exu_n1434), .B(exu_n6270), .Y(exu_n22597));
AND2X1 exu_U5818(.A(exu_n22601), .B(exu_n6271), .Y(bypass_rd_data_g[58]));
AND2X1 exu_U5819(.A(exu_n1435), .B(exu_n6272), .Y(exu_n22601));
AND2X1 exu_U5820(.A(exu_n22605), .B(exu_n6273), .Y(bypass_rd_data_g[57]));
AND2X1 exu_U5821(.A(exu_n1436), .B(exu_n6274), .Y(exu_n22605));
AND2X1 exu_U5822(.A(exu_n22609), .B(exu_n6275), .Y(bypass_rd_data_g[56]));
AND2X1 exu_U5823(.A(exu_n1437), .B(exu_n6276), .Y(exu_n22609));
AND2X1 exu_U5824(.A(exu_n22613), .B(exu_n6277), .Y(bypass_rd_data_g[55]));
AND2X1 exu_U5825(.A(exu_n1438), .B(exu_n6278), .Y(exu_n22613));
AND2X1 exu_U5826(.A(exu_n22617), .B(exu_n6279), .Y(bypass_rd_data_g[54]));
AND2X1 exu_U5827(.A(exu_n1439), .B(exu_n6280), .Y(exu_n22617));
AND2X1 exu_U5828(.A(exu_n22621), .B(exu_n6281), .Y(bypass_rd_data_g[53]));
AND2X1 exu_U5829(.A(exu_n1440), .B(exu_n6282), .Y(exu_n22621));
AND2X1 exu_U5830(.A(exu_n22625), .B(exu_n6283), .Y(bypass_rd_data_g[52]));
AND2X1 exu_U5831(.A(exu_n1441), .B(exu_n6284), .Y(exu_n22625));
AND2X1 exu_U5832(.A(exu_n22629), .B(exu_n6285), .Y(bypass_rd_data_g[51]));
AND2X1 exu_U5833(.A(exu_n1442), .B(exu_n6286), .Y(exu_n22629));
AND2X1 exu_U5834(.A(exu_n22633), .B(exu_n6287), .Y(bypass_rd_data_g[50]));
AND2X1 exu_U5835(.A(exu_n1443), .B(exu_n6288), .Y(exu_n22633));
AND2X1 exu_U5836(.A(exu_n22641), .B(exu_n6291), .Y(bypass_rd_data_g[49]));
AND2X1 exu_U5837(.A(exu_n1445), .B(exu_n6292), .Y(exu_n22641));
AND2X1 exu_U5838(.A(exu_n22645), .B(exu_n6293), .Y(bypass_rd_data_g[48]));
AND2X1 exu_U5839(.A(exu_n1446), .B(exu_n6294), .Y(exu_n22645));
AND2X1 exu_U5840(.A(exu_n22649), .B(exu_n6295), .Y(bypass_rd_data_g[47]));
AND2X1 exu_U5841(.A(exu_n1447), .B(exu_n6296), .Y(exu_n22649));
AND2X1 exu_U5842(.A(exu_n22653), .B(exu_n6297), .Y(bypass_rd_data_g[46]));
AND2X1 exu_U5843(.A(exu_n1448), .B(exu_n6298), .Y(exu_n22653));
AND2X1 exu_U5844(.A(exu_n22657), .B(exu_n6299), .Y(bypass_rd_data_g[45]));
AND2X1 exu_U5845(.A(exu_n1449), .B(exu_n6300), .Y(exu_n22657));
AND2X1 exu_U5846(.A(exu_n22661), .B(exu_n6301), .Y(bypass_rd_data_g[44]));
AND2X1 exu_U5847(.A(exu_n1450), .B(exu_n6302), .Y(exu_n22661));
AND2X1 exu_U5848(.A(exu_n22665), .B(exu_n6303), .Y(bypass_rd_data_g[43]));
AND2X1 exu_U5849(.A(exu_n1451), .B(exu_n6304), .Y(exu_n22665));
AND2X1 exu_U5850(.A(exu_n22669), .B(exu_n6305), .Y(bypass_rd_data_g[42]));
AND2X1 exu_U5851(.A(exu_n1452), .B(exu_n6306), .Y(exu_n22669));
AND2X1 exu_U5852(.A(exu_n22673), .B(exu_n6307), .Y(bypass_rd_data_g[41]));
AND2X1 exu_U5853(.A(exu_n1453), .B(exu_n6308), .Y(exu_n22673));
AND2X1 exu_U5854(.A(exu_n22677), .B(exu_n6309), .Y(bypass_rd_data_g[40]));
AND2X1 exu_U5855(.A(exu_n1454), .B(exu_n6310), .Y(exu_n22677));
AND2X1 exu_U5856(.A(exu_n22685), .B(exu_n6313), .Y(bypass_rd_data_g[39]));
AND2X1 exu_U5857(.A(exu_n1456), .B(exu_n6314), .Y(exu_n22685));
AND2X1 exu_U5858(.A(exu_n22689), .B(exu_n6315), .Y(bypass_rd_data_g[38]));
AND2X1 exu_U5859(.A(exu_n1457), .B(exu_n6316), .Y(exu_n22689));
AND2X1 exu_U5860(.A(exu_n22693), .B(exu_n6317), .Y(bypass_rd_data_g[37]));
AND2X1 exu_U5861(.A(exu_n1458), .B(exu_n6318), .Y(exu_n22693));
AND2X1 exu_U5862(.A(exu_n22697), .B(exu_n6319), .Y(bypass_rd_data_g[36]));
AND2X1 exu_U5863(.A(exu_n1459), .B(exu_n6320), .Y(exu_n22697));
AND2X1 exu_U5864(.A(exu_n22701), .B(exu_n6321), .Y(bypass_rd_data_g[35]));
AND2X1 exu_U5865(.A(exu_n1460), .B(exu_n6322), .Y(exu_n22701));
AND2X1 exu_U5866(.A(exu_n22705), .B(exu_n6323), .Y(bypass_rd_data_g[34]));
AND2X1 exu_U5867(.A(exu_n1461), .B(exu_n6324), .Y(exu_n22705));
AND2X1 exu_U5868(.A(exu_n22709), .B(exu_n6325), .Y(bypass_rd_data_g[33]));
AND2X1 exu_U5869(.A(exu_n1462), .B(exu_n6326), .Y(exu_n22709));
AND2X1 exu_U5870(.A(exu_n22713), .B(exu_n6327), .Y(bypass_rd_data_g[32]));
AND2X1 exu_U5871(.A(exu_n1463), .B(exu_n6328), .Y(exu_n22713));
AND2X1 exu_U5872(.A(exu_n22717), .B(exu_n6329), .Y(bypass_rd_data_g[31]));
AND2X1 exu_U5873(.A(exu_n1464), .B(exu_n6330), .Y(exu_n22717));
AND2X1 exu_U5874(.A(exu_n22721), .B(exu_n6331), .Y(bypass_rd_data_g[30]));
AND2X1 exu_U5875(.A(exu_n1465), .B(exu_n6332), .Y(exu_n22721));
AND2X1 exu_U5876(.A(exu_n22729), .B(exu_n6335), .Y(bypass_rd_data_g[29]));
AND2X1 exu_U5877(.A(exu_n1467), .B(exu_n6336), .Y(exu_n22729));
AND2X1 exu_U5878(.A(exu_n22733), .B(exu_n6337), .Y(bypass_rd_data_g[28]));
AND2X1 exu_U5879(.A(exu_n1468), .B(exu_n6338), .Y(exu_n22733));
AND2X1 exu_U5880(.A(exu_n22737), .B(exu_n6339), .Y(bypass_rd_data_g[27]));
AND2X1 exu_U5881(.A(exu_n1469), .B(exu_n6340), .Y(exu_n22737));
AND2X1 exu_U5882(.A(exu_n22741), .B(exu_n6341), .Y(bypass_rd_data_g[26]));
AND2X1 exu_U5883(.A(exu_n1470), .B(exu_n6342), .Y(exu_n22741));
AND2X1 exu_U5884(.A(exu_n22745), .B(exu_n6343), .Y(bypass_rd_data_g[25]));
AND2X1 exu_U5885(.A(exu_n1471), .B(exu_n6344), .Y(exu_n22745));
AND2X1 exu_U5886(.A(exu_n22749), .B(exu_n6345), .Y(bypass_rd_data_g[24]));
AND2X1 exu_U5887(.A(exu_n1472), .B(exu_n6346), .Y(exu_n22749));
AND2X1 exu_U5888(.A(exu_n22753), .B(exu_n6347), .Y(bypass_rd_data_g[23]));
AND2X1 exu_U5889(.A(exu_n1473), .B(exu_n6348), .Y(exu_n22753));
AND2X1 exu_U5890(.A(exu_n22757), .B(exu_n6349), .Y(bypass_rd_data_g[22]));
AND2X1 exu_U5891(.A(exu_n1474), .B(exu_n6350), .Y(exu_n22757));
AND2X1 exu_U5892(.A(exu_n22761), .B(exu_n6351), .Y(bypass_rd_data_g[21]));
AND2X1 exu_U5893(.A(exu_n1475), .B(exu_n6352), .Y(exu_n22761));
AND2X1 exu_U5894(.A(exu_n22765), .B(exu_n6353), .Y(bypass_rd_data_g[20]));
AND2X1 exu_U5895(.A(exu_n1476), .B(exu_n6354), .Y(exu_n22765));
AND2X1 exu_U5896(.A(exu_n22773), .B(exu_n6357), .Y(bypass_rd_data_g[19]));
AND2X1 exu_U5897(.A(exu_n1478), .B(exu_n6358), .Y(exu_n22773));
AND2X1 exu_U5898(.A(exu_n22777), .B(exu_n6359), .Y(bypass_rd_data_g[18]));
AND2X1 exu_U5899(.A(exu_n1479), .B(exu_n6360), .Y(exu_n22777));
AND2X1 exu_U5900(.A(exu_n22781), .B(exu_n6361), .Y(bypass_rd_data_g[17]));
AND2X1 exu_U5901(.A(exu_n1480), .B(exu_n6362), .Y(exu_n22781));
AND2X1 exu_U5902(.A(exu_n22785), .B(exu_n6363), .Y(bypass_rd_data_g[16]));
AND2X1 exu_U5903(.A(exu_n1481), .B(exu_n6364), .Y(exu_n22785));
AND2X1 exu_U5904(.A(exu_n22789), .B(exu_n6365), .Y(bypass_rd_data_g[15]));
AND2X1 exu_U5905(.A(exu_n1482), .B(exu_n6366), .Y(exu_n22789));
AND2X1 exu_U5906(.A(exu_n22793), .B(exu_n6367), .Y(bypass_rd_data_g[14]));
AND2X1 exu_U5907(.A(exu_n1483), .B(exu_n6368), .Y(exu_n22793));
AND2X1 exu_U5908(.A(exu_n22797), .B(exu_n6369), .Y(bypass_rd_data_g[13]));
AND2X1 exu_U5909(.A(exu_n1484), .B(exu_n6370), .Y(exu_n22797));
AND2X1 exu_U5910(.A(exu_n22801), .B(exu_n6371), .Y(bypass_rd_data_g[12]));
AND2X1 exu_U5911(.A(exu_n1485), .B(exu_n6372), .Y(exu_n22801));
AND2X1 exu_U5912(.A(exu_n22805), .B(exu_n6373), .Y(bypass_rd_data_g[11]));
AND2X1 exu_U5913(.A(exu_n1486), .B(exu_n6374), .Y(exu_n22805));
AND2X1 exu_U5914(.A(exu_n22809), .B(exu_n6375), .Y(bypass_rd_data_g[10]));
AND2X1 exu_U5915(.A(exu_n1487), .B(exu_n6376), .Y(exu_n22809));
AND2X1 exu_U5916(.A(exu_n22561), .B(exu_n6251), .Y(bypass_rd_data_g[9]));
AND2X1 exu_U5917(.A(exu_n1425), .B(exu_n6252), .Y(exu_n22561));
AND2X1 exu_U5918(.A(exu_n22565), .B(exu_n6253), .Y(bypass_rd_data_g[8]));
AND2X1 exu_U5919(.A(exu_n1426), .B(exu_n6254), .Y(exu_n22565));
AND2X1 exu_U5920(.A(exu_n22569), .B(exu_n6255), .Y(bypass_rd_data_g[7]));
AND2X1 exu_U5921(.A(exu_n1427), .B(exu_n6256), .Y(exu_n22569));
INVX1 exu_U5922(.A(exu_n16053), .Y(exu_n16047));
AND2X1 exu_U5923(.A(exu_n22573), .B(exu_n6257), .Y(bypass_rd_data_g[6]));
AND2X1 exu_U5924(.A(exu_n1428), .B(exu_n6258), .Y(exu_n22573));
AND2X1 exu_U5925(.A(exu_n22593), .B(exu_n6267), .Y(bypass_rd_data_g[5]));
AND2X1 exu_U5926(.A(exu_n1433), .B(exu_n6268), .Y(exu_n22593));
AND2X1 exu_U5927(.A(exu_n22637), .B(exu_n6289), .Y(bypass_rd_data_g[4]));
AND2X1 exu_U5928(.A(exu_n1444), .B(exu_n6290), .Y(exu_n22637));
AND2X1 exu_U5929(.A(exu_n22681), .B(exu_n6311), .Y(bypass_rd_data_g[3]));
AND2X1 exu_U5930(.A(exu_n1455), .B(exu_n6312), .Y(exu_n22681));
INVX1 exu_U5931(.A(exu_n16052), .Y(exu_n16051));
AND2X1 exu_U5932(.A(exu_n22725), .B(exu_n6333), .Y(bypass_rd_data_g[2]));
AND2X1 exu_U5933(.A(exu_n1466), .B(exu_n6334), .Y(exu_n22725));
INVX1 exu_U5934(.A(exu_n16052), .Y(exu_n16050));
AND2X1 exu_U5935(.A(exu_n22769), .B(exu_n6355), .Y(bypass_rd_data_g[1]));
AND2X1 exu_U5936(.A(exu_n1477), .B(exu_n6356), .Y(exu_n22769));
INVX1 exu_U5937(.A(exu_n16052), .Y(exu_n16049));
AND2X1 exu_U5938(.A(exu_n22813), .B(exu_n6377), .Y(bypass_rd_data_g[0]));
AND2X1 exu_U5939(.A(exu_n1488), .B(exu_n6378), .Y(exu_n22813));
INVX1 exu_U5940(.A(exu_n16053), .Y(exu_n16048));
AND2X1 exu_U5941(.A(exu_n1805), .B(exu_n6835), .Y(exu_n23978));
AND2X1 exu_U5942(.A(exu_n1806), .B(exu_n6836), .Y(exu_n23977));
AND2X1 exu_U5943(.A(exu_n1807), .B(exu_n6837), .Y(exu_n23984));
AND2X1 exu_U5944(.A(exu_n1808), .B(exu_n6838), .Y(exu_n23983));
AND2X1 exu_U5945(.A(exu_n1809), .B(exu_n6839), .Y(exu_n23990));
AND2X1 exu_U5946(.A(exu_n1810), .B(exu_n6840), .Y(exu_n23989));
AND2X1 exu_U5947(.A(exu_n1811), .B(exu_n6841), .Y(exu_n23996));
AND2X1 exu_U5948(.A(exu_n1812), .B(exu_n6842), .Y(exu_n23995));
AND2X1 exu_U5949(.A(exu_n1815), .B(exu_n6845), .Y(exu_n24008));
AND2X1 exu_U5950(.A(exu_n1816), .B(exu_n6846), .Y(exu_n24007));
AND2X1 exu_U5951(.A(exu_n1817), .B(exu_n6847), .Y(exu_n24014));
AND2X1 exu_U5952(.A(exu_n1818), .B(exu_n6848), .Y(exu_n24013));
AND2X1 exu_U5953(.A(exu_n1819), .B(exu_n6849), .Y(exu_n24020));
AND2X1 exu_U5954(.A(exu_n1820), .B(exu_n6850), .Y(exu_n24019));
AND2X1 exu_U5955(.A(exu_n1821), .B(exu_n6851), .Y(exu_n24026));
AND2X1 exu_U5956(.A(exu_n1822), .B(exu_n6852), .Y(exu_n24025));
AND2X1 exu_U5957(.A(exu_n1823), .B(exu_n6853), .Y(exu_n24032));
AND2X1 exu_U5958(.A(exu_n1824), .B(exu_n6854), .Y(exu_n24031));
AND2X1 exu_U5959(.A(exu_n1825), .B(exu_n6855), .Y(exu_n24038));
AND2X1 exu_U5960(.A(exu_n1826), .B(exu_n6856), .Y(exu_n24037));
AND2X1 exu_U5961(.A(exu_n1827), .B(exu_n6857), .Y(exu_n24044));
AND2X1 exu_U5962(.A(exu_n1828), .B(exu_n6858), .Y(exu_n24043));
AND2X1 exu_U5963(.A(exu_n1829), .B(exu_n6859), .Y(exu_n24050));
AND2X1 exu_U5964(.A(exu_n1830), .B(exu_n6860), .Y(exu_n24049));
AND2X1 exu_U5965(.A(exu_n1831), .B(exu_n6861), .Y(exu_n24056));
AND2X1 exu_U5966(.A(exu_n1832), .B(exu_n6862), .Y(exu_n24055));
AND2X1 exu_U5967(.A(exu_n1833), .B(exu_n6863), .Y(exu_n24062));
AND2X1 exu_U5968(.A(exu_n1834), .B(exu_n6864), .Y(exu_n24061));
AND2X1 exu_U5969(.A(exu_n1837), .B(exu_n6867), .Y(exu_n24074));
AND2X1 exu_U5970(.A(exu_n1838), .B(exu_n6868), .Y(exu_n24073));
AND2X1 exu_U5971(.A(exu_n1839), .B(exu_n6869), .Y(exu_n24080));
AND2X1 exu_U5972(.A(exu_n1840), .B(exu_n6870), .Y(exu_n24079));
AND2X1 exu_U5973(.A(exu_n1841), .B(exu_n6871), .Y(exu_n24086));
AND2X1 exu_U5974(.A(exu_n1842), .B(exu_n6872), .Y(exu_n24085));
AND2X1 exu_U5975(.A(exu_n1843), .B(exu_n6873), .Y(exu_n24092));
AND2X1 exu_U5976(.A(exu_n1844), .B(exu_n6874), .Y(exu_n24091));
AND2X1 exu_U5977(.A(exu_n1845), .B(exu_n6875), .Y(exu_n24098));
AND2X1 exu_U5978(.A(exu_n1846), .B(exu_n6876), .Y(exu_n24097));
AND2X1 exu_U5979(.A(exu_n1847), .B(exu_n6877), .Y(exu_n24104));
AND2X1 exu_U5980(.A(exu_n1848), .B(exu_n6878), .Y(exu_n24103));
AND2X1 exu_U5981(.A(exu_n1849), .B(exu_n6879), .Y(exu_n24110));
AND2X1 exu_U5982(.A(exu_n1850), .B(exu_n6880), .Y(exu_n24109));
AND2X1 exu_U5983(.A(exu_n1851), .B(exu_n6881), .Y(exu_n24116));
AND2X1 exu_U5984(.A(exu_n1852), .B(exu_n6882), .Y(exu_n24115));
AND2X1 exu_U5985(.A(exu_n1853), .B(exu_n6883), .Y(exu_n24122));
AND2X1 exu_U5986(.A(exu_n1854), .B(exu_n6884), .Y(exu_n24121));
AND2X1 exu_U5987(.A(exu_n1855), .B(exu_n6885), .Y(exu_n24128));
AND2X1 exu_U5988(.A(exu_n1856), .B(exu_n6886), .Y(exu_n24127));
AND2X1 exu_U5989(.A(exu_n1859), .B(exu_n6889), .Y(exu_n24140));
AND2X1 exu_U5990(.A(exu_n1860), .B(exu_n6890), .Y(exu_n24139));
AND2X1 exu_U5991(.A(exu_n1861), .B(exu_n6891), .Y(exu_n24146));
AND2X1 exu_U5992(.A(exu_n1862), .B(exu_n6892), .Y(exu_n24145));
AND2X1 exu_U5993(.A(exu_n1863), .B(exu_n6893), .Y(exu_n24152));
AND2X1 exu_U5994(.A(exu_n1864), .B(exu_n6894), .Y(exu_n24151));
AND2X1 exu_U5995(.A(exu_n1865), .B(exu_n6895), .Y(exu_n24158));
AND2X1 exu_U5996(.A(exu_n1866), .B(exu_n6896), .Y(exu_n24157));
AND2X1 exu_U5997(.A(exu_n1867), .B(exu_n6897), .Y(exu_n24164));
AND2X1 exu_U5998(.A(exu_n1868), .B(exu_n6898), .Y(exu_n24163));
AND2X1 exu_U5999(.A(exu_n1869), .B(exu_n6899), .Y(exu_n24170));
AND2X1 exu_U6000(.A(exu_n1870), .B(exu_n6900), .Y(exu_n24169));
AND2X1 exu_U6001(.A(exu_n1871), .B(exu_n6901), .Y(exu_n24176));
AND2X1 exu_U6002(.A(exu_n1872), .B(exu_n6902), .Y(exu_n24175));
AND2X1 exu_U6003(.A(exu_n1873), .B(exu_n6903), .Y(exu_n24182));
AND2X1 exu_U6004(.A(exu_n1874), .B(exu_n6904), .Y(exu_n24181));
AND2X1 exu_U6005(.A(exu_n1875), .B(exu_n6905), .Y(exu_n24188));
AND2X1 exu_U6006(.A(exu_n1876), .B(exu_n6906), .Y(exu_n24187));
AND2X1 exu_U6007(.A(exu_n1877), .B(exu_n6907), .Y(exu_n24194));
AND2X1 exu_U6008(.A(exu_n1878), .B(exu_n6908), .Y(exu_n24193));
AND2X1 exu_U6009(.A(exu_n1881), .B(exu_n6911), .Y(exu_n24206));
AND2X1 exu_U6010(.A(exu_n1882), .B(exu_n6912), .Y(exu_n24205));
AND2X1 exu_U6011(.A(exu_n1883), .B(exu_n6913), .Y(exu_n24212));
AND2X1 exu_U6012(.A(exu_n1884), .B(exu_n6914), .Y(exu_n24211));
AND2X1 exu_U6013(.A(exu_n1885), .B(exu_n6915), .Y(exu_n24218));
AND2X1 exu_U6014(.A(exu_n1886), .B(exu_n6916), .Y(exu_n24217));
AND2X1 exu_U6015(.A(exu_n1887), .B(exu_n6917), .Y(exu_n24224));
AND2X1 exu_U6016(.A(exu_n1888), .B(exu_n6918), .Y(exu_n24223));
AND2X1 exu_U6017(.A(exu_n1889), .B(exu_n6919), .Y(exu_n24230));
AND2X1 exu_U6018(.A(exu_n1890), .B(exu_n6920), .Y(exu_n24229));
AND2X1 exu_U6019(.A(exu_n1891), .B(exu_n6921), .Y(exu_n24236));
AND2X1 exu_U6020(.A(exu_n1892), .B(exu_n6922), .Y(exu_n24235));
AND2X1 exu_U6021(.A(exu_n1893), .B(exu_n6923), .Y(exu_n24242));
AND2X1 exu_U6022(.A(exu_n1894), .B(exu_n6924), .Y(exu_n24241));
AND2X1 exu_U6023(.A(exu_n1895), .B(exu_n6925), .Y(exu_n24248));
AND2X1 exu_U6024(.A(exu_n1896), .B(exu_n6926), .Y(exu_n24247));
AND2X1 exu_U6025(.A(exu_n1897), .B(exu_n6927), .Y(exu_n24254));
AND2X1 exu_U6026(.A(exu_n1898), .B(exu_n6928), .Y(exu_n24253));
AND2X1 exu_U6027(.A(exu_n1899), .B(exu_n6929), .Y(exu_n24260));
AND2X1 exu_U6028(.A(exu_n1900), .B(exu_n6930), .Y(exu_n24259));
AND2X1 exu_U6029(.A(exu_n1903), .B(exu_n6933), .Y(exu_n24272));
AND2X1 exu_U6030(.A(exu_n1904), .B(exu_n6934), .Y(exu_n24271));
AND2X1 exu_U6031(.A(exu_n1905), .B(exu_n6935), .Y(exu_n24278));
AND2X1 exu_U6032(.A(exu_n1906), .B(exu_n6936), .Y(exu_n24277));
AND2X1 exu_U6033(.A(exu_n1907), .B(exu_n6937), .Y(exu_n24284));
AND2X1 exu_U6034(.A(exu_n1908), .B(exu_n6938), .Y(exu_n24283));
AND2X1 exu_U6035(.A(exu_n1909), .B(exu_n6939), .Y(exu_n24290));
AND2X1 exu_U6036(.A(exu_n1910), .B(exu_n6940), .Y(exu_n24289));
AND2X1 exu_U6037(.A(exu_n1911), .B(exu_n6941), .Y(exu_n24296));
AND2X1 exu_U6038(.A(exu_n1912), .B(exu_n6942), .Y(exu_n24295));
AND2X1 exu_U6039(.A(exu_n1913), .B(exu_n6943), .Y(exu_n24302));
AND2X1 exu_U6040(.A(exu_n1914), .B(exu_n6944), .Y(exu_n24301));
AND2X1 exu_U6041(.A(exu_n1915), .B(exu_n6945), .Y(exu_n24308));
AND2X1 exu_U6042(.A(exu_n1916), .B(exu_n6946), .Y(exu_n24307));
AND2X1 exu_U6043(.A(exu_n1917), .B(exu_n6947), .Y(exu_n24314));
AND2X1 exu_U6044(.A(exu_n1918), .B(exu_n6948), .Y(exu_n24313));
AND2X1 exu_U6045(.A(exu_n1919), .B(exu_n6949), .Y(exu_n24320));
AND2X1 exu_U6046(.A(exu_n1920), .B(exu_n6950), .Y(exu_n24319));
AND2X1 exu_U6047(.A(exu_n1921), .B(exu_n6951), .Y(exu_n24326));
AND2X1 exu_U6048(.A(exu_n1922), .B(exu_n6952), .Y(exu_n24325));
AND2X1 exu_U6049(.A(exu_n1797), .B(exu_n6827), .Y(exu_n23954));
AND2X1 exu_U6050(.A(exu_n1798), .B(exu_n6828), .Y(exu_n23953));
AND2X1 exu_U6051(.A(exu_n1799), .B(exu_n6829), .Y(exu_n23960));
AND2X1 exu_U6052(.A(exu_n1800), .B(exu_n6830), .Y(exu_n23959));
AND2X1 exu_U6053(.A(exu_n1801), .B(exu_n6831), .Y(exu_n23966));
AND2X1 exu_U6054(.A(exu_n1802), .B(exu_n6832), .Y(exu_n23965));
INVX1 exu_U6055(.A(exu_n16060), .Y(exu_n16054));
AND2X1 exu_U6056(.A(exu_n1803), .B(exu_n6833), .Y(exu_n23972));
AND2X1 exu_U6057(.A(exu_n1804), .B(exu_n6834), .Y(exu_n23971));
AND2X1 exu_U6058(.A(exu_n1813), .B(exu_n6843), .Y(exu_n24002));
AND2X1 exu_U6059(.A(exu_n1814), .B(exu_n6844), .Y(exu_n24001));
AND2X1 exu_U6060(.A(exu_n1835), .B(exu_n6865), .Y(exu_n24068));
AND2X1 exu_U6061(.A(exu_n1836), .B(exu_n6866), .Y(exu_n24067));
AND2X1 exu_U6062(.A(exu_n1857), .B(exu_n6887), .Y(exu_n24134));
AND2X1 exu_U6063(.A(exu_n1858), .B(exu_n6888), .Y(exu_n24133));
INVX1 exu_U6064(.A(exu_n16059), .Y(exu_n16058));
AND2X1 exu_U6065(.A(exu_n1879), .B(exu_n6909), .Y(exu_n24200));
AND2X1 exu_U6066(.A(exu_n1880), .B(exu_n6910), .Y(exu_n24199));
INVX1 exu_U6067(.A(exu_n16059), .Y(exu_n16057));
AND2X1 exu_U6068(.A(exu_n1901), .B(exu_n6931), .Y(exu_n24266));
AND2X1 exu_U6069(.A(exu_n1902), .B(exu_n6932), .Y(exu_n24265));
INVX1 exu_U6070(.A(exu_n16059), .Y(exu_n16056));
AND2X1 exu_U6071(.A(exu_n1923), .B(exu_n6953), .Y(exu_n24332));
AND2X1 exu_U6072(.A(exu_n1924), .B(exu_n6954), .Y(exu_n24331));
INVX1 exu_U6073(.A(exu_n16060), .Y(exu_n16055));
AND2X1 exu_U6074(.A(exu_n2255), .B(exu_n7283), .Y(exu_n25354));
AND2X1 exu_U6075(.A(exu_n2256), .B(exu_n7284), .Y(exu_n25353));
AND2X1 exu_U6076(.A(exu_n2257), .B(exu_n7285), .Y(exu_n25360));
AND2X1 exu_U6077(.A(exu_n2258), .B(exu_n7286), .Y(exu_n25359));
AND2X1 exu_U6078(.A(exu_n2259), .B(exu_n7287), .Y(exu_n25366));
AND2X1 exu_U6079(.A(exu_n2260), .B(exu_n7288), .Y(exu_n25365));
AND2X1 exu_U6080(.A(exu_n2261), .B(exu_n7289), .Y(exu_n25372));
AND2X1 exu_U6081(.A(exu_n2262), .B(exu_n7290), .Y(exu_n25371));
AND2X1 exu_U6082(.A(exu_n2265), .B(exu_n7293), .Y(exu_n25384));
AND2X1 exu_U6083(.A(exu_n2266), .B(exu_n7294), .Y(exu_n25383));
AND2X1 exu_U6084(.A(exu_n2267), .B(exu_n7295), .Y(exu_n25390));
AND2X1 exu_U6085(.A(exu_n2268), .B(exu_n7296), .Y(exu_n25389));
AND2X1 exu_U6086(.A(exu_n2269), .B(exu_n7297), .Y(exu_n25396));
AND2X1 exu_U6087(.A(exu_n2270), .B(exu_n7298), .Y(exu_n25395));
AND2X1 exu_U6088(.A(exu_n2271), .B(exu_n7299), .Y(exu_n25402));
AND2X1 exu_U6089(.A(exu_n2272), .B(exu_n7300), .Y(exu_n25401));
AND2X1 exu_U6090(.A(exu_n2273), .B(exu_n7301), .Y(exu_n25408));
AND2X1 exu_U6091(.A(exu_n2274), .B(exu_n7302), .Y(exu_n25407));
AND2X1 exu_U6092(.A(exu_n2275), .B(exu_n7303), .Y(exu_n25414));
AND2X1 exu_U6093(.A(exu_n2276), .B(exu_n7304), .Y(exu_n25413));
AND2X1 exu_U6094(.A(exu_n2277), .B(exu_n7305), .Y(exu_n25420));
AND2X1 exu_U6095(.A(exu_n2278), .B(exu_n7306), .Y(exu_n25419));
AND2X1 exu_U6096(.A(exu_n2279), .B(exu_n7307), .Y(exu_n25426));
AND2X1 exu_U6097(.A(exu_n2280), .B(exu_n7308), .Y(exu_n25425));
AND2X1 exu_U6098(.A(exu_n2281), .B(exu_n7309), .Y(exu_n25432));
AND2X1 exu_U6099(.A(exu_n2282), .B(exu_n7310), .Y(exu_n25431));
AND2X1 exu_U6100(.A(exu_n2283), .B(exu_n7311), .Y(exu_n25438));
AND2X1 exu_U6101(.A(exu_n2284), .B(exu_n7312), .Y(exu_n25437));
AND2X1 exu_U6102(.A(exu_n2287), .B(exu_n7315), .Y(exu_n25450));
AND2X1 exu_U6103(.A(exu_n2288), .B(exu_n7316), .Y(exu_n25449));
AND2X1 exu_U6104(.A(exu_n2289), .B(exu_n7317), .Y(exu_n25456));
AND2X1 exu_U6105(.A(exu_n2290), .B(exu_n7318), .Y(exu_n25455));
AND2X1 exu_U6106(.A(exu_n2291), .B(exu_n7319), .Y(exu_n25462));
AND2X1 exu_U6107(.A(exu_n2292), .B(exu_n7320), .Y(exu_n25461));
AND2X1 exu_U6108(.A(exu_n2293), .B(exu_n7321), .Y(exu_n25468));
AND2X1 exu_U6109(.A(exu_n2294), .B(exu_n7322), .Y(exu_n25467));
AND2X1 exu_U6110(.A(exu_n2295), .B(exu_n7323), .Y(exu_n25474));
AND2X1 exu_U6111(.A(exu_n2296), .B(exu_n7324), .Y(exu_n25473));
AND2X1 exu_U6112(.A(exu_n2297), .B(exu_n7325), .Y(exu_n25480));
AND2X1 exu_U6113(.A(exu_n2298), .B(exu_n7326), .Y(exu_n25479));
AND2X1 exu_U6114(.A(exu_n2299), .B(exu_n7327), .Y(exu_n25486));
AND2X1 exu_U6115(.A(exu_n2300), .B(exu_n7328), .Y(exu_n25485));
AND2X1 exu_U6116(.A(exu_n2301), .B(exu_n7329), .Y(exu_n25492));
AND2X1 exu_U6117(.A(exu_n2302), .B(exu_n7330), .Y(exu_n25491));
AND2X1 exu_U6118(.A(exu_n2303), .B(exu_n7331), .Y(exu_n25498));
AND2X1 exu_U6119(.A(exu_n2304), .B(exu_n7332), .Y(exu_n25497));
AND2X1 exu_U6120(.A(exu_n2305), .B(exu_n7333), .Y(exu_n25504));
AND2X1 exu_U6121(.A(exu_n2306), .B(exu_n7334), .Y(exu_n25503));
AND2X1 exu_U6122(.A(exu_n2309), .B(exu_n7337), .Y(exu_n25516));
AND2X1 exu_U6123(.A(exu_n2310), .B(exu_n7338), .Y(exu_n25515));
AND2X1 exu_U6124(.A(exu_n2311), .B(exu_n7339), .Y(exu_n25522));
AND2X1 exu_U6125(.A(exu_n2312), .B(exu_n7340), .Y(exu_n25521));
AND2X1 exu_U6126(.A(exu_n2313), .B(exu_n7341), .Y(exu_n25528));
AND2X1 exu_U6127(.A(exu_n2314), .B(exu_n7342), .Y(exu_n25527));
AND2X1 exu_U6128(.A(exu_n2315), .B(exu_n7343), .Y(exu_n25534));
AND2X1 exu_U6129(.A(exu_n2316), .B(exu_n7344), .Y(exu_n25533));
AND2X1 exu_U6130(.A(exu_n2317), .B(exu_n7345), .Y(exu_n25540));
AND2X1 exu_U6131(.A(exu_n2318), .B(exu_n7346), .Y(exu_n25539));
AND2X1 exu_U6132(.A(exu_n2319), .B(exu_n7347), .Y(exu_n25546));
AND2X1 exu_U6133(.A(exu_n2320), .B(exu_n7348), .Y(exu_n25545));
AND2X1 exu_U6134(.A(exu_n2321), .B(exu_n7349), .Y(exu_n25552));
AND2X1 exu_U6135(.A(exu_n2322), .B(exu_n7350), .Y(exu_n25551));
AND2X1 exu_U6136(.A(exu_n2323), .B(exu_n7351), .Y(exu_n25558));
AND2X1 exu_U6137(.A(exu_n2324), .B(exu_n7352), .Y(exu_n25557));
AND2X1 exu_U6138(.A(exu_n2325), .B(exu_n7353), .Y(exu_n25564));
AND2X1 exu_U6139(.A(exu_n2326), .B(exu_n7354), .Y(exu_n25563));
AND2X1 exu_U6140(.A(exu_n2327), .B(exu_n7355), .Y(exu_n25570));
AND2X1 exu_U6141(.A(exu_n2328), .B(exu_n7356), .Y(exu_n25569));
AND2X1 exu_U6142(.A(exu_n2331), .B(exu_n7359), .Y(exu_n25582));
AND2X1 exu_U6143(.A(exu_n2332), .B(exu_n7360), .Y(exu_n25581));
AND2X1 exu_U6144(.A(exu_n2333), .B(exu_n7361), .Y(exu_n25588));
AND2X1 exu_U6145(.A(exu_n2334), .B(exu_n7362), .Y(exu_n25587));
AND2X1 exu_U6146(.A(exu_n2335), .B(exu_n7363), .Y(exu_n25594));
AND2X1 exu_U6147(.A(exu_n2336), .B(exu_n7364), .Y(exu_n25593));
AND2X1 exu_U6148(.A(exu_n2337), .B(exu_n7365), .Y(exu_n25600));
AND2X1 exu_U6149(.A(exu_n2338), .B(exu_n7366), .Y(exu_n25599));
AND2X1 exu_U6150(.A(exu_n2339), .B(exu_n7367), .Y(exu_n25606));
AND2X1 exu_U6151(.A(exu_n2340), .B(exu_n7368), .Y(exu_n25605));
AND2X1 exu_U6152(.A(exu_n2341), .B(exu_n7369), .Y(exu_n25612));
AND2X1 exu_U6153(.A(exu_n2342), .B(exu_n7370), .Y(exu_n25611));
AND2X1 exu_U6154(.A(exu_n2343), .B(exu_n7371), .Y(exu_n25618));
AND2X1 exu_U6155(.A(exu_n2344), .B(exu_n7372), .Y(exu_n25617));
AND2X1 exu_U6156(.A(exu_n2345), .B(exu_n7373), .Y(exu_n25624));
AND2X1 exu_U6157(.A(exu_n2346), .B(exu_n7374), .Y(exu_n25623));
AND2X1 exu_U6158(.A(exu_n2347), .B(exu_n7375), .Y(exu_n25630));
AND2X1 exu_U6159(.A(exu_n2348), .B(exu_n7376), .Y(exu_n25629));
AND2X1 exu_U6160(.A(exu_n2349), .B(exu_n7377), .Y(exu_n25636));
AND2X1 exu_U6161(.A(exu_n2350), .B(exu_n7378), .Y(exu_n25635));
AND2X1 exu_U6162(.A(exu_n2353), .B(exu_n7381), .Y(exu_n25648));
AND2X1 exu_U6163(.A(exu_n2354), .B(exu_n7382), .Y(exu_n25647));
AND2X1 exu_U6164(.A(exu_n2355), .B(exu_n7383), .Y(exu_n25654));
AND2X1 exu_U6165(.A(exu_n2356), .B(exu_n7384), .Y(exu_n25653));
AND2X1 exu_U6166(.A(exu_n2357), .B(exu_n7385), .Y(exu_n25660));
AND2X1 exu_U6167(.A(exu_n2358), .B(exu_n7386), .Y(exu_n25659));
AND2X1 exu_U6168(.A(exu_n2359), .B(exu_n7387), .Y(exu_n25666));
AND2X1 exu_U6169(.A(exu_n2360), .B(exu_n7388), .Y(exu_n25665));
AND2X1 exu_U6170(.A(exu_n2361), .B(exu_n7389), .Y(exu_n25672));
AND2X1 exu_U6171(.A(exu_n2362), .B(exu_n7390), .Y(exu_n25671));
AND2X1 exu_U6172(.A(exu_n2363), .B(exu_n7391), .Y(exu_n25678));
AND2X1 exu_U6173(.A(exu_n2364), .B(exu_n7392), .Y(exu_n25677));
AND2X1 exu_U6174(.A(exu_n2365), .B(exu_n7393), .Y(exu_n25684));
AND2X1 exu_U6175(.A(exu_n2366), .B(exu_n7394), .Y(exu_n25683));
AND2X1 exu_U6176(.A(exu_n2367), .B(exu_n7395), .Y(exu_n25690));
AND2X1 exu_U6177(.A(exu_n2368), .B(exu_n7396), .Y(exu_n25689));
AND2X1 exu_U6178(.A(exu_n2369), .B(exu_n7397), .Y(exu_n25696));
AND2X1 exu_U6179(.A(exu_n2370), .B(exu_n7398), .Y(exu_n25695));
AND2X1 exu_U6180(.A(exu_n2371), .B(exu_n7399), .Y(exu_n25702));
AND2X1 exu_U6181(.A(exu_n2372), .B(exu_n7400), .Y(exu_n25701));
AND2X1 exu_U6182(.A(exu_n2247), .B(exu_n7275), .Y(exu_n25330));
AND2X1 exu_U6183(.A(exu_n2248), .B(exu_n7276), .Y(exu_n25329));
AND2X1 exu_U6184(.A(exu_n2249), .B(exu_n7277), .Y(exu_n25336));
AND2X1 exu_U6185(.A(exu_n2250), .B(exu_n7278), .Y(exu_n25335));
AND2X1 exu_U6186(.A(exu_n2251), .B(exu_n7279), .Y(exu_n25342));
AND2X1 exu_U6187(.A(exu_n2252), .B(exu_n7280), .Y(exu_n25341));
INVX1 exu_U6188(.A(exu_n16067), .Y(exu_n16061));
AND2X1 exu_U6189(.A(exu_n2253), .B(exu_n7281), .Y(exu_n25348));
AND2X1 exu_U6190(.A(exu_n2254), .B(exu_n7282), .Y(exu_n25347));
AND2X1 exu_U6191(.A(exu_n2263), .B(exu_n7291), .Y(exu_n25378));
AND2X1 exu_U6192(.A(exu_n2264), .B(exu_n7292), .Y(exu_n25377));
AND2X1 exu_U6193(.A(exu_n2285), .B(exu_n7313), .Y(exu_n25444));
AND2X1 exu_U6194(.A(exu_n2286), .B(exu_n7314), .Y(exu_n25443));
AND2X1 exu_U6195(.A(exu_n2307), .B(exu_n7335), .Y(exu_n25510));
AND2X1 exu_U6196(.A(exu_n2308), .B(exu_n7336), .Y(exu_n25509));
INVX1 exu_U6197(.A(exu_n16066), .Y(exu_n16065));
AND2X1 exu_U6198(.A(exu_n2329), .B(exu_n7357), .Y(exu_n25576));
AND2X1 exu_U6199(.A(exu_n2330), .B(exu_n7358), .Y(exu_n25575));
INVX1 exu_U6200(.A(exu_n16066), .Y(exu_n16064));
AND2X1 exu_U6201(.A(exu_n2351), .B(exu_n7379), .Y(exu_n25642));
AND2X1 exu_U6202(.A(exu_n2352), .B(exu_n7380), .Y(exu_n25641));
INVX1 exu_U6203(.A(exu_n16066), .Y(exu_n16063));
AND2X1 exu_U6204(.A(exu_n2373), .B(exu_n7401), .Y(exu_n25708));
AND2X1 exu_U6205(.A(exu_n2374), .B(exu_n7402), .Y(exu_n25707));
INVX1 exu_U6206(.A(exu_n16067), .Y(exu_n16062));
AND2X1 exu_U6207(.A(exu_n2447), .B(exu_n7475), .Y(exu_n25994));
AND2X1 exu_U6208(.A(exu_n2448), .B(exu_n7476), .Y(exu_n25993));
AND2X1 exu_U6209(.A(exu_n2449), .B(exu_n7477), .Y(exu_n26000));
AND2X1 exu_U6210(.A(exu_n2450), .B(exu_n7478), .Y(exu_n25999));
AND2X1 exu_U6211(.A(exu_n2451), .B(exu_n7479), .Y(exu_n26006));
AND2X1 exu_U6212(.A(exu_n2452), .B(exu_n7480), .Y(exu_n26005));
AND2X1 exu_U6213(.A(exu_n2453), .B(exu_n7481), .Y(exu_n26012));
AND2X1 exu_U6214(.A(exu_n2454), .B(exu_n7482), .Y(exu_n26011));
AND2X1 exu_U6215(.A(exu_n2457), .B(exu_n7485), .Y(exu_n26024));
AND2X1 exu_U6216(.A(exu_n2458), .B(exu_n7486), .Y(exu_n26023));
AND2X1 exu_U6217(.A(exu_n2459), .B(exu_n7487), .Y(exu_n26030));
AND2X1 exu_U6218(.A(exu_n2460), .B(exu_n7488), .Y(exu_n26029));
AND2X1 exu_U6219(.A(exu_n2461), .B(exu_n7489), .Y(exu_n26036));
AND2X1 exu_U6220(.A(exu_n2462), .B(exu_n7490), .Y(exu_n26035));
AND2X1 exu_U6221(.A(exu_n2463), .B(exu_n7491), .Y(exu_n26042));
AND2X1 exu_U6222(.A(exu_n2464), .B(exu_n7492), .Y(exu_n26041));
AND2X1 exu_U6223(.A(exu_n2465), .B(exu_n7493), .Y(exu_n26048));
AND2X1 exu_U6224(.A(exu_n2466), .B(exu_n7494), .Y(exu_n26047));
AND2X1 exu_U6225(.A(exu_n2467), .B(exu_n7495), .Y(exu_n26054));
AND2X1 exu_U6226(.A(exu_n2468), .B(exu_n7496), .Y(exu_n26053));
AND2X1 exu_U6227(.A(exu_n2469), .B(exu_n7497), .Y(exu_n26060));
AND2X1 exu_U6228(.A(exu_n2470), .B(exu_n7498), .Y(exu_n26059));
AND2X1 exu_U6229(.A(exu_n2471), .B(exu_n7499), .Y(exu_n26066));
AND2X1 exu_U6230(.A(exu_n2472), .B(exu_n7500), .Y(exu_n26065));
AND2X1 exu_U6231(.A(exu_n2473), .B(exu_n7501), .Y(exu_n26072));
AND2X1 exu_U6232(.A(exu_n2474), .B(exu_n7502), .Y(exu_n26071));
AND2X1 exu_U6233(.A(exu_n2475), .B(exu_n7503), .Y(exu_n26078));
AND2X1 exu_U6234(.A(exu_n2476), .B(exu_n7504), .Y(exu_n26077));
AND2X1 exu_U6235(.A(exu_n2479), .B(exu_n7507), .Y(exu_n26090));
AND2X1 exu_U6236(.A(exu_n2480), .B(exu_n7508), .Y(exu_n26089));
AND2X1 exu_U6237(.A(exu_n2481), .B(exu_n7509), .Y(exu_n26096));
AND2X1 exu_U6238(.A(exu_n2482), .B(exu_n7510), .Y(exu_n26095));
AND2X1 exu_U6239(.A(exu_n2483), .B(exu_n7511), .Y(exu_n26102));
AND2X1 exu_U6240(.A(exu_n2484), .B(exu_n7512), .Y(exu_n26101));
AND2X1 exu_U6241(.A(exu_n2485), .B(exu_n7513), .Y(exu_n26108));
AND2X1 exu_U6242(.A(exu_n2486), .B(exu_n7514), .Y(exu_n26107));
AND2X1 exu_U6243(.A(exu_n2487), .B(exu_n7515), .Y(exu_n26114));
AND2X1 exu_U6244(.A(exu_n2488), .B(exu_n7516), .Y(exu_n26113));
AND2X1 exu_U6245(.A(exu_n2489), .B(exu_n7517), .Y(exu_n26120));
AND2X1 exu_U6246(.A(exu_n2490), .B(exu_n7518), .Y(exu_n26119));
AND2X1 exu_U6247(.A(exu_n2491), .B(exu_n7519), .Y(exu_n26126));
AND2X1 exu_U6248(.A(exu_n2492), .B(exu_n7520), .Y(exu_n26125));
AND2X1 exu_U6249(.A(exu_n2493), .B(exu_n7521), .Y(exu_n26132));
AND2X1 exu_U6250(.A(exu_n2494), .B(exu_n7522), .Y(exu_n26131));
AND2X1 exu_U6251(.A(exu_n2495), .B(exu_n7523), .Y(exu_n26138));
AND2X1 exu_U6252(.A(exu_n2496), .B(exu_n7524), .Y(exu_n26137));
AND2X1 exu_U6253(.A(exu_n2497), .B(exu_n7525), .Y(exu_n26144));
AND2X1 exu_U6254(.A(exu_n2498), .B(exu_n7526), .Y(exu_n26143));
AND2X1 exu_U6255(.A(exu_n2501), .B(exu_n7529), .Y(exu_n26156));
AND2X1 exu_U6256(.A(exu_n2502), .B(exu_n7530), .Y(exu_n26155));
AND2X1 exu_U6257(.A(exu_n2503), .B(exu_n7531), .Y(exu_n26162));
AND2X1 exu_U6258(.A(exu_n2504), .B(exu_n7532), .Y(exu_n26161));
AND2X1 exu_U6259(.A(exu_n2505), .B(exu_n7533), .Y(exu_n26168));
AND2X1 exu_U6260(.A(exu_n2506), .B(exu_n7534), .Y(exu_n26167));
AND2X1 exu_U6261(.A(exu_n2507), .B(exu_n7535), .Y(exu_n26174));
AND2X1 exu_U6262(.A(exu_n2508), .B(exu_n7536), .Y(exu_n26173));
AND2X1 exu_U6263(.A(exu_n2509), .B(exu_n7537), .Y(exu_n26180));
AND2X1 exu_U6264(.A(exu_n2510), .B(exu_n7538), .Y(exu_n26179));
AND2X1 exu_U6265(.A(exu_n2511), .B(exu_n7539), .Y(exu_n26186));
AND2X1 exu_U6266(.A(exu_n2512), .B(exu_n7540), .Y(exu_n26185));
AND2X1 exu_U6267(.A(exu_n2513), .B(exu_n7541), .Y(exu_n26192));
AND2X1 exu_U6268(.A(exu_n2514), .B(exu_n7542), .Y(exu_n26191));
AND2X1 exu_U6269(.A(exu_n2515), .B(exu_n7543), .Y(exu_n26198));
AND2X1 exu_U6270(.A(exu_n2516), .B(exu_n7544), .Y(exu_n26197));
AND2X1 exu_U6271(.A(exu_n2517), .B(exu_n7545), .Y(exu_n26204));
AND2X1 exu_U6272(.A(exu_n2518), .B(exu_n7546), .Y(exu_n26203));
AND2X1 exu_U6273(.A(exu_n2519), .B(exu_n7547), .Y(exu_n26210));
AND2X1 exu_U6274(.A(exu_n2520), .B(exu_n7548), .Y(exu_n26209));
AND2X1 exu_U6275(.A(exu_n2523), .B(exu_n7551), .Y(exu_n26222));
AND2X1 exu_U6276(.A(exu_n2524), .B(exu_n7552), .Y(exu_n26221));
AND2X1 exu_U6277(.A(exu_n2525), .B(exu_n7553), .Y(exu_n26228));
AND2X1 exu_U6278(.A(exu_n2526), .B(exu_n7554), .Y(exu_n26227));
AND2X1 exu_U6279(.A(exu_n2527), .B(exu_n7555), .Y(exu_n26234));
AND2X1 exu_U6280(.A(exu_n2528), .B(exu_n7556), .Y(exu_n26233));
AND2X1 exu_U6281(.A(exu_n2529), .B(exu_n7557), .Y(exu_n26240));
AND2X1 exu_U6282(.A(exu_n2530), .B(exu_n7558), .Y(exu_n26239));
AND2X1 exu_U6283(.A(exu_n2531), .B(exu_n7559), .Y(exu_n26246));
AND2X1 exu_U6284(.A(exu_n2532), .B(exu_n7560), .Y(exu_n26245));
AND2X1 exu_U6285(.A(exu_n2533), .B(exu_n7561), .Y(exu_n26252));
AND2X1 exu_U6286(.A(exu_n2534), .B(exu_n7562), .Y(exu_n26251));
AND2X1 exu_U6287(.A(exu_n2535), .B(exu_n7563), .Y(exu_n26258));
AND2X1 exu_U6288(.A(exu_n2536), .B(exu_n7564), .Y(exu_n26257));
AND2X1 exu_U6289(.A(exu_n2537), .B(exu_n7565), .Y(exu_n26264));
AND2X1 exu_U6290(.A(exu_n2538), .B(exu_n7566), .Y(exu_n26263));
AND2X1 exu_U6291(.A(exu_n2539), .B(exu_n7567), .Y(exu_n26270));
AND2X1 exu_U6292(.A(exu_n2540), .B(exu_n7568), .Y(exu_n26269));
AND2X1 exu_U6293(.A(exu_n2541), .B(exu_n7569), .Y(exu_n26276));
AND2X1 exu_U6294(.A(exu_n2542), .B(exu_n7570), .Y(exu_n26275));
AND2X1 exu_U6295(.A(exu_n2545), .B(exu_n7573), .Y(exu_n26288));
AND2X1 exu_U6296(.A(exu_n2546), .B(exu_n7574), .Y(exu_n26287));
AND2X1 exu_U6297(.A(exu_n2547), .B(exu_n7575), .Y(exu_n26294));
AND2X1 exu_U6298(.A(exu_n2548), .B(exu_n7576), .Y(exu_n26293));
AND2X1 exu_U6299(.A(exu_n2549), .B(exu_n7577), .Y(exu_n26300));
AND2X1 exu_U6300(.A(exu_n2550), .B(exu_n7578), .Y(exu_n26299));
AND2X1 exu_U6301(.A(exu_n2551), .B(exu_n7579), .Y(exu_n26306));
AND2X1 exu_U6302(.A(exu_n2552), .B(exu_n7580), .Y(exu_n26305));
AND2X1 exu_U6303(.A(exu_n2553), .B(exu_n7581), .Y(exu_n26312));
AND2X1 exu_U6304(.A(exu_n2554), .B(exu_n7582), .Y(exu_n26311));
AND2X1 exu_U6305(.A(exu_n2555), .B(exu_n7583), .Y(exu_n26318));
AND2X1 exu_U6306(.A(exu_n2556), .B(exu_n7584), .Y(exu_n26317));
AND2X1 exu_U6307(.A(exu_n2557), .B(exu_n7585), .Y(exu_n26324));
AND2X1 exu_U6308(.A(exu_n2558), .B(exu_n7586), .Y(exu_n26323));
AND2X1 exu_U6309(.A(exu_n2559), .B(exu_n7587), .Y(exu_n26330));
AND2X1 exu_U6310(.A(exu_n2560), .B(exu_n7588), .Y(exu_n26329));
AND2X1 exu_U6311(.A(exu_n2561), .B(exu_n7589), .Y(exu_n26336));
AND2X1 exu_U6312(.A(exu_n2562), .B(exu_n7590), .Y(exu_n26335));
AND2X1 exu_U6313(.A(exu_n2563), .B(exu_n7591), .Y(exu_n26342));
AND2X1 exu_U6314(.A(exu_n2564), .B(exu_n7592), .Y(exu_n26341));
AND2X1 exu_U6315(.A(exu_n2439), .B(exu_n7467), .Y(exu_n25970));
AND2X1 exu_U6316(.A(exu_n2440), .B(exu_n7468), .Y(exu_n25969));
AND2X1 exu_U6317(.A(exu_n2441), .B(exu_n7469), .Y(exu_n25976));
AND2X1 exu_U6318(.A(exu_n2442), .B(exu_n7470), .Y(exu_n25975));
AND2X1 exu_U6319(.A(exu_n2443), .B(exu_n7471), .Y(exu_n25982));
AND2X1 exu_U6320(.A(exu_n2444), .B(exu_n7472), .Y(exu_n25981));
INVX1 exu_U6321(.A(exu_n16074), .Y(exu_n16068));
AND2X1 exu_U6322(.A(exu_n2445), .B(exu_n7473), .Y(exu_n25988));
AND2X1 exu_U6323(.A(exu_n2446), .B(exu_n7474), .Y(exu_n25987));
AND2X1 exu_U6324(.A(exu_n2455), .B(exu_n7483), .Y(exu_n26018));
AND2X1 exu_U6325(.A(exu_n2456), .B(exu_n7484), .Y(exu_n26017));
AND2X1 exu_U6326(.A(exu_n2477), .B(exu_n7505), .Y(exu_n26084));
AND2X1 exu_U6327(.A(exu_n2478), .B(exu_n7506), .Y(exu_n26083));
AND2X1 exu_U6328(.A(exu_n2499), .B(exu_n7527), .Y(exu_n26150));
AND2X1 exu_U6329(.A(exu_n2500), .B(exu_n7528), .Y(exu_n26149));
INVX1 exu_U6330(.A(exu_n16073), .Y(exu_n16072));
AND2X1 exu_U6331(.A(exu_n2521), .B(exu_n7549), .Y(exu_n26216));
AND2X1 exu_U6332(.A(exu_n2522), .B(exu_n7550), .Y(exu_n26215));
INVX1 exu_U6333(.A(exu_n16073), .Y(exu_n16071));
AND2X1 exu_U6334(.A(exu_n2543), .B(exu_n7571), .Y(exu_n26282));
AND2X1 exu_U6335(.A(exu_n2544), .B(exu_n7572), .Y(exu_n26281));
INVX1 exu_U6336(.A(exu_n16073), .Y(exu_n16070));
AND2X1 exu_U6337(.A(exu_n2565), .B(exu_n7593), .Y(exu_n26348));
AND2X1 exu_U6338(.A(exu_n2566), .B(exu_n7594), .Y(exu_n26347));
INVX1 exu_U6339(.A(exu_n16074), .Y(exu_n16069));
AND2X1 exu_U6340(.A(exu_n1997), .B(exu_n7027), .Y(exu_n24618));
AND2X1 exu_U6341(.A(exu_n1998), .B(exu_n7028), .Y(exu_n24617));
AND2X1 exu_U6342(.A(exu_n1999), .B(exu_n7029), .Y(exu_n24624));
AND2X1 exu_U6343(.A(exu_n2000), .B(exu_n7030), .Y(exu_n24623));
AND2X1 exu_U6344(.A(exu_n2001), .B(exu_n7031), .Y(exu_n24630));
AND2X1 exu_U6345(.A(exu_n2002), .B(exu_n7032), .Y(exu_n24629));
AND2X1 exu_U6346(.A(exu_n2003), .B(exu_n7033), .Y(exu_n24636));
AND2X1 exu_U6347(.A(exu_n2004), .B(exu_n7034), .Y(exu_n24635));
AND2X1 exu_U6348(.A(exu_n2007), .B(exu_n7037), .Y(exu_n24648));
AND2X1 exu_U6349(.A(exu_n2008), .B(exu_n7038), .Y(exu_n24647));
AND2X1 exu_U6350(.A(exu_n2009), .B(exu_n7039), .Y(exu_n24654));
AND2X1 exu_U6351(.A(exu_n2010), .B(exu_n7040), .Y(exu_n24653));
AND2X1 exu_U6352(.A(exu_n2011), .B(exu_n7041), .Y(exu_n24660));
AND2X1 exu_U6353(.A(exu_n2012), .B(exu_n7042), .Y(exu_n24659));
AND2X1 exu_U6354(.A(exu_n2013), .B(exu_n7043), .Y(exu_n24666));
AND2X1 exu_U6355(.A(exu_n2014), .B(exu_n7044), .Y(exu_n24665));
AND2X1 exu_U6356(.A(exu_n2015), .B(exu_n7045), .Y(exu_n24672));
AND2X1 exu_U6357(.A(exu_n2016), .B(exu_n7046), .Y(exu_n24671));
AND2X1 exu_U6358(.A(exu_n2017), .B(exu_n7047), .Y(exu_n24678));
AND2X1 exu_U6359(.A(exu_n2018), .B(exu_n7048), .Y(exu_n24677));
AND2X1 exu_U6360(.A(exu_n2019), .B(exu_n7049), .Y(exu_n24684));
AND2X1 exu_U6361(.A(exu_n2020), .B(exu_n7050), .Y(exu_n24683));
AND2X1 exu_U6362(.A(exu_n2021), .B(exu_n7051), .Y(exu_n24690));
AND2X1 exu_U6363(.A(exu_n2022), .B(exu_n7052), .Y(exu_n24689));
AND2X1 exu_U6364(.A(exu_n2023), .B(exu_n7053), .Y(exu_n24696));
AND2X1 exu_U6365(.A(exu_n2024), .B(exu_n7054), .Y(exu_n24695));
AND2X1 exu_U6366(.A(exu_n2025), .B(exu_n7055), .Y(exu_n24702));
AND2X1 exu_U6367(.A(exu_n2026), .B(exu_n7056), .Y(exu_n24701));
AND2X1 exu_U6368(.A(exu_n2029), .B(exu_n7059), .Y(exu_n24714));
AND2X1 exu_U6369(.A(exu_n2030), .B(exu_n7060), .Y(exu_n24713));
AND2X1 exu_U6370(.A(exu_n2031), .B(exu_n7061), .Y(exu_n24720));
AND2X1 exu_U6371(.A(exu_n2032), .B(exu_n7062), .Y(exu_n24719));
AND2X1 exu_U6372(.A(exu_n2033), .B(exu_n7063), .Y(exu_n24726));
AND2X1 exu_U6373(.A(exu_n2034), .B(exu_n7064), .Y(exu_n24725));
AND2X1 exu_U6374(.A(exu_n2035), .B(exu_n7065), .Y(exu_n24732));
AND2X1 exu_U6375(.A(exu_n2036), .B(exu_n7066), .Y(exu_n24731));
AND2X1 exu_U6376(.A(exu_n2037), .B(exu_n7067), .Y(exu_n24738));
AND2X1 exu_U6377(.A(exu_n2038), .B(exu_n7068), .Y(exu_n24737));
AND2X1 exu_U6378(.A(exu_n2039), .B(exu_n7069), .Y(exu_n24744));
AND2X1 exu_U6379(.A(exu_n2040), .B(exu_n7070), .Y(exu_n24743));
AND2X1 exu_U6380(.A(exu_n2041), .B(exu_n7071), .Y(exu_n24750));
AND2X1 exu_U6381(.A(exu_n2042), .B(exu_n7072), .Y(exu_n24749));
AND2X1 exu_U6382(.A(exu_n2043), .B(exu_n7073), .Y(exu_n24756));
AND2X1 exu_U6383(.A(exu_n2044), .B(exu_n7074), .Y(exu_n24755));
AND2X1 exu_U6384(.A(exu_n2045), .B(exu_n7075), .Y(exu_n24762));
AND2X1 exu_U6385(.A(exu_n2046), .B(exu_n7076), .Y(exu_n24761));
AND2X1 exu_U6386(.A(exu_n2047), .B(exu_n7077), .Y(exu_n24768));
AND2X1 exu_U6387(.A(exu_n2048), .B(exu_n7078), .Y(exu_n24767));
AND2X1 exu_U6388(.A(exu_n2051), .B(exu_n7081), .Y(exu_n24780));
AND2X1 exu_U6389(.A(exu_n2052), .B(exu_n7082), .Y(exu_n24779));
AND2X1 exu_U6390(.A(exu_n2053), .B(exu_n7083), .Y(exu_n24786));
AND2X1 exu_U6391(.A(exu_n2054), .B(exu_n7084), .Y(exu_n24785));
AND2X1 exu_U6392(.A(exu_n2055), .B(exu_n7085), .Y(exu_n24792));
AND2X1 exu_U6393(.A(exu_n2056), .B(exu_n7086), .Y(exu_n24791));
AND2X1 exu_U6394(.A(exu_n2057), .B(exu_n7087), .Y(exu_n24798));
AND2X1 exu_U6395(.A(exu_n2058), .B(exu_n7088), .Y(exu_n24797));
AND2X1 exu_U6396(.A(exu_n2059), .B(exu_n7089), .Y(exu_n24804));
AND2X1 exu_U6397(.A(exu_n2060), .B(exu_n7090), .Y(exu_n24803));
AND2X1 exu_U6398(.A(exu_n2061), .B(exu_n7091), .Y(exu_n24810));
AND2X1 exu_U6399(.A(exu_n2062), .B(exu_n7092), .Y(exu_n24809));
AND2X1 exu_U6400(.A(exu_n2063), .B(exu_n7093), .Y(exu_n24816));
AND2X1 exu_U6401(.A(exu_n2064), .B(exu_n7094), .Y(exu_n24815));
AND2X1 exu_U6402(.A(exu_n2065), .B(exu_n7095), .Y(exu_n24822));
AND2X1 exu_U6403(.A(exu_n2066), .B(exu_n7096), .Y(exu_n24821));
AND2X1 exu_U6404(.A(exu_n2067), .B(exu_n7097), .Y(exu_n24828));
AND2X1 exu_U6405(.A(exu_n2068), .B(exu_n7098), .Y(exu_n24827));
AND2X1 exu_U6406(.A(exu_n2069), .B(exu_n7099), .Y(exu_n24834));
AND2X1 exu_U6407(.A(exu_n2070), .B(exu_n7100), .Y(exu_n24833));
AND2X1 exu_U6408(.A(exu_n2073), .B(exu_n7103), .Y(exu_n24846));
AND2X1 exu_U6409(.A(exu_n2074), .B(exu_n7104), .Y(exu_n24845));
AND2X1 exu_U6410(.A(exu_n2075), .B(exu_n7105), .Y(exu_n24852));
AND2X1 exu_U6411(.A(exu_n2076), .B(exu_n7106), .Y(exu_n24851));
AND2X1 exu_U6412(.A(exu_n2077), .B(exu_n7107), .Y(exu_n24858));
AND2X1 exu_U6413(.A(exu_n2078), .B(exu_n7108), .Y(exu_n24857));
AND2X1 exu_U6414(.A(exu_n2079), .B(exu_n7109), .Y(exu_n24864));
AND2X1 exu_U6415(.A(exu_n2080), .B(exu_n7110), .Y(exu_n24863));
AND2X1 exu_U6416(.A(exu_n2081), .B(exu_n7111), .Y(exu_n24870));
AND2X1 exu_U6417(.A(exu_n2082), .B(exu_n7112), .Y(exu_n24869));
AND2X1 exu_U6418(.A(exu_n2083), .B(exu_n7113), .Y(exu_n24876));
AND2X1 exu_U6419(.A(exu_n2084), .B(exu_n7114), .Y(exu_n24875));
AND2X1 exu_U6420(.A(exu_n2085), .B(exu_n7115), .Y(exu_n24882));
AND2X1 exu_U6421(.A(exu_n2086), .B(exu_n7116), .Y(exu_n24881));
AND2X1 exu_U6422(.A(exu_n2087), .B(exu_n7117), .Y(exu_n24888));
AND2X1 exu_U6423(.A(exu_n2088), .B(exu_n7118), .Y(exu_n24887));
AND2X1 exu_U6424(.A(exu_n2089), .B(exu_n7119), .Y(exu_n24894));
AND2X1 exu_U6425(.A(exu_n2090), .B(exu_n7120), .Y(exu_n24893));
AND2X1 exu_U6426(.A(exu_n2091), .B(exu_n7121), .Y(exu_n24900));
AND2X1 exu_U6427(.A(exu_n2092), .B(exu_n7122), .Y(exu_n24899));
AND2X1 exu_U6428(.A(exu_n2095), .B(exu_n7125), .Y(exu_n24912));
AND2X1 exu_U6429(.A(exu_n2096), .B(exu_n7126), .Y(exu_n24911));
AND2X1 exu_U6430(.A(exu_n2097), .B(exu_n7127), .Y(exu_n24918));
AND2X1 exu_U6431(.A(exu_n2098), .B(exu_n7128), .Y(exu_n24917));
AND2X1 exu_U6432(.A(exu_n2099), .B(exu_n7129), .Y(exu_n24924));
AND2X1 exu_U6433(.A(exu_n2100), .B(exu_n7130), .Y(exu_n24923));
AND2X1 exu_U6434(.A(exu_n2101), .B(exu_n7131), .Y(exu_n24930));
AND2X1 exu_U6435(.A(exu_n2102), .B(exu_n7132), .Y(exu_n24929));
AND2X1 exu_U6436(.A(exu_n2103), .B(exu_n7133), .Y(exu_n24936));
AND2X1 exu_U6437(.A(exu_n2104), .B(exu_n7134), .Y(exu_n24935));
AND2X1 exu_U6438(.A(exu_n2105), .B(exu_n7135), .Y(exu_n24942));
AND2X1 exu_U6439(.A(exu_n2106), .B(exu_n7136), .Y(exu_n24941));
AND2X1 exu_U6440(.A(exu_n2107), .B(exu_n7137), .Y(exu_n24948));
AND2X1 exu_U6441(.A(exu_n2108), .B(exu_n7138), .Y(exu_n24947));
AND2X1 exu_U6442(.A(exu_n2109), .B(exu_n7139), .Y(exu_n24954));
AND2X1 exu_U6443(.A(exu_n2110), .B(exu_n7140), .Y(exu_n24953));
AND2X1 exu_U6444(.A(exu_n2111), .B(exu_n7141), .Y(exu_n24960));
AND2X1 exu_U6445(.A(exu_n2112), .B(exu_n7142), .Y(exu_n24959));
AND2X1 exu_U6446(.A(exu_n2113), .B(exu_n7143), .Y(exu_n24966));
AND2X1 exu_U6447(.A(exu_n2114), .B(exu_n7144), .Y(exu_n24965));
AND2X1 exu_U6448(.A(exu_n1989), .B(exu_n7019), .Y(exu_n24594));
AND2X1 exu_U6449(.A(exu_n1990), .B(exu_n7020), .Y(exu_n24593));
AND2X1 exu_U6450(.A(exu_n1991), .B(exu_n7021), .Y(exu_n24600));
AND2X1 exu_U6451(.A(exu_n1992), .B(exu_n7022), .Y(exu_n24599));
AND2X1 exu_U6452(.A(exu_n1993), .B(exu_n7023), .Y(exu_n24606));
AND2X1 exu_U6453(.A(exu_n1994), .B(exu_n7024), .Y(exu_n24605));
INVX1 exu_U6454(.A(exu_n16081), .Y(exu_n16075));
AND2X1 exu_U6455(.A(exu_n1995), .B(exu_n7025), .Y(exu_n24612));
AND2X1 exu_U6456(.A(exu_n1996), .B(exu_n7026), .Y(exu_n24611));
AND2X1 exu_U6457(.A(exu_n2005), .B(exu_n7035), .Y(exu_n24642));
AND2X1 exu_U6458(.A(exu_n2006), .B(exu_n7036), .Y(exu_n24641));
AND2X1 exu_U6459(.A(exu_n2027), .B(exu_n7057), .Y(exu_n24708));
AND2X1 exu_U6460(.A(exu_n2028), .B(exu_n7058), .Y(exu_n24707));
AND2X1 exu_U6461(.A(exu_n2049), .B(exu_n7079), .Y(exu_n24774));
AND2X1 exu_U6462(.A(exu_n2050), .B(exu_n7080), .Y(exu_n24773));
INVX1 exu_U6463(.A(exu_n16080), .Y(exu_n16079));
AND2X1 exu_U6464(.A(exu_n2071), .B(exu_n7101), .Y(exu_n24840));
AND2X1 exu_U6465(.A(exu_n2072), .B(exu_n7102), .Y(exu_n24839));
INVX1 exu_U6466(.A(exu_n16080), .Y(exu_n16078));
AND2X1 exu_U6467(.A(exu_n2093), .B(exu_n7123), .Y(exu_n24906));
AND2X1 exu_U6468(.A(exu_n2094), .B(exu_n7124), .Y(exu_n24905));
INVX1 exu_U6469(.A(exu_n16080), .Y(exu_n16077));
AND2X1 exu_U6470(.A(exu_n2115), .B(exu_n7145), .Y(exu_n24972));
AND2X1 exu_U6471(.A(exu_n2116), .B(exu_n7146), .Y(exu_n24971));
INVX1 exu_U6472(.A(exu_n16081), .Y(exu_n16076));
INVX1 exu_U6473(.A(exu_n16088), .Y(exu_n16082));
INVX1 exu_U6474(.A(exu_n16087), .Y(exu_n16086));
INVX1 exu_U6475(.A(exu_n16087), .Y(exu_n16085));
INVX1 exu_U6476(.A(exu_n16087), .Y(exu_n16084));
INVX1 exu_U6477(.A(exu_n16088), .Y(exu_n16083));
INVX1 exu_U6478(.A(exu_n16095), .Y(exu_n16089));
INVX1 exu_U6479(.A(exu_n16094), .Y(exu_n16093));
INVX1 exu_U6480(.A(exu_n16094), .Y(exu_n16092));
INVX1 exu_U6481(.A(exu_n16094), .Y(exu_n16091));
INVX1 exu_U6482(.A(exu_n16095), .Y(exu_n16090));
INVX1 exu_U6483(.A(exu_n16102), .Y(exu_n16096));
INVX1 exu_U6484(.A(exu_n16101), .Y(exu_n16100));
INVX1 exu_U6485(.A(exu_n16101), .Y(exu_n16099));
INVX1 exu_U6486(.A(exu_n16101), .Y(exu_n16098));
INVX1 exu_U6487(.A(exu_n16102), .Y(exu_n16097));
AND2X1 exu_U6488(.A(exu_n748), .B(exu_n5509), .Y(div_xin[62]));
AND2X1 exu_U6489(.A(exu_n750), .B(exu_n5513), .Y(div_xin[61]));
AND2X1 exu_U6490(.A(exu_n751), .B(exu_n5515), .Y(div_xin[60]));
AND2X1 exu_U6491(.A(exu_n752), .B(exu_n5517), .Y(div_xin[59]));
AND2X1 exu_U6492(.A(exu_n753), .B(exu_n5519), .Y(div_xin[58]));
AND2X1 exu_U6493(.A(exu_n754), .B(exu_n5521), .Y(div_xin[57]));
AND2X1 exu_U6494(.A(exu_n755), .B(exu_n5523), .Y(div_xin[56]));
AND2X1 exu_U6495(.A(exu_n756), .B(exu_n5525), .Y(div_xin[55]));
AND2X1 exu_U6496(.A(exu_n757), .B(exu_n5527), .Y(div_xin[54]));
AND2X1 exu_U6497(.A(exu_n758), .B(exu_n5529), .Y(div_xin[53]));
AND2X1 exu_U6498(.A(exu_n759), .B(exu_n5530), .Y(div_xin[52]));
AND2X1 exu_U6499(.A(exu_n761), .B(exu_n5530), .Y(div_xin[51]));
AND2X1 exu_U6500(.A(exu_n762), .B(exu_n5530), .Y(div_xin[50]));
AND2X1 exu_U6501(.A(exu_n763), .B(exu_n5530), .Y(div_xin[49]));
AND2X1 exu_U6502(.A(exu_n764), .B(exu_n5530), .Y(div_xin[48]));
AND2X1 exu_U6503(.A(exu_n765), .B(exu_n5530), .Y(div_xin[47]));
AND2X1 exu_U6504(.A(exu_n766), .B(exu_n5530), .Y(div_xin[46]));
AND2X1 exu_U6505(.A(exu_n767), .B(exu_n5530), .Y(div_xin[45]));
AND2X1 exu_U6506(.A(exu_n768), .B(exu_n5530), .Y(div_xin[44]));
AND2X1 exu_U6507(.A(exu_n769), .B(exu_n5530), .Y(div_xin[43]));
AND2X1 exu_U6508(.A(exu_n770), .B(exu_n5530), .Y(div_xin[42]));
AND2X1 exu_U6509(.A(exu_n740), .B(exu_n5497), .Y(div_xin[41]));
AND2X1 exu_U6510(.A(exu_n741), .B(exu_n5497), .Y(div_xin[40]));
AND2X1 exu_U6511(.A(exu_n742), .B(exu_n5499), .Y(div_xin[39]));
AND2X1 exu_U6512(.A(exu_n743), .B(exu_n5501), .Y(div_xin[38]));
AND2X1 exu_U6513(.A(exu_n744), .B(exu_n5503), .Y(div_xin[37]));
AND2X1 exu_U6514(.A(exu_n745), .B(exu_n5505), .Y(div_xin[36]));
AND2X1 exu_U6515(.A(exu_n746), .B(exu_n5507), .Y(div_xin[35]));
AND2X1 exu_U6516(.A(exu_n749), .B(exu_n5511), .Y(div_xin[34]));
AND2X1 exu_U6517(.A(exu_n760), .B(exu_n5530), .Y(div_xin[33]));
AND2X1 exu_U6518(.A(exu_n771), .B(exu_n5530), .Y(div_xin[32]));
AND2X1 exu_U6519(.A(div_input_data_e[95]), .B(exu_n16613), .Y(div_xin[31]));
AND2X1 exu_U6520(.A(div_input_data_e[94]), .B(exu_n16613), .Y(div_xin[30]));
AND2X1 exu_U6521(.A(div_input_data_e[93]), .B(exu_n16613), .Y(div_xin[29]));
AND2X1 exu_U6522(.A(div_input_data_e[92]), .B(exu_n16613), .Y(div_xin[28]));
AND2X1 exu_U6523(.A(div_input_data_e[91]), .B(exu_n16613), .Y(div_xin[27]));
AND2X1 exu_U6524(.A(div_input_data_e[90]), .B(exu_n16613), .Y(div_xin[26]));
AND2X1 exu_U6525(.A(div_input_data_e[89]), .B(exu_n16613), .Y(div_xin[25]));
AND2X1 exu_U6526(.A(div_input_data_e[88]), .B(exu_n16613), .Y(div_xin[24]));
AND2X1 exu_U6527(.A(div_input_data_e[87]), .B(exu_n16613), .Y(div_xin[23]));
AND2X1 exu_U6528(.A(div_input_data_e[86]), .B(exu_n16613), .Y(div_xin[22]));
AND2X1 exu_U6529(.A(div_input_data_e[85]), .B(exu_n16613), .Y(div_xin[21]));
AND2X1 exu_U6530(.A(div_input_data_e[84]), .B(exu_n16613), .Y(div_xin[20]));
AND2X1 exu_U6531(.A(div_input_data_e[83]), .B(exu_n16613), .Y(div_xin[19]));
AND2X1 exu_U6532(.A(div_input_data_e[82]), .B(exu_n16613), .Y(div_xin[18]));
AND2X1 exu_U6533(.A(div_input_data_e[81]), .B(exu_n16613), .Y(div_xin[17]));
AND2X1 exu_U6534(.A(div_input_data_e[80]), .B(exu_n16613), .Y(div_xin[16]));
AND2X1 exu_U6535(.A(div_input_data_e[79]), .B(exu_n16613), .Y(div_xin[15]));
AND2X1 exu_U6536(.A(div_input_data_e[78]), .B(exu_n16613), .Y(div_xin[14]));
AND2X1 exu_U6537(.A(div_input_data_e[77]), .B(exu_n16613), .Y(div_xin[13]));
AND2X1 exu_U6538(.A(div_input_data_e[76]), .B(exu_n16613), .Y(div_xin[12]));
AND2X1 exu_U6539(.A(div_input_data_e[75]), .B(exu_n16613), .Y(div_xin[11]));
AND2X1 exu_U6540(.A(div_input_data_e[74]), .B(exu_n16613), .Y(div_xin[10]));
AND2X1 exu_U6541(.A(div_input_data_e[73]), .B(exu_n16613), .Y(div_xin[9]));
AND2X1 exu_U6542(.A(div_input_data_e[72]), .B(exu_n16613), .Y(div_xin[8]));
AND2X1 exu_U6543(.A(div_input_data_e[71]), .B(exu_n16613), .Y(div_xin[7]));
INVX1 exu_U6544(.A(exu_n16109), .Y(exu_n16103));
AND2X1 exu_U6545(.A(div_input_data_e[70]), .B(exu_n16613), .Y(div_xin[6]));
AND2X1 exu_U6546(.A(div_input_data_e[69]), .B(exu_n16613), .Y(div_xin[5]));
AND2X1 exu_U6547(.A(div_input_data_e[68]), .B(exu_n16613), .Y(div_xin[4]));
AND2X1 exu_U6548(.A(div_input_data_e[67]), .B(exu_n16613), .Y(div_xin[3]));
INVX1 exu_U6549(.A(exu_n16108), .Y(exu_n16107));
AND2X1 exu_U6550(.A(div_input_data_e[66]), .B(exu_n16613), .Y(div_xin[2]));
INVX1 exu_U6551(.A(exu_n16108), .Y(exu_n16106));
AND2X1 exu_U6552(.A(div_input_data_e[65]), .B(exu_n16613), .Y(div_xin[1]));
INVX1 exu_U6553(.A(exu_n16108), .Y(exu_n16105));
AND2X1 exu_U6554(.A(div_input_data_e[64]), .B(exu_n16613), .Y(div_xin[0]));
INVX1 exu_U6555(.A(exu_n16109), .Y(exu_n16104));
INVX1 exu_U6556(.A(exu_n16116), .Y(exu_n16110));
INVX1 exu_U6557(.A(exu_n16115), .Y(exu_n16114));
INVX1 exu_U6558(.A(exu_n16115), .Y(exu_n16113));
INVX1 exu_U6559(.A(exu_n16115), .Y(exu_n16112));
INVX1 exu_U6560(.A(exu_n16116), .Y(exu_n16111));
AND2X1 exu_U6561(.A(rml_cwp_swap_slot0_state[1]), .B(exu_n9120), .Y(rml_cwp_swap_slot0_state_valid[1]));
AND2X1 exu_U6562(.A(rml_cwp_swap_thr[0]), .B(rml_cwp_n45), .Y(rml_cwp_swap_next_state[0]));
AND2X1 exu_U6563(.A(exu_n15026), .B(rml_cwp_N99), .Y(rml_cwp_n45));
AND2X1 exu_U6564(.A(exu_n15026), .B(exu_n9121), .Y(rml_cwp_swap_keep_state[0]));
AND2X1 exu_U6565(.A(exu_n15960), .B(rml_cwp_n73), .Y(rml_cwp_swap_sel_tlu[0]));
AND2X1 exu_U6566(.A(rml_cwp_cwpccr_update_w), .B(exu_n15410), .Y(rml_cwp_n73));
AND2X1 exu_U6567(.A(exu_n4148), .B(rml_cwp_cwpccr_update_w), .Y(rml_cwp_valid_tlu_swap_w));
INVX1 exu_U6568(.A(rml_cwp_swap_sel_tlu[0]), .Y(exu_n16393));
INVX1 exu_U6569(.A(se), .Y(ecl_mdqctl_mul_data_dff_n1));
OR2X1 exu_U6570(.A(ecl_div_zero_m), .B(exu_n15363), .Y(ecl_mdqctl_n54));
INVX1 exu_U6571(.A(ecl_mdqctl_new_div_vld), .Y(exu_n16387));
AND2X1 exu_U6572(.A(div_input_data_e[95]), .B(exu_n15814), .Y(ecl_divcntl_inputs_neg_d));
INVX1 exu_U6573(.A(ecl_divcntl_inputs_neg_dff_n6), .Y(exu_n16370));
OR2X1 exu_U6574(.A(exu_n16505), .B(exu_n15398), .Y(ecl_divcntl_n26));
INVX1 exu_U6575(.A(ecl_divcntl_div_state[4]), .Y(exu_n16504));
INVX1 exu_U6576(.A(ecl_divcntl_div_state[3]), .Y(exu_n16503));
OR2X1 exu_U6577(.A(exu_n15471), .B(exu_n14749), .Y(ecl_divcntl_n33));
INVX1 exu_U6578(.A(se), .Y(ecl_divcntl_divstate_dff_n1));
AND2X1 exu_U6579(.A(exu_n4528), .B(ecl_bypass_m), .Y(ecl_writeback_valid_m));
INVX1 exu_U6580(.A(se), .Y(rml_oddwin_dff_n1));
AND2X1 exu_U6581(.A(exu_n10942), .B(exu_n5475), .Y(div_din[94]));
AND2X1 exu_U6582(.A(exu_n10944), .B(exu_n5477), .Y(div_din[93]));
AND2X1 exu_U6583(.A(exu_n10948), .B(exu_n5481), .Y(div_din[92]));
AND2X1 exu_U6584(.A(exu_n10950), .B(exu_n5483), .Y(div_din[91]));
AND2X1 exu_U6585(.A(exu_n10952), .B(exu_n5485), .Y(div_din[90]));
AND2X1 exu_U6586(.A(exu_n10954), .B(exu_n5487), .Y(div_din[89]));
AND2X1 exu_U6587(.A(exu_n10956), .B(exu_n5489), .Y(div_din[88]));
AND2X1 exu_U6588(.A(exu_n10958), .B(exu_n5491), .Y(div_din[87]));
AND2X1 exu_U6589(.A(exu_n10960), .B(exu_n5493), .Y(div_din[86]));
AND2X1 exu_U6590(.A(exu_n10962), .B(exu_n5494), .Y(div_din[85]));
AND2X1 exu_U6591(.A(exu_n10964), .B(exu_n5494), .Y(div_din[84]));
AND2X1 exu_U6592(.A(exu_n10966), .B(exu_n5494), .Y(div_din[83]));
AND2X1 exu_U6593(.A(exu_n10970), .B(exu_n5494), .Y(div_din[82]));
AND2X1 exu_U6594(.A(exu_n10972), .B(exu_n5494), .Y(div_din[81]));
AND2X1 exu_U6595(.A(exu_n10974), .B(exu_n5494), .Y(div_din[80]));
AND2X1 exu_U6596(.A(exu_n10976), .B(exu_n5494), .Y(div_din[79]));
AND2X1 exu_U6597(.A(exu_n10978), .B(exu_n5494), .Y(div_din[78]));
AND2X1 exu_U6598(.A(exu_n10980), .B(exu_n5494), .Y(div_din[77]));
AND2X1 exu_U6599(.A(exu_n10982), .B(exu_n5494), .Y(div_din[76]));
AND2X1 exu_U6600(.A(exu_n10984), .B(exu_n5494), .Y(div_din[75]));
AND2X1 exu_U6601(.A(exu_n10986), .B(exu_n5494), .Y(div_din[74]));
AND2X1 exu_U6602(.A(exu_n10988), .B(exu_n5494), .Y(div_din[73]));
AND2X1 exu_U6603(.A(exu_n10928), .B(exu_n5463), .Y(div_din[72]));
AND2X1 exu_U6604(.A(exu_n10930), .B(exu_n5463), .Y(div_din[71]));
AND2X1 exu_U6605(.A(exu_n10932), .B(exu_n5465), .Y(div_din[70]));
AND2X1 exu_U6606(.A(exu_n10934), .B(exu_n5467), .Y(div_din[69]));
AND2X1 exu_U6607(.A(exu_n10936), .B(exu_n5469), .Y(div_din[68]));
AND2X1 exu_U6608(.A(exu_n10938), .B(exu_n5471), .Y(div_din[67]));
AND2X1 exu_U6609(.A(exu_n10940), .B(exu_n5473), .Y(div_din[66]));
AND2X1 exu_U6610(.A(exu_n10946), .B(exu_n5479), .Y(div_din[65]));
AND2X1 exu_U6611(.A(exu_n10968), .B(exu_n5494), .Y(div_din[64]));
OR2X1 exu_U6612(.A(exu_n28720), .B(exu_n16248), .Y(div_out64[63]));
AND2X1 exu_U6613(.A(exu_n10990), .B(exu_n5495), .Y(div_din[63]));
OR2X1 exu_U6614(.A(exu_n28721), .B(exu_n16248), .Y(div_out64[62]));
AND2X1 exu_U6615(.A(exu_n10880), .B(exu_n5438), .Y(div_dividend[62]));
OR2X1 exu_U6616(.A(exu_n28722), .B(ecl_div_sel_neg32), .Y(div_out64[61]));
AND2X1 exu_U6617(.A(exu_n10884), .B(exu_n5440), .Y(div_dividend[61]));
OR2X1 exu_U6618(.A(exu_n28723), .B(ecl_div_sel_neg32), .Y(div_out64[60]));
AND2X1 exu_U6619(.A(exu_n10886), .B(exu_n5441), .Y(div_dividend[60]));
OR2X1 exu_U6620(.A(exu_n28730), .B(exu_n16248), .Y(div_out64[59]));
AND2X1 exu_U6621(.A(exu_n10888), .B(exu_n5442), .Y(div_dividend[59]));
OR2X1 exu_U6622(.A(exu_n28731), .B(ecl_div_sel_neg32), .Y(div_out64[58]));
AND2X1 exu_U6623(.A(exu_n10890), .B(exu_n5443), .Y(div_dividend[58]));
OR2X1 exu_U6624(.A(exu_n28732), .B(ecl_div_sel_neg32), .Y(div_out64[57]));
AND2X1 exu_U6625(.A(exu_n10892), .B(exu_n5444), .Y(div_dividend[57]));
OR2X1 exu_U6626(.A(exu_n28733), .B(exu_n16248), .Y(div_out64[56]));
AND2X1 exu_U6627(.A(exu_n10894), .B(exu_n5445), .Y(div_dividend[56]));
OR2X1 exu_U6628(.A(exu_n28734), .B(exu_n16248), .Y(div_out64[55]));
AND2X1 exu_U6629(.A(exu_n10896), .B(exu_n5446), .Y(div_dividend[55]));
OR2X1 exu_U6630(.A(exu_n28735), .B(exu_n16248), .Y(div_out64[54]));
AND2X1 exu_U6631(.A(exu_n10898), .B(exu_n5447), .Y(div_dividend[54]));
OR2X1 exu_U6632(.A(exu_n28736), .B(ecl_div_sel_neg32), .Y(div_out64[53]));
AND2X1 exu_U6633(.A(exu_n10900), .B(exu_n5448), .Y(div_dividend[53]));
OR2X1 exu_U6634(.A(exu_n28737), .B(ecl_div_sel_neg32), .Y(div_out64[52]));
AND2X1 exu_U6635(.A(exu_n10902), .B(exu_n5449), .Y(div_dividend[52]));
OR2X1 exu_U6636(.A(exu_n28738), .B(ecl_div_sel_neg32), .Y(div_out64[51]));
AND2X1 exu_U6637(.A(exu_n10906), .B(exu_n5451), .Y(div_dividend[51]));
OR2X1 exu_U6638(.A(exu_n28739), .B(exu_n16248), .Y(div_out64[50]));
AND2X1 exu_U6639(.A(exu_n10908), .B(exu_n5452), .Y(div_dividend[50]));
OR2X1 exu_U6640(.A(exu_n28746), .B(ecl_div_sel_neg32), .Y(div_out64[49]));
AND2X1 exu_U6641(.A(exu_n10910), .B(exu_n5453), .Y(div_dividend[49]));
OR2X1 exu_U6642(.A(exu_n28747), .B(exu_n16248), .Y(div_out64[48]));
AND2X1 exu_U6643(.A(exu_n10912), .B(exu_n5454), .Y(div_dividend[48]));
OR2X1 exu_U6644(.A(exu_n28748), .B(ecl_div_sel_neg32), .Y(div_out64[47]));
AND2X1 exu_U6645(.A(exu_n10914), .B(exu_n5455), .Y(div_dividend[47]));
OR2X1 exu_U6646(.A(exu_n28749), .B(ecl_div_sel_neg32), .Y(div_out64[46]));
AND2X1 exu_U6647(.A(exu_n10916), .B(exu_n5456), .Y(div_dividend[46]));
OR2X1 exu_U6648(.A(exu_n28750), .B(ecl_div_sel_neg32), .Y(div_out64[45]));
AND2X1 exu_U6649(.A(exu_n10918), .B(exu_n5457), .Y(div_dividend[45]));
OR2X1 exu_U6650(.A(exu_n28751), .B(ecl_div_sel_neg32), .Y(div_out64[44]));
AND2X1 exu_U6651(.A(exu_n10920), .B(exu_n5458), .Y(div_dividend[44]));
OR2X1 exu_U6652(.A(exu_n28752), .B(ecl_div_sel_neg32), .Y(div_out64[43]));
AND2X1 exu_U6653(.A(exu_n10922), .B(exu_n5459), .Y(div_dividend[43]));
OR2X1 exu_U6654(.A(exu_n28753), .B(ecl_div_sel_neg32), .Y(div_out64[42]));
AND2X1 exu_U6655(.A(exu_n10924), .B(exu_n5460), .Y(div_dividend[42]));
OR2X1 exu_U6656(.A(exu_n28754), .B(ecl_div_sel_neg32), .Y(div_out64[41]));
AND2X1 exu_U6657(.A(exu_n10866), .B(exu_n5430), .Y(div_dividend[41]));
OR2X1 exu_U6658(.A(exu_n28755), .B(ecl_div_sel_neg32), .Y(div_out64[40]));
AND2X1 exu_U6659(.A(exu_n10868), .B(exu_n5431), .Y(div_dividend[40]));
OR2X1 exu_U6660(.A(exu_n28762), .B(ecl_div_sel_neg32), .Y(div_out64[39]));
AND2X1 exu_U6661(.A(exu_n10870), .B(exu_n5432), .Y(div_dividend[39]));
OR2X1 exu_U6662(.A(exu_n28763), .B(ecl_div_sel_neg32), .Y(div_out64[38]));
AND2X1 exu_U6663(.A(exu_n10872), .B(exu_n5433), .Y(div_dividend[38]));
OR2X1 exu_U6664(.A(exu_n28764), .B(exu_n16248), .Y(div_out64[37]));
AND2X1 exu_U6665(.A(exu_n10874), .B(exu_n5434), .Y(div_dividend[37]));
OR2X1 exu_U6666(.A(exu_n28765), .B(ecl_div_sel_neg32), .Y(div_out64[36]));
AND2X1 exu_U6667(.A(exu_n10876), .B(exu_n5435), .Y(div_dividend[36]));
OR2X1 exu_U6668(.A(exu_n28766), .B(exu_n16248), .Y(div_out64[35]));
AND2X1 exu_U6669(.A(exu_n10878), .B(exu_n5436), .Y(div_dividend[35]));
OR2X1 exu_U6670(.A(exu_n28767), .B(ecl_div_sel_neg32), .Y(div_out64[34]));
AND2X1 exu_U6671(.A(exu_n10882), .B(exu_n5439), .Y(div_dividend[34]));
OR2X1 exu_U6672(.A(exu_n28768), .B(exu_n16248), .Y(div_out64[33]));
AND2X1 exu_U6673(.A(exu_n10904), .B(exu_n5450), .Y(div_dividend[33]));
OR2X1 exu_U6674(.A(exu_n28769), .B(ecl_div_sel_neg32), .Y(div_out64[32]));
AND2X1 exu_U6675(.A(exu_n10926), .B(exu_n5461), .Y(div_dividend[32]));
OR2X1 exu_U6676(.A(exu_n13303), .B(ecl_div_sel_neg32), .Y(div_out64[31]));
OR2X1 exu_U6677(.A(exu_n13304), .B(exu_n14611), .Y(div_out64[30]));
OR2X1 exu_U6678(.A(exu_n13306), .B(exu_n14613), .Y(div_out64[29]));
OR2X1 exu_U6679(.A(exu_n13307), .B(exu_n14614), .Y(div_out64[28]));
OR2X1 exu_U6680(.A(exu_n13308), .B(exu_n14615), .Y(div_out64[27]));
OR2X1 exu_U6681(.A(exu_n13309), .B(exu_n14616), .Y(div_out64[26]));
OR2X1 exu_U6682(.A(exu_n13310), .B(exu_n14617), .Y(div_out64[25]));
OR2X1 exu_U6683(.A(exu_n13311), .B(exu_n14618), .Y(div_out64[24]));
OR2X1 exu_U6684(.A(exu_n13312), .B(exu_n14619), .Y(div_out64[23]));
OR2X1 exu_U6685(.A(exu_n13313), .B(exu_n14620), .Y(div_out64[22]));
OR2X1 exu_U6686(.A(exu_n13314), .B(exu_n14621), .Y(div_out64[21]));
OR2X1 exu_U6687(.A(exu_n13315), .B(exu_n14622), .Y(div_out64[20]));
OR2X1 exu_U6688(.A(exu_n13317), .B(exu_n14624), .Y(div_out64[19]));
OR2X1 exu_U6689(.A(exu_n13318), .B(exu_n14625), .Y(div_out64[18]));
OR2X1 exu_U6690(.A(exu_n13319), .B(exu_n14626), .Y(div_out64[17]));
OR2X1 exu_U6691(.A(exu_n13320), .B(exu_n14627), .Y(div_out64[16]));
OR2X1 exu_U6692(.A(exu_n13321), .B(exu_n14628), .Y(div_out64[15]));
OR2X1 exu_U6693(.A(exu_n13322), .B(exu_n14629), .Y(div_out64[14]));
OR2X1 exu_U6694(.A(exu_n13323), .B(exu_n14630), .Y(div_out64[13]));
OR2X1 exu_U6695(.A(exu_n13324), .B(exu_n14631), .Y(div_out64[12]));
OR2X1 exu_U6696(.A(exu_n13325), .B(exu_n14632), .Y(div_out64[11]));
OR2X1 exu_U6697(.A(exu_n13326), .B(exu_n14633), .Y(div_out64[10]));
INVX1 exu_U6698(.A(exu_n16129), .Y(exu_n16119));
OR2X1 exu_U6699(.A(exu_n13296), .B(exu_n14604), .Y(div_out64[9]));
INVX1 exu_U6700(.A(exu_n16129), .Y(exu_n16118));
OR2X1 exu_U6701(.A(exu_n13297), .B(exu_n14605), .Y(div_out64[8]));
OR2X1 exu_U6702(.A(exu_n13298), .B(exu_n14606), .Y(div_out64[7]));
INVX1 exu_U6703(.A(exu_n16130), .Y(exu_n16117));
INVX1 exu_U6704(.A(div_d_dff_n1), .Y(exu_n16130));
OR2X1 exu_U6705(.A(exu_n13299), .B(exu_n14607), .Y(div_out64[6]));
INVX1 exu_U6706(.A(exu_n16127), .Y(exu_n16126));
OR2X1 exu_U6707(.A(exu_n13300), .B(exu_n14608), .Y(div_out64[5]));
INVX1 exu_U6708(.A(exu_n16127), .Y(exu_n16125));
OR2X1 exu_U6709(.A(exu_n13301), .B(exu_n14609), .Y(div_out64[4]));
INVX1 exu_U6710(.A(exu_n16127), .Y(exu_n16124));
OR2X1 exu_U6711(.A(exu_n13302), .B(exu_n14610), .Y(div_out64[3]));
INVX1 exu_U6712(.A(exu_n16128), .Y(exu_n16123));
OR2X1 exu_U6713(.A(exu_n13305), .B(exu_n14612), .Y(div_out64[2]));
INVX1 exu_U6714(.A(exu_n16128), .Y(exu_n16122));
OR2X1 exu_U6715(.A(exu_n13316), .B(exu_n14623), .Y(div_out64[1]));
INVX1 exu_U6716(.A(exu_n16128), .Y(exu_n16121));
OR2X1 exu_U6717(.A(exu_n13327), .B(exu_n14634), .Y(div_out64[0]));
INVX1 exu_U6718(.A(exu_n16129), .Y(exu_n16120));
AND2X1 exu_U6719(.A(exu_n11929), .B(exu_n9669), .Y(ecl_early1_ttype_e[5]));
AND2X1 exu_U6720(.A(rml_ecl_wtype_e[2]), .B(exu_n15030), .Y(ecl_early1_ttype_e[4]));
AND2X1 exu_U6721(.A(exu_n11932), .B(exu_n9670), .Y(ecl_early1_ttype_e[3]));
AND2X1 exu_U6722(.A(exu_n11934), .B(exu_n9671), .Y(ecl_early1_ttype_e[2]));
OR2X1 exu_U6723(.A(exu_n15239), .B(exu_n15362), .Y(ecl_early1_ttype_e[1]));
INVX1 exu_U6724(.A(se), .Y(ecl_ttype_e2m_n1));
INVX1 exu_U6725(.A(se), .Y(ecl_dff_aluop_d2e_n1));
INVX1 exu_U6726(.A(se), .Y(ecl_dff_ld_tid_m2g_n1));
INVX1 exu_U6727(.A(se), .Y(ecl_dff_rs1_s2d_n1));
INVX1 exu_U6728(.A(se), .Y(ecc_rs1_err_e2m_n1));
INVX1 exu_U6729(.A(se), .Y(ecc_rs1_ecc_d2e_n1));
AND2X1 exu_U6730(.A(exu_n800), .B(exu_n5561), .Y(exu_n20519));
AND2X1 exu_U6731(.A(exu_n801), .B(exu_n5562), .Y(exu_n20518));
AND2X1 exu_U6732(.A(exu_n802), .B(exu_n5563), .Y(exu_n20525));
AND2X1 exu_U6733(.A(exu_n803), .B(exu_n5564), .Y(exu_n20524));
AND2X1 exu_U6734(.A(exu_n806), .B(exu_n5567), .Y(exu_n20537));
AND2X1 exu_U6735(.A(exu_n807), .B(exu_n5568), .Y(exu_n20536));
AND2X1 exu_U6736(.A(exu_n808), .B(exu_n5569), .Y(exu_n20543));
AND2X1 exu_U6737(.A(exu_n809), .B(exu_n5570), .Y(exu_n20542));
AND2X1 exu_U6738(.A(exu_n810), .B(exu_n5571), .Y(exu_n20549));
AND2X1 exu_U6739(.A(exu_n811), .B(exu_n5572), .Y(exu_n20548));
AND2X1 exu_U6740(.A(exu_n812), .B(exu_n5573), .Y(exu_n20555));
AND2X1 exu_U6741(.A(exu_n813), .B(exu_n5574), .Y(exu_n20554));
AND2X1 exu_U6742(.A(exu_n814), .B(exu_n5575), .Y(exu_n20561));
AND2X1 exu_U6743(.A(exu_n815), .B(exu_n5576), .Y(exu_n20560));
AND2X1 exu_U6744(.A(exu_n816), .B(exu_n5577), .Y(exu_n20567));
AND2X1 exu_U6745(.A(exu_n817), .B(exu_n5578), .Y(exu_n20566));
AND2X1 exu_U6746(.A(exu_n818), .B(exu_n5579), .Y(exu_n20573));
AND2X1 exu_U6747(.A(exu_n819), .B(exu_n5580), .Y(exu_n20572));
AND2X1 exu_U6748(.A(exu_n820), .B(exu_n5581), .Y(exu_n20579));
AND2X1 exu_U6749(.A(exu_n821), .B(exu_n5582), .Y(exu_n20578));
AND2X1 exu_U6750(.A(exu_n822), .B(exu_n5583), .Y(exu_n20585));
AND2X1 exu_U6751(.A(exu_n823), .B(exu_n5584), .Y(exu_n20584));
AND2X1 exu_U6752(.A(exu_n824), .B(exu_n5585), .Y(exu_n20591));
AND2X1 exu_U6753(.A(exu_n825), .B(exu_n5586), .Y(exu_n20590));
AND2X1 exu_U6754(.A(exu_n828), .B(exu_n5589), .Y(exu_n20603));
AND2X1 exu_U6755(.A(exu_n829), .B(exu_n5590), .Y(exu_n20602));
AND2X1 exu_U6756(.A(exu_n830), .B(exu_n5591), .Y(exu_n20609));
AND2X1 exu_U6757(.A(exu_n831), .B(exu_n5592), .Y(exu_n20608));
AND2X1 exu_U6758(.A(exu_n832), .B(exu_n5593), .Y(exu_n20615));
AND2X1 exu_U6759(.A(exu_n833), .B(exu_n5594), .Y(exu_n20614));
AND2X1 exu_U6760(.A(exu_n834), .B(exu_n5595), .Y(exu_n20621));
AND2X1 exu_U6761(.A(exu_n835), .B(exu_n5596), .Y(exu_n20620));
AND2X1 exu_U6762(.A(exu_n836), .B(exu_n5597), .Y(exu_n20627));
AND2X1 exu_U6763(.A(exu_n837), .B(exu_n5598), .Y(exu_n20626));
AND2X1 exu_U6764(.A(exu_n838), .B(exu_n5599), .Y(exu_n20633));
AND2X1 exu_U6765(.A(exu_n839), .B(exu_n5600), .Y(exu_n20632));
AND2X1 exu_U6766(.A(exu_n840), .B(exu_n5601), .Y(exu_n20639));
AND2X1 exu_U6767(.A(exu_n841), .B(exu_n5602), .Y(exu_n20638));
AND2X1 exu_U6768(.A(exu_n842), .B(exu_n5603), .Y(exu_n20645));
AND2X1 exu_U6769(.A(exu_n843), .B(exu_n5604), .Y(exu_n20644));
AND2X1 exu_U6770(.A(exu_n844), .B(exu_n5605), .Y(exu_n20651));
AND2X1 exu_U6771(.A(exu_n845), .B(exu_n5606), .Y(exu_n20650));
AND2X1 exu_U6772(.A(exu_n846), .B(exu_n5607), .Y(exu_n20657));
AND2X1 exu_U6773(.A(exu_n847), .B(exu_n5608), .Y(exu_n20656));
AND2X1 exu_U6774(.A(exu_n786), .B(exu_n5547), .Y(exu_n20477));
AND2X1 exu_U6775(.A(exu_n787), .B(exu_n5548), .Y(exu_n20476));
AND2X1 exu_U6776(.A(exu_n788), .B(exu_n5549), .Y(exu_n20483));
AND2X1 exu_U6777(.A(exu_n789), .B(exu_n5550), .Y(exu_n20482));
AND2X1 exu_U6778(.A(exu_n790), .B(exu_n5551), .Y(exu_n20489));
AND2X1 exu_U6779(.A(exu_n791), .B(exu_n5552), .Y(exu_n20488));
INVX1 exu_U6780(.A(exu_n16134), .Y(exu_n16131));
AND2X1 exu_U6781(.A(exu_n792), .B(exu_n5553), .Y(exu_n20495));
AND2X1 exu_U6782(.A(exu_n793), .B(exu_n5554), .Y(exu_n20494));
AND2X1 exu_U6783(.A(exu_n794), .B(exu_n5555), .Y(exu_n20501));
AND2X1 exu_U6784(.A(exu_n795), .B(exu_n5556), .Y(exu_n20500));
AND2X1 exu_U6785(.A(exu_n796), .B(exu_n5557), .Y(exu_n20507));
AND2X1 exu_U6786(.A(exu_n797), .B(exu_n5558), .Y(exu_n20506));
AND2X1 exu_U6787(.A(exu_n798), .B(exu_n5559), .Y(exu_n20513));
AND2X1 exu_U6788(.A(exu_n799), .B(exu_n5560), .Y(exu_n20512));
AND2X1 exu_U6789(.A(exu_n804), .B(exu_n5565), .Y(exu_n20531));
AND2X1 exu_U6790(.A(exu_n805), .B(exu_n5566), .Y(exu_n20530));
AND2X1 exu_U6791(.A(exu_n826), .B(exu_n5587), .Y(exu_n20597));
AND2X1 exu_U6792(.A(exu_n827), .B(exu_n5588), .Y(exu_n20596));
INVX1 exu_U6793(.A(exu_n16134), .Y(exu_n16133));
AND2X1 exu_U6794(.A(exu_n848), .B(exu_n5609), .Y(exu_n20663));
AND2X1 exu_U6795(.A(exu_n849), .B(exu_n5610), .Y(exu_n20662));
INVX1 exu_U6796(.A(exu_n16134), .Y(exu_n16132));
INVX1 exu_U6797(.A(exu_n16141), .Y(exu_n16135));
INVX1 exu_U6798(.A(exu_n16140), .Y(exu_n16139));
INVX1 exu_U6799(.A(exu_n16140), .Y(exu_n16138));
INVX1 exu_U6800(.A(exu_n16140), .Y(exu_n16137));
INVX1 exu_U6801(.A(exu_n16141), .Y(exu_n16136));
AND2X1 exu_U6802(.A(exu_n781), .B(exu_n5544), .Y(exu_n19946));
AND2X1 exu_U6803(.A(exu_n780), .B(exu_n5543), .Y(exu_n19942));
AND2X1 exu_U6804(.A(exu_n779), .B(exu_n5542), .Y(exu_n19938));
AND2X1 exu_U6805(.A(exu_n778), .B(exu_n5541), .Y(exu_n19934));
AND2X1 exu_U6806(.A(exu_n777), .B(exu_n5540), .Y(exu_n19930));
AND2X1 exu_U6807(.A(exu_n776), .B(exu_n5539), .Y(exu_n19926));
AND2X1 exu_U6808(.A(exu_n775), .B(exu_n5538), .Y(exu_n19922));
AND2X1 exu_U6809(.A(exu_n4073), .B(exu_n9064), .Y(ecl_eccctl_ecc_synd7_mux_n1));
AND2X1 exu_U6810(.A(exu_n4566), .B(exu_n9351), .Y(exu_n31748));
AND2X1 exu_U6811(.A(exu_n4565), .B(exu_n9350), .Y(exu_n31747));
AND2X1 exu_U6812(.A(exu_n4564), .B(exu_n9349), .Y(exu_n31746));
AND2X1 exu_U6813(.A(exu_n4563), .B(exu_n9348), .Y(exu_n31745));
AND2X1 exu_U6814(.A(exu_n4562), .B(exu_n9347), .Y(exu_n31744));
AND2X1 exu_U6815(.A(exu_n4561), .B(exu_n9346), .Y(exu_n31743));
AND2X1 exu_U6816(.A(exu_n4560), .B(exu_n9345), .Y(exu_n31742));
AND2X1 exu_U6817(.A(exu_n4559), .B(exu_n9344), .Y(exu_n31741));
AND2X1 exu_U6818(.A(exu_n227), .B(exu_n5154), .Y(exu_n17724));
AND2X1 exu_U6819(.A(exu_n226), .B(exu_n5153), .Y(exu_n17720));
AND2X1 exu_U6820(.A(exu_n225), .B(exu_n5152), .Y(exu_n17716));
AND2X1 exu_U6821(.A(exu_n17712), .B(exu_n5150), .Y(exu_n31740));
AND2X1 exu_U6822(.A(exu_n224), .B(exu_n5151), .Y(exu_n17712));
AND2X1 exu_U6823(.A(exu_n17708), .B(exu_n5148), .Y(exu_n31739));
AND2X1 exu_U6824(.A(exu_n223), .B(exu_n5149), .Y(exu_n17708));
AND2X1 exu_U6825(.A(ecl_eccctl_cwp_m[2]), .B(ecl_eccctl_n25), .Y(exu_ifu_err_reg_m[7]));
AND2X1 exu_U6826(.A(exu_n4538), .B(exu_n9336), .Y(ecl_writeback_n118));
AND2X1 exu_U6827(.A(exu_n4535), .B(exu_n9333), .Y(ecl_writeback_n111));
AND2X1 exu_U6828(.A(exu_n4534), .B(exu_n9332), .Y(ecl_writeback_n103));
AND2X1 exu_U6829(.A(exu_n4533), .B(exu_n9331), .Y(ecl_writeback_n92));
INVX1 exu_U6830(.A(ecl_alu_ecl_mem_addr_invalid_m_l), .Y(exu_ifu_va_oor_m));
AND2X1 exu_U6831(.A(exu_n3642), .B(exu_n8659), .Y(exu_n31737));
OR2X1 exu_U6832(.A(exu_tlu_ue_trap_m), .B(ecl_fill_trap_m), .Y(exu_lsu_priority_trap_m));
AND2X1 exu_U6833(.A(exu_n3625), .B(exu_n8642), .Y(exu_n31736));
AND2X1 exu_U6834(.A(exu_n3614), .B(exu_n8631), .Y(exu_n31735));
AND2X1 exu_U6835(.A(exu_n3603), .B(exu_n8620), .Y(exu_n31734));
AND2X1 exu_U6836(.A(exu_n3600), .B(exu_n8617), .Y(exu_n31733));
AND2X1 exu_U6837(.A(exu_n3599), .B(exu_n8616), .Y(exu_n31732));
AND2X1 exu_U6838(.A(exu_n3598), .B(exu_n8615), .Y(exu_n31731));
AND2X1 exu_U6839(.A(exu_n3597), .B(exu_n8614), .Y(exu_n31730));
AND2X1 exu_U6840(.A(exu_n3596), .B(exu_n8613), .Y(exu_n31729));
AND2X1 exu_U6841(.A(exu_n3595), .B(exu_n8612), .Y(exu_n31728));
AND2X1 exu_U6842(.A(exu_n3594), .B(exu_n8611), .Y(exu_n31727));
AND2X1 exu_U6843(.A(exu_n3624), .B(exu_n8641), .Y(exu_n31726));
AND2X1 exu_U6844(.A(exu_n3623), .B(exu_n8640), .Y(exu_n31725));
AND2X1 exu_U6845(.A(exu_n3622), .B(exu_n8639), .Y(exu_n31724));
AND2X1 exu_U6846(.A(exu_n3621), .B(exu_n8638), .Y(exu_n31723));
AND2X1 exu_U6847(.A(exu_n3620), .B(exu_n8637), .Y(exu_n31722));
AND2X1 exu_U6848(.A(exu_n3619), .B(exu_n8636), .Y(exu_n31721));
AND2X1 exu_U6849(.A(exu_n3618), .B(exu_n8635), .Y(exu_n31720));
AND2X1 exu_U6850(.A(exu_n3617), .B(exu_n8634), .Y(exu_n31719));
AND2X1 exu_U6851(.A(exu_n3616), .B(exu_n8633), .Y(exu_n31718));
AND2X1 exu_U6852(.A(exu_n3615), .B(exu_n8632), .Y(exu_n31717));
AND2X1 exu_U6853(.A(exu_n3613), .B(exu_n8630), .Y(exu_n31716));
AND2X1 exu_U6854(.A(exu_n3612), .B(exu_n8629), .Y(exu_n31715));
AND2X1 exu_U6855(.A(exu_n3611), .B(exu_n8628), .Y(exu_n31714));
AND2X1 exu_U6856(.A(exu_n3610), .B(exu_n8627), .Y(exu_n31713));
AND2X1 exu_U6857(.A(exu_n3609), .B(exu_n8626), .Y(exu_n31712));
AND2X1 exu_U6858(.A(exu_n3608), .B(exu_n8625), .Y(exu_n31711));
AND2X1 exu_U6859(.A(exu_n3607), .B(exu_n8624), .Y(exu_n31710));
AND2X1 exu_U6860(.A(exu_n3606), .B(exu_n8623), .Y(exu_n31709));
AND2X1 exu_U6861(.A(exu_n3605), .B(exu_n8622), .Y(exu_n31708));
AND2X1 exu_U6862(.A(exu_n3604), .B(exu_n8621), .Y(exu_n31707));
AND2X1 exu_U6863(.A(exu_n3602), .B(exu_n8619), .Y(exu_n31706));
AND2X1 exu_U6864(.A(exu_n3601), .B(exu_n8618), .Y(exu_n31705));
OR2X1 exu_U6865(.A(ecl_early_ttype_m[0]), .B(exu_tlu_ue_trap_m), .Y(exu_tlu_ttype_m[0]));
AND2X1 exu_U6866(.A(ecl_early_ttype_m[1]), .B(exu_n16595), .Y(exu_tlu_ttype_m[1]));
AND2X1 exu_U6867(.A(ecl_early_ttype_m[2]), .B(exu_n16595), .Y(exu_tlu_ttype_m[2]));
OR2X1 exu_U6868(.A(ecl_early_ttype_m[3]), .B(exu_tlu_ue_trap_m), .Y(exu_tlu_ttype_m[3]));
AND2X1 exu_U6869(.A(ecl_early_ttype_m[4]), .B(exu_n16595), .Y(exu_tlu_ttype_m[4]));
OR2X1 exu_U6870(.A(ecl_early_ttype_m[5]), .B(exu_tlu_ue_trap_m), .Y(exu_tlu_ttype_m[5]));
AND2X1 exu_U6871(.A(ecl_early_ttype_m[6]), .B(exu_n16595), .Y(exu_tlu_ttype_m[6]));
AND2X1 exu_U6872(.A(ecl_early_ttype_m[8]), .B(exu_n16595), .Y(exu_tlu_ttype_m[8]));
OR2X1 exu_U6873(.A(ecl_div_zero_m), .B(ecl_n102), .Y(exu_tlu_ttype_vld_m));
OR2X1 exu_U6874(.A(exu_tlu_ue_trap_m), .B(ecl_early_ttype_vld_m), .Y(ecl_n102));
AND2X1 exu_U6875(.A(ecl_eccctl_nceen_m), .B(exu_ifu_ecc_ue_m), .Y(exu_tlu_ue_trap_m));
AND2X1 exu_U6876(.A(ecl_ifu_exu_range_check_jlret_m), .B(exu_ifu_va_oor_m), .Y(exu_tlu_va_oor_jl_ret_m));
AND2X1 exu_U6877(.A(ecl_ifu_exu_range_check_other_m), .B(exu_ifu_va_oor_m), .Y(exu_tlu_va_oor_m));
OR2X1 exu_U6878(.A(exu_n13429), .B(exu_n14742), .Y(rml_irf_old_agp[0]));
AND2X1 exu_U6879(.A(exu_n4139), .B(exu_n9115), .Y(rml_mux_agp_out1_n7));
OR2X1 exu_U6880(.A(exu_n13428), .B(exu_n14741), .Y(rml_irf_old_agp[1]));
AND2X1 exu_U6881(.A(exu_n4137), .B(exu_n9113), .Y(rml_mux_agp_out1_n1));
OR2X1 exu_U6882(.A(rml_n59), .B(rml_kill_restore_w), .Y(rml_irf_kill_restore_w));
AND2X1 exu_U6883(.A(rml_did_restore_w), .B(exu_n15740), .Y(rml_n59));
OR2X1 exu_U6884(.A(exu_n15346), .B(rml_swap_locals_ins), .Y(rml_irf_swap_local_e));
OR2X1 exu_U6885(.A(exu_n13393), .B(exu_n14700), .Y(ecl_irf_tid_g[0]));
AND2X1 exu_U6886(.A(exu_n3966), .B(exu_n8981), .Y(exu_n31463));
OR2X1 exu_U6887(.A(exu_n13392), .B(exu_n14699), .Y(ecl_irf_tid_g[1]));
AND2X1 exu_U6888(.A(exu_n3964), .B(exu_n8979), .Y(exu_n31457));
INVX1 exu_U6889(.A(bypass_rd_synd_w2_l[0]), .Y(byp_irf_rd_data_w2[64]));
INVX1 exu_U6890(.A(bypass_rd_synd_w2_l[1]), .Y(byp_irf_rd_data_w2[65]));
INVX1 exu_U6891(.A(bypass_rd_synd_w2_l[2]), .Y(byp_irf_rd_data_w2[66]));
INVX1 exu_U6892(.A(bypass_rd_synd_w2_l[3]), .Y(byp_irf_rd_data_w2[67]));
INVX1 exu_U6893(.A(bypass_rd_synd_w2_l[4]), .Y(byp_irf_rd_data_w2[68]));
INVX1 exu_U6894(.A(bypass_rd_synd_w2_l[5]), .Y(byp_irf_rd_data_w2[69]));
INVX1 exu_U6895(.A(bypass_rd_synd_w2_l[6]), .Y(byp_irf_rd_data_w2[70]));
INVX1 exu_U6896(.A(bypass_rd_synd_w2_l[7]), .Y(byp_irf_rd_data_w2[71]));
INVX1 exu_U6897(.A(bypass_rd_synd_w_l[0]), .Y(byp_irf_rd_data_w[64]));
INVX1 exu_U6898(.A(bypass_rd_synd_w_l[1]), .Y(byp_irf_rd_data_w[65]));
INVX1 exu_U6899(.A(bypass_rd_synd_w_l[2]), .Y(byp_irf_rd_data_w[66]));
INVX1 exu_U6900(.A(bypass_rd_synd_w_l[3]), .Y(byp_irf_rd_data_w[67]));
INVX1 exu_U6901(.A(bypass_rd_synd_w_l[4]), .Y(byp_irf_rd_data_w[68]));
INVX1 exu_U6902(.A(bypass_rd_synd_w_l[5]), .Y(byp_irf_rd_data_w[69]));
INVX1 exu_U6903(.A(bypass_rd_synd_w_l[6]), .Y(byp_irf_rd_data_w[70]));
INVX1 exu_U6904(.A(bypass_rd_synd_w_l[7]), .Y(byp_irf_rd_data_w[71]));
OR2X1 exu_U6905(.A(exu_n13419), .B(exu_n14732), .Y(ecl_irf_rd_g[0]));
AND2X1 exu_U6906(.A(exu_n4095), .B(exu_n9089), .Y(ecl_writeback_rd_g_mux_n25));
OR2X1 exu_U6907(.A(exu_n13418), .B(exu_n14731), .Y(ecl_irf_rd_g[1]));
AND2X1 exu_U6908(.A(exu_n4093), .B(exu_n9087), .Y(ecl_writeback_rd_g_mux_n19));
OR2X1 exu_U6909(.A(exu_n13417), .B(exu_n14730), .Y(ecl_irf_rd_g[2]));
AND2X1 exu_U6910(.A(exu_n4091), .B(exu_n9085), .Y(ecl_writeback_rd_g_mux_n13));
OR2X1 exu_U6911(.A(exu_n13416), .B(exu_n14729), .Y(ecl_irf_rd_g[3]));
AND2X1 exu_U6912(.A(exu_n4089), .B(exu_n9083), .Y(ecl_writeback_rd_g_mux_n7));
OR2X1 exu_U6913(.A(exu_n13415), .B(exu_n14728), .Y(ecl_irf_rd_g[4]));
AND2X1 exu_U6914(.A(exu_n4087), .B(exu_n9081), .Y(ecl_writeback_rd_g_mux_n1));
OR2X1 exu_U6915(.A(exu_n12136), .B(exu_n13552), .Y(ecl_irf_rd_m[0]));
AND2X1 exu_U6916(.A(exu_n321), .B(exu_n5248), .Y(exu_n18005));
OR2X1 exu_U6917(.A(exu_n12135), .B(exu_n13551), .Y(ecl_irf_rd_m[1]));
AND2X1 exu_U6918(.A(exu_n319), .B(exu_n5246), .Y(exu_n17999));
OR2X1 exu_U6919(.A(exu_n12134), .B(exu_n13550), .Y(ecl_irf_rd_m[2]));
AND2X1 exu_U6920(.A(exu_n317), .B(exu_n5244), .Y(exu_n17993));
OR2X1 exu_U6921(.A(exu_n12133), .B(exu_n13549), .Y(ecl_irf_rd_m[3]));
AND2X1 exu_U6922(.A(exu_n315), .B(exu_n5242), .Y(exu_n17987));
OR2X1 exu_U6923(.A(exu_n12132), .B(exu_n13548), .Y(ecl_irf_rd_m[4]));
AND2X1 exu_U6924(.A(exu_n313), .B(exu_n5240), .Y(exu_n17981));
OR2X1 exu_U6925(.A(rml_cwp_n37), .B(exu_n14702), .Y(rml_cwp_next_slot1_state[1]));
AND2X1 exu_U6926(.A(exu_n3968), .B(exu_n8983), .Y(exu_n31474));
OR2X1 exu_U6927(.A(exu_n31478), .B(exu_n31477), .Y(rml_cwp_next_slot1_state[0]));
AND2X1 exu_U6928(.A(exu_n163), .B(exu_n5123), .Y(exu_n17513));
AND2X1 exu_U6929(.A(exu_n165), .B(exu_n5124), .Y(exu_n17517));
AND2X1 exu_U6930(.A(exu_n167), .B(exu_n5125), .Y(exu_n17521));
AND2X1 exu_U6931(.A(exu_n169), .B(exu_n5126), .Y(exu_n17525));
AND2X1 exu_U6932(.A(exu_n171), .B(exu_n5127), .Y(exu_n17529));
AND2X1 exu_U6933(.A(exu_n176), .B(exu_n5128), .Y(exu_n17539));
OR2X1 exu_U6934(.A(rml_cwp_n36), .B(exu_n14703), .Y(rml_cwp_next_slot2_state[1]));
AND2X1 exu_U6935(.A(exu_n3969), .B(exu_n8984), .Y(exu_n31479));
OR2X1 exu_U6936(.A(exu_n31483), .B(exu_n31482), .Y(rml_cwp_next_slot2_state[0]));
AND2X1 exu_U6937(.A(exu_n182), .B(exu_n5129), .Y(exu_n17550));
AND2X1 exu_U6938(.A(exu_n184), .B(exu_n5130), .Y(exu_n17554));
AND2X1 exu_U6939(.A(exu_n186), .B(exu_n5131), .Y(exu_n17558));
AND2X1 exu_U6940(.A(exu_n188), .B(exu_n5132), .Y(exu_n17562));
AND2X1 exu_U6941(.A(exu_n190), .B(exu_n5133), .Y(exu_n17566));
AND2X1 exu_U6942(.A(exu_n195), .B(exu_n5134), .Y(exu_n17576));
OR2X1 exu_U6943(.A(rml_cwp_n35), .B(exu_n14704), .Y(rml_cwp_next_slot3_state[1]));
AND2X1 exu_U6944(.A(exu_n3970), .B(exu_n8985), .Y(exu_n31484));
OR2X1 exu_U6945(.A(exu_n31488), .B(exu_n31487), .Y(rml_cwp_next_slot3_state[0]));
AND2X1 exu_U6946(.A(exu_n201), .B(exu_n5135), .Y(exu_n17587));
AND2X1 exu_U6947(.A(exu_n203), .B(exu_n5136), .Y(exu_n17591));
AND2X1 exu_U6948(.A(exu_n205), .B(exu_n5137), .Y(exu_n17595));
AND2X1 exu_U6949(.A(exu_n207), .B(exu_n5138), .Y(exu_n17599));
AND2X1 exu_U6950(.A(exu_n209), .B(exu_n5139), .Y(exu_n17603));
AND2X1 exu_U6951(.A(exu_n214), .B(exu_n5140), .Y(exu_n17613));
OR2X1 exu_U6952(.A(ecl_divcntl_cnt6_n16), .B(exu_n14723), .Y(ecl_divcntl_cnt6_n15));
OR2X1 exu_U6953(.A(exu_n15387), .B(exu_n14724), .Y(ecl_divcntl_cnt6_n22));
AND2X1 exu_U6954(.A(ecl_divcntl_cnt6_n32), .B(ecl_divcntl_div_state_1), .Y(ecl_divcntl_cnt6_next_cntr[1]));
AND2X1 exu_U6955(.A(rml_cwp_swap_data[7]), .B(rml_cwp_n96), .Y(rml_cwp_cwp_cmplt_next));
OR2X1 exu_U6956(.A(exu_n13408), .B(exu_n14719), .Y(rml_cwp_swap_data_12));
AND2X1 exu_U6957(.A(exu_n678), .B(exu_n5399), .Y(exu_n18956));
AND2X1 exu_U6958(.A(exu_n681), .B(exu_n5400), .Y(exu_n18959));
AND2X1 exu_U6959(.A(exu_n684), .B(exu_n5401), .Y(exu_n18962));
AND2X1 exu_U6960(.A(exu_n687), .B(exu_n5402), .Y(exu_n18965));
AND2X1 exu_U6961(.A(exu_n690), .B(exu_n5403), .Y(exu_n18968));
AND2X1 exu_U6962(.A(exu_n693), .B(exu_n5404), .Y(exu_n18971));
AND2X1 exu_U6963(.A(exu_n696), .B(exu_n5405), .Y(exu_n18974));
AND2X1 exu_U6964(.A(exu_n699), .B(exu_n5406), .Y(exu_n18977));
AND2X1 exu_U6965(.A(exu_n704), .B(exu_n5408), .Y(exu_n18984));
AND2X1 exu_U6966(.A(exu_n707), .B(exu_n5409), .Y(exu_n18987));
AND2X1 exu_U6967(.A(exu_n710), .B(exu_n5410), .Y(exu_n18990));
AND2X1 exu_U6968(.A(exu_n713), .B(exu_n5411), .Y(exu_n18993));
AND2X1 exu_U6969(.A(exu_n716), .B(exu_n5412), .Y(exu_n18996));
AND2X1 exu_U6970(.A(exu_n719), .B(exu_n5413), .Y(exu_n18999));
AND2X1 exu_U6971(.A(exu_n480), .B(exu_n5303), .Y(exu_n18607));
AND2X1 exu_U6972(.A(exu_n480), .B(exu_n5304), .Y(exu_n18610));
AND2X1 exu_U6973(.A(exu_n483), .B(exu_n5305), .Y(exu_n18613));
AND2X1 exu_U6974(.A(exu_n486), .B(exu_n5306), .Y(exu_n18616));
AND2X1 exu_U6975(.A(exu_n488), .B(exu_n5307), .Y(exu_n18619));
AND2X1 exu_U6976(.A(exu_n490), .B(exu_n5308), .Y(exu_n18623));
AND2X1 exu_U6977(.A(exu_n492), .B(exu_n5309), .Y(exu_n18627));
AND2X1 exu_U6978(.A(exu_n494), .B(exu_n5310), .Y(exu_n18631));
AND2X1 exu_U6979(.A(exu_n496), .B(exu_n5311), .Y(exu_n18635));
AND2X1 exu_U6980(.A(exu_n498), .B(exu_n5312), .Y(exu_n18639));
AND2X1 exu_U6981(.A(exu_n502), .B(exu_n5314), .Y(exu_n18647));
AND2X1 exu_U6982(.A(exu_n504), .B(exu_n5315), .Y(exu_n18651));
AND2X1 exu_U6983(.A(exu_n506), .B(exu_n5316), .Y(exu_n18655));
AND2X1 exu_U6984(.A(exu_n508), .B(exu_n5317), .Y(exu_n18659));
AND2X1 exu_U6985(.A(exu_n510), .B(exu_n5318), .Y(exu_n18663));
AND2X1 exu_U6986(.A(exu_n512), .B(exu_n5319), .Y(exu_n18667));
AND2X1 exu_U6987(.A(exu_n514), .B(exu_n5320), .Y(exu_n18671));
AND2X1 exu_U6988(.A(exu_n516), .B(exu_n5321), .Y(exu_n18675));
AND2X1 exu_U6989(.A(exu_n518), .B(exu_n5322), .Y(exu_n18679));
AND2X1 exu_U6990(.A(exu_n520), .B(exu_n5323), .Y(exu_n18683));
AND2X1 exu_U6991(.A(exu_n524), .B(exu_n5325), .Y(exu_n18691));
AND2X1 exu_U6992(.A(exu_n526), .B(exu_n5326), .Y(exu_n18695));
AND2X1 exu_U6993(.A(exu_n528), .B(exu_n5327), .Y(exu_n18699));
AND2X1 exu_U6994(.A(exu_n530), .B(exu_n5328), .Y(exu_n18703));
AND2X1 exu_U6995(.A(exu_n532), .B(exu_n5329), .Y(exu_n18707));
AND2X1 exu_U6996(.A(exu_n534), .B(exu_n5330), .Y(exu_n18711));
AND2X1 exu_U6997(.A(exu_n536), .B(exu_n5331), .Y(exu_n18715));
AND2X1 exu_U6998(.A(exu_n538), .B(exu_n5332), .Y(exu_n18719));
AND2X1 exu_U6999(.A(exu_n540), .B(exu_n5333), .Y(exu_n18723));
AND2X1 exu_U7000(.A(exu_n542), .B(exu_n5334), .Y(exu_n18727));
AND2X1 exu_U7001(.A(exu_n546), .B(exu_n5336), .Y(exu_n18735));
AND2X1 exu_U7002(.A(exu_n548), .B(exu_n5337), .Y(exu_n18739));
AND2X1 exu_U7003(.A(exu_n550), .B(exu_n5338), .Y(exu_n18743));
AND2X1 exu_U7004(.A(exu_n552), .B(exu_n5339), .Y(exu_n18747));
AND2X1 exu_U7005(.A(exu_n554), .B(exu_n5340), .Y(exu_n18751));
AND2X1 exu_U7006(.A(exu_n556), .B(exu_n5341), .Y(exu_n18755));
AND2X1 exu_U7007(.A(exu_n560), .B(exu_n5342), .Y(exu_n18759));
AND2X1 exu_U7008(.A(exu_n560), .B(exu_n5343), .Y(exu_n18762));
AND2X1 exu_U7009(.A(exu_n563), .B(exu_n5344), .Y(exu_n18765));
AND2X1 exu_U7010(.A(exu_n566), .B(exu_n5345), .Y(exu_n18768));
AND2X1 exu_U7011(.A(exu_n571), .B(exu_n5347), .Y(exu_n18775));
AND2X1 exu_U7012(.A(exu_n574), .B(exu_n5348), .Y(exu_n18778));
AND2X1 exu_U7013(.A(exu_n577), .B(exu_n5349), .Y(exu_n18781));
AND2X1 exu_U7014(.A(exu_n580), .B(exu_n5350), .Y(exu_n18784));
AND2X1 exu_U7015(.A(exu_n583), .B(exu_n5351), .Y(exu_n18787));
AND2X1 exu_U7016(.A(exu_n586), .B(exu_n5352), .Y(exu_n18790));
AND2X1 exu_U7017(.A(exu_n589), .B(exu_n5353), .Y(exu_n18793));
AND2X1 exu_U7018(.A(exu_n592), .B(exu_n5354), .Y(exu_n18796));
AND2X1 exu_U7019(.A(exu_n595), .B(exu_n5355), .Y(exu_n18799));
AND2X1 exu_U7020(.A(exu_n598), .B(exu_n5356), .Y(exu_n18802));
AND2X1 exu_U7021(.A(exu_n603), .B(exu_n5358), .Y(exu_n18809));
AND2X1 exu_U7022(.A(exu_n606), .B(exu_n5359), .Y(exu_n18812));
AND2X1 exu_U7023(.A(exu_n609), .B(exu_n5360), .Y(exu_n18815));
AND2X1 exu_U7024(.A(exu_n612), .B(exu_n5361), .Y(exu_n18818));
AND2X1 exu_U7025(.A(exu_n615), .B(exu_n5362), .Y(exu_n18821));
AND2X1 exu_U7026(.A(exu_n633), .B(exu_n5377), .Y(exu_n18868));
AND2X1 exu_U7027(.A(exu_n635), .B(exu_n5378), .Y(exu_n18872));
AND2X1 exu_U7028(.A(exu_n639), .B(exu_n5380), .Y(exu_n18880));
AND2X1 exu_U7029(.A(exu_n641), .B(exu_n5381), .Y(exu_n18884));
AND2X1 exu_U7030(.A(exu_n643), .B(exu_n5382), .Y(exu_n18888));
AND2X1 exu_U7031(.A(exu_n645), .B(exu_n5383), .Y(exu_n18892));
AND2X1 exu_U7032(.A(exu_n647), .B(exu_n5384), .Y(exu_n18896));
AND2X1 exu_U7033(.A(exu_n649), .B(exu_n5385), .Y(exu_n18900));
AND2X1 exu_U7034(.A(exu_n651), .B(exu_n5386), .Y(exu_n18904));
AND2X1 exu_U7035(.A(exu_n653), .B(exu_n5387), .Y(exu_n18908));
AND2X1 exu_U7036(.A(exu_n655), .B(exu_n5388), .Y(exu_n18912));
AND2X1 exu_U7037(.A(exu_n657), .B(exu_n5389), .Y(exu_n18916));
AND2X1 exu_U7038(.A(exu_n661), .B(exu_n5391), .Y(exu_n18924));
AND2X1 exu_U7039(.A(exu_n663), .B(exu_n5392), .Y(exu_n18928));
AND2X1 exu_U7040(.A(exu_n665), .B(exu_n5393), .Y(exu_n18932));
AND2X1 exu_U7041(.A(exu_n667), .B(exu_n5394), .Y(exu_n18936));
AND2X1 exu_U7042(.A(exu_n669), .B(exu_n5395), .Y(exu_n18940));
AND2X1 exu_U7043(.A(exu_n671), .B(exu_n5396), .Y(exu_n18944));
AND2X1 exu_U7044(.A(exu_n673), .B(exu_n5397), .Y(exu_n18948));
AND2X1 exu_U7045(.A(exu_n675), .B(exu_n5398), .Y(exu_n18952));
AND2X1 exu_U7046(.A(exu_n701), .B(exu_n5407), .Y(exu_n18980));
AND2X1 exu_U7047(.A(exu_n725), .B(exu_n5418), .Y(exu_n19014));
AND2X1 exu_U7048(.A(exu_n476), .B(exu_n5302), .Y(exu_n18603));
AND2X1 exu_U7049(.A(exu_n500), .B(exu_n5313), .Y(exu_n18643));
AND2X1 exu_U7050(.A(exu_n522), .B(exu_n5324), .Y(exu_n18687));
AND2X1 exu_U7051(.A(exu_n544), .B(exu_n5335), .Y(exu_n18731));
AND2X1 exu_U7052(.A(exu_n568), .B(exu_n5346), .Y(exu_n18771));
AND2X1 exu_U7053(.A(exu_n600), .B(exu_n5357), .Y(exu_n18805));
AND2X1 exu_U7054(.A(exu_n622), .B(exu_n5368), .Y(exu_n18839));
AND2X1 exu_U7055(.A(exu_n637), .B(exu_n5379), .Y(exu_n18876));
AND2X1 exu_U7056(.A(exu_n659), .B(exu_n5390), .Y(exu_n18920));
AND2X1 exu_U7057(.A(exu_n738), .B(exu_n5429), .Y(exu_n19049));
AND2X1 exu_U7058(.A(exu_n4961), .B(exu_n9661), .Y(ecl_dff_sel_sum_d2e_din[0]));
OR2X1 exu_U7059(.A(ifu_exu_rs3o_vld_d), .B(ifu_exu_rs3e_vld_d), .Y(ecl_rs3_vld_d));
INVX1 exu_U7060(.A(se), .Y(exu_n19283));
INVX1 exu_U7061(.A(ifu_exu_muls_d), .Y(exu_n16386));
INVX1 exu_U7062(.A(se), .Y(exu_n19287));
INVX1 exu_U7063(.A(se), .Y(exu_n19295));
INVX1 exu_U7064(.A(se), .Y(exu_n19297));
INVX1 exu_U7065(.A(se), .Y(exu_n19299));
INVX1 exu_U7066(.A(se), .Y(exu_n19301));
INVX1 exu_U7067(.A(se), .Y(exu_n19303));
INVX1 exu_U7068(.A(se), .Y(exu_n19305));
INVX1 exu_U7069(.A(se), .Y(exu_n19307));
INVX1 exu_U7070(.A(se), .Y(exu_n19309));
INVX1 exu_U7071(.A(se), .Y(exu_n19311));
INVX1 exu_U7072(.A(se), .Y(exu_n19313));
INVX1 exu_U7073(.A(se), .Y(exu_n19315));
INVX1 exu_U7074(.A(se), .Y(exu_n19317));
OR2X1 exu_U7075(.A(ecl_ifu_tlu_flush_w), .B(lsu_exu_flush_pipe_w), .Y(ecl_flush_w));
INVX1 exu_U7076(.A(se), .Y(exu_n19319));
INVX1 exu_U7077(.A(se), .Y(exu_n19321));
INVX1 exu_U7078(.A(se), .Y(exu_n19323));
AND2X1 exu_U7079(.A(ifu_exu_rs3o_vld_d), .B(ifu_exu_rs3e_vld_d), .Y(ecl_std_d));
INVX1 exu_U7080(.A(se), .Y(exu_n19325));
OR2X1 exu_U7081(.A(exu_n13501), .B(ecl_n111), .Y(ecl_early_ttype_vld_e));
OR2X1 exu_U7082(.A(exu_n15493), .B(ecl_misalign_addr_e), .Y(ecl_n111));
INVX1 exu_U7083(.A(se), .Y(exu_n19327));
INVX1 exu_U7084(.A(se), .Y(exu_n19329));
INVX1 exu_U7085(.A(se), .Y(exu_n19331));
INVX1 exu_U7086(.A(se), .Y(exu_n19333));
INVX1 exu_U7087(.A(se), .Y(exu_n19335));
INVX1 exu_U7088(.A(se), .Y(exu_n19291));
INVX1 exu_U7089(.A(se), .Y(exu_n19339));
INVX1 exu_U7090(.A(se), .Y(exu_n19293));
INVX1 exu_U7091(.A(se), .Y(exu_n19341));
OR2X1 exu_U7092(.A(rml_ecl_clean_window_e), .B(rml_rml_ecl_kill_e), .Y(rml_win_trap_e));
INVX1 exu_U7093(.A(se), .Y(exu_n19343));
INVX1 exu_U7094(.A(se), .Y(exu_n19345));
INVX1 exu_U7095(.A(se), .Y(exu_n19347));
INVX1 exu_U7096(.A(se), .Y(exu_n19349));
INVX1 exu_U7097(.A(se), .Y(exu_n19351));
INVX1 exu_U7098(.A(se), .Y(exu_n19353));
INVX1 exu_U7099(.A(se), .Y(exu_n19355));
INVX1 exu_U7100(.A(se), .Y(exu_n19357));
INVX1 exu_U7101(.A(se), .Y(exu_n19359));
INVX1 exu_U7102(.A(se), .Y(exu_n19361));
INVX1 exu_U7103(.A(se), .Y(exu_n19363));
INVX1 exu_U7104(.A(se), .Y(exu_n19365));
INVX1 exu_U7105(.A(se), .Y(exu_n19367));
INVX1 exu_U7106(.A(se), .Y(exu_n19369));
INVX1 exu_U7107(.A(se), .Y(exu_n19371));
INVX1 exu_U7108(.A(se), .Y(exu_n19373));
INVX1 exu_U7109(.A(se), .Y(exu_n19375));
INVX1 exu_U7110(.A(se), .Y(exu_n19381));
INVX1 exu_U7111(.A(se), .Y(exu_n19383));
INVX1 exu_U7112(.A(se), .Y(exu_n19385));
INVX1 exu_U7113(.A(se), .Y(exu_n19387));
INVX1 exu_U7114(.A(se), .Y(exu_n19389));
INVX1 exu_U7115(.A(se), .Y(exu_n19391));
INVX1 exu_U7116(.A(se), .Y(exu_n19393));
INVX1 exu_U7117(.A(se), .Y(exu_n19395));
INVX1 exu_U7118(.A(se), .Y(exu_n19397));
INVX1 exu_U7119(.A(se), .Y(exu_n19399));
INVX1 exu_U7120(.A(exu_n16171), .Y(exu_n16172));
INVX1 exu_U7121(.A(se), .Y(exu_n19401));
INVX1 exu_U7122(.A(se), .Y(exu_n19403));
INVX1 exu_U7123(.A(se), .Y(exu_n19405));
INVX1 exu_U7124(.A(se), .Y(exu_n19407));
INVX1 exu_U7125(.A(se), .Y(exu_n19409));
INVX1 exu_U7126(.A(se), .Y(exu_n19411));
INVX1 exu_U7127(.A(se), .Y(exu_n19413));
INVX1 exu_U7128(.A(se), .Y(exu_n19415));
INVX1 exu_U7129(.A(se), .Y(exu_n19417));
INVX1 exu_U7130(.A(se), .Y(exu_n19419));
INVX1 exu_U7131(.A(se), .Y(exu_n19421));
INVX1 exu_U7132(.A(se), .Y(exu_n19423));
INVX1 exu_U7133(.A(se), .Y(exu_n19425));
INVX1 exu_U7134(.A(exu_n16171), .Y(exu_n16173));
INVX1 exu_U7135(.A(se), .Y(exu_n19427));
INVX1 exu_U7136(.A(se), .Y(exu_n19429));
INVX1 exu_U7137(.A(se), .Y(exu_n19431));
INVX1 exu_U7138(.A(se), .Y(exu_n19433));
INVX1 exu_U7139(.A(se), .Y(exu_n19435));
INVX1 exu_U7140(.A(se), .Y(exu_n19437));
INVX1 exu_U7141(.A(se), .Y(exu_n19439));
INVX1 exu_U7142(.A(se), .Y(exu_n19441));
INVX1 exu_U7143(.A(se), .Y(exu_n19443));
INVX1 exu_U7144(.A(se), .Y(exu_n19445));
INVX1 exu_U7145(.A(se), .Y(exu_n19447));
INVX1 exu_U7146(.A(se), .Y(exu_n19449));
INVX1 exu_U7147(.A(se), .Y(exu_n19451));
INVX1 exu_U7148(.A(exu_n16171), .Y(exu_n16174));
INVX1 exu_U7149(.A(se), .Y(exu_n19453));
INVX1 exu_U7150(.A(se), .Y(exu_n19455));
INVX1 exu_U7151(.A(se), .Y(exu_n19457));
INVX1 exu_U7152(.A(se), .Y(exu_n19459));
INVX1 exu_U7153(.A(se), .Y(exu_n19461));
INVX1 exu_U7154(.A(se), .Y(exu_n19463));
INVX1 exu_U7155(.A(se), .Y(exu_n19465));
INVX1 exu_U7156(.A(se), .Y(exu_n19467));
INVX1 exu_U7157(.A(se), .Y(exu_n19469));
INVX1 exu_U7158(.A(se), .Y(exu_n19471));
INVX1 exu_U7159(.A(se), .Y(exu_n19473));
INVX1 exu_U7160(.A(se), .Y(exu_n19475));
INVX1 exu_U7161(.A(se), .Y(exu_n19377));
INVX1 exu_U7162(.A(exu_n16171), .Y(exu_n16175));
INVX1 exu_U7163(.A(se), .Y(exu_n19379));
INVX1 exu_U7164(.A(se), .Y(exu_n19477));
INVX1 exu_U7165(.A(se), .Y(exu_n19479));
INVX1 exu_U7166(.A(se), .Y(exu_n19481));
INVX1 exu_U7167(.A(se), .Y(exu_n19483));
INVX1 exu_U7168(.A(se), .Y(exu_n19485));
INVX1 exu_U7169(.A(se), .Y(exu_n19487));
INVX1 exu_U7170(.A(se), .Y(exu_n19489));
INVX1 exu_U7171(.A(se), .Y(exu_n19491));
INVX1 exu_U7172(.A(se), .Y(exu_n19493));
INVX1 exu_U7173(.A(se), .Y(exu_n19495));
INVX1 exu_U7174(.A(se), .Y(exu_n19497));
INVX1 exu_U7175(.A(se), .Y(exu_n19499));
INVX1 exu_U7176(.A(exu_n16171), .Y(exu_n16176));
INVX1 exu_U7177(.A(se), .Y(exu_n19501));
INVX1 exu_U7178(.A(se), .Y(exu_n19503));
INVX1 exu_U7179(.A(se), .Y(exu_n19505));
INVX1 exu_U7180(.A(se), .Y(exu_n19507));
INVX1 exu_U7181(.A(se), .Y(exu_n19509));
INVX1 exu_U7182(.A(se), .Y(exu_n19511));
INVX1 exu_U7183(.A(se), .Y(exu_n19513));
INVX1 exu_U7184(.A(se), .Y(exu_n19515));
INVX1 exu_U7185(.A(se), .Y(exu_n19517));
INVX1 exu_U7186(.A(se), .Y(exu_n19519));
INVX1 exu_U7187(.A(se), .Y(exu_n19521));
INVX1 exu_U7188(.A(se), .Y(exu_n19523));
INVX1 exu_U7189(.A(se), .Y(exu_n19525));
INVX1 exu_U7190(.A(exu_n16171), .Y(exu_n16177));
INVX1 exu_U7191(.A(se), .Y(exu_n19527));
INVX1 exu_U7192(.A(se), .Y(exu_n19529));
INVX1 exu_U7193(.A(se), .Y(exu_n19531));
INVX1 exu_U7194(.A(se), .Y(exu_n19533));
INVX1 exu_U7195(.A(se), .Y(exu_n19535));
INVX1 exu_U7196(.A(se), .Y(exu_n19537));
INVX1 exu_U7197(.A(se), .Y(exu_n19539));
INVX1 exu_U7198(.A(se), .Y(exu_n19541));
INVX1 exu_U7199(.A(se), .Y(exu_n19543));
INVX1 exu_U7200(.A(se), .Y(exu_n19545));
INVX1 exu_U7201(.A(se), .Y(exu_n19547));
INVX1 exu_U7202(.A(se), .Y(exu_n19549));
INVX1 exu_U7203(.A(se), .Y(exu_n19551));
INVX1 exu_U7204(.A(exu_n16171), .Y(exu_n16178));
INVX1 exu_U7205(.A(se), .Y(exu_n19553));
INVX1 exu_U7206(.A(se), .Y(exu_n19555));
INVX1 exu_U7207(.A(se), .Y(exu_n19557));
INVX1 exu_U7208(.A(se), .Y(exu_n19559));
INVX1 exu_U7209(.A(se), .Y(exu_n19561));
INVX1 exu_U7210(.A(se), .Y(exu_n19563));
INVX1 exu_U7211(.A(se), .Y(exu_n19565));
INVX1 exu_U7212(.A(se), .Y(exu_n19567));
INVX1 exu_U7213(.A(se), .Y(exu_n19569));
INVX1 exu_U7214(.A(se), .Y(exu_n19571));
INVX1 exu_U7215(.A(se), .Y(exu_n19573));
INVX1 exu_U7216(.A(se), .Y(exu_n19575));
INVX1 exu_U7217(.A(se), .Y(exu_n19577));
OR2X1 exu_U7218(.A(tlu_exu_cwpccr_update_m), .B(ecl_ccr_setcc_m), .Y(ecl_ccr_valid_setcc_m));
INVX1 exu_U7219(.A(se), .Y(exu_n19579));
OR2X1 exu_U7220(.A(exu_n16269), .B(lsu_exu_dfill_vld_g), .Y(ecl_writeback_ld_g));
INVX1 exu_U7221(.A(se), .Y(exu_n19581));
INVX1 exu_U7222(.A(se), .Y(exu_n19583));
INVX1 exu_U7223(.A(se), .Y(exu_n19585));
INVX1 exu_U7224(.A(se), .Y(exu_n19587));
INVX1 exu_U7225(.A(se), .Y(exu_n19589));
INVX1 exu_U7226(.A(se), .Y(exu_n19591));
INVX1 exu_U7227(.A(se), .Y(exu_n19593));
INVX1 exu_U7228(.A(se), .Y(exu_n19595));
INVX1 exu_U7229(.A(se), .Y(exu_n19597));
AND2X1 exu_U7230(.A(ifu_exu_inst_vld_w), .B(exu_n9327), .Y(ecl_writeback_yreg_wen_w));
INVX1 exu_U7231(.A(se), .Y(exu_n19599));
INVX1 exu_U7232(.A(se), .Y(exu_n19601));
INVX1 exu_U7233(.A(se), .Y(exu_n19603));
INVX1 exu_U7234(.A(se), .Y(exu_n19605));
INVX1 exu_U7235(.A(se), .Y(exu_n19607));
AND2X1 exu_U7236(.A(ifu_exu_inst_vld_e), .B(ecl_writeback_n65), .Y(ecl_writeback_short_longop_done_e));
AND2X1 exu_U7237(.A(ecl_writeback_n66), .B(exu_n16389), .Y(ecl_writeback_n65));
INVX1 exu_U7238(.A(se), .Y(exu_n19609));
INVX1 exu_U7239(.A(se), .Y(exu_n19611));
INVX1 exu_U7240(.A(se), .Y(exu_n19613));
INVX1 exu_U7241(.A(se), .Y(exu_n19615));
INVX1 exu_U7242(.A(se), .Y(exu_n19617));
INVX1 exu_U7243(.A(se), .Y(exu_n19619));
INVX1 exu_U7244(.A(se), .Y(exu_n19623));
AND2X1 exu_U7245(.A(exu_n16391), .B(ecc_ecl_rs2_ce), .Y(ecl_eccctl_sel_rs2_e));
INVX1 exu_U7246(.A(ecc_ecl_rs1_ce), .Y(exu_n16391));
INVX1 exu_U7247(.A(se), .Y(exu_n19625));
INVX1 exu_U7248(.A(se), .Y(exu_n19627));
INVX1 exu_U7249(.A(se), .Y(exu_n19629));
INVX1 exu_U7250(.A(se), .Y(exu_n19621));
INVX1 exu_U7251(.A(se), .Y(exu_n19631));
INVX1 exu_U7252(.A(se), .Y(exu_n19633));
INVX1 exu_U7253(.A(se), .Y(exu_n19635));
INVX1 exu_U7254(.A(se), .Y(exu_n19637));
INVX1 exu_U7255(.A(se), .Y(exu_n19640));
INVX1 exu_U7256(.A(se), .Y(exu_n19642));
INVX1 exu_U7257(.A(se), .Y(exu_n19644));
INVX1 exu_U7258(.A(se), .Y(exu_n19646));
INVX1 exu_U7259(.A(se), .Y(exu_n19648));
INVX1 exu_U7260(.A(se), .Y(exu_n19650));
INVX1 exu_U7261(.A(se), .Y(exu_n19652));
AND2X1 exu_U7262(.A(ecl_mdqctl_n51), .B(exu_n16213), .Y(ecl_mdqctl_isdiv_e_valid));
INVX1 exu_U7263(.A(se), .Y(exu_n19654));
AND2X1 exu_U7264(.A(ecl_mdqctl_n51), .B(ecl_mdqctl_isdiv_m), .Y(ecl_mdqctl_isdiv_m_valid));
INVX1 exu_U7265(.A(se), .Y(exu_n19656));
AND2X1 exu_U7266(.A(ecl_mdqctl_ismul_m), .B(ecl_mdqctl_n22), .Y(ecl_mdqctl_ismul_m_valid));
OR2X1 exu_U7267(.A(exu_n13431), .B(exu_n14748), .Y(ecl_mdqctl_n17));
AND2X1 exu_U7268(.A(ecl_mdqctl_n23), .B(ecl_mdqctl_mul_done_c0), .Y(ecl_mdqctl_mul_done_valid_c0));
AND2X1 exu_U7269(.A(ecl_mdqctl_n22), .B(exu_n15425), .Y(ecl_mdqctl_n23));
AND2X1 exu_U7270(.A(ecl_mdqctl_mul_done_c1), .B(ecl_mdqctl_n22), .Y(ecl_mdqctl_mul_done_valid_c1));
AND2X1 exu_U7271(.A(exu_n4487), .B(exu_n15458), .Y(ecl_mdqctl_next_mul_done));
AND2X1 exu_U7272(.A(ifu_exu_shiftop_d[2]), .B(ifu_exu_enshift_d), .Y(ecl_shiftop_d[2]));
AND2X1 exu_U7273(.A(ifu_exu_shiftop_d[1]), .B(ifu_exu_enshift_d), .Y(ecl_shiftop_d[1]));
AND2X1 exu_U7274(.A(ifu_exu_shiftop_d[0]), .B(ifu_exu_enshift_d), .Y(ecl_shiftop_d[0]));
AND2X1 exu_U7275(.A(exu_n4085), .B(ecl_mdqctl_n63), .Y(ecl_wb_ccr_setcc_g));
INVX1 exu_U7276(.A(ecl_muls_rs1_31_m_l), .Y(exu_n16612));
OR2X1 exu_U7277(.A(exu_n12102), .B(exu_n13518), .Y(rml_cwp_cwp_thr0_next[2]));
OR2X1 exu_U7278(.A(exu_n12103), .B(exu_n13519), .Y(rml_cwp_cwp_thr0_next[1]));
OR2X1 exu_U7279(.A(exu_n12105), .B(exu_n13521), .Y(rml_cwp_cwp_thr1_next[2]));
OR2X1 exu_U7280(.A(exu_n12106), .B(exu_n13522), .Y(rml_cwp_cwp_thr1_next[1]));
OR2X1 exu_U7281(.A(exu_n12108), .B(exu_n13524), .Y(rml_cwp_cwp_thr2_next[2]));
OR2X1 exu_U7282(.A(exu_n12109), .B(exu_n13525), .Y(rml_cwp_cwp_thr2_next[1]));
OR2X1 exu_U7283(.A(exu_n12111), .B(exu_n13527), .Y(rml_cwp_cwp_thr3_next[2]));
OR2X1 exu_U7284(.A(exu_n12112), .B(exu_n13528), .Y(rml_cwp_cwp_thr3_next[1]));
AND2X1 exu_U7285(.A(exu_n16265), .B(ifu_exu_rd_ffusr_e), .Y(ecl_read_ffusr_e));
AND2X1 exu_U7286(.A(exu_n4949), .B(exu_n15420), .Y(ecl_read_tlusr_e));
OR2X1 exu_U7287(.A(exu_n13495), .B(exu_n14810), .Y(rml_ecl_gl_e[1]));
OR2X1 exu_U7288(.A(exu_n13496), .B(exu_n14811), .Y(rml_ecl_gl_e[0]));
INVX1 exu_U7289(.A(div_u32eql_notequal), .Y(exu_n16436));
OR2X1 exu_U7290(.A(exu_n13396), .B(exu_n14707), .Y(div_u32eql_notequal));
OR2X1 exu_U7291(.A(exu_n13430), .B(exu_n14747), .Y(div_ecl_low32_nonzero));
OR2X1 exu_U7292(.A(exu_n13398), .B(exu_n14709), .Y(rml_cwp_swap_data[8]));
OR2X1 exu_U7293(.A(exu_n13409), .B(exu_n14720), .Y(rml_cwp_spill_wtype_next[2]));
OR2X1 exu_U7294(.A(exu_n13410), .B(exu_n14721), .Y(rml_cwp_spill_wtype_next[1]));
OR2X1 exu_U7295(.A(exu_n13397), .B(exu_n14708), .Y(rml_cwp_spill_wtype_next[0]));
INVX1 exu_U7296(.A(irf_byp_rs2_data_d_l[71]), .Y(byp_ecc_rs2_synd_d[7]));
INVX1 exu_U7297(.A(irf_byp_rs2_data_d_l[70]), .Y(byp_ecc_rs2_synd_d[6]));
INVX1 exu_U7298(.A(irf_byp_rs2_data_d_l[69]), .Y(byp_ecc_rs2_synd_d[5]));
INVX1 exu_U7299(.A(irf_byp_rs2_data_d_l[68]), .Y(byp_ecc_rs2_synd_d[4]));
INVX1 exu_U7300(.A(irf_byp_rs2_data_d_l[67]), .Y(byp_ecc_rs2_synd_d[3]));
INVX1 exu_U7301(.A(irf_byp_rs2_data_d_l[66]), .Y(byp_ecc_rs2_synd_d[2]));
INVX1 exu_U7302(.A(irf_byp_rs2_data_d_l[65]), .Y(byp_ecc_rs2_synd_d[1]));
INVX1 exu_U7303(.A(irf_byp_rs2_data_d_l[64]), .Y(byp_ecc_rs2_synd_d[0]));
INVX1 exu_U7304(.A(irf_byp_rs3_data_d_l[71]), .Y(byp_ecc_rs3_synd_d[7]));
INVX1 exu_U7305(.A(irf_byp_rs3_data_d_l[70]), .Y(byp_ecc_rs3_synd_d[6]));
INVX1 exu_U7306(.A(irf_byp_rs3_data_d_l[69]), .Y(byp_ecc_rs3_synd_d[5]));
INVX1 exu_U7307(.A(irf_byp_rs3_data_d_l[68]), .Y(byp_ecc_rs3_synd_d[4]));
INVX1 exu_U7308(.A(irf_byp_rs3_data_d_l[67]), .Y(byp_ecc_rs3_synd_d[3]));
INVX1 exu_U7309(.A(irf_byp_rs3_data_d_l[66]), .Y(byp_ecc_rs3_synd_d[2]));
INVX1 exu_U7310(.A(irf_byp_rs3_data_d_l[65]), .Y(byp_ecc_rs3_synd_d[1]));
INVX1 exu_U7311(.A(irf_byp_rs3_data_d_l[64]), .Y(byp_ecc_rs3_synd_d[0]));
AND2X1 exu_U7312(.A(exu_n4113), .B(exu_n9106), .Y(ecl_ccr_mux_ccrin0_n1));
AND2X1 exu_U7313(.A(exu_n4115), .B(exu_n9107), .Y(ecl_ccr_mux_ccrin0_n5));
AND2X1 exu_U7314(.A(exu_n4119), .B(exu_n9108), .Y(ecl_ccr_mux_ccrin0_n17));
AND2X1 exu_U7315(.A(exu_n4121), .B(exu_n9109), .Y(ecl_ccr_mux_ccrin0_n21));
AND2X1 exu_U7316(.A(exu_n4123), .B(exu_n9110), .Y(ecl_ccr_mux_ccrin0_n25));
AND2X1 exu_U7317(.A(exu_n4125), .B(exu_n9111), .Y(ecl_ccr_mux_ccrin0_n29));
AND2X1 exu_U7318(.A(exu_n329), .B(exu_n5255), .Y(exu_n18037));
AND2X1 exu_U7319(.A(exu_n331), .B(exu_n5256), .Y(exu_n18041));
AND2X1 exu_U7320(.A(exu_n335), .B(exu_n5257), .Y(exu_n18049));
AND2X1 exu_U7321(.A(exu_n337), .B(exu_n5258), .Y(exu_n18053));
AND2X1 exu_U7322(.A(exu_n339), .B(exu_n5259), .Y(exu_n18057));
AND2X1 exu_U7323(.A(exu_n341), .B(exu_n5260), .Y(exu_n18061));
AND2X1 exu_U7324(.A(exu_n343), .B(exu_n5261), .Y(exu_n18065));
AND2X1 exu_U7325(.A(exu_n345), .B(exu_n5262), .Y(exu_n18069));
AND2X1 exu_U7326(.A(exu_n349), .B(exu_n5263), .Y(exu_n18077));
AND2X1 exu_U7327(.A(exu_n351), .B(exu_n5264), .Y(exu_n18081));
AND2X1 exu_U7328(.A(exu_n353), .B(exu_n5265), .Y(exu_n18085));
AND2X1 exu_U7329(.A(exu_n355), .B(exu_n5266), .Y(exu_n18089));
AND2X1 exu_U7330(.A(exu_n357), .B(exu_n5267), .Y(exu_n18093));
AND2X1 exu_U7331(.A(exu_n359), .B(exu_n5268), .Y(exu_n18097));
AND2X1 exu_U7332(.A(exu_n363), .B(exu_n5269), .Y(exu_n18105));
AND2X1 exu_U7333(.A(exu_n365), .B(exu_n5270), .Y(exu_n18109));
AND2X1 exu_U7334(.A(exu_n367), .B(exu_n5271), .Y(exu_n18113));
AND2X1 exu_U7335(.A(exu_n369), .B(exu_n5272), .Y(exu_n18117));
OR2X1 exu_U7336(.A(exu_n18014), .B(exu_n18013), .Y(ecl_writeback_rdpr_mux2_out[5]));
OR2X1 exu_U7337(.A(exu_n18016), .B(exu_n18015), .Y(ecl_writeback_rdpr_mux2_out[4]));
OR2X1 exu_U7338(.A(exu_n18018), .B(exu_n18017), .Y(ecl_writeback_rdpr_mux2_out[3]));
OR2X1 exu_U7339(.A(exu_n12137), .B(exu_n13553), .Y(ecl_writeback_rdpr_mux2_out[2]));
OR2X1 exu_U7340(.A(exu_n12138), .B(exu_n13554), .Y(ecl_writeback_rdpr_mux2_out[1]));
OR2X1 exu_U7341(.A(exu_n12139), .B(exu_n13555), .Y(ecl_writeback_rdpr_mux2_out[0]));
OR2X1 exu_U7342(.A(exu_n12217), .B(exu_n13629), .Y(div_yreg_next_yreg_thr0[31]));
OR2X1 exu_U7343(.A(exu_n12218), .B(exu_n13630), .Y(div_yreg_next_yreg_thr0[30]));
OR2X1 exu_U7344(.A(exu_n12220), .B(exu_n13632), .Y(div_yreg_next_yreg_thr0[29]));
OR2X1 exu_U7345(.A(exu_n12221), .B(exu_n13633), .Y(div_yreg_next_yreg_thr0[28]));
OR2X1 exu_U7346(.A(exu_n12222), .B(exu_n13634), .Y(div_yreg_next_yreg_thr0[27]));
OR2X1 exu_U7347(.A(exu_n12223), .B(exu_n13635), .Y(div_yreg_next_yreg_thr0[26]));
OR2X1 exu_U7348(.A(exu_n12224), .B(exu_n13636), .Y(div_yreg_next_yreg_thr0[25]));
OR2X1 exu_U7349(.A(exu_n12225), .B(exu_n13637), .Y(div_yreg_next_yreg_thr0[24]));
OR2X1 exu_U7350(.A(exu_n12226), .B(exu_n13638), .Y(div_yreg_next_yreg_thr0[23]));
OR2X1 exu_U7351(.A(exu_n12227), .B(exu_n13639), .Y(div_yreg_next_yreg_thr0[22]));
OR2X1 exu_U7352(.A(exu_n12228), .B(exu_n13640), .Y(div_yreg_next_yreg_thr0[21]));
OR2X1 exu_U7353(.A(exu_n12229), .B(exu_n13641), .Y(div_yreg_next_yreg_thr0[20]));
OR2X1 exu_U7354(.A(exu_n12231), .B(exu_n13643), .Y(div_yreg_next_yreg_thr0[19]));
OR2X1 exu_U7355(.A(exu_n12232), .B(exu_n13644), .Y(div_yreg_next_yreg_thr0[18]));
OR2X1 exu_U7356(.A(exu_n12233), .B(exu_n13645), .Y(div_yreg_next_yreg_thr0[17]));
OR2X1 exu_U7357(.A(exu_n12234), .B(exu_n13646), .Y(div_yreg_next_yreg_thr0[16]));
OR2X1 exu_U7358(.A(exu_n12235), .B(exu_n13647), .Y(div_yreg_next_yreg_thr0[15]));
OR2X1 exu_U7359(.A(exu_n12236), .B(exu_n13648), .Y(div_yreg_next_yreg_thr0[14]));
OR2X1 exu_U7360(.A(exu_n12237), .B(exu_n13649), .Y(div_yreg_next_yreg_thr0[13]));
OR2X1 exu_U7361(.A(exu_n12238), .B(exu_n13650), .Y(div_yreg_next_yreg_thr0[12]));
OR2X1 exu_U7362(.A(exu_n12239), .B(exu_n13651), .Y(div_yreg_next_yreg_thr0[11]));
OR2X1 exu_U7363(.A(exu_n12240), .B(exu_n13652), .Y(div_yreg_next_yreg_thr0[10]));
OR2X1 exu_U7364(.A(exu_n12210), .B(exu_n13622), .Y(div_yreg_next_yreg_thr0[9]));
OR2X1 exu_U7365(.A(exu_n12211), .B(exu_n13623), .Y(div_yreg_next_yreg_thr0[8]));
OR2X1 exu_U7366(.A(exu_n12212), .B(exu_n13624), .Y(div_yreg_next_yreg_thr0[7]));
OR2X1 exu_U7367(.A(exu_n12213), .B(exu_n13625), .Y(div_yreg_next_yreg_thr0[6]));
OR2X1 exu_U7368(.A(exu_n12214), .B(exu_n13626), .Y(div_yreg_next_yreg_thr0[5]));
OR2X1 exu_U7369(.A(exu_n12215), .B(exu_n13627), .Y(div_yreg_next_yreg_thr0[4]));
OR2X1 exu_U7370(.A(exu_n12216), .B(exu_n13628), .Y(div_yreg_next_yreg_thr0[3]));
OR2X1 exu_U7371(.A(exu_n12219), .B(exu_n13631), .Y(div_yreg_next_yreg_thr0[2]));
OR2X1 exu_U7372(.A(exu_n12230), .B(exu_n13642), .Y(div_yreg_next_yreg_thr0[1]));
OR2X1 exu_U7373(.A(exu_n12241), .B(exu_n13653), .Y(div_yreg_next_yreg_thr0[0]));
OR2X1 exu_U7374(.A(exu_n12249), .B(exu_n13661), .Y(div_yreg_next_yreg_thr1[31]));
OR2X1 exu_U7375(.A(exu_n12250), .B(exu_n13662), .Y(div_yreg_next_yreg_thr1[30]));
OR2X1 exu_U7376(.A(exu_n12252), .B(exu_n13664), .Y(div_yreg_next_yreg_thr1[29]));
OR2X1 exu_U7377(.A(exu_n12253), .B(exu_n13665), .Y(div_yreg_next_yreg_thr1[28]));
OR2X1 exu_U7378(.A(exu_n12254), .B(exu_n13666), .Y(div_yreg_next_yreg_thr1[27]));
OR2X1 exu_U7379(.A(exu_n12255), .B(exu_n13667), .Y(div_yreg_next_yreg_thr1[26]));
OR2X1 exu_U7380(.A(exu_n12256), .B(exu_n13668), .Y(div_yreg_next_yreg_thr1[25]));
OR2X1 exu_U7381(.A(exu_n12257), .B(exu_n13669), .Y(div_yreg_next_yreg_thr1[24]));
OR2X1 exu_U7382(.A(exu_n12258), .B(exu_n13670), .Y(div_yreg_next_yreg_thr1[23]));
OR2X1 exu_U7383(.A(exu_n12259), .B(exu_n13671), .Y(div_yreg_next_yreg_thr1[22]));
OR2X1 exu_U7384(.A(exu_n12260), .B(exu_n13672), .Y(div_yreg_next_yreg_thr1[21]));
OR2X1 exu_U7385(.A(exu_n12261), .B(exu_n13673), .Y(div_yreg_next_yreg_thr1[20]));
OR2X1 exu_U7386(.A(exu_n12263), .B(exu_n13675), .Y(div_yreg_next_yreg_thr1[19]));
OR2X1 exu_U7387(.A(exu_n12264), .B(exu_n13676), .Y(div_yreg_next_yreg_thr1[18]));
OR2X1 exu_U7388(.A(exu_n12265), .B(exu_n13677), .Y(div_yreg_next_yreg_thr1[17]));
OR2X1 exu_U7389(.A(exu_n12266), .B(exu_n13678), .Y(div_yreg_next_yreg_thr1[16]));
OR2X1 exu_U7390(.A(exu_n12267), .B(exu_n13679), .Y(div_yreg_next_yreg_thr1[15]));
OR2X1 exu_U7391(.A(exu_n12268), .B(exu_n13680), .Y(div_yreg_next_yreg_thr1[14]));
OR2X1 exu_U7392(.A(exu_n12269), .B(exu_n13681), .Y(div_yreg_next_yreg_thr1[13]));
OR2X1 exu_U7393(.A(exu_n12270), .B(exu_n13682), .Y(div_yreg_next_yreg_thr1[12]));
OR2X1 exu_U7394(.A(exu_n12271), .B(exu_n13683), .Y(div_yreg_next_yreg_thr1[11]));
OR2X1 exu_U7395(.A(exu_n12272), .B(exu_n13684), .Y(div_yreg_next_yreg_thr1[10]));
OR2X1 exu_U7396(.A(exu_n12242), .B(exu_n13654), .Y(div_yreg_next_yreg_thr1[9]));
OR2X1 exu_U7397(.A(exu_n12243), .B(exu_n13655), .Y(div_yreg_next_yreg_thr1[8]));
OR2X1 exu_U7398(.A(exu_n12244), .B(exu_n13656), .Y(div_yreg_next_yreg_thr1[7]));
OR2X1 exu_U7399(.A(exu_n12245), .B(exu_n13657), .Y(div_yreg_next_yreg_thr1[6]));
OR2X1 exu_U7400(.A(exu_n12246), .B(exu_n13658), .Y(div_yreg_next_yreg_thr1[5]));
OR2X1 exu_U7401(.A(exu_n12247), .B(exu_n13659), .Y(div_yreg_next_yreg_thr1[4]));
OR2X1 exu_U7402(.A(exu_n12248), .B(exu_n13660), .Y(div_yreg_next_yreg_thr1[3]));
OR2X1 exu_U7403(.A(exu_n12251), .B(exu_n13663), .Y(div_yreg_next_yreg_thr1[2]));
OR2X1 exu_U7404(.A(exu_n12262), .B(exu_n13674), .Y(div_yreg_next_yreg_thr1[1]));
OR2X1 exu_U7405(.A(exu_n12273), .B(exu_n13685), .Y(div_yreg_next_yreg_thr1[0]));
OR2X1 exu_U7406(.A(exu_n12281), .B(exu_n13693), .Y(div_yreg_next_yreg_thr2[31]));
OR2X1 exu_U7407(.A(exu_n12282), .B(exu_n13694), .Y(div_yreg_next_yreg_thr2[30]));
OR2X1 exu_U7408(.A(exu_n12284), .B(exu_n13696), .Y(div_yreg_next_yreg_thr2[29]));
OR2X1 exu_U7409(.A(exu_n12285), .B(exu_n13697), .Y(div_yreg_next_yreg_thr2[28]));
OR2X1 exu_U7410(.A(exu_n12286), .B(exu_n13698), .Y(div_yreg_next_yreg_thr2[27]));
OR2X1 exu_U7411(.A(exu_n12287), .B(exu_n13699), .Y(div_yreg_next_yreg_thr2[26]));
OR2X1 exu_U7412(.A(exu_n12288), .B(exu_n13700), .Y(div_yreg_next_yreg_thr2[25]));
OR2X1 exu_U7413(.A(exu_n12289), .B(exu_n13701), .Y(div_yreg_next_yreg_thr2[24]));
OR2X1 exu_U7414(.A(exu_n12290), .B(exu_n13702), .Y(div_yreg_next_yreg_thr2[23]));
OR2X1 exu_U7415(.A(exu_n12291), .B(exu_n13703), .Y(div_yreg_next_yreg_thr2[22]));
OR2X1 exu_U7416(.A(exu_n12292), .B(exu_n13704), .Y(div_yreg_next_yreg_thr2[21]));
OR2X1 exu_U7417(.A(exu_n12293), .B(exu_n13705), .Y(div_yreg_next_yreg_thr2[20]));
OR2X1 exu_U7418(.A(exu_n12295), .B(exu_n13707), .Y(div_yreg_next_yreg_thr2[19]));
OR2X1 exu_U7419(.A(exu_n12296), .B(exu_n13708), .Y(div_yreg_next_yreg_thr2[18]));
OR2X1 exu_U7420(.A(exu_n12297), .B(exu_n13709), .Y(div_yreg_next_yreg_thr2[17]));
OR2X1 exu_U7421(.A(exu_n12298), .B(exu_n13710), .Y(div_yreg_next_yreg_thr2[16]));
OR2X1 exu_U7422(.A(exu_n12299), .B(exu_n13711), .Y(div_yreg_next_yreg_thr2[15]));
OR2X1 exu_U7423(.A(exu_n12300), .B(exu_n13712), .Y(div_yreg_next_yreg_thr2[14]));
OR2X1 exu_U7424(.A(exu_n12301), .B(exu_n13713), .Y(div_yreg_next_yreg_thr2[13]));
OR2X1 exu_U7425(.A(exu_n12302), .B(exu_n13714), .Y(div_yreg_next_yreg_thr2[12]));
OR2X1 exu_U7426(.A(exu_n12303), .B(exu_n13715), .Y(div_yreg_next_yreg_thr2[11]));
OR2X1 exu_U7427(.A(exu_n12304), .B(exu_n13716), .Y(div_yreg_next_yreg_thr2[10]));
OR2X1 exu_U7428(.A(exu_n12274), .B(exu_n13686), .Y(div_yreg_next_yreg_thr2[9]));
OR2X1 exu_U7429(.A(exu_n12275), .B(exu_n13687), .Y(div_yreg_next_yreg_thr2[8]));
OR2X1 exu_U7430(.A(exu_n12276), .B(exu_n13688), .Y(div_yreg_next_yreg_thr2[7]));
OR2X1 exu_U7431(.A(exu_n12277), .B(exu_n13689), .Y(div_yreg_next_yreg_thr2[6]));
OR2X1 exu_U7432(.A(exu_n12278), .B(exu_n13690), .Y(div_yreg_next_yreg_thr2[5]));
OR2X1 exu_U7433(.A(exu_n12279), .B(exu_n13691), .Y(div_yreg_next_yreg_thr2[4]));
OR2X1 exu_U7434(.A(exu_n12280), .B(exu_n13692), .Y(div_yreg_next_yreg_thr2[3]));
OR2X1 exu_U7435(.A(exu_n12283), .B(exu_n13695), .Y(div_yreg_next_yreg_thr2[2]));
OR2X1 exu_U7436(.A(exu_n12294), .B(exu_n13706), .Y(div_yreg_next_yreg_thr2[1]));
OR2X1 exu_U7437(.A(exu_n12305), .B(exu_n13717), .Y(div_yreg_next_yreg_thr2[0]));
OR2X1 exu_U7438(.A(exu_n12313), .B(exu_n13725), .Y(div_yreg_next_yreg_thr3[31]));
OR2X1 exu_U7439(.A(exu_n12314), .B(exu_n13726), .Y(div_yreg_next_yreg_thr3[30]));
OR2X1 exu_U7440(.A(exu_n12316), .B(exu_n13728), .Y(div_yreg_next_yreg_thr3[29]));
OR2X1 exu_U7441(.A(exu_n12317), .B(exu_n13729), .Y(div_yreg_next_yreg_thr3[28]));
OR2X1 exu_U7442(.A(exu_n12318), .B(exu_n13730), .Y(div_yreg_next_yreg_thr3[27]));
OR2X1 exu_U7443(.A(exu_n12319), .B(exu_n13731), .Y(div_yreg_next_yreg_thr3[26]));
OR2X1 exu_U7444(.A(exu_n12320), .B(exu_n13732), .Y(div_yreg_next_yreg_thr3[25]));
OR2X1 exu_U7445(.A(exu_n12321), .B(exu_n13733), .Y(div_yreg_next_yreg_thr3[24]));
OR2X1 exu_U7446(.A(exu_n12322), .B(exu_n13734), .Y(div_yreg_next_yreg_thr3[23]));
OR2X1 exu_U7447(.A(exu_n12323), .B(exu_n13735), .Y(div_yreg_next_yreg_thr3[22]));
OR2X1 exu_U7448(.A(exu_n12324), .B(exu_n13736), .Y(div_yreg_next_yreg_thr3[21]));
OR2X1 exu_U7449(.A(exu_n12325), .B(exu_n13737), .Y(div_yreg_next_yreg_thr3[20]));
OR2X1 exu_U7450(.A(exu_n12327), .B(exu_n13739), .Y(div_yreg_next_yreg_thr3[19]));
OR2X1 exu_U7451(.A(exu_n12328), .B(exu_n13740), .Y(div_yreg_next_yreg_thr3[18]));
OR2X1 exu_U7452(.A(exu_n12329), .B(exu_n13741), .Y(div_yreg_next_yreg_thr3[17]));
OR2X1 exu_U7453(.A(exu_n12330), .B(exu_n13742), .Y(div_yreg_next_yreg_thr3[16]));
OR2X1 exu_U7454(.A(exu_n12331), .B(exu_n13743), .Y(div_yreg_next_yreg_thr3[15]));
OR2X1 exu_U7455(.A(exu_n12332), .B(exu_n13744), .Y(div_yreg_next_yreg_thr3[14]));
OR2X1 exu_U7456(.A(exu_n12333), .B(exu_n13745), .Y(div_yreg_next_yreg_thr3[13]));
OR2X1 exu_U7457(.A(exu_n12334), .B(exu_n13746), .Y(div_yreg_next_yreg_thr3[12]));
OR2X1 exu_U7458(.A(exu_n12335), .B(exu_n13747), .Y(div_yreg_next_yreg_thr3[11]));
OR2X1 exu_U7459(.A(exu_n12336), .B(exu_n13748), .Y(div_yreg_next_yreg_thr3[10]));
OR2X1 exu_U7460(.A(exu_n12306), .B(exu_n13718), .Y(div_yreg_next_yreg_thr3[9]));
OR2X1 exu_U7461(.A(exu_n12307), .B(exu_n13719), .Y(div_yreg_next_yreg_thr3[8]));
OR2X1 exu_U7462(.A(exu_n12308), .B(exu_n13720), .Y(div_yreg_next_yreg_thr3[7]));
OR2X1 exu_U7463(.A(exu_n12309), .B(exu_n13721), .Y(div_yreg_next_yreg_thr3[6]));
OR2X1 exu_U7464(.A(exu_n12310), .B(exu_n13722), .Y(div_yreg_next_yreg_thr3[5]));
OR2X1 exu_U7465(.A(exu_n12311), .B(exu_n13723), .Y(div_yreg_next_yreg_thr3[4]));
OR2X1 exu_U7466(.A(exu_n12312), .B(exu_n13724), .Y(div_yreg_next_yreg_thr3[3]));
OR2X1 exu_U7467(.A(exu_n12315), .B(exu_n13727), .Y(div_yreg_next_yreg_thr3[2]));
OR2X1 exu_U7468(.A(exu_n12326), .B(exu_n13738), .Y(div_yreg_next_yreg_thr3[1]));
OR2X1 exu_U7469(.A(exu_n12337), .B(exu_n13749), .Y(div_yreg_next_yreg_thr3[0]));
OR2X1 exu_U7470(.A(bypass_ifu_exu_sr_mux_n240), .B(exu_n14783), .Y(bypass_rd_data_e[31]));
OR2X1 exu_U7471(.A(bypass_ifu_exu_sr_mux_n246), .B(exu_n14784), .Y(bypass_rd_data_e[30]));
OR2X1 exu_U7472(.A(bypass_ifu_exu_sr_mux_n258), .B(exu_n14786), .Y(bypass_rd_data_e[29]));
OR2X1 exu_U7473(.A(bypass_ifu_exu_sr_mux_n264), .B(exu_n14787), .Y(bypass_rd_data_e[28]));
OR2X1 exu_U7474(.A(bypass_ifu_exu_sr_mux_n270), .B(exu_n14788), .Y(bypass_rd_data_e[27]));
OR2X1 exu_U7475(.A(bypass_ifu_exu_sr_mux_n276), .B(exu_n14789), .Y(bypass_rd_data_e[26]));
OR2X1 exu_U7476(.A(bypass_ifu_exu_sr_mux_n282), .B(exu_n14790), .Y(bypass_rd_data_e[25]));
OR2X1 exu_U7477(.A(bypass_ifu_exu_sr_mux_n288), .B(exu_n14791), .Y(bypass_rd_data_e[24]));
OR2X1 exu_U7478(.A(bypass_ifu_exu_sr_mux_n294), .B(exu_n14792), .Y(bypass_rd_data_e[23]));
OR2X1 exu_U7479(.A(bypass_ifu_exu_sr_mux_n300), .B(exu_n14793), .Y(bypass_rd_data_e[22]));
OR2X1 exu_U7480(.A(bypass_ifu_exu_sr_mux_n306), .B(exu_n14794), .Y(bypass_rd_data_e[21]));
OR2X1 exu_U7481(.A(bypass_ifu_exu_sr_mux_n312), .B(exu_n14795), .Y(bypass_rd_data_e[20]));
OR2X1 exu_U7482(.A(bypass_ifu_exu_sr_mux_n324), .B(exu_n14797), .Y(bypass_rd_data_e[19]));
OR2X1 exu_U7483(.A(bypass_ifu_exu_sr_mux_n330), .B(exu_n14798), .Y(bypass_rd_data_e[18]));
OR2X1 exu_U7484(.A(bypass_ifu_exu_sr_mux_n336), .B(exu_n14799), .Y(bypass_rd_data_e[17]));
OR2X1 exu_U7485(.A(bypass_ifu_exu_sr_mux_n342), .B(exu_n14800), .Y(bypass_rd_data_e[16]));
OR2X1 exu_U7486(.A(bypass_ifu_exu_sr_mux_n348), .B(exu_n14801), .Y(bypass_rd_data_e[15]));
OR2X1 exu_U7487(.A(bypass_ifu_exu_sr_mux_n354), .B(exu_n14802), .Y(bypass_rd_data_e[14]));
OR2X1 exu_U7488(.A(bypass_ifu_exu_sr_mux_n360), .B(exu_n14803), .Y(bypass_rd_data_e[13]));
OR2X1 exu_U7489(.A(bypass_ifu_exu_sr_mux_n366), .B(exu_n14804), .Y(bypass_rd_data_e[12]));
OR2X1 exu_U7490(.A(bypass_ifu_exu_sr_mux_n372), .B(exu_n14805), .Y(bypass_rd_data_e[11]));
OR2X1 exu_U7491(.A(bypass_ifu_exu_sr_mux_n378), .B(exu_n14806), .Y(bypass_rd_data_e[10]));
OR2X1 exu_U7492(.A(bypass_ifu_exu_sr_mux_n6), .B(exu_n14776), .Y(bypass_rd_data_e[9]));
OR2X1 exu_U7493(.A(bypass_ifu_exu_sr_mux_n12), .B(exu_n14777), .Y(bypass_rd_data_e[8]));
OR2X1 exu_U7494(.A(exu_n13487), .B(exu_n14778), .Y(bypass_rd_data_e[7]));
OR2X1 exu_U7495(.A(exu_n13488), .B(exu_n14779), .Y(bypass_rd_data_e[6]));
OR2X1 exu_U7496(.A(exu_n13489), .B(exu_n14780), .Y(bypass_rd_data_e[5]));
OR2X1 exu_U7497(.A(exu_n13490), .B(exu_n14781), .Y(bypass_rd_data_e[4]));
OR2X1 exu_U7498(.A(exu_n13491), .B(exu_n14782), .Y(bypass_rd_data_e[3]));
OR2X1 exu_U7499(.A(exu_n13492), .B(exu_n14785), .Y(bypass_rd_data_e[2]));
OR2X1 exu_U7500(.A(exu_n13493), .B(exu_n14796), .Y(bypass_rd_data_e[1]));
OR2X1 exu_U7501(.A(exu_n13494), .B(exu_n14807), .Y(bypass_rd_data_e[0]));
INVX1 exu_U7502(.A(exu_n16171), .Y(exu_n16179));
INVX1 exu_U7503(.A(exu_n16171), .Y(exu_n16180));
INVX1 exu_U7504(.A(exu_n16171), .Y(exu_n16181));
INVX1 exu_U7505(.A(exu_n16171), .Y(exu_n16182));
INVX1 exu_U7506(.A(exu_n16171), .Y(exu_n16183));
INVX1 exu_U7507(.A(exu_n16171), .Y(exu_n16184));
OR2X1 exu_U7508(.A(exu_n12470), .B(exu_n13882), .Y(bypass_byp_alu_rs1_data_d[63]));
OR2X1 exu_U7509(.A(exu_n12471), .B(exu_n13883), .Y(bypass_byp_alu_rs1_data_d[62]));
OR2X1 exu_U7510(.A(exu_n12472), .B(exu_n13884), .Y(bypass_byp_alu_rs1_data_d[61]));
OR2X1 exu_U7511(.A(exu_n12473), .B(exu_n13885), .Y(bypass_byp_alu_rs1_data_d[60]));
OR2X1 exu_U7512(.A(exu_n12475), .B(exu_n13887), .Y(bypass_byp_alu_rs1_data_d[59]));
OR2X1 exu_U7513(.A(exu_n12476), .B(exu_n13888), .Y(bypass_byp_alu_rs1_data_d[58]));
OR2X1 exu_U7514(.A(exu_n12477), .B(exu_n13889), .Y(bypass_byp_alu_rs1_data_d[57]));
OR2X1 exu_U7515(.A(exu_n12478), .B(exu_n13890), .Y(bypass_byp_alu_rs1_data_d[56]));
OR2X1 exu_U7516(.A(exu_n12479), .B(exu_n13891), .Y(bypass_byp_alu_rs1_data_d[55]));
OR2X1 exu_U7517(.A(exu_n12480), .B(exu_n13892), .Y(bypass_byp_alu_rs1_data_d[54]));
OR2X1 exu_U7518(.A(exu_n12481), .B(exu_n13893), .Y(bypass_byp_alu_rs1_data_d[53]));
OR2X1 exu_U7519(.A(exu_n12482), .B(exu_n13894), .Y(bypass_byp_alu_rs1_data_d[52]));
OR2X1 exu_U7520(.A(exu_n12483), .B(exu_n13895), .Y(bypass_byp_alu_rs1_data_d[51]));
OR2X1 exu_U7521(.A(exu_n12484), .B(exu_n13896), .Y(bypass_byp_alu_rs1_data_d[50]));
OR2X1 exu_U7522(.A(exu_n12486), .B(exu_n13898), .Y(bypass_byp_alu_rs1_data_d[49]));
OR2X1 exu_U7523(.A(exu_n12487), .B(exu_n13899), .Y(bypass_byp_alu_rs1_data_d[48]));
OR2X1 exu_U7524(.A(exu_n12488), .B(exu_n13900), .Y(bypass_byp_alu_rs1_data_d[47]));
OR2X1 exu_U7525(.A(exu_n12489), .B(exu_n13901), .Y(bypass_byp_alu_rs1_data_d[46]));
OR2X1 exu_U7526(.A(exu_n12490), .B(exu_n13902), .Y(bypass_byp_alu_rs1_data_d[45]));
OR2X1 exu_U7527(.A(exu_n12491), .B(exu_n13903), .Y(bypass_byp_alu_rs1_data_d[44]));
OR2X1 exu_U7528(.A(exu_n12492), .B(exu_n13904), .Y(bypass_byp_alu_rs1_data_d[43]));
OR2X1 exu_U7529(.A(exu_n12493), .B(exu_n13905), .Y(bypass_byp_alu_rs1_data_d[42]));
OR2X1 exu_U7530(.A(exu_n12494), .B(exu_n13906), .Y(bypass_byp_alu_rs1_data_d[41]));
OR2X1 exu_U7531(.A(exu_n12495), .B(exu_n13907), .Y(bypass_byp_alu_rs1_data_d[40]));
OR2X1 exu_U7532(.A(exu_n12497), .B(exu_n13909), .Y(bypass_byp_alu_rs1_data_d[39]));
OR2X1 exu_U7533(.A(exu_n12498), .B(exu_n13910), .Y(bypass_byp_alu_rs1_data_d[38]));
OR2X1 exu_U7534(.A(exu_n12499), .B(exu_n13911), .Y(bypass_byp_alu_rs1_data_d[37]));
OR2X1 exu_U7535(.A(exu_n12500), .B(exu_n13912), .Y(bypass_byp_alu_rs1_data_d[36]));
OR2X1 exu_U7536(.A(exu_n12501), .B(exu_n13913), .Y(bypass_byp_alu_rs1_data_d[35]));
OR2X1 exu_U7537(.A(exu_n12502), .B(exu_n13914), .Y(bypass_byp_alu_rs1_data_d[34]));
OR2X1 exu_U7538(.A(exu_n12503), .B(exu_n13915), .Y(bypass_byp_alu_rs1_data_d[33]));
OR2X1 exu_U7539(.A(exu_n12504), .B(exu_n13916), .Y(bypass_byp_alu_rs1_data_d[32]));
OR2X1 exu_U7540(.A(exu_n12505), .B(exu_n13917), .Y(bypass_byp_alu_rs1_data_d[31]));
OR2X1 exu_U7541(.A(exu_n12506), .B(exu_n13918), .Y(bypass_byp_alu_rs1_data_d[30]));
OR2X1 exu_U7542(.A(exu_n12508), .B(exu_n13920), .Y(bypass_byp_alu_rs1_data_d[29]));
OR2X1 exu_U7543(.A(exu_n12509), .B(exu_n13921), .Y(bypass_byp_alu_rs1_data_d[28]));
OR2X1 exu_U7544(.A(exu_n12510), .B(exu_n13922), .Y(bypass_byp_alu_rs1_data_d[27]));
OR2X1 exu_U7545(.A(exu_n12511), .B(exu_n13923), .Y(bypass_byp_alu_rs1_data_d[26]));
OR2X1 exu_U7546(.A(exu_n12512), .B(exu_n13924), .Y(bypass_byp_alu_rs1_data_d[25]));
OR2X1 exu_U7547(.A(exu_n12513), .B(exu_n13925), .Y(bypass_byp_alu_rs1_data_d[24]));
OR2X1 exu_U7548(.A(exu_n12514), .B(exu_n13926), .Y(bypass_byp_alu_rs1_data_d[23]));
OR2X1 exu_U7549(.A(exu_n12515), .B(exu_n13927), .Y(bypass_byp_alu_rs1_data_d[22]));
OR2X1 exu_U7550(.A(exu_n12516), .B(exu_n13928), .Y(bypass_byp_alu_rs1_data_d[21]));
OR2X1 exu_U7551(.A(exu_n12517), .B(exu_n13929), .Y(bypass_byp_alu_rs1_data_d[20]));
OR2X1 exu_U7552(.A(exu_n12519), .B(exu_n13931), .Y(bypass_byp_alu_rs1_data_d[19]));
OR2X1 exu_U7553(.A(exu_n12520), .B(exu_n13932), .Y(bypass_byp_alu_rs1_data_d[18]));
OR2X1 exu_U7554(.A(exu_n12521), .B(exu_n13933), .Y(bypass_byp_alu_rs1_data_d[17]));
OR2X1 exu_U7555(.A(exu_n12522), .B(exu_n13934), .Y(bypass_byp_alu_rs1_data_d[16]));
OR2X1 exu_U7556(.A(exu_n12523), .B(exu_n13935), .Y(bypass_byp_alu_rs1_data_d[15]));
OR2X1 exu_U7557(.A(exu_n12524), .B(exu_n13936), .Y(bypass_byp_alu_rs1_data_d[14]));
OR2X1 exu_U7558(.A(exu_n12525), .B(exu_n13937), .Y(bypass_byp_alu_rs1_data_d[13]));
OR2X1 exu_U7559(.A(exu_n12526), .B(exu_n13938), .Y(bypass_byp_alu_rs1_data_d[12]));
OR2X1 exu_U7560(.A(exu_n12527), .B(exu_n13939), .Y(bypass_byp_alu_rs1_data_d[11]));
OR2X1 exu_U7561(.A(exu_n12528), .B(exu_n13940), .Y(bypass_byp_alu_rs1_data_d[10]));
OR2X1 exu_U7562(.A(exu_n12466), .B(exu_n13878), .Y(bypass_byp_alu_rs1_data_d[9]));
OR2X1 exu_U7563(.A(exu_n12467), .B(exu_n13879), .Y(bypass_byp_alu_rs1_data_d[8]));
OR2X1 exu_U7564(.A(exu_n12468), .B(exu_n13880), .Y(bypass_byp_alu_rs1_data_d[7]));
OR2X1 exu_U7565(.A(exu_n12469), .B(exu_n13881), .Y(bypass_byp_alu_rs1_data_d[6]));
OR2X1 exu_U7566(.A(exu_n12474), .B(exu_n13886), .Y(bypass_byp_alu_rs1_data_d[5]));
OR2X1 exu_U7567(.A(exu_n12485), .B(exu_n13897), .Y(bypass_byp_alu_rs1_data_d[4]));
OR2X1 exu_U7568(.A(exu_n12496), .B(exu_n13908), .Y(bypass_byp_alu_rs1_data_d[3]));
OR2X1 exu_U7569(.A(exu_n12507), .B(exu_n13919), .Y(bypass_byp_alu_rs1_data_d[2]));
OR2X1 exu_U7570(.A(exu_n12518), .B(exu_n13930), .Y(bypass_byp_alu_rs1_data_d[1]));
OR2X1 exu_U7571(.A(exu_n12529), .B(exu_n13941), .Y(bypass_byp_alu_rs1_data_d[0]));
OR2X1 exu_U7572(.A(exu_n12726), .B(exu_n14074), .Y(bypass_byp_alu_rs2_data_d[63]));
OR2X1 exu_U7573(.A(exu_n12727), .B(exu_n14075), .Y(bypass_byp_alu_rs2_data_d[62]));
OR2X1 exu_U7574(.A(exu_n12728), .B(exu_n14076), .Y(bypass_byp_alu_rs2_data_d[61]));
OR2X1 exu_U7575(.A(exu_n12729), .B(exu_n14077), .Y(bypass_byp_alu_rs2_data_d[60]));
OR2X1 exu_U7576(.A(exu_n12731), .B(exu_n14079), .Y(bypass_byp_alu_rs2_data_d[59]));
OR2X1 exu_U7577(.A(exu_n12732), .B(exu_n14080), .Y(bypass_byp_alu_rs2_data_d[58]));
OR2X1 exu_U7578(.A(exu_n12733), .B(exu_n14081), .Y(bypass_byp_alu_rs2_data_d[57]));
OR2X1 exu_U7579(.A(exu_n12734), .B(exu_n14082), .Y(bypass_byp_alu_rs2_data_d[56]));
OR2X1 exu_U7580(.A(exu_n12735), .B(exu_n14083), .Y(bypass_byp_alu_rs2_data_d[55]));
OR2X1 exu_U7581(.A(exu_n12736), .B(exu_n14084), .Y(bypass_byp_alu_rs2_data_d[54]));
OR2X1 exu_U7582(.A(exu_n12737), .B(exu_n14085), .Y(bypass_byp_alu_rs2_data_d[53]));
OR2X1 exu_U7583(.A(exu_n12738), .B(exu_n14086), .Y(bypass_byp_alu_rs2_data_d[52]));
OR2X1 exu_U7584(.A(exu_n12739), .B(exu_n14087), .Y(bypass_byp_alu_rs2_data_d[51]));
OR2X1 exu_U7585(.A(exu_n12740), .B(exu_n14088), .Y(bypass_byp_alu_rs2_data_d[50]));
OR2X1 exu_U7586(.A(exu_n12742), .B(exu_n14090), .Y(bypass_byp_alu_rs2_data_d[49]));
OR2X1 exu_U7587(.A(exu_n12743), .B(exu_n14091), .Y(bypass_byp_alu_rs2_data_d[48]));
OR2X1 exu_U7588(.A(exu_n12744), .B(exu_n14092), .Y(bypass_byp_alu_rs2_data_d[47]));
OR2X1 exu_U7589(.A(exu_n12745), .B(exu_n14093), .Y(bypass_byp_alu_rs2_data_d[46]));
OR2X1 exu_U7590(.A(exu_n12746), .B(exu_n14094), .Y(bypass_byp_alu_rs2_data_d[45]));
OR2X1 exu_U7591(.A(exu_n12747), .B(exu_n14095), .Y(bypass_byp_alu_rs2_data_d[44]));
OR2X1 exu_U7592(.A(exu_n12748), .B(exu_n14096), .Y(bypass_byp_alu_rs2_data_d[43]));
OR2X1 exu_U7593(.A(exu_n12749), .B(exu_n14097), .Y(bypass_byp_alu_rs2_data_d[42]));
OR2X1 exu_U7594(.A(exu_n12750), .B(exu_n14098), .Y(bypass_byp_alu_rs2_data_d[41]));
OR2X1 exu_U7595(.A(exu_n12751), .B(exu_n14099), .Y(bypass_byp_alu_rs2_data_d[40]));
OR2X1 exu_U7596(.A(exu_n12753), .B(exu_n14101), .Y(bypass_byp_alu_rs2_data_d[39]));
OR2X1 exu_U7597(.A(exu_n12754), .B(exu_n14102), .Y(bypass_byp_alu_rs2_data_d[38]));
OR2X1 exu_U7598(.A(exu_n12755), .B(exu_n14103), .Y(bypass_byp_alu_rs2_data_d[37]));
OR2X1 exu_U7599(.A(exu_n12756), .B(exu_n14104), .Y(bypass_byp_alu_rs2_data_d[36]));
OR2X1 exu_U7600(.A(exu_n12757), .B(exu_n14105), .Y(bypass_byp_alu_rs2_data_d[35]));
OR2X1 exu_U7601(.A(exu_n12758), .B(exu_n14106), .Y(bypass_byp_alu_rs2_data_d[34]));
OR2X1 exu_U7602(.A(exu_n12759), .B(exu_n14107), .Y(bypass_byp_alu_rs2_data_d[33]));
OR2X1 exu_U7603(.A(exu_n12760), .B(exu_n14108), .Y(bypass_byp_alu_rs2_data_d[32]));
OR2X1 exu_U7604(.A(exu_n12761), .B(exu_n14109), .Y(bypass_byp_alu_rs2_data_d[31]));
OR2X1 exu_U7605(.A(exu_n12762), .B(exu_n14110), .Y(bypass_byp_alu_rs2_data_d[30]));
OR2X1 exu_U7606(.A(exu_n12764), .B(exu_n14112), .Y(bypass_byp_alu_rs2_data_d[29]));
OR2X1 exu_U7607(.A(exu_n12765), .B(exu_n14113), .Y(bypass_byp_alu_rs2_data_d[28]));
OR2X1 exu_U7608(.A(exu_n12766), .B(exu_n14114), .Y(bypass_byp_alu_rs2_data_d[27]));
OR2X1 exu_U7609(.A(exu_n12767), .B(exu_n14115), .Y(bypass_byp_alu_rs2_data_d[26]));
OR2X1 exu_U7610(.A(exu_n12768), .B(exu_n14116), .Y(bypass_byp_alu_rs2_data_d[25]));
OR2X1 exu_U7611(.A(exu_n12769), .B(exu_n14117), .Y(bypass_byp_alu_rs2_data_d[24]));
OR2X1 exu_U7612(.A(exu_n12770), .B(exu_n14118), .Y(bypass_byp_alu_rs2_data_d[23]));
OR2X1 exu_U7613(.A(exu_n12771), .B(exu_n14119), .Y(bypass_byp_alu_rs2_data_d[22]));
OR2X1 exu_U7614(.A(exu_n12772), .B(exu_n14120), .Y(bypass_byp_alu_rs2_data_d[21]));
OR2X1 exu_U7615(.A(exu_n12773), .B(exu_n14121), .Y(bypass_byp_alu_rs2_data_d[20]));
OR2X1 exu_U7616(.A(exu_n12775), .B(exu_n14123), .Y(bypass_byp_alu_rs2_data_d[19]));
OR2X1 exu_U7617(.A(exu_n12776), .B(exu_n14124), .Y(bypass_byp_alu_rs2_data_d[18]));
OR2X1 exu_U7618(.A(exu_n12777), .B(exu_n14125), .Y(bypass_byp_alu_rs2_data_d[17]));
OR2X1 exu_U7619(.A(exu_n12778), .B(exu_n14126), .Y(bypass_byp_alu_rs2_data_d[16]));
OR2X1 exu_U7620(.A(exu_n12779), .B(exu_n14127), .Y(bypass_byp_alu_rs2_data_d[15]));
OR2X1 exu_U7621(.A(exu_n12780), .B(exu_n14128), .Y(bypass_byp_alu_rs2_data_d[14]));
OR2X1 exu_U7622(.A(exu_n12781), .B(exu_n14129), .Y(bypass_byp_alu_rs2_data_d[13]));
OR2X1 exu_U7623(.A(exu_n12782), .B(exu_n14130), .Y(bypass_byp_alu_rs2_data_d[12]));
OR2X1 exu_U7624(.A(exu_n12783), .B(exu_n14131), .Y(bypass_byp_alu_rs2_data_d[11]));
OR2X1 exu_U7625(.A(exu_n12784), .B(exu_n14132), .Y(bypass_byp_alu_rs2_data_d[10]));
OR2X1 exu_U7626(.A(exu_n12722), .B(exu_n14070), .Y(bypass_byp_alu_rs2_data_d[9]));
OR2X1 exu_U7627(.A(exu_n12723), .B(exu_n14071), .Y(bypass_byp_alu_rs2_data_d[8]));
OR2X1 exu_U7628(.A(exu_n12724), .B(exu_n14072), .Y(bypass_byp_alu_rs2_data_d[7]));
OR2X1 exu_U7629(.A(exu_n12725), .B(exu_n14073), .Y(bypass_byp_alu_rs2_data_d[6]));
OR2X1 exu_U7630(.A(exu_n12730), .B(exu_n14078), .Y(bypass_byp_alu_rs2_data_d[5]));
OR2X1 exu_U7631(.A(exu_n12741), .B(exu_n14089), .Y(bypass_byp_alu_rs2_data_d[4]));
OR2X1 exu_U7632(.A(exu_n12752), .B(exu_n14100), .Y(bypass_byp_alu_rs2_data_d[3]));
OR2X1 exu_U7633(.A(exu_n12763), .B(exu_n14111), .Y(bypass_byp_alu_rs2_data_d[2]));
OR2X1 exu_U7634(.A(exu_n12774), .B(exu_n14122), .Y(bypass_byp_alu_rs2_data_d[1]));
OR2X1 exu_U7635(.A(exu_n12785), .B(exu_n14133), .Y(bypass_byp_alu_rs2_data_d[0]));
OR2X1 exu_U7636(.A(exu_n12854), .B(exu_n14138), .Y(bypass_rs3_data_d[63]));
OR2X1 exu_U7637(.A(exu_n12855), .B(exu_n14139), .Y(bypass_rs3_data_d[62]));
OR2X1 exu_U7638(.A(exu_n12856), .B(exu_n14140), .Y(bypass_rs3_data_d[61]));
OR2X1 exu_U7639(.A(exu_n12857), .B(exu_n14141), .Y(bypass_rs3_data_d[60]));
OR2X1 exu_U7640(.A(exu_n12859), .B(exu_n14143), .Y(bypass_rs3_data_d[59]));
OR2X1 exu_U7641(.A(exu_n12860), .B(exu_n14144), .Y(bypass_rs3_data_d[58]));
OR2X1 exu_U7642(.A(exu_n12861), .B(exu_n14145), .Y(bypass_rs3_data_d[57]));
OR2X1 exu_U7643(.A(exu_n12862), .B(exu_n14146), .Y(bypass_rs3_data_d[56]));
OR2X1 exu_U7644(.A(exu_n12863), .B(exu_n14147), .Y(bypass_rs3_data_d[55]));
OR2X1 exu_U7645(.A(exu_n12864), .B(exu_n14148), .Y(bypass_rs3_data_d[54]));
OR2X1 exu_U7646(.A(exu_n12865), .B(exu_n14149), .Y(bypass_rs3_data_d[53]));
OR2X1 exu_U7647(.A(exu_n12866), .B(exu_n14150), .Y(bypass_rs3_data_d[52]));
OR2X1 exu_U7648(.A(exu_n12867), .B(exu_n14151), .Y(bypass_rs3_data_d[51]));
OR2X1 exu_U7649(.A(exu_n12868), .B(exu_n14152), .Y(bypass_rs3_data_d[50]));
OR2X1 exu_U7650(.A(exu_n12870), .B(exu_n14154), .Y(bypass_rs3_data_d[49]));
OR2X1 exu_U7651(.A(exu_n12871), .B(exu_n14155), .Y(bypass_rs3_data_d[48]));
OR2X1 exu_U7652(.A(exu_n12872), .B(exu_n14156), .Y(bypass_rs3_data_d[47]));
OR2X1 exu_U7653(.A(exu_n12873), .B(exu_n14157), .Y(bypass_rs3_data_d[46]));
OR2X1 exu_U7654(.A(exu_n12874), .B(exu_n14158), .Y(bypass_rs3_data_d[45]));
OR2X1 exu_U7655(.A(exu_n12875), .B(exu_n14159), .Y(bypass_rs3_data_d[44]));
OR2X1 exu_U7656(.A(exu_n12876), .B(exu_n14160), .Y(bypass_rs3_data_d[43]));
OR2X1 exu_U7657(.A(exu_n12877), .B(exu_n14161), .Y(bypass_rs3_data_d[42]));
OR2X1 exu_U7658(.A(exu_n12878), .B(exu_n14162), .Y(bypass_rs3_data_d[41]));
OR2X1 exu_U7659(.A(exu_n12879), .B(exu_n14163), .Y(bypass_rs3_data_d[40]));
OR2X1 exu_U7660(.A(exu_n12881), .B(exu_n14165), .Y(bypass_rs3_data_d[39]));
OR2X1 exu_U7661(.A(exu_n12882), .B(exu_n14166), .Y(bypass_rs3_data_d[38]));
OR2X1 exu_U7662(.A(exu_n12883), .B(exu_n14167), .Y(bypass_rs3_data_d[37]));
OR2X1 exu_U7663(.A(exu_n12884), .B(exu_n14168), .Y(bypass_rs3_data_d[36]));
OR2X1 exu_U7664(.A(exu_n12885), .B(exu_n14169), .Y(bypass_rs3_data_d[35]));
OR2X1 exu_U7665(.A(exu_n12886), .B(exu_n14170), .Y(bypass_rs3_data_d[34]));
OR2X1 exu_U7666(.A(exu_n12887), .B(exu_n14171), .Y(bypass_rs3_data_d[33]));
OR2X1 exu_U7667(.A(exu_n12888), .B(exu_n14172), .Y(bypass_rs3_data_d[32]));
OR2X1 exu_U7668(.A(exu_n12889), .B(exu_n14173), .Y(bypass_rs3_data_d[31]));
OR2X1 exu_U7669(.A(exu_n12890), .B(exu_n14174), .Y(bypass_rs3_data_d[30]));
OR2X1 exu_U7670(.A(exu_n12892), .B(exu_n14176), .Y(bypass_rs3_data_d[29]));
OR2X1 exu_U7671(.A(exu_n12893), .B(exu_n14177), .Y(bypass_rs3_data_d[28]));
OR2X1 exu_U7672(.A(exu_n12894), .B(exu_n14178), .Y(bypass_rs3_data_d[27]));
OR2X1 exu_U7673(.A(exu_n12895), .B(exu_n14179), .Y(bypass_rs3_data_d[26]));
OR2X1 exu_U7674(.A(exu_n12896), .B(exu_n14180), .Y(bypass_rs3_data_d[25]));
OR2X1 exu_U7675(.A(exu_n12897), .B(exu_n14181), .Y(bypass_rs3_data_d[24]));
OR2X1 exu_U7676(.A(exu_n12898), .B(exu_n14182), .Y(bypass_rs3_data_d[23]));
OR2X1 exu_U7677(.A(exu_n12899), .B(exu_n14183), .Y(bypass_rs3_data_d[22]));
OR2X1 exu_U7678(.A(exu_n12900), .B(exu_n14184), .Y(bypass_rs3_data_d[21]));
OR2X1 exu_U7679(.A(exu_n12901), .B(exu_n14185), .Y(bypass_rs3_data_d[20]));
OR2X1 exu_U7680(.A(exu_n12903), .B(exu_n14187), .Y(bypass_rs3_data_d[19]));
OR2X1 exu_U7681(.A(exu_n12904), .B(exu_n14188), .Y(bypass_rs3_data_d[18]));
OR2X1 exu_U7682(.A(exu_n12905), .B(exu_n14189), .Y(bypass_rs3_data_d[17]));
OR2X1 exu_U7683(.A(exu_n12906), .B(exu_n14190), .Y(bypass_rs3_data_d[16]));
OR2X1 exu_U7684(.A(exu_n12907), .B(exu_n14191), .Y(bypass_rs3_data_d[15]));
OR2X1 exu_U7685(.A(exu_n12908), .B(exu_n14192), .Y(bypass_rs3_data_d[14]));
OR2X1 exu_U7686(.A(exu_n12909), .B(exu_n14193), .Y(bypass_rs3_data_d[13]));
OR2X1 exu_U7687(.A(exu_n12910), .B(exu_n14194), .Y(bypass_rs3_data_d[12]));
OR2X1 exu_U7688(.A(exu_n12911), .B(exu_n14195), .Y(bypass_rs3_data_d[11]));
OR2X1 exu_U7689(.A(exu_n12912), .B(exu_n14196), .Y(bypass_rs3_data_d[10]));
OR2X1 exu_U7690(.A(exu_n12850), .B(exu_n14134), .Y(bypass_rs3_data_d[9]));
OR2X1 exu_U7691(.A(exu_n12851), .B(exu_n14135), .Y(bypass_rs3_data_d[8]));
OR2X1 exu_U7692(.A(exu_n12852), .B(exu_n14136), .Y(bypass_rs3_data_d[7]));
OR2X1 exu_U7693(.A(exu_n12853), .B(exu_n14137), .Y(bypass_rs3_data_d[6]));
OR2X1 exu_U7694(.A(exu_n12858), .B(exu_n14142), .Y(bypass_rs3_data_d[5]));
OR2X1 exu_U7695(.A(exu_n12869), .B(exu_n14153), .Y(bypass_rs3_data_d[4]));
OR2X1 exu_U7696(.A(exu_n12880), .B(exu_n14164), .Y(bypass_rs3_data_d[3]));
OR2X1 exu_U7697(.A(exu_n12891), .B(exu_n14175), .Y(bypass_rs3_data_d[2]));
OR2X1 exu_U7698(.A(exu_n12902), .B(exu_n14186), .Y(bypass_rs3_data_d[1]));
OR2X1 exu_U7699(.A(exu_n12913), .B(exu_n14197), .Y(bypass_rs3_data_d[0]));
OR2X1 exu_U7700(.A(exu_n12598), .B(exu_n13946), .Y(bypass_byp_alu_rcc_data_d[63]));
OR2X1 exu_U7701(.A(exu_n12599), .B(exu_n13947), .Y(bypass_byp_alu_rcc_data_d[62]));
OR2X1 exu_U7702(.A(exu_n12600), .B(exu_n13948), .Y(bypass_byp_alu_rcc_data_d[61]));
OR2X1 exu_U7703(.A(exu_n12601), .B(exu_n13949), .Y(bypass_byp_alu_rcc_data_d[60]));
OR2X1 exu_U7704(.A(exu_n12603), .B(exu_n13951), .Y(bypass_byp_alu_rcc_data_d[59]));
OR2X1 exu_U7705(.A(exu_n12604), .B(exu_n13952), .Y(bypass_byp_alu_rcc_data_d[58]));
OR2X1 exu_U7706(.A(exu_n12605), .B(exu_n13953), .Y(bypass_byp_alu_rcc_data_d[57]));
OR2X1 exu_U7707(.A(exu_n12606), .B(exu_n13954), .Y(bypass_byp_alu_rcc_data_d[56]));
OR2X1 exu_U7708(.A(exu_n12607), .B(exu_n13955), .Y(bypass_byp_alu_rcc_data_d[55]));
OR2X1 exu_U7709(.A(exu_n12608), .B(exu_n13956), .Y(bypass_byp_alu_rcc_data_d[54]));
OR2X1 exu_U7710(.A(exu_n12609), .B(exu_n13957), .Y(bypass_byp_alu_rcc_data_d[53]));
OR2X1 exu_U7711(.A(exu_n12610), .B(exu_n13958), .Y(bypass_byp_alu_rcc_data_d[52]));
OR2X1 exu_U7712(.A(exu_n12611), .B(exu_n13959), .Y(bypass_byp_alu_rcc_data_d[51]));
OR2X1 exu_U7713(.A(exu_n12612), .B(exu_n13960), .Y(bypass_byp_alu_rcc_data_d[50]));
OR2X1 exu_U7714(.A(exu_n12614), .B(exu_n13962), .Y(bypass_byp_alu_rcc_data_d[49]));
OR2X1 exu_U7715(.A(exu_n12615), .B(exu_n13963), .Y(bypass_byp_alu_rcc_data_d[48]));
OR2X1 exu_U7716(.A(exu_n12616), .B(exu_n13964), .Y(bypass_byp_alu_rcc_data_d[47]));
OR2X1 exu_U7717(.A(exu_n12617), .B(exu_n13965), .Y(bypass_byp_alu_rcc_data_d[46]));
OR2X1 exu_U7718(.A(exu_n12618), .B(exu_n13966), .Y(bypass_byp_alu_rcc_data_d[45]));
OR2X1 exu_U7719(.A(exu_n12619), .B(exu_n13967), .Y(bypass_byp_alu_rcc_data_d[44]));
OR2X1 exu_U7720(.A(exu_n12620), .B(exu_n13968), .Y(bypass_byp_alu_rcc_data_d[43]));
OR2X1 exu_U7721(.A(exu_n12621), .B(exu_n13969), .Y(bypass_byp_alu_rcc_data_d[42]));
OR2X1 exu_U7722(.A(exu_n12622), .B(exu_n13970), .Y(bypass_byp_alu_rcc_data_d[41]));
OR2X1 exu_U7723(.A(exu_n12623), .B(exu_n13971), .Y(bypass_byp_alu_rcc_data_d[40]));
OR2X1 exu_U7724(.A(exu_n12625), .B(exu_n13973), .Y(bypass_byp_alu_rcc_data_d[39]));
OR2X1 exu_U7725(.A(exu_n12626), .B(exu_n13974), .Y(bypass_byp_alu_rcc_data_d[38]));
OR2X1 exu_U7726(.A(exu_n12627), .B(exu_n13975), .Y(bypass_byp_alu_rcc_data_d[37]));
OR2X1 exu_U7727(.A(exu_n12628), .B(exu_n13976), .Y(bypass_byp_alu_rcc_data_d[36]));
OR2X1 exu_U7728(.A(exu_n12629), .B(exu_n13977), .Y(bypass_byp_alu_rcc_data_d[35]));
OR2X1 exu_U7729(.A(exu_n12630), .B(exu_n13978), .Y(bypass_byp_alu_rcc_data_d[34]));
OR2X1 exu_U7730(.A(exu_n12631), .B(exu_n13979), .Y(bypass_byp_alu_rcc_data_d[33]));
OR2X1 exu_U7731(.A(exu_n12632), .B(exu_n13980), .Y(bypass_byp_alu_rcc_data_d[32]));
OR2X1 exu_U7732(.A(exu_n12633), .B(exu_n13981), .Y(bypass_byp_alu_rcc_data_d[31]));
OR2X1 exu_U7733(.A(exu_n12634), .B(exu_n13982), .Y(bypass_byp_alu_rcc_data_d[30]));
OR2X1 exu_U7734(.A(exu_n12636), .B(exu_n13984), .Y(bypass_byp_alu_rcc_data_d[29]));
OR2X1 exu_U7735(.A(exu_n12637), .B(exu_n13985), .Y(bypass_byp_alu_rcc_data_d[28]));
OR2X1 exu_U7736(.A(exu_n12638), .B(exu_n13986), .Y(bypass_byp_alu_rcc_data_d[27]));
OR2X1 exu_U7737(.A(exu_n12639), .B(exu_n13987), .Y(bypass_byp_alu_rcc_data_d[26]));
OR2X1 exu_U7738(.A(exu_n12640), .B(exu_n13988), .Y(bypass_byp_alu_rcc_data_d[25]));
OR2X1 exu_U7739(.A(exu_n12641), .B(exu_n13989), .Y(bypass_byp_alu_rcc_data_d[24]));
OR2X1 exu_U7740(.A(exu_n12642), .B(exu_n13990), .Y(bypass_byp_alu_rcc_data_d[23]));
OR2X1 exu_U7741(.A(exu_n12643), .B(exu_n13991), .Y(bypass_byp_alu_rcc_data_d[22]));
OR2X1 exu_U7742(.A(exu_n12644), .B(exu_n13992), .Y(bypass_byp_alu_rcc_data_d[21]));
OR2X1 exu_U7743(.A(exu_n12645), .B(exu_n13993), .Y(bypass_byp_alu_rcc_data_d[20]));
OR2X1 exu_U7744(.A(exu_n12647), .B(exu_n13995), .Y(bypass_byp_alu_rcc_data_d[19]));
OR2X1 exu_U7745(.A(exu_n12648), .B(exu_n13996), .Y(bypass_byp_alu_rcc_data_d[18]));
OR2X1 exu_U7746(.A(exu_n12649), .B(exu_n13997), .Y(bypass_byp_alu_rcc_data_d[17]));
OR2X1 exu_U7747(.A(exu_n12650), .B(exu_n13998), .Y(bypass_byp_alu_rcc_data_d[16]));
OR2X1 exu_U7748(.A(exu_n12651), .B(exu_n13999), .Y(bypass_byp_alu_rcc_data_d[15]));
OR2X1 exu_U7749(.A(exu_n12652), .B(exu_n14000), .Y(bypass_byp_alu_rcc_data_d[14]));
OR2X1 exu_U7750(.A(exu_n12653), .B(exu_n14001), .Y(bypass_byp_alu_rcc_data_d[13]));
OR2X1 exu_U7751(.A(exu_n12654), .B(exu_n14002), .Y(bypass_byp_alu_rcc_data_d[12]));
OR2X1 exu_U7752(.A(exu_n12655), .B(exu_n14003), .Y(bypass_byp_alu_rcc_data_d[11]));
OR2X1 exu_U7753(.A(exu_n12656), .B(exu_n14004), .Y(bypass_byp_alu_rcc_data_d[10]));
OR2X1 exu_U7754(.A(exu_n12594), .B(exu_n13942), .Y(bypass_byp_alu_rcc_data_d[9]));
OR2X1 exu_U7755(.A(exu_n12595), .B(exu_n13943), .Y(bypass_byp_alu_rcc_data_d[8]));
OR2X1 exu_U7756(.A(exu_n12596), .B(exu_n13944), .Y(bypass_byp_alu_rcc_data_d[7]));
OR2X1 exu_U7757(.A(exu_n12597), .B(exu_n13945), .Y(bypass_byp_alu_rcc_data_d[6]));
OR2X1 exu_U7758(.A(exu_n12602), .B(exu_n13950), .Y(bypass_byp_alu_rcc_data_d[5]));
OR2X1 exu_U7759(.A(exu_n12613), .B(exu_n13961), .Y(bypass_byp_alu_rcc_data_d[4]));
OR2X1 exu_U7760(.A(exu_n12624), .B(exu_n13972), .Y(bypass_byp_alu_rcc_data_d[3]));
OR2X1 exu_U7761(.A(exu_n12635), .B(exu_n13983), .Y(bypass_byp_alu_rcc_data_d[2]));
OR2X1 exu_U7762(.A(exu_n12646), .B(exu_n13994), .Y(bypass_byp_alu_rcc_data_d[1]));
OR2X1 exu_U7763(.A(exu_n12657), .B(exu_n14005), .Y(bypass_byp_alu_rcc_data_d[0]));
INVX1 exu_U7764(.A(se), .Y(exu_n19289));
INVX1 exu_U7765(.A(exu_n23081), .Y(exu_n16443));
AND2X1 exu_U7766(.A(exu_n3839), .B(exu_n6511), .Y(exu_n23081));
INVX1 exu_U7767(.A(exu_n23083), .Y(exu_n16444));
AND2X1 exu_U7768(.A(exu_n3840), .B(exu_n6512), .Y(exu_n23083));
INVX1 exu_U7769(.A(exu_n23085), .Y(exu_n16445));
AND2X1 exu_U7770(.A(exu_n3841), .B(exu_n6513), .Y(exu_n23085));
INVX1 exu_U7771(.A(exu_n23087), .Y(exu_n16446));
AND2X1 exu_U7772(.A(exu_n3842), .B(exu_n6514), .Y(exu_n23087));
INVX1 exu_U7773(.A(exu_n23091), .Y(exu_n16448));
AND2X1 exu_U7774(.A(exu_n3844), .B(exu_n6516), .Y(exu_n23091));
INVX1 exu_U7775(.A(exu_n23093), .Y(exu_n16449));
AND2X1 exu_U7776(.A(exu_n3845), .B(exu_n6517), .Y(exu_n23093));
INVX1 exu_U7777(.A(exu_n23095), .Y(exu_n16450));
AND2X1 exu_U7778(.A(exu_n3846), .B(exu_n6518), .Y(exu_n23095));
INVX1 exu_U7779(.A(exu_n23097), .Y(exu_n16451));
AND2X1 exu_U7780(.A(exu_n3847), .B(exu_n6519), .Y(exu_n23097));
INVX1 exu_U7781(.A(exu_n23099), .Y(exu_n16452));
AND2X1 exu_U7782(.A(exu_n3848), .B(exu_n6520), .Y(exu_n23099));
INVX1 exu_U7783(.A(exu_n23101), .Y(exu_n16453));
AND2X1 exu_U7784(.A(exu_n3849), .B(exu_n6521), .Y(exu_n23101));
INVX1 exu_U7785(.A(exu_n23103), .Y(exu_n16454));
AND2X1 exu_U7786(.A(exu_n3850), .B(exu_n6522), .Y(exu_n23103));
INVX1 exu_U7787(.A(exu_n23105), .Y(exu_n16455));
AND2X1 exu_U7788(.A(exu_n3851), .B(exu_n6523), .Y(exu_n23105));
INVX1 exu_U7789(.A(exu_n23107), .Y(exu_n16456));
AND2X1 exu_U7790(.A(exu_n3852), .B(exu_n6524), .Y(exu_n23107));
INVX1 exu_U7791(.A(exu_n23109), .Y(exu_n16457));
AND2X1 exu_U7792(.A(exu_n3853), .B(exu_n6525), .Y(exu_n23109));
INVX1 exu_U7793(.A(exu_n23113), .Y(exu_n16459));
AND2X1 exu_U7794(.A(exu_n3855), .B(exu_n6527), .Y(exu_n23113));
INVX1 exu_U7795(.A(exu_n23115), .Y(exu_n16460));
AND2X1 exu_U7796(.A(exu_n3856), .B(exu_n6528), .Y(exu_n23115));
INVX1 exu_U7797(.A(exu_n23117), .Y(exu_n16461));
AND2X1 exu_U7798(.A(exu_n3857), .B(exu_n6529), .Y(exu_n23117));
INVX1 exu_U7799(.A(exu_n23119), .Y(exu_n16462));
AND2X1 exu_U7800(.A(exu_n3858), .B(exu_n6530), .Y(exu_n23119));
INVX1 exu_U7801(.A(exu_n23121), .Y(exu_n16463));
AND2X1 exu_U7802(.A(exu_n3859), .B(exu_n6531), .Y(exu_n23121));
INVX1 exu_U7803(.A(exu_n23123), .Y(exu_n16464));
AND2X1 exu_U7804(.A(exu_n3860), .B(exu_n6532), .Y(exu_n23123));
INVX1 exu_U7805(.A(exu_n23125), .Y(exu_n16465));
AND2X1 exu_U7806(.A(exu_n3861), .B(exu_n6533), .Y(exu_n23125));
INVX1 exu_U7807(.A(exu_n23127), .Y(exu_n16466));
AND2X1 exu_U7808(.A(exu_n3862), .B(exu_n6534), .Y(exu_n23127));
INVX1 exu_U7809(.A(exu_n23129), .Y(exu_n16467));
AND2X1 exu_U7810(.A(exu_n3863), .B(exu_n6535), .Y(exu_n23129));
INVX1 exu_U7811(.A(exu_n23131), .Y(exu_n16468));
AND2X1 exu_U7812(.A(exu_n3864), .B(exu_n6536), .Y(exu_n23131));
INVX1 exu_U7813(.A(exu_n23135), .Y(exu_n16470));
AND2X1 exu_U7814(.A(exu_n3866), .B(exu_n6538), .Y(exu_n23135));
INVX1 exu_U7815(.A(exu_n23137), .Y(exu_n16471));
AND2X1 exu_U7816(.A(exu_n3867), .B(exu_n6539), .Y(exu_n23137));
INVX1 exu_U7817(.A(exu_n23139), .Y(exu_n16472));
AND2X1 exu_U7818(.A(exu_n3868), .B(exu_n6540), .Y(exu_n23139));
INVX1 exu_U7819(.A(exu_n23141), .Y(exu_n16473));
AND2X1 exu_U7820(.A(exu_n3869), .B(exu_n6541), .Y(exu_n23141));
INVX1 exu_U7821(.A(exu_n23143), .Y(exu_n16474));
AND2X1 exu_U7822(.A(exu_n3870), .B(exu_n6542), .Y(exu_n23143));
INVX1 exu_U7823(.A(exu_n23145), .Y(exu_n16475));
AND2X1 exu_U7824(.A(exu_n3871), .B(exu_n6543), .Y(exu_n23145));
INVX1 exu_U7825(.A(exu_n23147), .Y(exu_n16476));
AND2X1 exu_U7826(.A(exu_n3872), .B(exu_n6544), .Y(exu_n23147));
INVX1 exu_U7827(.A(exu_n23149), .Y(exu_n16477));
AND2X1 exu_U7828(.A(exu_n3873), .B(exu_n6545), .Y(exu_n23149));
INVX1 exu_U7829(.A(exu_n23151), .Y(exu_n16478));
AND2X1 exu_U7830(.A(exu_n3874), .B(exu_n6546), .Y(exu_n23151));
INVX1 exu_U7831(.A(exu_n23153), .Y(exu_n16479));
AND2X1 exu_U7832(.A(exu_n3875), .B(exu_n6547), .Y(exu_n23153));
INVX1 exu_U7833(.A(exu_n23157), .Y(exu_n16481));
AND2X1 exu_U7834(.A(exu_n3877), .B(exu_n6549), .Y(exu_n23157));
INVX1 exu_U7835(.A(exu_n23159), .Y(exu_n16482));
AND2X1 exu_U7836(.A(exu_n3878), .B(exu_n6550), .Y(exu_n23159));
INVX1 exu_U7837(.A(exu_n23161), .Y(exu_n16483));
AND2X1 exu_U7838(.A(exu_n3879), .B(exu_n6551), .Y(exu_n23161));
INVX1 exu_U7839(.A(exu_n23163), .Y(exu_n16484));
AND2X1 exu_U7840(.A(exu_n3880), .B(exu_n6552), .Y(exu_n23163));
INVX1 exu_U7841(.A(exu_n23165), .Y(exu_n16485));
AND2X1 exu_U7842(.A(exu_n3881), .B(exu_n6553), .Y(exu_n23165));
INVX1 exu_U7843(.A(exu_n23167), .Y(exu_n16486));
AND2X1 exu_U7844(.A(exu_n3882), .B(exu_n6554), .Y(exu_n23167));
INVX1 exu_U7845(.A(exu_n23169), .Y(exu_n16487));
AND2X1 exu_U7846(.A(exu_n3883), .B(exu_n6555), .Y(exu_n23169));
INVX1 exu_U7847(.A(exu_n23171), .Y(exu_n16488));
AND2X1 exu_U7848(.A(exu_n3884), .B(exu_n6556), .Y(exu_n23171));
INVX1 exu_U7849(.A(exu_n23173), .Y(exu_n16489));
AND2X1 exu_U7850(.A(exu_n3885), .B(exu_n6557), .Y(exu_n23173));
INVX1 exu_U7851(.A(exu_n23175), .Y(exu_n16490));
AND2X1 exu_U7852(.A(exu_n3886), .B(exu_n6558), .Y(exu_n23175));
INVX1 exu_U7853(.A(exu_n23179), .Y(exu_n16492));
AND2X1 exu_U7854(.A(exu_n3888), .B(exu_n6560), .Y(exu_n23179));
INVX1 exu_U7855(.A(exu_n23181), .Y(exu_n16493));
AND2X1 exu_U7856(.A(exu_n3889), .B(exu_n6561), .Y(exu_n23181));
INVX1 exu_U7857(.A(exu_n23183), .Y(exu_n16494));
AND2X1 exu_U7858(.A(exu_n3890), .B(exu_n6562), .Y(exu_n23183));
INVX1 exu_U7859(.A(exu_n23185), .Y(exu_n16495));
AND2X1 exu_U7860(.A(exu_n3891), .B(exu_n6563), .Y(exu_n23185));
INVX1 exu_U7861(.A(exu_n23187), .Y(exu_n16496));
AND2X1 exu_U7862(.A(exu_n3892), .B(exu_n6564), .Y(exu_n23187));
INVX1 exu_U7863(.A(exu_n23189), .Y(exu_n16497));
AND2X1 exu_U7864(.A(exu_n3893), .B(exu_n6565), .Y(exu_n23189));
INVX1 exu_U7865(.A(exu_n23191), .Y(exu_n16498));
AND2X1 exu_U7866(.A(exu_n3894), .B(exu_n6566), .Y(exu_n23191));
INVX1 exu_U7867(.A(exu_n23193), .Y(exu_n16499));
AND2X1 exu_U7868(.A(exu_n3895), .B(exu_n6567), .Y(exu_n23193));
INVX1 exu_U7869(.A(exu_n23195), .Y(exu_n16500));
AND2X1 exu_U7870(.A(exu_n3896), .B(exu_n6568), .Y(exu_n23195));
INVX1 exu_U7871(.A(exu_n23197), .Y(exu_n16501));
AND2X1 exu_U7872(.A(exu_n3897), .B(exu_n6569), .Y(exu_n23197));
INVX1 exu_U7873(.A(exu_n23073), .Y(exu_n16439));
AND2X1 exu_U7874(.A(exu_n3835), .B(exu_n6507), .Y(exu_n23073));
INVX1 exu_U7875(.A(exu_n23075), .Y(exu_n16440));
AND2X1 exu_U7876(.A(exu_n3836), .B(exu_n6508), .Y(exu_n23075));
INVX1 exu_U7877(.A(exu_n23077), .Y(exu_n16441));
AND2X1 exu_U7878(.A(exu_n3837), .B(exu_n6509), .Y(exu_n23077));
INVX1 exu_U7879(.A(exu_n23079), .Y(exu_n16442));
AND2X1 exu_U7880(.A(exu_n3838), .B(exu_n6510), .Y(exu_n23079));
INVX1 exu_U7881(.A(exu_n23089), .Y(exu_n16447));
AND2X1 exu_U7882(.A(exu_n3843), .B(exu_n6515), .Y(exu_n23089));
INVX1 exu_U7883(.A(exu_n23111), .Y(exu_n16458));
AND2X1 exu_U7884(.A(exu_n3854), .B(exu_n6526), .Y(exu_n23111));
INVX1 exu_U7885(.A(exu_n23133), .Y(exu_n16469));
AND2X1 exu_U7886(.A(exu_n3865), .B(exu_n6537), .Y(exu_n23133));
INVX1 exu_U7887(.A(exu_n23155), .Y(exu_n16480));
AND2X1 exu_U7888(.A(exu_n3876), .B(exu_n6548), .Y(exu_n23155));
INVX1 exu_U7889(.A(exu_n23177), .Y(exu_n16491));
AND2X1 exu_U7890(.A(exu_n3887), .B(exu_n6559), .Y(exu_n23177));
INVX1 exu_U7891(.A(exu_n23199), .Y(exu_n16502));
AND2X1 exu_U7892(.A(exu_n3898), .B(exu_n6570), .Y(exu_n23199));
INVX1 exu_U7893(.A(se), .Y(exu_n19337));
OR2X1 exu_U7894(.A(rml_cwp_n74), .B(exu_n14701), .Y(rml_cwp_next_slot0_state[1]));
AND2X1 exu_U7895(.A(exu_n3967), .B(exu_n8982), .Y(exu_n31469));
OR2X1 exu_U7896(.A(exu_n31473), .B(exu_n31472), .Y(rml_cwp_next_slot0_state[0]));
AND2X1 exu_U7897(.A(exu_n4040), .B(exu_n9054), .Y(rml_cwp_slot0_data_mux_n17));
AND2X1 exu_U7898(.A(exu_n4042), .B(exu_n9055), .Y(rml_cwp_slot0_data_mux_n21));
AND2X1 exu_U7899(.A(exu_n4044), .B(exu_n9056), .Y(rml_cwp_slot0_data_mux_n25));
AND2X1 exu_U7900(.A(exu_n4046), .B(exu_n9057), .Y(rml_cwp_slot0_data_mux_n29));
AND2X1 exu_U7901(.A(exu_n4048), .B(exu_n9058), .Y(rml_cwp_slot0_data_mux_n33));
AND2X1 exu_U7902(.A(exu_n4053), .B(exu_n9059), .Y(rml_cwp_slot0_data_mux_n49));
AND2X1 exu_U7903(.A(exu_n15815), .B(exu_n9308), .Y(ecl_divcntl_next_state[5]));
AND2X1 exu_U7904(.A(exu_n15815), .B(exu_n9309), .Y(ecl_divcntl_next_state[4]));
AND2X1 exu_U7905(.A(exu_n15815), .B(exu_n9310), .Y(ecl_divcntl_next_state[1]));
AND2X1 exu_U7906(.A(exu_n4505), .B(exu_n9311), .Y(ecl_divcntl_n35));
AND2X1 exu_U7907(.A(exu_n4354), .B(exu_n9231), .Y(div_d_mux_n389));
AND2X1 exu_U7908(.A(exu_n4356), .B(exu_n9232), .Y(div_d_mux_n393));
AND2X1 exu_U7909(.A(exu_n4358), .B(exu_n9233), .Y(div_d_mux_n397));
AND2X1 exu_U7910(.A(exu_n4360), .B(exu_n9234), .Y(div_d_mux_n401));
AND2X1 exu_U7911(.A(exu_n4362), .B(exu_n9235), .Y(div_d_mux_n405));
AND2X1 exu_U7912(.A(exu_n4364), .B(exu_n9236), .Y(div_d_mux_n409));
AND2X1 exu_U7913(.A(exu_n4366), .B(exu_n9237), .Y(div_d_mux_n413));
AND2X1 exu_U7914(.A(exu_n4368), .B(exu_n9238), .Y(div_d_mux_n417));
AND2X1 exu_U7915(.A(exu_n4372), .B(exu_n9240), .Y(div_d_mux_n425));
AND2X1 exu_U7916(.A(exu_n4374), .B(exu_n9241), .Y(div_d_mux_n429));
AND2X1 exu_U7917(.A(exu_n4376), .B(exu_n9242), .Y(div_d_mux_n433));
AND2X1 exu_U7918(.A(exu_n4378), .B(exu_n9243), .Y(div_d_mux_n437));
AND2X1 exu_U7919(.A(exu_n4380), .B(exu_n9244), .Y(div_d_mux_n441));
AND2X1 exu_U7920(.A(exu_n4382), .B(exu_n9245), .Y(div_d_mux_n445));
AND2X1 exu_U7921(.A(exu_n4384), .B(exu_n9246), .Y(div_d_mux_n449));
AND2X1 exu_U7922(.A(exu_n4386), .B(exu_n9247), .Y(div_d_mux_n453));
AND2X1 exu_U7923(.A(exu_n4388), .B(exu_n9248), .Y(div_d_mux_n457));
AND2X1 exu_U7924(.A(exu_n4390), .B(exu_n9249), .Y(div_d_mux_n461));
AND2X1 exu_U7925(.A(exu_n4394), .B(exu_n9251), .Y(div_d_mux_n469));
AND2X1 exu_U7926(.A(exu_n4396), .B(exu_n9252), .Y(div_d_mux_n473));
AND2X1 exu_U7927(.A(exu_n4398), .B(exu_n9253), .Y(div_d_mux_n477));
AND2X1 exu_U7928(.A(exu_n4400), .B(exu_n9254), .Y(div_d_mux_n481));
AND2X1 exu_U7929(.A(exu_n4402), .B(exu_n9255), .Y(div_d_mux_n485));
AND2X1 exu_U7930(.A(exu_n4404), .B(exu_n9256), .Y(div_d_mux_n489));
AND2X1 exu_U7931(.A(exu_n4406), .B(exu_n9257), .Y(div_d_mux_n493));
AND2X1 exu_U7932(.A(exu_n4408), .B(exu_n9258), .Y(div_d_mux_n497));
AND2X1 exu_U7933(.A(exu_n4410), .B(exu_n9259), .Y(div_d_mux_n501));
AND2X1 exu_U7934(.A(exu_n4412), .B(exu_n9260), .Y(div_d_mux_n505));
AND2X1 exu_U7935(.A(exu_n4162), .B(exu_n9135), .Y(div_d_mux_n5));
AND2X1 exu_U7936(.A(exu_n4164), .B(exu_n9136), .Y(div_d_mux_n9));
AND2X1 exu_U7937(.A(exu_n4166), .B(exu_n9137), .Y(div_d_mux_n13));
AND2X1 exu_U7938(.A(exu_n4168), .B(exu_n9138), .Y(div_d_mux_n17));
AND2X1 exu_U7939(.A(exu_n4170), .B(exu_n9139), .Y(div_d_mux_n21));
AND2X1 exu_U7940(.A(exu_n4172), .B(exu_n9140), .Y(div_d_mux_n25));
AND2X1 exu_U7941(.A(exu_n4174), .B(exu_n9141), .Y(div_d_mux_n29));
AND2X1 exu_U7942(.A(exu_n4176), .B(exu_n9142), .Y(div_d_mux_n33));
AND2X1 exu_U7943(.A(exu_n4178), .B(exu_n9143), .Y(div_d_mux_n37));
AND2X1 exu_U7944(.A(exu_n4180), .B(exu_n9144), .Y(div_d_mux_n41));
AND2X1 exu_U7945(.A(exu_n4184), .B(exu_n9146), .Y(div_d_mux_n49));
AND2X1 exu_U7946(.A(exu_n4186), .B(exu_n9147), .Y(div_d_mux_n53));
AND2X1 exu_U7947(.A(exu_n4188), .B(exu_n9148), .Y(div_d_mux_n57));
AND2X1 exu_U7948(.A(exu_n4190), .B(exu_n9149), .Y(div_d_mux_n61));
AND2X1 exu_U7949(.A(exu_n4192), .B(exu_n9150), .Y(div_d_mux_n65));
AND2X1 exu_U7950(.A(exu_n4194), .B(exu_n9151), .Y(div_d_mux_n69));
AND2X1 exu_U7951(.A(exu_n4196), .B(exu_n9152), .Y(div_d_mux_n73));
AND2X1 exu_U7952(.A(exu_n4198), .B(exu_n9153), .Y(div_d_mux_n77));
AND2X1 exu_U7953(.A(exu_n4200), .B(exu_n9154), .Y(div_d_mux_n81));
AND2X1 exu_U7954(.A(exu_n4202), .B(exu_n9155), .Y(div_d_mux_n85));
AND2X1 exu_U7955(.A(exu_n4206), .B(exu_n9157), .Y(div_d_mux_n93));
AND2X1 exu_U7956(.A(exu_n4208), .B(exu_n9158), .Y(div_d_mux_n97));
AND2X1 exu_U7957(.A(exu_n4210), .B(exu_n9159), .Y(div_d_mux_n101));
AND2X1 exu_U7958(.A(exu_n4212), .B(exu_n9160), .Y(div_d_mux_n105));
AND2X1 exu_U7959(.A(exu_n4214), .B(exu_n9161), .Y(div_d_mux_n109));
AND2X1 exu_U7960(.A(exu_n4216), .B(exu_n9162), .Y(div_d_mux_n113));
AND2X1 exu_U7961(.A(exu_n4218), .B(exu_n9163), .Y(div_d_mux_n117));
AND2X1 exu_U7962(.A(exu_n4220), .B(exu_n9164), .Y(div_d_mux_n121));
AND2X1 exu_U7963(.A(exu_n4222), .B(exu_n9165), .Y(div_d_mux_n125));
AND2X1 exu_U7964(.A(exu_n4224), .B(exu_n9166), .Y(div_d_mux_n129));
AND2X1 exu_U7965(.A(exu_n4228), .B(exu_n9168), .Y(div_d_mux_n137));
AND2X1 exu_U7966(.A(exu_n4230), .B(exu_n9169), .Y(div_d_mux_n141));
AND2X1 exu_U7967(.A(exu_n4232), .B(exu_n9170), .Y(div_d_mux_n145));
AND2X1 exu_U7968(.A(exu_n4234), .B(exu_n9171), .Y(div_d_mux_n149));
AND2X1 exu_U7969(.A(exu_n4236), .B(exu_n9172), .Y(div_d_mux_n153));
AND2X1 exu_U7970(.A(exu_n4238), .B(exu_n9173), .Y(div_d_mux_n157));
AND2X1 exu_U7971(.A(exu_n4240), .B(exu_n9174), .Y(div_d_mux_n161));
AND2X1 exu_U7972(.A(exu_n4242), .B(exu_n9175), .Y(div_d_mux_n165));
AND2X1 exu_U7973(.A(exu_n4244), .B(exu_n9176), .Y(div_d_mux_n169));
AND2X1 exu_U7974(.A(exu_n4246), .B(exu_n9177), .Y(div_d_mux_n173));
AND2X1 exu_U7975(.A(exu_n4250), .B(exu_n9179), .Y(div_d_mux_n181));
AND2X1 exu_U7976(.A(exu_n4252), .B(exu_n9180), .Y(div_d_mux_n185));
AND2X1 exu_U7977(.A(exu_n4254), .B(exu_n9181), .Y(div_d_mux_n189));
AND2X1 exu_U7978(.A(exu_n4256), .B(exu_n9182), .Y(div_d_mux_n193));
AND2X1 exu_U7979(.A(exu_n4258), .B(exu_n9183), .Y(div_d_mux_n197));
AND2X1 exu_U7980(.A(exu_n4260), .B(exu_n9184), .Y(div_d_mux_n201));
AND2X1 exu_U7981(.A(exu_n4262), .B(exu_n9185), .Y(div_d_mux_n205));
AND2X1 exu_U7982(.A(exu_n4264), .B(exu_n9186), .Y(div_d_mux_n209));
AND2X1 exu_U7983(.A(exu_n4266), .B(exu_n9187), .Y(div_d_mux_n213));
AND2X1 exu_U7984(.A(exu_n4268), .B(exu_n9188), .Y(div_d_mux_n217));
AND2X1 exu_U7985(.A(exu_n4272), .B(exu_n9190), .Y(div_d_mux_n225));
AND2X1 exu_U7986(.A(exu_n4274), .B(exu_n9191), .Y(div_d_mux_n229));
AND2X1 exu_U7987(.A(exu_n4276), .B(exu_n9192), .Y(div_d_mux_n233));
AND2X1 exu_U7988(.A(exu_n4278), .B(exu_n9193), .Y(div_d_mux_n237));
AND2X1 exu_U7989(.A(exu_n4280), .B(exu_n9194), .Y(div_d_mux_n241));
AND2X1 exu_U7990(.A(exu_n4282), .B(exu_n9195), .Y(div_d_mux_n245));
AND2X1 exu_U7991(.A(exu_n4284), .B(exu_n9196), .Y(div_d_mux_n249));
AND2X1 exu_U7992(.A(exu_n4286), .B(exu_n9197), .Y(div_d_mux_n253));
AND2X1 exu_U7993(.A(exu_n4288), .B(exu_n9198), .Y(div_d_mux_n257));
AND2X1 exu_U7994(.A(exu_n4290), .B(exu_n9199), .Y(div_d_mux_n261));
AND2X1 exu_U7995(.A(exu_n4294), .B(exu_n9201), .Y(div_d_mux_n269));
AND2X1 exu_U7996(.A(exu_n4296), .B(exu_n9202), .Y(div_d_mux_n273));
AND2X1 exu_U7997(.A(exu_n4298), .B(exu_n9203), .Y(div_d_mux_n277));
AND2X1 exu_U7998(.A(exu_n4300), .B(exu_n9204), .Y(div_d_mux_n281));
AND2X1 exu_U7999(.A(exu_n4302), .B(exu_n9205), .Y(div_d_mux_n285));
AND2X1 exu_U8000(.A(exu_n4304), .B(exu_n9206), .Y(div_d_mux_n289));
AND2X1 exu_U8001(.A(exu_n4306), .B(exu_n9207), .Y(div_d_mux_n293));
AND2X1 exu_U8002(.A(exu_n4308), .B(exu_n9208), .Y(div_d_mux_n297));
AND2X1 exu_U8003(.A(exu_n4310), .B(exu_n9209), .Y(div_d_mux_n301));
AND2X1 exu_U8004(.A(exu_n4312), .B(exu_n9210), .Y(div_d_mux_n305));
AND2X1 exu_U8005(.A(exu_n4316), .B(exu_n9212), .Y(div_d_mux_n313));
AND2X1 exu_U8006(.A(exu_n4318), .B(exu_n9213), .Y(div_d_mux_n317));
AND2X1 exu_U8007(.A(exu_n4320), .B(exu_n9214), .Y(div_d_mux_n321));
AND2X1 exu_U8008(.A(exu_n4322), .B(exu_n9215), .Y(div_d_mux_n325));
AND2X1 exu_U8009(.A(exu_n4324), .B(exu_n9216), .Y(div_d_mux_n329));
AND2X1 exu_U8010(.A(exu_n4326), .B(exu_n9217), .Y(div_d_mux_n333));
AND2X1 exu_U8011(.A(exu_n4328), .B(exu_n9218), .Y(div_d_mux_n337));
AND2X1 exu_U8012(.A(exu_n4330), .B(exu_n9219), .Y(div_d_mux_n341));
AND2X1 exu_U8013(.A(exu_n4332), .B(exu_n9220), .Y(div_d_mux_n345));
AND2X1 exu_U8014(.A(exu_n4334), .B(exu_n9221), .Y(div_d_mux_n349));
AND2X1 exu_U8015(.A(exu_n4338), .B(exu_n9223), .Y(div_d_mux_n357));
AND2X1 exu_U8016(.A(exu_n4340), .B(exu_n9224), .Y(div_d_mux_n361));
AND2X1 exu_U8017(.A(exu_n4342), .B(exu_n9225), .Y(div_d_mux_n365));
AND2X1 exu_U8018(.A(exu_n4344), .B(exu_n9226), .Y(div_d_mux_n369));
AND2X1 exu_U8019(.A(exu_n4346), .B(exu_n9227), .Y(div_d_mux_n373));
AND2X1 exu_U8020(.A(exu_n4348), .B(exu_n9228), .Y(div_d_mux_n377));
AND2X1 exu_U8021(.A(exu_n4350), .B(exu_n9229), .Y(div_d_mux_n381));
AND2X1 exu_U8022(.A(exu_n4352), .B(exu_n9230), .Y(div_d_mux_n385));
AND2X1 exu_U8023(.A(exu_n4370), .B(exu_n9239), .Y(div_d_mux_n421));
AND2X1 exu_U8024(.A(exu_n4392), .B(exu_n9250), .Y(div_d_mux_n465));
AND2X1 exu_U8025(.A(exu_n4160), .B(exu_n9134), .Y(div_d_mux_n1));
AND2X1 exu_U8026(.A(exu_n4182), .B(exu_n9145), .Y(div_d_mux_n45));
AND2X1 exu_U8027(.A(exu_n4204), .B(exu_n9156), .Y(div_d_mux_n89));
AND2X1 exu_U8028(.A(exu_n4226), .B(exu_n9167), .Y(div_d_mux_n133));
AND2X1 exu_U8029(.A(exu_n4248), .B(exu_n9178), .Y(div_d_mux_n177));
AND2X1 exu_U8030(.A(exu_n4270), .B(exu_n9189), .Y(div_d_mux_n221));
AND2X1 exu_U8031(.A(exu_n4292), .B(exu_n9200), .Y(div_d_mux_n265));
AND2X1 exu_U8032(.A(exu_n4314), .B(exu_n9211), .Y(div_d_mux_n309));
AND2X1 exu_U8033(.A(exu_n4336), .B(exu_n9222), .Y(div_d_mux_n353));
AND2X1 exu_U8034(.A(exu_n4414), .B(exu_n9261), .Y(div_d_mux_n509));
INVX1 exu_U8035(.A(ecl_ttype_mux_n5), .Y(exu_n16380));
AND2X1 exu_U8036(.A(exu_n4567), .B(exu_n9352), .Y(ecl_ttype_mux_n5));
INVX1 exu_U8037(.A(ecl_ttype_mux_n9), .Y(exu_n16379));
AND2X1 exu_U8038(.A(exu_n4568), .B(exu_n9352), .Y(ecl_ttype_mux_n9));
AND2X1 exu_U8039(.A(exu_n4570), .B(exu_n9353), .Y(ecl_ttype_mux_n13));
AND2X1 exu_U8040(.A(exu_n4572), .B(exu_n9354), .Y(ecl_ttype_mux_n17));
INVX1 exu_U8041(.A(ecl_ttype_mux_n21), .Y(exu_n16378));
AND2X1 exu_U8042(.A(exu_n4573), .B(exu_n9355), .Y(ecl_ttype_mux_n21));
AND2X1 exu_U8043(.A(exu_n4575), .B(exu_n9356), .Y(ecl_ttype_mux_n25));
INVX1 exu_U8044(.A(ecl_ttype_mux_n29), .Y(exu_n16377));
AND2X1 exu_U8045(.A(exu_n4576), .B(exu_n9357), .Y(ecl_ttype_mux_n29));
INVX1 exu_U8046(.A(ecl_ttype_mux_n33), .Y(exu_n16376));
AND2X1 exu_U8047(.A(exu_n4577), .B(exu_n9357), .Y(ecl_ttype_mux_n33));
INVX1 exu_U8048(.A(irf_byp_rs1_data_d_l[71]), .Y(byp_ecc_rs1_synd_d[7]));
INVX1 exu_U8049(.A(irf_byp_rs1_data_d_l[70]), .Y(byp_ecc_rs1_synd_d[6]));
INVX1 exu_U8050(.A(irf_byp_rs1_data_d_l[69]), .Y(byp_ecc_rs1_synd_d[5]));
INVX1 exu_U8051(.A(irf_byp_rs1_data_d_l[68]), .Y(byp_ecc_rs1_synd_d[4]));
INVX1 exu_U8052(.A(irf_byp_rs1_data_d_l[67]), .Y(byp_ecc_rs1_synd_d[3]));
INVX1 exu_U8053(.A(irf_byp_rs1_data_d_l[66]), .Y(byp_ecc_rs1_synd_d[2]));
INVX1 exu_U8054(.A(irf_byp_rs1_data_d_l[65]), .Y(byp_ecc_rs1_synd_d[1]));
INVX1 exu_U8055(.A(irf_byp_rs1_data_d_l[64]), .Y(byp_ecc_rs1_synd_d[0]));
OR2X1 exu_U8056(.A(exu_n12153), .B(exu_n13565), .Y(bypass_rs3h_data_d[31]));
OR2X1 exu_U8057(.A(exu_n12154), .B(exu_n13566), .Y(bypass_rs3h_data_d[30]));
OR2X1 exu_U8058(.A(exu_n12156), .B(exu_n13568), .Y(bypass_rs3h_data_d[29]));
OR2X1 exu_U8059(.A(exu_n12157), .B(exu_n13569), .Y(bypass_rs3h_data_d[28]));
OR2X1 exu_U8060(.A(exu_n12158), .B(exu_n13570), .Y(bypass_rs3h_data_d[27]));
OR2X1 exu_U8061(.A(exu_n12159), .B(exu_n13571), .Y(bypass_rs3h_data_d[26]));
OR2X1 exu_U8062(.A(exu_n12160), .B(exu_n13572), .Y(bypass_rs3h_data_d[25]));
OR2X1 exu_U8063(.A(exu_n12161), .B(exu_n13573), .Y(bypass_rs3h_data_d[24]));
OR2X1 exu_U8064(.A(exu_n12162), .B(exu_n13574), .Y(bypass_rs3h_data_d[23]));
OR2X1 exu_U8065(.A(exu_n12163), .B(exu_n13575), .Y(bypass_rs3h_data_d[22]));
OR2X1 exu_U8066(.A(exu_n12164), .B(exu_n13576), .Y(bypass_rs3h_data_d[21]));
OR2X1 exu_U8067(.A(exu_n12165), .B(exu_n13577), .Y(bypass_rs3h_data_d[20]));
OR2X1 exu_U8068(.A(exu_n12167), .B(exu_n13579), .Y(bypass_rs3h_data_d[19]));
OR2X1 exu_U8069(.A(exu_n12168), .B(exu_n13580), .Y(bypass_rs3h_data_d[18]));
OR2X1 exu_U8070(.A(exu_n12169), .B(exu_n13581), .Y(bypass_rs3h_data_d[17]));
OR2X1 exu_U8071(.A(exu_n12170), .B(exu_n13582), .Y(bypass_rs3h_data_d[16]));
OR2X1 exu_U8072(.A(exu_n12171), .B(exu_n13583), .Y(bypass_rs3h_data_d[15]));
OR2X1 exu_U8073(.A(exu_n12172), .B(exu_n13584), .Y(bypass_rs3h_data_d[14]));
OR2X1 exu_U8074(.A(exu_n12173), .B(exu_n13585), .Y(bypass_rs3h_data_d[13]));
OR2X1 exu_U8075(.A(exu_n12174), .B(exu_n13586), .Y(bypass_rs3h_data_d[12]));
OR2X1 exu_U8076(.A(exu_n12175), .B(exu_n13587), .Y(bypass_rs3h_data_d[11]));
OR2X1 exu_U8077(.A(exu_n12176), .B(exu_n13588), .Y(bypass_rs3h_data_d[10]));
OR2X1 exu_U8078(.A(exu_n12146), .B(exu_n13558), .Y(bypass_rs3h_data_d[9]));
OR2X1 exu_U8079(.A(exu_n12147), .B(exu_n13559), .Y(bypass_rs3h_data_d[8]));
OR2X1 exu_U8080(.A(exu_n12148), .B(exu_n13560), .Y(bypass_rs3h_data_d[7]));
OR2X1 exu_U8081(.A(exu_n12149), .B(exu_n13561), .Y(bypass_rs3h_data_d[6]));
OR2X1 exu_U8082(.A(exu_n12150), .B(exu_n13562), .Y(bypass_rs3h_data_d[5]));
OR2X1 exu_U8083(.A(exu_n12151), .B(exu_n13563), .Y(bypass_rs3h_data_d[4]));
OR2X1 exu_U8084(.A(exu_n12152), .B(exu_n13564), .Y(bypass_rs3h_data_d[3]));
OR2X1 exu_U8085(.A(exu_n12155), .B(exu_n13567), .Y(bypass_rs3h_data_d[2]));
OR2X1 exu_U8086(.A(exu_n12166), .B(exu_n13578), .Y(bypass_rs3h_data_d[1]));
OR2X1 exu_U8087(.A(exu_n12177), .B(exu_n13589), .Y(bypass_rs3h_data_d[0]));
INVX1 exu_U8088(.A(rclk), .Y(bypass_irf_write_clkbuf_n1));
INVX1 exu_U8089(.A(se), .Y(exu_n19281));
INVX1 exu_U8090(.A(se), .Y(exu_n19279));
INVX1 exu_U8091(.A(se), .Y(exu_n19275));
INVX1 exu_U8092(.A(se), .Y(exu_n19273));
INVX1 exu_U8093(.A(se), .Y(exu_n19271));
INVX1 exu_U8094(.A(se), .Y(exu_n19269));
INVX1 exu_U8095(.A(exu_n16159), .Y(exu_n16157));
INVX1 exu_U8096(.A(se), .Y(exu_n19267));
AND2X1 exu_U8097(.A(exu_n15968), .B(exu_n15203), .Y(ecl_byp_rcc_mux1_sel_w2));
INVX1 exu_U8098(.A(shft_shift16_e[3]), .Y(exu_n16142));
INVX1 exu_U8099(.A(ecl_shft_extendbit_e), .Y(exu_n16190));
INVX1 exu_U8100(.A(se), .Y(exu_n19265));
INVX1 exu_U8101(.A(exu_n16270), .Y(exu_n16269));
INVX1 exu_U8102(.A(exu_n16165), .Y(exu_n16170));
INVX1 exu_U8103(.A(exu_n16165), .Y(exu_n16169));
INVX1 exu_U8104(.A(exu_n15380), .Y(exu_n15964));
AND2X1 exu_U8105(.A(exu_n4517), .B(exu_n9320), .Y(ecl_byplog_rs2_n29));
INVX1 exu_U8106(.A(exu_n16204), .Y(exu_n16217));
INVX1 exu_U8107(.A(se), .Y(exu_n19263));
INVX1 exu_U8108(.A(ecl_div_mul_get_new_data), .Y(exu_n16255));
INVX1 exu_U8109(.A(exu_n15979), .Y(exu_n15978));
INVX1 exu_U8110(.A(ecl_div_sel_adder), .Y(exu_n16251));
INVX1 exu_U8111(.A(shft_shift16_e[2]), .Y(exu_n16145));
AND2X1 exu_U8112(.A(exu_n773), .B(exu_n5534), .Y(exu_n19199));
OR2X1 exu_U8113(.A(exu_n13441), .B(exu_n14760), .Y(ecl_byplog_rs1_n17));
INVX1 exu_U8114(.A(ecl_shft_shift4_e[2]), .Y(exu_n16232));
INVX1 exu_U8115(.A(exu_n16203), .Y(exu_n16215));
INVX1 exu_U8116(.A(se), .Y(exu_n19261));
INVX1 exu_U8117(.A(ecl_byp_rcc_mux1_sel_w2), .Y(exu_n16300));
INVX1 exu_U8118(.A(exu_n15968), .Y(exu_n15967));
INVX1 exu_U8119(.A(exu_n15818), .Y(exu_n15965));
INVX1 exu_U8120(.A(ecl_byp_rcc_mux1_sel_w), .Y(exu_n16301));
INVX1 exu_U8121(.A(ecl_mdqctl_ismul_e), .Y(exu_n15985));
INVX1 exu_U8122(.A(exu_n16255), .Y(exu_n16254));
INVX1 exu_U8123(.A(exu_n15381), .Y(exu_n15963));
INVX1 exu_U8124(.A(exu_n15820), .Y(exu_n15966));
INVX1 exu_U8125(.A(exu_n15382), .Y(exu_n15988));
INVX1 exu_U8126(.A(exu_n16196), .Y(exu_n16195));
AND2X1 exu_U8127(.A(ecl_divcntl_cnt6_n26), .B(exu_n9062), .Y(ecl_divcntl_cnt6_n20));
INVX1 exu_U8128(.A(ecl_shft_extendbit_e), .Y(exu_n16191));
OR2X1 exu_U8129(.A(ecl_byplog_rs1_n26), .B(exu_n14756), .Y(ecl_byp_rcc_mux2_sel_usemux1));
AND2X1 exu_U8130(.A(exu_n15201), .B(exu_n9316), .Y(ecl_byp_rs2_mux2_sel_usemux1));
INVX1 exu_U8131(.A(se), .Y(exu_n19259));
INVX1 exu_U8132(.A(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n16315));
INVX1 exu_U8133(.A(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n16298));
AND2X1 exu_U8134(.A(exu_n4151), .B(exu_n9126), .Y(rml_cwp_N99));
INVX1 exu_U8135(.A(ecl_shft_lshift_e_l), .Y(exu_n16236));
INVX1 exu_U8136(.A(ecl_alu_casa_e), .Y(exu_n16262));
INVX1 exu_U8137(.A(exu_n15962), .Y(exu_n15961));
INVX1 exu_U8138(.A(exu_n15972), .Y(exu_n15971));
INVX1 exu_U8139(.A(ecl_byp_rcc_mux2_sel_rf), .Y(exu_n16305));
INVX1 exu_U8140(.A(exu_n19187), .Y(exu_n16004));
AND2X1 exu_U8141(.A(exu_n4519), .B(exu_n15476), .Y(ecl_byplog_rs1_n20));
INVX1 exu_U8142(.A(exu_n16167), .Y(exu_n16165));
INVX1 exu_U8143(.A(exu_n16167), .Y(exu_n16164));
INVX1 exu_U8144(.A(ecl_alu_out_sel_shift_e_l), .Y(exu_n15977));
INVX1 exu_U8145(.A(ecl_shft_shift1_e[0]), .Y(exu_n16223));
INVX1 exu_U8146(.A(ecl_shft_shift1_e[1]), .Y(exu_n16225));
INVX1 exu_U8147(.A(ecl_shft_shift4_e[0]), .Y(exu_n16230));
INVX1 exu_U8148(.A(ecl_div_keep_d), .Y(exu_n16258));
AND2X1 exu_U8149(.A(exu_n747), .B(exu_n5509), .Y(div_xin[63]));
INVX1 exu_U8150(.A(exu_n15976), .Y(exu_n15975));
INVX1 exu_U8151(.A(exu_n15761), .Y(exu_n15989));
INVX1 exu_U8152(.A(ecl_byp_rcc_mux2_sel_e), .Y(exu_n16306));
INVX1 exu_U8153(.A(ecl_byp_rs2_mux1_sel_m), .Y(exu_n16294));
INVX1 exu_U8154(.A(ecl_byp_rs3_mux1_sel_m), .Y(exu_n16290));
INVX1 exu_U8155(.A(exu_n16193), .Y(exu_n16198));
INVX1 exu_U8156(.A(exu_n16196), .Y(exu_n16194));
INVX1 exu_U8157(.A(exu_n16199), .Y(exu_n16193));
AND2X1 exu_U8158(.A(exu_n11662), .B(ifu_exu_inst_vld_w), .Y(ecl_writeback_n149));
INVX1 exu_U8159(.A(ecl_div_ld_inputs), .Y(exu_n16205));
OR2X1 exu_U8160(.A(exu_n15359), .B(exu_n15435), .Y(ecl_byp_rs2_mux1_sel_w));
OR2X1 exu_U8161(.A(ecl_byplog_rs2_n21), .B(exu_n14755), .Y(ecl_byp_rs2_mux2_sel_ld));
OR2X1 exu_U8162(.A(exu_n15357), .B(exu_n15433), .Y(ecl_byp_rs3_mux1_sel_w));
OR2X1 exu_U8163(.A(exu_n19192), .B(exu_n13556), .Y(ecl_byp_rs3_mux2_sel_ld));
AND2X1 exu_U8164(.A(exu_n16402), .B(exu_n9668), .Y(ecl_alu_log_sel_move_e));
OR2X1 exu_U8165(.A(exu_n16401), .B(exu_n14820), .Y(ecl_alu_log_sel_or_e));
AND2X1 exu_U8166(.A(ecl_byplog_rs1_n14), .B(exu_n9321), .Y(ecl_byp_rs1_mux2_sel_usemux1));
OR2X1 exu_U8167(.A(exu_n16401), .B(exu_n14819), .Y(ecl_alu_log_sel_xor_e));
OR2X1 exu_U8168(.A(exu_n16400), .B(exu_n14821), .Y(ecl_alu_log_sel_and_e));
INVX1 exu_U8169(.A(se), .Y(exu_n19257));
AND2X1 exu_U8170(.A(exu_n19235), .B(exu_n5535), .Y(exu_n19223));
OR2X1 exu_U8171(.A(exu_n13451), .B(exu_n14770), .Y(ecl_writeback_n85));
OR2X1 exu_U8172(.A(exu_n13450), .B(exu_n15364), .Y(ecl_writeback_n81));
OR2X1 exu_U8173(.A(exu_n13449), .B(exu_n15364), .Y(ecl_writeback_n77));
OR2X1 exu_U8174(.A(exu_n15358), .B(exu_n15434), .Y(ecl_byp_rs3h_mux1_sel_w));
OR2X1 exu_U8175(.A(exu_n15219), .B(exu_n14765), .Y(ecl_div_yreg_wen_l[1]));
OR2X1 exu_U8176(.A(exu_n15218), .B(exu_n14764), .Y(ecl_div_yreg_wen_l[2]));
OR2X1 exu_U8177(.A(exu_n15217), .B(exu_n14763), .Y(ecl_div_yreg_wen_l[3]));
OR2X1 exu_U8178(.A(exu_n13452), .B(exu_n14771), .Y(ecl_div_yreg_wen_g[0]));
INVX1 exu_U8179(.A(ecl_div_sel_neg32), .Y(exu_n16249));
INVX1 exu_U8180(.A(shft_shift16_e[0]), .Y(exu_n16149));
INVX1 exu_U8181(.A(exu_n16280), .Y(exu_n16279));
INVX1 exu_U8182(.A(alu_invert_e), .Y(exu_n16151));
INVX1 exu_U8183(.A(ecl_byp_sel_pipe_m), .Y(exu_n16274));
INVX1 exu_U8184(.A(ecl_div_yreg_wen_g[0]), .Y(exu_n16245));
INVX1 exu_U8185(.A(exu_n19223), .Y(exu_n16005));
INVX1 exu_U8186(.A(ecl_div_yreg_wen_l[1]), .Y(exu_n16242));
INVX1 exu_U8187(.A(ecl_div_yreg_wen_l[2]), .Y(exu_n16243));
INVX1 exu_U8188(.A(ecl_div_yreg_wen_l[3]), .Y(exu_n16244));
INVX1 exu_U8189(.A(ecl_byp_rs3h_mux1_sel_w), .Y(exu_n16285));
INVX1 exu_U8190(.A(ecl_writeback_n85), .Y(exu_n15980));
INVX1 exu_U8191(.A(ecl_writeback_n81), .Y(exu_n15981));
INVX1 exu_U8192(.A(ecl_writeback_n77), .Y(exu_n15982));
AND2X1 exu_U8193(.A(exu_n15349), .B(exu_n15685), .Y(rml_exu_tlu_spill_e));
INVX1 exu_U8194(.A(exu_n15970), .Y(exu_n15969));
INVX1 exu_U8195(.A(exu_n15023), .Y(exu_n15973));
INVX1 exu_U8196(.A(ecl_div_last_cycle), .Y(exu_n16257));
INVX1 exu_U8197(.A(ecl_byp_rcc_mux1_sel_m), .Y(exu_n16302));
INVX1 exu_U8198(.A(exu_n16229), .Y(exu_n16228));
INVX1 exu_U8199(.A(ecl_shft_shift1_e[2]), .Y(exu_n16227));
INVX1 exu_U8200(.A(exu_n16235), .Y(exu_n16234));
AND2X1 exu_U8201(.A(ifu_exu_restored_e), .B(exu_n9616), .Y(rml_n131));
INVX1 exu_U8202(.A(exu_n15022), .Y(exu_n15974));
INVX1 exu_U8203(.A(exu_n16167), .Y(exu_n16166));
INVX1 exu_U8204(.A(ecl_byp_sel_ifex_m), .Y(exu_n16264));
AND2X1 exu_U8205(.A(exu_n3711), .B(exu_n8790), .Y(div_gencc_in[63]));
INVX1 exu_U8206(.A(exu_n16155), .Y(exu_n16161));
AND2X1 exu_U8207(.A(exu_n15375), .B(exu_n6186), .Y(exu_n25714));
AND2X1 exu_U8208(.A(exu_n1299), .B(exu_n15375), .Y(exu_n25718));
AND2X1 exu_U8209(.A(exu_n1301), .B(exu_n19200), .Y(exu_n25722));
AND2X1 exu_U8210(.A(exu_n1303), .B(exu_n15375), .Y(exu_n25726));
AND2X1 exu_U8211(.A(exu_n1305), .B(exu_n19200), .Y(exu_n25730));
AND2X1 exu_U8212(.A(exu_n1307), .B(exu_n15375), .Y(exu_n25734));
AND2X1 exu_U8213(.A(exu_n1309), .B(exu_n19200), .Y(exu_n25738));
AND2X1 exu_U8214(.A(exu_n1311), .B(exu_n15375), .Y(exu_n25742));
AND2X1 exu_U8215(.A(exu_n1313), .B(exu_n19200), .Y(exu_n25746));
AND2X1 exu_U8216(.A(exu_n1315), .B(exu_n15375), .Y(exu_n25750));
AND2X1 exu_U8217(.A(exu_n1317), .B(exu_n19200), .Y(exu_n25754));
AND2X1 exu_U8218(.A(exu_n1319), .B(exu_n15375), .Y(exu_n25758));
AND2X1 exu_U8219(.A(exu_n1321), .B(exu_n19200), .Y(exu_n25762));
AND2X1 exu_U8220(.A(exu_n4672), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n160));
AND2X1 exu_U8221(.A(exu_n4674), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n166));
AND2X1 exu_U8222(.A(exu_n4676), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n172));
AND2X1 exu_U8223(.A(exu_n4678), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n178));
AND2X1 exu_U8224(.A(exu_n4680), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n184));
AND2X1 exu_U8225(.A(exu_n4682), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n190));
AND2X1 exu_U8226(.A(exu_n15205), .B(exu_n9325), .Y(ecl_eccctl_n21));
AND2X1 exu_U8227(.A(exu_n16618), .B(exu_n9053), .Y(rml_cwp_cwp_output_queue_n22));
AND2X1 exu_U8228(.A(exu_n215), .B(exu_n19285), .Y(exu_n19639));
AND2X1 exu_U8229(.A(exu_n15351), .B(exu_n9667), .Y(ecl_shft_extendbit_e));
INVX1 exu_U8230(.A(exu_n16205), .Y(exu_n16204));
INVX1 exu_U8231(.A(exu_n16203), .Y(exu_n16216));
INVX1 exu_U8232(.A(shft_shift16_e[1]), .Y(exu_n16147));
INVX1 exu_U8233(.A(se), .Y(exu_n19255));
OR2X1 exu_U8234(.A(exu_n19228), .B(exu_n13557), .Y(ecl_byp_rs3h_mux2_sel_ld));
OR2X1 exu_U8235(.A(exu_n15386), .B(exu_n19222), .Y(ecl_byp_rs3h_mux2_sel_e));
INVX1 exu_U8236(.A(exu_n16309), .Y(exu_n16308));
INVX1 exu_U8237(.A(ecl_byp_rs3h_mux1_sel_m), .Y(exu_n16286));
INVX1 exu_U8238(.A(ecl_div_sel_u32), .Y(exu_n16247));
INVX1 exu_U8239(.A(ecl_div_yreg_wen_w[0]), .Y(exu_n16241));
INVX1 exu_U8240(.A(ecl_div_thr_e[0]), .Y(exu_n16220));
OR2X1 exu_U8241(.A(exu_n15356), .B(exu_n16554), .Y(ecl_wb_ccr_wrccr_w));
INVX1 exu_U8242(.A(ecl_byp_restore_m), .Y(exu_n16268));
INVX1 exu_U8243(.A(exu_n16283), .Y(exu_n16282));
INVX1 exu_U8244(.A(exu_n16277), .Y(exu_n16276));
INVX1 exu_U8245(.A(exu_n16317), .Y(exu_n16316));
INVX1 exu_U8246(.A(ecl_byp_rs3h_mux2_sel_ld), .Y(exu_n16287));
INVX1 exu_U8247(.A(ecl_byp_rs3h_mux2_sel_e), .Y(exu_n16288));
OR2X1 exu_U8248(.A(exu_n15436), .B(exu_n16155), .Y(ecl_alu_out_sel_shift_e_l));
AND2X1 exu_U8249(.A(exu_n4557), .B(ecl_ccr_setcc_w2), .Y(ecl_ccr_n19));
AND2X1 exu_U8250(.A(exu_n4555), .B(ecl_ccr_thr_w2[0]), .Y(ecl_ccr_n17));
AND2X1 exu_U8251(.A(exu_n4553), .B(ecl_ccr_thr_w2[1]), .Y(ecl_ccr_n15));
INVX1 exu_U8252(.A(ecl_byp_ldxa_g), .Y(exu_n16270));
AND2X1 exu_U8253(.A(exu_n149), .B(exu_n5116), .Y(alu_addsub_cout64_e));
AND2X1 exu_U8254(.A(exu_n4510), .B(exu_n16205), .Y(ecl_div_sel_adder));
INVX1 exu_U8255(.A(exu_n16251), .Y(exu_n16250));
AND2X1 U8256 ( .A(n773), .B(1'b1), .Y(n19235) );
AND2X1 exu_U8257(.A(exu_n16597), .B(exu_n9339), .Y(ecl_writeback_n50));
XNOR2X1 exu_U8258(.A(exu_n15525), .B(exu_n15526), .Y(exu_n1));
INVX1 exu_U8259(.A(ecl_shiftop_e[2]), .Y(exu_n16154));
INVX1 exu_U8260(.A(ecl_div_muls), .Y(exu_n16185));
INVX1 exu_U8261(.A(exu_n16155), .Y(exu_n16159));
INVX1 exu_U8262(.A(exu_n16156), .Y(exu_n16155));
AND2X1 exu_U8263(.A(exu_n4520), .B(exu_n9322), .Y(ecl_byplog_rs1_n26));
AND2X1 exu_U8264(.A(exu_n1401), .B(exu_n19200), .Y(exu_n25922));
AND2X1 exu_U8265(.A(exu_n1403), .B(exu_n19200), .Y(exu_n25926));
AND2X1 exu_U8266(.A(exu_n1405), .B(exu_n15375), .Y(exu_n25930));
AND2X1 exu_U8267(.A(exu_n1407), .B(exu_n15375), .Y(exu_n25934));
AND2X1 exu_U8268(.A(exu_n1409), .B(exu_n19200), .Y(exu_n25938));
AND2X1 exu_U8269(.A(exu_n1411), .B(exu_n19200), .Y(exu_n25942));
AND2X1 exu_U8270(.A(exu_n1413), .B(exu_n15375), .Y(exu_n25946));
AND2X1 exu_U8271(.A(exu_n1415), .B(exu_n19200), .Y(exu_n25950));
AND2X1 exu_U8272(.A(exu_n1417), .B(exu_n15375), .Y(exu_n25954));
AND2X1 exu_U8273(.A(exu_n1419), .B(exu_n15375), .Y(exu_n25958));
AND2X1 exu_U8274(.A(exu_n1421), .B(exu_n19200), .Y(exu_n25962));
AND2X1 exu_U8275(.A(exu_n1423), .B(exu_n19200), .Y(exu_n25966));
INVX1 exu_U8276(.A(exu_n16169), .Y(exu_n16163));
INVX1 exu_U8277(.A(ecl_std_e), .Y(exu_n16167));
AND2X1 exu_U8278(.A(ecl_byplog_rs2_n29), .B(exu_n9318), .Y(ecl_byplog_rs2_n30));
INVX1 exu_U8279(.A(exu_n19184), .Y(exu_n15962));
AND2X1 exu_U8280(.A(exu_n772), .B(exu_n19186), .Y(exu_n19184));
OR2X1 exu_U8281(.A(exu_n13432), .B(exu_n14751), .Y(ecl_div_sel_div));
AND2X1 exu_U8282(.A(exu_n15424), .B(exu_n16219), .Y(ecl_divcntl_N56));
OR2X1 exu_U8283(.A(ecl_divcntl_div_state_1), .B(exu_n14750), .Y(ecl_div_keep_d));
INVX1 exu_U8284(.A(exu_n16204), .Y(exu_n16219));
OR2X1 exu_U8285(.A(ecl_byp_sel_ecc_m), .B(exu_n15237), .Y(ecl_byp_sel_pipe_m));
OR2X1 exu_U8286(.A(exu_n15358), .B(exu_n19238), .Y(ecl_byp_rs3h_mux1_sel_m));
OR2X1 exu_U8287(.A(exu_n15220), .B(ecl_writeback_n182), .Y(ecl_div_yreg_wen_w[0]));
INVX1 exu_U8288(.A(ecl_div_upper33_zero), .Y(exu_n16246));
INVX1 exu_U8289(.A(ecl_byp_rs3h_longmux_sel_g2), .Y(exu_n16275));
INVX1 exu_U8290(.A(ecl_div_thr_e[1]), .Y(exu_n16221));
AND2X1 exu_U8291(.A(exu_n15689), .B(exu_n15460), .Y(ecc_decode_n27));
INVX1 exu_U8292(.A(ecl_shft_shift4_e[3]), .Y(exu_n16235));
INVX1 exu_U8293(.A(ecl_divcntl_subtract), .Y(exu_n15987));
AND2X1 exu_U8294(.A(exu_n15689), .B(ecc_err_m[3]), .Y(ecc_decode_n35));
INVX1 exu_U8295(.A(bypass_sehold_clk), .Y(exu_n16171));
AND2X1 exu_U8296(.A(div_input_data_e[65]), .B(div_input_data_e[64]), .Y(ecl_shft_shift1_e[3]));
INVX1 exu_U8297(.A(ecl_byp_sel_load_g), .Y(exu_n16272));
INVX1 exu_U8298(.A(exu_n16272), .Y(exu_n16271));
INVX1 exu_U8299(.A(ecl_div_sel_64b), .Y(exu_n16253));
INVX1 exu_U8300(.A(ecl_byp_rs1_mux2_sel_e), .Y(exu_n16317));
INVX1 exu_U8301(.A(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n16283));
INVX1 exu_U8302(.A(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n16280));
INVX1 exu_U8303(.A(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n16277));
INVX1 exu_U8304(.A(ecl_byp_sel_ifusr_e), .Y(exu_n16267));
AND2X1 exu_U8305(.A(exu_n4898), .B(exu_n15817), .Y(rml_rml_kill_w));
INVX1 exu_U8306(.A(ecl_byp_sel_ecc_m), .Y(exu_n16273));
OR2X1 exu_U8307(.A(exu_n15359), .B(ecl_byplog_rs2_n32), .Y(ecl_byp_rs2_mux1_sel_m));
OR2X1 exu_U8308(.A(exu_n15389), .B(ecl_byplog_rs2_n15), .Y(ecl_byp_rs2_mux2_sel_e));
OR2X1 exu_U8309(.A(exu_n15357), .B(exu_n19202), .Y(ecl_byp_rs3_mux1_sel_m));
OR2X1 exu_U8310(.A(exu_n15385), .B(exu_n19186), .Y(ecl_byp_rs3_mux2_sel_e));
OR2X1 exu_U8311(.A(exu_n13445), .B(ecl_writeback_n135), .Y(ecl_rml_cwp_wen_e));
AND2X1 exu_U8312(.A(rml_ecl_other_e), .B(exu_n9614), .Y(rml_n130));
INVX1 exu_U8313(.A(exu_n16170), .Y(exu_n16162));
INVX1 exu_U8314(.A(ecl_alu_out_sel_rs3_e_l), .Y(exu_n15972));
AND2X1 exu_U8315(.A(exu_n4957), .B(exu_n15436), .Y(ecl_alu_out_sel_rs3_e_l));
AND2X1 exu_U8316(.A(ecl_byplog_rs1_n30), .B(exu_n15437), .Y(ecl_byplog_rs1_n24));
AND2X1 exu_U8317(.A(exu_n15690), .B(exu_n16519), .Y(shft_shift16_e[0]));
AND2X1 exu_U8318(.A(exu_n15441), .B(ecc_err_m[1]), .Y(ecc_decode_n21));
AND2X1 exu_U8319(.A(div_input_data_e[68]), .B(exu_n15690), .Y(shft_shift16_e[1]));
AND2X1 exu_U8320(.A(exu_n4516), .B(exu_n15201), .Y(ecl_byp_rs2_mux2_sel_rf));
INVX1 exu_U8321(.A(exu_n16298), .Y(exu_n16297));
AND2X1 exu_U8322(.A(exu_n4518), .B(exu_n16395), .Y(ecl_byp_rs1_mux2_sel_rf));
INVX1 exu_U8323(.A(exu_n16315), .Y(exu_n16314));
AND2X1 exu_U8324(.A(exu_n15236), .B(exu_n15398), .Y(ecl_mdqctl_n63));
INVX1 exu_U8325(.A(ecl_byp_rs1_mux1_sel_w2), .Y(exu_n16307));
AND2X1 exu_U8326(.A(ecl_ldxa_g), .B(ifu_exu_inst_vld_w), .Y(ecl_byp_ldxa_g));
AND2X1 exu_U8327(.A(exu_n4512), .B(exu_n15221), .Y(ecl_div_sel_neg32));
INVX1 exu_U8328(.A(exu_n16249), .Y(exu_n16248));
AND2X1 exu_U8329(.A(ecc_syn_mux_n25), .B(exu_n9372), .Y(ecc_err_m[0]));
AND2X1 exu_U8330(.A(exu_n1323), .B(exu_n19200), .Y(exu_n25766));
AND2X1 exu_U8331(.A(exu_n1325), .B(exu_n15375), .Y(exu_n25770));
AND2X1 exu_U8332(.A(exu_n1327), .B(exu_n19200), .Y(exu_n25774));
AND2X1 exu_U8333(.A(exu_n1329), .B(exu_n15375), .Y(exu_n25778));
AND2X1 exu_U8334(.A(exu_n1331), .B(exu_n19200), .Y(exu_n25782));
AND2X1 exu_U8335(.A(exu_n1333), .B(exu_n15375), .Y(exu_n25786));
AND2X1 exu_U8336(.A(exu_n1335), .B(exu_n15375), .Y(exu_n25790));
AND2X1 exu_U8337(.A(exu_n1337), .B(exu_n19200), .Y(exu_n25794));
AND2X1 exu_U8338(.A(exu_n1339), .B(exu_n15375), .Y(exu_n25798));
AND2X1 exu_U8339(.A(exu_n1341), .B(exu_n19200), .Y(exu_n25802));
AND2X1 exu_U8340(.A(exu_n1343), .B(exu_n19200), .Y(exu_n25806));
AND2X1 exu_U8341(.A(exu_n1345), .B(exu_n15375), .Y(exu_n25810));
AND2X1 exu_U8342(.A(exu_n1347), .B(exu_n15375), .Y(exu_n25814));
AND2X1 exu_U8343(.A(exu_n1349), .B(exu_n15375), .Y(exu_n25818));
AND2X1 exu_U8344(.A(exu_n1351), .B(exu_n15375), .Y(exu_n25822));
AND2X1 exu_U8345(.A(exu_n1353), .B(exu_n19200), .Y(exu_n25826));
AND2X1 exu_U8346(.A(exu_n1355), .B(exu_n15375), .Y(exu_n25830));
AND2X1 exu_U8347(.A(exu_n1357), .B(exu_n19200), .Y(exu_n25834));
AND2X1 exu_U8348(.A(exu_n1359), .B(exu_n19200), .Y(exu_n25838));
AND2X1 exu_U8349(.A(exu_n1361), .B(exu_n15375), .Y(exu_n25842));
AND2X1 exu_U8350(.A(exu_n1363), .B(exu_n15375), .Y(exu_n25846));
AND2X1 exu_U8351(.A(exu_n1365), .B(exu_n19200), .Y(exu_n25850));
AND2X1 exu_U8352(.A(exu_n1367), .B(exu_n15375), .Y(exu_n25854));
AND2X1 exu_U8353(.A(exu_n1369), .B(exu_n19200), .Y(exu_n25858));
AND2X1 exu_U8354(.A(exu_n1371), .B(exu_n19200), .Y(exu_n25862));
AND2X1 exu_U8355(.A(exu_n1373), .B(exu_n15375), .Y(exu_n25866));
AND2X1 exu_U8356(.A(exu_n1375), .B(exu_n19200), .Y(exu_n25870));
AND2X1 exu_U8357(.A(exu_n1377), .B(exu_n15375), .Y(exu_n25874));
AND2X1 exu_U8358(.A(exu_n1379), .B(exu_n15375), .Y(exu_n25878));
AND2X1 exu_U8359(.A(exu_n1381), .B(exu_n15375), .Y(exu_n25882));
AND2X1 exu_U8360(.A(exu_n1383), .B(exu_n19200), .Y(exu_n25886));
AND2X1 exu_U8361(.A(exu_n1385), .B(exu_n15375), .Y(exu_n25890));
AND2X1 exu_U8362(.A(exu_n1387), .B(exu_n19200), .Y(exu_n25894));
AND2X1 exu_U8363(.A(exu_n1389), .B(exu_n19200), .Y(exu_n25898));
AND2X1 exu_U8364(.A(exu_n1391), .B(exu_n19200), .Y(exu_n25902));
AND2X1 exu_U8365(.A(exu_n1393), .B(exu_n15375), .Y(exu_n25906));
AND2X1 exu_U8366(.A(exu_n1395), .B(exu_n19200), .Y(exu_n25910));
AND2X1 exu_U8367(.A(exu_n1397), .B(exu_n15375), .Y(exu_n25914));
AND2X1 exu_U8368(.A(exu_n1399), .B(exu_n19200), .Y(exu_n25918));
AND2X1 exu_U8369(.A(exu_n19236), .B(exu_n9407), .Y(bypass_mux_rs3h_data_1_n4));
AND2X1 exu_U8370(.A(exu_n4622), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n10));
AND2X1 exu_U8371(.A(exu_n4624), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n16));
AND2X1 exu_U8372(.A(exu_n4626), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n22));
AND2X1 exu_U8373(.A(exu_n4628), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n28));
AND2X1 exu_U8374(.A(exu_n4630), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n34));
AND2X1 exu_U8375(.A(exu_n4632), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n40));
AND2X1 exu_U8376(.A(exu_n4634), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n46));
AND2X1 exu_U8377(.A(exu_n4636), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n52));
AND2X1 exu_U8378(.A(exu_n4638), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n58));
AND2X1 exu_U8379(.A(exu_n4640), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n64));
AND2X1 exu_U8380(.A(exu_n4642), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n70));
AND2X1 exu_U8381(.A(exu_n4644), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n76));
AND2X1 exu_U8382(.A(exu_n4646), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n82));
AND2X1 exu_U8383(.A(exu_n4648), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n88));
AND2X1 exu_U8384(.A(exu_n4650), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n94));
AND2X1 exu_U8385(.A(exu_n4652), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n100));
AND2X1 exu_U8386(.A(exu_n4654), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n106));
AND2X1 exu_U8387(.A(exu_n4656), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n112));
AND2X1 exu_U8388(.A(exu_n4658), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n118));
AND2X1 exu_U8389(.A(exu_n4660), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n124));
AND2X1 exu_U8390(.A(exu_n4662), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n130));
AND2X1 exu_U8391(.A(exu_n4664), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n136));
AND2X1 exu_U8392(.A(exu_n4666), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n142));
AND2X1 exu_U8393(.A(exu_n4668), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n148));
AND2X1 exu_U8394(.A(exu_n4670), .B(exu_n19236), .Y(bypass_mux_rs3h_data_1_n154));
OR2X1 exu_U8395(.A(exu_n16398), .B(exu_n15363), .Y(ecl_divcntl_n24));
INVX1 exu_U8396(.A(ecl_alu_out_sel_logic_e_l), .Y(exu_n15970));
AND2X1 exu_U8397(.A(rml_save_e), .B(exu_n15343), .Y(exu_ifu_spill_e));
INVX1 exu_U8398(.A(ecl_shft_shift4_e[2]), .Y(exu_n16233));
AND2X1 exu_U8399(.A(ecc_syn_mux_n9), .B(exu_n9364), .Y(ecc_err_m[4]));
AND2X1 exu_U8400(.A(exu_n4947), .B(exu_n19285), .Y(exu_n19286));
AND2X1 exu_U8401(.A(exu_n4526), .B(exu_n19601), .Y(exu_n19602));
AND2X1 exu_U8402(.A(exu_n4150), .B(exu_n19277), .Y(exu_n19669));
AND2X1 exu_U8403(.A(exu_n4063), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n7));
INVX1 exu_U8404(.A(ecl_div_keep_d), .Y(exu_n16259));
INVX1 exu_U8405(.A(shft_shift16_e[3]), .Y(exu_n16143));
INVX1 exu_U8406(.A(shft_shift16_e[3]), .Y(exu_n16144));
AND2X1 exu_U8407(.A(ecc_syn_mux_n17), .B(exu_n9368), .Y(ecc_err_m[2]));
INVX1 exu_U8408(.A(exu_n16204), .Y(exu_n16218));
INVX1 exu_U8409(.A(exu_n16218), .Y(exu_n16213));
INVX1 exu_U8410(.A(ecl_shft_extendbit_e), .Y(exu_n16189));
AND2X1 exu_U8411(.A(exu_n15381), .B(exu_n9317), .Y(ecl_byplog_rs2_n14));
INVX1 exu_U8412(.A(se), .Y(exu_n19285));
INVX1 exu_U8413(.A(ecl_byp_sel_alu_e), .Y(exu_n16265));
INVX1 exu_U8414(.A(ecl_div_thr_e[2]), .Y(exu_n16222));
AND2X1 exu_U8415(.A(exu_n15460), .B(ecc_err_m[0]), .Y(ecc_decode_n29));
INVX1 exu_U8416(.A(exu_n16151), .Y(exu_n16150));
AND2X1 exu_U8417(.A(exu_n16301), .B(ecl_byplog_rs1_n20), .Y(ecl_byp_rs1_mux1_sel_w));
INVX1 exu_U8418(.A(ecl_byp_rs1_mux1_sel_w), .Y(exu_n16309));
AND2X1 exu_U8419(.A(div_input_data_e[67]), .B(div_input_data_e[66]), .Y(ecl_shft_shift4_e[3]));
INVX1 exu_U8420(.A(ecl_shft_shift1_e[3]), .Y(exu_n16229));
INVX1 exu_U8421(.A(ecl_ecc_sel_rs1_m_l), .Y(exu_n15976));
AND2X1 exu_U8422(.A(exu_n15441), .B(exu_n15461), .Y(ecc_decode_n18));
AND2X1 exu_U8423(.A(exu_n15461), .B(ecc_err_m[2]), .Y(ecc_decode_n22));
OR2X1 exu_U8424(.A(ecl_div_div64), .B(ecl_div_muls), .Y(ecl_div_sel_64b));
INVX1 exu_U8425(.A(exu_n16253), .Y(exu_n16252));
AND2X1 exu_U8426(.A(ecl_byplog_rs1_n20), .B(exu_n15769), .Y(ecl_byp_rs1_mux2_sel_e));
AND2X1 exu_U8427(.A(exu_n15968), .B(exu_n15465), .Y(ecl_byp_rs1_longmux_sel_w2));
AND2X1 exu_U8428(.A(exu_n15820), .B(exu_n15464), .Y(ecl_byp_rs2_longmux_sel_w2));
AND2X1 exu_U8429(.A(exu_n15818), .B(exu_n15462), .Y(ecl_byp_rs3_longmux_sel_w2));
AND2X1 exu_U8430(.A(exu_n16265), .B(ifu_exu_rd_ifusr_e), .Y(ecl_byp_sel_ifusr_e));
INVX1 exu_U8431(.A(exu_n16267), .Y(exu_n16266));
INVX1 exu_U8432(.A(ecl_byp_rs1_mux1_sel_m), .Y(exu_n16311));
AND2X1 exu_U8433(.A(exu_n16302), .B(ecl_byplog_rs1_n20), .Y(ecl_byp_rs1_mux1_sel_m));
INVX1 exu_U8434(.A(exu_n16311), .Y(exu_n16310));
OR2X1 exu_U8435(.A(exu_ifu_err_reg_m[4]), .B(exu_ifu_err_reg_m[3]), .Y(ecl_eccctl_n25));
AND2X1 exu_U8436(.A(ecc_syn_mux_n13), .B(exu_n9366), .Y(ecc_err_m[3]));
INVX1 exu_U8437(.A(ecl_shft_shift1_e[0]), .Y(exu_n16224));
OR2X1 exu_U8438(.A(exu_n15362), .B(exu_n14817), .Y(ecl_pick_not_aligned));
AND2X1 exu_U8439(.A(exu_n19199), .B(exu_n5532), .Y(exu_n19200));
INVX1 exu_U8440(.A(ecl_byplog_rs1_n22), .Y(exu_n15968));
AND2X1 exu_U8441(.A(exu_n172), .B(exu_n15941), .Y(exu_n17462));
AND2X1 exu_U8442(.A(exu_n173), .B(exu_n15941), .Y(exu_n17463));
AND2X1 exu_U8443(.A(exu_n174), .B(exu_n15941), .Y(exu_n17464));
AND2X1 exu_U8444(.A(exu_n158), .B(exu_n15941), .Y(exu_n17465));
AND2X1 exu_U8445(.A(exu_n159), .B(exu_n15941), .Y(exu_n17466));
AND2X1 exu_U8446(.A(exu_n160), .B(exu_n15941), .Y(exu_n17467));
AND2X1 exu_U8447(.A(exu_n161), .B(exu_n15941), .Y(exu_n17468));
AND2X1 exu_U8448(.A(exu_n162), .B(exu_n15941), .Y(exu_n17469));
AND2X1 exu_U8449(.A(exu_n164), .B(exu_n15941), .Y(exu_n17470));
AND2X1 exu_U8450(.A(exu_n166), .B(exu_n15941), .Y(exu_n17471));
AND2X1 exu_U8451(.A(exu_n168), .B(exu_n15941), .Y(exu_n17472));
AND2X1 exu_U8452(.A(exu_n170), .B(exu_n15941), .Y(exu_n17473));
AND2X1 exu_U8453(.A(exu_n175), .B(exu_n15941), .Y(exu_n17474));
AND2X1 exu_U8454(.A(exu_n191), .B(exu_n15942), .Y(exu_n17478));
AND2X1 exu_U8455(.A(exu_n192), .B(exu_n15942), .Y(exu_n17479));
AND2X1 exu_U8456(.A(exu_n193), .B(exu_n15942), .Y(exu_n17480));
AND2X1 exu_U8457(.A(exu_n177), .B(exu_n15942), .Y(exu_n17481));
AND2X1 exu_U8458(.A(exu_n178), .B(exu_n15942), .Y(exu_n17482));
AND2X1 exu_U8459(.A(exu_n179), .B(exu_n15942), .Y(exu_n17483));
AND2X1 exu_U8460(.A(exu_n180), .B(exu_n15942), .Y(exu_n17484));
AND2X1 exu_U8461(.A(exu_n181), .B(exu_n15942), .Y(exu_n17485));
AND2X1 exu_U8462(.A(exu_n183), .B(exu_n15942), .Y(exu_n17486));
AND2X1 exu_U8463(.A(exu_n185), .B(exu_n15942), .Y(exu_n17487));
AND2X1 exu_U8464(.A(exu_n187), .B(exu_n15942), .Y(exu_n17488));
AND2X1 exu_U8465(.A(exu_n189), .B(exu_n15942), .Y(exu_n17489));
AND2X1 exu_U8466(.A(exu_n194), .B(exu_n15942), .Y(exu_n17490));
AND2X1 exu_U8467(.A(exu_n210), .B(exu_n15943), .Y(exu_n17493));
AND2X1 exu_U8468(.A(exu_n211), .B(exu_n15943), .Y(exu_n17494));
AND2X1 exu_U8469(.A(exu_n212), .B(exu_n15943), .Y(exu_n17495));
AND2X1 exu_U8470(.A(exu_n196), .B(exu_n15943), .Y(exu_n17496));
AND2X1 exu_U8471(.A(exu_n197), .B(exu_n15943), .Y(exu_n17497));
AND2X1 exu_U8472(.A(exu_n198), .B(exu_n15943), .Y(exu_n17498));
AND2X1 exu_U8473(.A(exu_n199), .B(exu_n15943), .Y(exu_n17499));
AND2X1 exu_U8474(.A(exu_n200), .B(exu_n15943), .Y(exu_n17500));
AND2X1 exu_U8475(.A(exu_n202), .B(exu_n15943), .Y(exu_n17501));
AND2X1 exu_U8476(.A(exu_n204), .B(exu_n15943), .Y(exu_n17502));
AND2X1 exu_U8477(.A(exu_n206), .B(exu_n15943), .Y(exu_n17503));
AND2X1 exu_U8478(.A(exu_n208), .B(exu_n15943), .Y(exu_n17504));
AND2X1 exu_U8479(.A(exu_n213), .B(exu_n15943), .Y(exu_n17505));
AND2X1 exu_U8480(.A(exu_n4067), .B(exu_n17619), .Y(exu_n17620));
AND2X1 exu_U8481(.A(exu_n4068), .B(exu_n17619), .Y(exu_n17621));
AND2X1 exu_U8482(.A(exu_n4069), .B(exu_n17619), .Y(exu_n17622));
AND2X1 exu_U8483(.A(exu_n4070), .B(exu_n17619), .Y(exu_n17623));
AND2X1 exu_U8484(.A(exu_n15024), .B(exu_n9116), .Y(exu_n17980));
AND2X1 exu_U8485(.A(exu_n394), .B(exu_n18198), .Y(exu_n18195));
AND2X1 exu_U8486(.A(exu_n393), .B(exu_n18198), .Y(exu_n18196));
AND2X1 exu_U8487(.A(exu_n392), .B(exu_n18198), .Y(exu_n18197));
AND2X1 exu_U8488(.A(exu_n397), .B(exu_n18202), .Y(exu_n18199));
AND2X1 exu_U8489(.A(exu_n396), .B(exu_n18202), .Y(exu_n18200));
AND2X1 exu_U8490(.A(exu_n395), .B(exu_n18202), .Y(exu_n18201));
AND2X1 exu_U8491(.A(exu_n400), .B(exu_n18206), .Y(exu_n18203));
AND2X1 exu_U8492(.A(exu_n399), .B(exu_n18206), .Y(exu_n18204));
AND2X1 exu_U8493(.A(exu_n398), .B(exu_n18206), .Y(exu_n18205));
AND2X1 exu_U8494(.A(exu_n403), .B(exu_n18210), .Y(exu_n18207));
AND2X1 exu_U8495(.A(exu_n402), .B(exu_n18210), .Y(exu_n18208));
AND2X1 exu_U8496(.A(exu_n401), .B(exu_n18210), .Y(exu_n18209));
AND2X1 exu_U8497(.A(exu_n406), .B(exu_n18242), .Y(exu_n18239));
AND2X1 exu_U8498(.A(exu_n405), .B(exu_n18242), .Y(exu_n18240));
AND2X1 exu_U8499(.A(exu_n404), .B(exu_n18242), .Y(exu_n18241));
AND2X1 exu_U8500(.A(exu_n409), .B(exu_n18246), .Y(exu_n18243));
AND2X1 exu_U8501(.A(exu_n408), .B(exu_n18246), .Y(exu_n18244));
AND2X1 exu_U8502(.A(exu_n407), .B(exu_n18246), .Y(exu_n18245));
AND2X1 exu_U8503(.A(exu_n412), .B(exu_n18250), .Y(exu_n18247));
AND2X1 exu_U8504(.A(exu_n411), .B(exu_n18250), .Y(exu_n18248));
AND2X1 exu_U8505(.A(exu_n410), .B(exu_n18250), .Y(exu_n18249));
AND2X1 exu_U8506(.A(exu_n415), .B(exu_n18254), .Y(exu_n18251));
AND2X1 exu_U8507(.A(exu_n414), .B(exu_n18254), .Y(exu_n18252));
AND2X1 exu_U8508(.A(exu_n413), .B(exu_n18254), .Y(exu_n18253));
AND2X1 exu_U8509(.A(exu_n418), .B(exu_n18286), .Y(exu_n18283));
AND2X1 exu_U8510(.A(exu_n417), .B(exu_n18286), .Y(exu_n18284));
AND2X1 exu_U8511(.A(exu_n416), .B(exu_n18286), .Y(exu_n18285));
AND2X1 exu_U8512(.A(exu_n421), .B(exu_n18290), .Y(exu_n18287));
AND2X1 exu_U8513(.A(exu_n420), .B(exu_n18290), .Y(exu_n18288));
AND2X1 exu_U8514(.A(exu_n419), .B(exu_n18290), .Y(exu_n18289));
AND2X1 exu_U8515(.A(exu_n424), .B(exu_n18294), .Y(exu_n18291));
AND2X1 exu_U8516(.A(exu_n423), .B(exu_n18294), .Y(exu_n18292));
AND2X1 exu_U8517(.A(exu_n422), .B(exu_n18294), .Y(exu_n18293));
AND2X1 exu_U8518(.A(exu_n427), .B(exu_n18298), .Y(exu_n18295));
AND2X1 exu_U8519(.A(exu_n426), .B(exu_n18298), .Y(exu_n18296));
AND2X1 exu_U8520(.A(exu_n425), .B(exu_n18298), .Y(exu_n18297));
AND2X1 exu_U8521(.A(exu_n430), .B(exu_n18330), .Y(exu_n18327));
AND2X1 exu_U8522(.A(exu_n429), .B(exu_n18330), .Y(exu_n18328));
AND2X1 exu_U8523(.A(exu_n428), .B(exu_n18330), .Y(exu_n18329));
AND2X1 exu_U8524(.A(exu_n433), .B(exu_n18334), .Y(exu_n18331));
AND2X1 exu_U8525(.A(exu_n432), .B(exu_n18334), .Y(exu_n18332));
AND2X1 exu_U8526(.A(exu_n431), .B(exu_n18334), .Y(exu_n18333));
AND2X1 exu_U8527(.A(exu_n436), .B(exu_n18338), .Y(exu_n18335));
AND2X1 exu_U8528(.A(exu_n435), .B(exu_n18338), .Y(exu_n18336));
AND2X1 exu_U8529(.A(exu_n434), .B(exu_n18338), .Y(exu_n18337));
AND2X1 exu_U8530(.A(exu_n439), .B(exu_n18342), .Y(exu_n18339));
AND2X1 exu_U8531(.A(exu_n438), .B(exu_n18342), .Y(exu_n18340));
AND2X1 exu_U8532(.A(exu_n437), .B(exu_n18342), .Y(exu_n18341));
AND2X1 exu_U8533(.A(exu_n442), .B(exu_n18370), .Y(exu_n18367));
AND2X1 exu_U8534(.A(exu_n441), .B(exu_n18370), .Y(exu_n18368));
AND2X1 exu_U8535(.A(exu_n440), .B(exu_n18370), .Y(exu_n18369));
AND2X1 exu_U8536(.A(exu_n445), .B(exu_n18374), .Y(exu_n18371));
AND2X1 exu_U8537(.A(exu_n444), .B(exu_n18374), .Y(exu_n18372));
AND2X1 exu_U8538(.A(exu_n443), .B(exu_n18374), .Y(exu_n18373));
AND2X1 exu_U8539(.A(exu_n448), .B(exu_n18378), .Y(exu_n18375));
AND2X1 exu_U8540(.A(exu_n447), .B(exu_n18378), .Y(exu_n18376));
AND2X1 exu_U8541(.A(exu_n446), .B(exu_n18378), .Y(exu_n18377));
AND2X1 exu_U8542(.A(exu_n451), .B(exu_n18382), .Y(exu_n18379));
AND2X1 exu_U8543(.A(exu_n450), .B(exu_n18382), .Y(exu_n18380));
AND2X1 exu_U8544(.A(exu_n449), .B(exu_n18382), .Y(exu_n18381));
AND2X1 exu_U8545(.A(exu_n4143), .B(exu_n18412), .Y(exu_n18413));
AND2X1 exu_U8546(.A(exu_n4144), .B(exu_n18412), .Y(exu_n18414));
AND2X1 exu_U8547(.A(exu_n4145), .B(exu_n18412), .Y(exu_n18415));
AND2X1 exu_U8548(.A(exu_n4146), .B(exu_n18412), .Y(exu_n18416));
AND2X1 exu_U8549(.A(exu_n676), .B(exu_n15992), .Y(exu_n18568));
AND2X1 exu_U8550(.A(exu_n679), .B(exu_n15992), .Y(exu_n18570));
AND2X1 exu_U8551(.A(exu_n682), .B(exu_n15992), .Y(exu_n18571));
AND2X1 exu_U8552(.A(exu_n685), .B(exu_n15992), .Y(exu_n18572));
AND2X1 exu_U8553(.A(exu_n688), .B(exu_n15992), .Y(exu_n18573));
AND2X1 exu_U8554(.A(exu_n691), .B(exu_n15992), .Y(exu_n18574));
AND2X1 exu_U8555(.A(exu_n694), .B(exu_n15992), .Y(exu_n18575));
AND2X1 exu_U8556(.A(exu_n697), .B(exu_n15992), .Y(exu_n18576));
AND2X1 exu_U8557(.A(exu_n702), .B(exu_n15991), .Y(exu_n18577));
AND2X1 exu_U8558(.A(exu_n705), .B(exu_n15991), .Y(exu_n18578));
AND2X1 exu_U8559(.A(exu_n708), .B(exu_n15991), .Y(exu_n18579));
AND2X1 exu_U8560(.A(exu_n711), .B(exu_n15991), .Y(exu_n18581));
AND2X1 exu_U8561(.A(exu_n714), .B(exu_n15991), .Y(exu_n18582));
AND2X1 exu_U8562(.A(exu_n717), .B(exu_n15991), .Y(exu_n18583));
AND2X1 exu_U8563(.A(exu_n720), .B(exu_n15991), .Y(exu_n18584));
AND2X1 exu_U8564(.A(exu_n721), .B(exu_n15991), .Y(exu_n18585));
AND2X1 exu_U8565(.A(exu_n722), .B(exu_n15991), .Y(exu_n18586));
AND2X1 exu_U8566(.A(exu_n723), .B(exu_n15991), .Y(exu_n18587));
AND2X1 exu_U8567(.A(exu_n726), .B(exu_n15991), .Y(exu_n18588));
AND2X1 exu_U8568(.A(exu_n727), .B(exu_n15991), .Y(exu_n18589));
AND2X1 exu_U8569(.A(exu_n728), .B(exu_n15990), .Y(exu_n18590));
AND2X1 exu_U8570(.A(exu_n729), .B(exu_n15990), .Y(exu_n18592));
AND2X1 exu_U8571(.A(exu_n730), .B(exu_n15990), .Y(exu_n18593));
AND2X1 exu_U8572(.A(exu_n731), .B(exu_n15990), .Y(exu_n18594));
AND2X1 exu_U8573(.A(exu_n732), .B(exu_n15990), .Y(exu_n18595));
AND2X1 exu_U8574(.A(exu_n733), .B(exu_n15990), .Y(exu_n18596));
AND2X1 exu_U8575(.A(exu_n734), .B(exu_n15990), .Y(exu_n18597));
AND2X1 exu_U8576(.A(exu_n735), .B(exu_n15990), .Y(exu_n18598));
AND2X1 exu_U8577(.A(exu_n477), .B(exu_n15990), .Y(exu_n18599));
AND2X1 exu_U8578(.A(exu_n478), .B(exu_n15990), .Y(exu_n18600));
AND2X1 exu_U8579(.A(exu_n481), .B(exu_n15990), .Y(exu_n18601));
AND2X1 exu_U8580(.A(exu_n484), .B(exu_n15999), .Y(exu_n18475));
AND2X1 exu_U8581(.A(exu_n487), .B(exu_n15999), .Y(exu_n18476));
AND2X1 exu_U8582(.A(exu_n489), .B(exu_n15999), .Y(exu_n18477));
AND2X1 exu_U8583(.A(exu_n491), .B(exu_n15999), .Y(exu_n18478));
AND2X1 exu_U8584(.A(exu_n493), .B(exu_n15999), .Y(exu_n18479));
AND2X1 exu_U8585(.A(exu_n495), .B(exu_n15999), .Y(exu_n18480));
AND2X1 exu_U8586(.A(exu_n497), .B(exu_n15999), .Y(exu_n18481));
AND2X1 exu_U8587(.A(exu_n501), .B(exu_n15999), .Y(exu_n18482));
AND2X1 exu_U8588(.A(exu_n503), .B(exu_n15999), .Y(exu_n18483));
AND2X1 exu_U8589(.A(exu_n505), .B(exu_n15999), .Y(exu_n18484));
AND2X1 exu_U8590(.A(exu_n507), .B(exu_n15998), .Y(exu_n18486));
AND2X1 exu_U8591(.A(exu_n509), .B(exu_n15998), .Y(exu_n18487));
AND2X1 exu_U8592(.A(exu_n511), .B(exu_n15998), .Y(exu_n18488));
AND2X1 exu_U8593(.A(exu_n513), .B(exu_n15998), .Y(exu_n18489));
AND2X1 exu_U8594(.A(exu_n515), .B(exu_n15998), .Y(exu_n18490));
AND2X1 exu_U8595(.A(exu_n517), .B(exu_n15998), .Y(exu_n18491));
AND2X1 exu_U8596(.A(exu_n519), .B(exu_n15998), .Y(exu_n18492));
AND2X1 exu_U8597(.A(exu_n523), .B(exu_n15998), .Y(exu_n18493));
AND2X1 exu_U8598(.A(exu_n525), .B(exu_n15998), .Y(exu_n18494));
AND2X1 exu_U8599(.A(exu_n527), .B(exu_n15998), .Y(exu_n18495));
AND2X1 exu_U8600(.A(exu_n529), .B(exu_n15998), .Y(exu_n18497));
AND2X1 exu_U8601(.A(exu_n531), .B(exu_n15998), .Y(exu_n18498));
AND2X1 exu_U8602(.A(exu_n533), .B(exu_n15997), .Y(exu_n18499));
AND2X1 exu_U8603(.A(exu_n535), .B(exu_n15997), .Y(exu_n18500));
AND2X1 exu_U8604(.A(exu_n537), .B(exu_n15997), .Y(exu_n18501));
AND2X1 exu_U8605(.A(exu_n539), .B(exu_n15997), .Y(exu_n18502));
AND2X1 exu_U8606(.A(exu_n541), .B(exu_n15997), .Y(exu_n18503));
AND2X1 exu_U8607(.A(exu_n545), .B(exu_n15997), .Y(exu_n18504));
AND2X1 exu_U8608(.A(exu_n547), .B(exu_n15997), .Y(exu_n18505));
AND2X1 exu_U8609(.A(exu_n549), .B(exu_n15997), .Y(exu_n18506));
AND2X1 exu_U8610(.A(exu_n551), .B(exu_n15997), .Y(exu_n18508));
AND2X1 exu_U8611(.A(exu_n553), .B(exu_n15997), .Y(exu_n18509));
AND2X1 exu_U8612(.A(exu_n555), .B(exu_n15997), .Y(exu_n18510));
AND2X1 exu_U8613(.A(exu_n557), .B(exu_n15997), .Y(exu_n18511));
AND2X1 exu_U8614(.A(exu_n558), .B(exu_n15996), .Y(exu_n18512));
AND2X1 exu_U8615(.A(exu_n561), .B(exu_n15996), .Y(exu_n18513));
AND2X1 exu_U8616(.A(exu_n564), .B(exu_n15996), .Y(exu_n18514));
AND2X1 exu_U8617(.A(exu_n569), .B(exu_n15996), .Y(exu_n18515));
AND2X1 exu_U8618(.A(exu_n572), .B(exu_n15996), .Y(exu_n18516));
AND2X1 exu_U8619(.A(exu_n575), .B(exu_n15996), .Y(exu_n18517));
AND2X1 exu_U8620(.A(exu_n578), .B(exu_n15996), .Y(exu_n18519));
AND2X1 exu_U8621(.A(exu_n581), .B(exu_n15996), .Y(exu_n18520));
AND2X1 exu_U8622(.A(exu_n584), .B(exu_n15996), .Y(exu_n18521));
AND2X1 exu_U8623(.A(exu_n587), .B(exu_n15996), .Y(exu_n18522));
AND2X1 exu_U8624(.A(exu_n590), .B(exu_n15996), .Y(exu_n18523));
AND2X1 exu_U8625(.A(exu_n593), .B(exu_n15996), .Y(exu_n18524));
AND2X1 exu_U8626(.A(exu_n596), .B(exu_n15995), .Y(exu_n18525));
AND2X1 exu_U8627(.A(exu_n601), .B(exu_n15995), .Y(exu_n18526));
AND2X1 exu_U8628(.A(exu_n604), .B(exu_n15995), .Y(exu_n18527));
AND2X1 exu_U8629(.A(exu_n607), .B(exu_n15995), .Y(exu_n18528));
AND2X1 exu_U8630(.A(exu_n610), .B(exu_n15995), .Y(exu_n18530));
AND2X1 exu_U8631(.A(exu_n613), .B(exu_n15995), .Y(exu_n18531));
AND2X1 exu_U8632(.A(exu_n616), .B(exu_n15995), .Y(exu_n18532));
AND2X1 exu_U8633(.A(exu_n617), .B(exu_n15995), .Y(exu_n18533));
AND2X1 exu_U8634(.A(exu_n618), .B(exu_n15995), .Y(exu_n18534));
AND2X1 exu_U8635(.A(exu_n619), .B(exu_n15995), .Y(exu_n18535));
AND2X1 exu_U8636(.A(exu_n620), .B(exu_n15995), .Y(exu_n18536));
AND2X1 exu_U8637(.A(exu_n623), .B(exu_n15995), .Y(exu_n18537));
AND2X1 exu_U8638(.A(exu_n624), .B(exu_n15994), .Y(exu_n18538));
AND2X1 exu_U8639(.A(exu_n625), .B(exu_n15994), .Y(exu_n18539));
AND2X1 exu_U8640(.A(exu_n626), .B(exu_n15994), .Y(exu_n18541));
AND2X1 exu_U8641(.A(exu_n627), .B(exu_n15994), .Y(exu_n18542));
AND2X1 exu_U8642(.A(exu_n628), .B(exu_n15994), .Y(exu_n18543));
AND2X1 exu_U8643(.A(exu_n629), .B(exu_n15994), .Y(exu_n18544));
AND2X1 exu_U8644(.A(exu_n630), .B(exu_n15994), .Y(exu_n18545));
AND2X1 exu_U8645(.A(exu_n632), .B(exu_n15994), .Y(exu_n18546));
AND2X1 exu_U8646(.A(exu_n634), .B(exu_n15994), .Y(exu_n18547));
AND2X1 exu_U8647(.A(exu_n638), .B(exu_n15994), .Y(exu_n18548));
AND2X1 exu_U8648(.A(exu_n640), .B(exu_n15994), .Y(exu_n18549));
AND2X1 exu_U8649(.A(exu_n642), .B(exu_n15994), .Y(exu_n18550));
AND2X1 exu_U8650(.A(exu_n644), .B(exu_n15993), .Y(exu_n18552));
AND2X1 exu_U8651(.A(exu_n646), .B(exu_n15993), .Y(exu_n18553));
AND2X1 exu_U8652(.A(exu_n648), .B(exu_n15993), .Y(exu_n18554));
AND2X1 exu_U8653(.A(exu_n650), .B(exu_n15993), .Y(exu_n18555));
AND2X1 exu_U8654(.A(exu_n652), .B(exu_n15993), .Y(exu_n18556));
AND2X1 exu_U8655(.A(exu_n654), .B(exu_n15993), .Y(exu_n18557));
AND2X1 exu_U8656(.A(exu_n656), .B(exu_n15993), .Y(exu_n18558));
AND2X1 exu_U8657(.A(exu_n660), .B(exu_n15993), .Y(exu_n18559));
AND2X1 exu_U8658(.A(exu_n662), .B(exu_n15993), .Y(exu_n18560));
AND2X1 exu_U8659(.A(exu_n664), .B(exu_n15993), .Y(exu_n18561));
AND2X1 exu_U8660(.A(exu_n666), .B(exu_n15993), .Y(exu_n18562));
AND2X1 exu_U8661(.A(exu_n668), .B(exu_n15993), .Y(exu_n18563));
AND2X1 exu_U8662(.A(exu_n670), .B(exu_n15992), .Y(exu_n18564));
AND2X1 exu_U8663(.A(exu_n672), .B(exu_n15992), .Y(exu_n18565));
AND2X1 exu_U8664(.A(exu_n674), .B(exu_n15992), .Y(exu_n18566));
AND2X1 exu_U8665(.A(exu_n700), .B(exu_n15992), .Y(exu_n18567));
AND2X1 exu_U8666(.A(exu_n724), .B(exu_n15992), .Y(exu_n18569));
AND2X1 exu_U8667(.A(exu_n475), .B(exu_n15991), .Y(exu_n18580));
AND2X1 exu_U8668(.A(exu_n499), .B(exu_n15990), .Y(exu_n18591));
AND2X1 exu_U8669(.A(exu_n521), .B(exu_n15990), .Y(exu_n18602));
AND2X1 exu_U8670(.A(exu_n543), .B(exu_n15999), .Y(exu_n18485));
AND2X1 exu_U8671(.A(exu_n567), .B(exu_n15998), .Y(exu_n18496));
AND2X1 exu_U8672(.A(exu_n599), .B(exu_n15997), .Y(exu_n18507));
AND2X1 exu_U8673(.A(exu_n621), .B(exu_n15996), .Y(exu_n18518));
AND2X1 exu_U8674(.A(exu_n636), .B(exu_n15995), .Y(exu_n18529));
AND2X1 exu_U8675(.A(exu_n658), .B(exu_n15994), .Y(exu_n18540));
AND2X1 exu_U8676(.A(exu_n737), .B(exu_n15993), .Y(exu_n18551));
AND2X1 exu_U8677(.A(exu_n4030), .B(exu_n15024), .Y(exu_n19251));
AND2X1 exu_U8678(.A(exu_n4031), .B(exu_n15024), .Y(exu_n19252));
AND2X1 exu_U8679(.A(exu_n4032), .B(exu_n15024), .Y(exu_n19253));
AND2X1 exu_U8680(.A(exu_n4033), .B(exu_n15024), .Y(exu_n19254));
AND2X1 exu_U8681(.A(exu_n4955), .B(exu_n19277), .Y(exu_n19278));
AND2X1 exu_U8682(.A(exu_n4484), .B(exu_n19297), .Y(exu_n19298));
AND2X1 exu_U8683(.A(exu_n4948), .B(exu_n19303), .Y(exu_n19304));
AND2X1 exu_U8684(.A(exu_n4954), .B(exu_n19313), .Y(exu_n19314));
AND2X1 exu_U8685(.A(exu_n4963), .B(exu_n19319), .Y(exu_n19320));
AND2X1 exu_U8686(.A(exu_n4960), .B(exu_n19321), .Y(exu_n19322));
AND2X1 exu_U8687(.A(exu_n4958), .B(exu_n19329), .Y(exu_n19330));
AND2X1 exu_U8688(.A(exu_n4959), .B(exu_n19331), .Y(exu_n19332));
AND2X1 exu_U8689(.A(exu_n4962), .B(exu_n19333), .Y(exu_n19334));
AND2X1 exu_U8690(.A(exu_n4956), .B(exu_n19335), .Y(exu_n19336));
AND2X1 exu_U8691(.A(exu_n4895), .B(exu_n19355), .Y(exu_n19356));
AND2X1 exu_U8692(.A(exu_n4896), .B(exu_n19357), .Y(exu_n19358));
AND2X1 exu_U8693(.A(exu_n4542), .B(exu_n19581), .Y(exu_n19582));
AND2X1 exu_U8694(.A(exu_n4525), .B(exu_n19583), .Y(exu_n19584));
AND2X1 exu_U8695(.A(exu_n4532), .B(exu_n19585), .Y(exu_n19586));
AND2X1 exu_U8696(.A(exu_n4529), .B(exu_n19589), .Y(exu_n19590));
AND2X1 exu_U8697(.A(exu_n4530), .B(exu_n19605), .Y(exu_n19606));
AND2X1 exu_U8698(.A(exu_n4523), .B(exu_n19615), .Y(exu_n19616));
AND2X1 exu_U8699(.A(exu_n4521), .B(exu_n19617), .Y(exu_n19618));
AND2X1 exu_U8700(.A(exu_n4066), .B(exu_n19637), .Y(exu_n19638));
AND2X1 exu_U8701(.A(exu_n4508), .B(exu_n19642), .Y(exu_n19643));
AND2X1 exu_U8702(.A(exu_n4507), .B(exu_n19644), .Y(exu_n19645));
AND2X1 exu_U8703(.A(exu_n4506), .B(exu_n19646), .Y(exu_n19647));
AND2X1 exu_U8704(.A(exu_n4500), .B(exu_n19648), .Y(exu_n19649));
AND2X1 exu_U8705(.A(exu_n4488), .B(exu_n19275), .Y(exu_n19660));
AND2X1 exu_U8706(.A(exu_n4489), .B(exu_n19273), .Y(exu_n19661));
AND2X1 exu_U8707(.A(exu_n4158), .B(exu_n19674), .Y(exu_n19675));
AND2X1 exu_U8708(.A(exu_n4157), .B(exu_n19674), .Y(exu_n19676));
AND2X1 exu_U8709(.A(exu_n4156), .B(exu_n19674), .Y(exu_n19677));
AND2X1 exu_U8710(.A(exu_n4142), .B(exu_n19686), .Y(exu_n19687));
AND2X1 exu_U8711(.A(exu_n4141), .B(exu_n19686), .Y(exu_n19688));
AND2X1 exu_U8712(.A(exu_n4140), .B(exu_n19686), .Y(exu_n19689));
AND2X1 exu_U8713(.A(exu_n456), .B(exu_n19694), .Y(exu_n19695));
AND2X1 exu_U8714(.A(exu_n455), .B(exu_n19694), .Y(exu_n19696));
AND2X1 exu_U8715(.A(exu_n454), .B(exu_n19694), .Y(exu_n19697));
AND2X1 exu_U8716(.A(exu_n459), .B(exu_n19702), .Y(exu_n19703));
AND2X1 exu_U8717(.A(exu_n458), .B(exu_n19702), .Y(exu_n19704));
AND2X1 exu_U8718(.A(exu_n457), .B(exu_n19702), .Y(exu_n19705));
AND2X1 exu_U8719(.A(exu_n462), .B(exu_n19710), .Y(exu_n19711));
AND2X1 exu_U8720(.A(exu_n461), .B(exu_n19710), .Y(exu_n19712));
AND2X1 exu_U8721(.A(exu_n460), .B(exu_n19710), .Y(exu_n19713));
AND2X1 exu_U8722(.A(exu_n465), .B(exu_n19766), .Y(exu_n19767));
AND2X1 exu_U8723(.A(exu_n464), .B(exu_n19766), .Y(exu_n19768));
AND2X1 exu_U8724(.A(exu_n463), .B(exu_n19766), .Y(exu_n19769));
AND2X1 exu_U8725(.A(exu_n468), .B(exu_n19770), .Y(exu_n19771));
AND2X1 exu_U8726(.A(exu_n467), .B(exu_n19770), .Y(exu_n19772));
AND2X1 exu_U8727(.A(exu_n466), .B(exu_n19770), .Y(exu_n19773));
AND2X1 exu_U8728(.A(exu_n471), .B(exu_n19774), .Y(exu_n19775));
AND2X1 exu_U8729(.A(exu_n470), .B(exu_n19774), .Y(exu_n19776));
AND2X1 exu_U8730(.A(exu_n469), .B(exu_n19774), .Y(exu_n19777));
AND2X1 exu_U8731(.A(exu_n474), .B(exu_n19778), .Y(exu_n19779));
AND2X1 exu_U8732(.A(exu_n473), .B(exu_n19778), .Y(exu_n19780));
AND2X1 exu_U8733(.A(exu_n472), .B(exu_n19778), .Y(exu_n19781));
AND2X1 exu_U8734(.A(exu_n4135), .B(exu_n19806), .Y(exu_n19807));
AND2X1 exu_U8735(.A(exu_n4134), .B(exu_n19806), .Y(exu_n19808));
AND2X1 exu_U8736(.A(exu_n387), .B(exu_n19809), .Y(exu_n19810));
AND2X1 exu_U8737(.A(exu_n386), .B(exu_n19809), .Y(exu_n19811));
AND2X1 exu_U8738(.A(exu_n389), .B(exu_n19812), .Y(exu_n19813));
AND2X1 exu_U8739(.A(exu_n388), .B(exu_n19812), .Y(exu_n19814));
AND2X1 exu_U8740(.A(exu_n391), .B(exu_n19815), .Y(exu_n19816));
AND2X1 exu_U8741(.A(exu_n390), .B(exu_n19815), .Y(exu_n19817));
AND2X1 exu_U8742(.A(exu_n4133), .B(exu_n20295), .Y(exu_n20303));
AND2X1 exu_U8743(.A(exu_n4132), .B(exu_n20295), .Y(exu_n20296));
AND2X1 exu_U8744(.A(exu_n4131), .B(exu_n20295), .Y(exu_n20297));
AND2X1 exu_U8745(.A(exu_n4130), .B(exu_n20295), .Y(exu_n20298));
AND2X1 exu_U8746(.A(exu_n4129), .B(exu_n20295), .Y(exu_n20299));
AND2X1 exu_U8747(.A(exu_n4128), .B(exu_n20295), .Y(exu_n20300));
AND2X1 exu_U8748(.A(exu_n4127), .B(exu_n20295), .Y(exu_n20301));
AND2X1 exu_U8749(.A(exu_n4126), .B(exu_n20295), .Y(exu_n20302));
AND2X1 exu_U8750(.A(exu_n4112), .B(exu_n20304), .Y(exu_n20312));
AND2X1 exu_U8751(.A(exu_n4114), .B(exu_n20304), .Y(exu_n20305));
AND2X1 exu_U8752(.A(exu_n4116), .B(exu_n20304), .Y(exu_n20306));
AND2X1 exu_U8753(.A(exu_n4117), .B(exu_n20304), .Y(exu_n20307));
AND2X1 exu_U8754(.A(exu_n4118), .B(exu_n20304), .Y(exu_n20308));
AND2X1 exu_U8755(.A(exu_n4120), .B(exu_n20304), .Y(exu_n20309));
AND2X1 exu_U8756(.A(exu_n4122), .B(exu_n20304), .Y(exu_n20310));
AND2X1 exu_U8757(.A(exu_n4124), .B(exu_n20304), .Y(exu_n20311));
AND2X1 exu_U8758(.A(exu_n328), .B(exu_n20313), .Y(exu_n20321));
AND2X1 exu_U8759(.A(exu_n330), .B(exu_n20313), .Y(exu_n20314));
AND2X1 exu_U8760(.A(exu_n332), .B(exu_n20313), .Y(exu_n20315));
AND2X1 exu_U8761(.A(exu_n333), .B(exu_n20313), .Y(exu_n20316));
AND2X1 exu_U8762(.A(exu_n334), .B(exu_n20313), .Y(exu_n20317));
AND2X1 exu_U8763(.A(exu_n336), .B(exu_n20313), .Y(exu_n20318));
AND2X1 exu_U8764(.A(exu_n338), .B(exu_n20313), .Y(exu_n20319));
AND2X1 exu_U8765(.A(exu_n340), .B(exu_n20313), .Y(exu_n20320));
AND2X1 exu_U8766(.A(exu_n342), .B(exu_n20322), .Y(exu_n20330));
AND2X1 exu_U8767(.A(exu_n344), .B(exu_n20322), .Y(exu_n20323));
AND2X1 exu_U8768(.A(exu_n346), .B(exu_n20322), .Y(exu_n20324));
AND2X1 exu_U8769(.A(exu_n347), .B(exu_n20322), .Y(exu_n20325));
AND2X1 exu_U8770(.A(exu_n348), .B(exu_n20322), .Y(exu_n20326));
AND2X1 exu_U8771(.A(exu_n350), .B(exu_n20322), .Y(exu_n20327));
AND2X1 exu_U8772(.A(exu_n352), .B(exu_n20322), .Y(exu_n20328));
AND2X1 exu_U8773(.A(exu_n354), .B(exu_n20322), .Y(exu_n20329));
AND2X1 exu_U8774(.A(exu_n356), .B(exu_n20331), .Y(exu_n20339));
AND2X1 exu_U8775(.A(exu_n358), .B(exu_n20331), .Y(exu_n20332));
AND2X1 exu_U8776(.A(exu_n360), .B(exu_n20331), .Y(exu_n20333));
AND2X1 exu_U8777(.A(exu_n361), .B(exu_n20331), .Y(exu_n20334));
AND2X1 exu_U8778(.A(exu_n362), .B(exu_n20331), .Y(exu_n20335));
AND2X1 exu_U8779(.A(exu_n364), .B(exu_n20331), .Y(exu_n20336));
AND2X1 exu_U8780(.A(exu_n366), .B(exu_n20331), .Y(exu_n20337));
AND2X1 exu_U8781(.A(exu_n368), .B(exu_n20331), .Y(exu_n20338));
AND2X1 exu_U8782(.A(exu_n4754), .B(exu_n16030), .Y(exu_n29305));
AND2X1 exu_U8783(.A(exu_n4755), .B(exu_n16030), .Y(exu_n29306));
AND2X1 exu_U8784(.A(exu_n4756), .B(exu_n16030), .Y(exu_n29307));
AND2X1 exu_U8785(.A(exu_n4757), .B(exu_n16030), .Y(exu_n29308));
AND2X1 exu_U8786(.A(exu_n4760), .B(exu_n16030), .Y(exu_n29309));
AND2X1 exu_U8787(.A(exu_n4761), .B(exu_n16030), .Y(exu_n29310));
AND2X1 exu_U8788(.A(exu_n4762), .B(exu_n16030), .Y(exu_n29311));
AND2X1 exu_U8789(.A(exu_n4763), .B(exu_n16030), .Y(exu_n29313));
AND2X1 exu_U8790(.A(exu_n4764), .B(exu_n16029), .Y(exu_n29314));
AND2X1 exu_U8791(.A(exu_n4765), .B(exu_n16029), .Y(exu_n29315));
AND2X1 exu_U8792(.A(exu_n4766), .B(exu_n16029), .Y(exu_n29316));
AND2X1 exu_U8793(.A(exu_n4767), .B(exu_n16029), .Y(exu_n29317));
AND2X1 exu_U8794(.A(exu_n4768), .B(exu_n16029), .Y(exu_n29318));
AND2X1 exu_U8795(.A(exu_n4769), .B(exu_n16029), .Y(exu_n29319));
AND2X1 exu_U8796(.A(exu_n4772), .B(exu_n16029), .Y(exu_n29320));
AND2X1 exu_U8797(.A(exu_n4773), .B(exu_n16029), .Y(exu_n29321));
AND2X1 exu_U8798(.A(exu_n4774), .B(exu_n16029), .Y(exu_n29322));
AND2X1 exu_U8799(.A(exu_n4775), .B(exu_n16029), .Y(exu_n29324));
AND2X1 exu_U8800(.A(exu_n4776), .B(exu_n16029), .Y(exu_n29325));
AND2X1 exu_U8801(.A(exu_n4777), .B(exu_n16029), .Y(exu_n29326));
AND2X1 exu_U8802(.A(exu_n4778), .B(exu_n16028), .Y(exu_n29327));
AND2X1 exu_U8803(.A(exu_n4779), .B(exu_n16028), .Y(exu_n29328));
AND2X1 exu_U8804(.A(exu_n4780), .B(exu_n16028), .Y(exu_n29329));
AND2X1 exu_U8805(.A(exu_n4781), .B(exu_n16028), .Y(exu_n29330));
AND2X1 exu_U8806(.A(exu_n4784), .B(exu_n16028), .Y(exu_n29331));
AND2X1 exu_U8807(.A(exu_n4785), .B(exu_n16028), .Y(exu_n29332));
AND2X1 exu_U8808(.A(exu_n4786), .B(exu_n16028), .Y(exu_n29333));
AND2X1 exu_U8809(.A(exu_n4787), .B(exu_n16028), .Y(exu_n29335));
AND2X1 exu_U8810(.A(exu_n4788), .B(exu_n16028), .Y(exu_n29336));
AND2X1 exu_U8811(.A(exu_n4789), .B(exu_n16028), .Y(exu_n29337));
AND2X1 exu_U8812(.A(exu_n4790), .B(exu_n16028), .Y(exu_n29338));
AND2X1 exu_U8813(.A(exu_n4791), .B(exu_n16028), .Y(exu_n29339));
AND2X1 exu_U8814(.A(exu_n3534), .B(exu_n16037), .Y(exu_n29370));
AND2X1 exu_U8815(.A(exu_n3535), .B(exu_n16037), .Y(exu_n29371));
AND2X1 exu_U8816(.A(exu_n3536), .B(exu_n16037), .Y(exu_n29372));
AND2X1 exu_U8817(.A(exu_n3537), .B(exu_n16037), .Y(exu_n29373));
AND2X1 exu_U8818(.A(exu_n3539), .B(exu_n16037), .Y(exu_n29374));
AND2X1 exu_U8819(.A(exu_n3540), .B(exu_n16037), .Y(exu_n29375));
AND2X1 exu_U8820(.A(exu_n3541), .B(exu_n16037), .Y(exu_n29376));
AND2X1 exu_U8821(.A(exu_n3542), .B(exu_n16037), .Y(exu_n29378));
AND2X1 exu_U8822(.A(exu_n3543), .B(exu_n16036), .Y(exu_n29379));
AND2X1 exu_U8823(.A(exu_n3544), .B(exu_n16036), .Y(exu_n29380));
AND2X1 exu_U8824(.A(exu_n3545), .B(exu_n16036), .Y(exu_n29381));
AND2X1 exu_U8825(.A(exu_n3546), .B(exu_n16036), .Y(exu_n29382));
AND2X1 exu_U8826(.A(exu_n3547), .B(exu_n16036), .Y(exu_n29383));
AND2X1 exu_U8827(.A(exu_n3548), .B(exu_n16036), .Y(exu_n29384));
AND2X1 exu_U8828(.A(exu_n3550), .B(exu_n16036), .Y(exu_n29385));
AND2X1 exu_U8829(.A(exu_n3551), .B(exu_n16036), .Y(exu_n29386));
AND2X1 exu_U8830(.A(exu_n3552), .B(exu_n16036), .Y(exu_n29387));
AND2X1 exu_U8831(.A(exu_n3553), .B(exu_n16036), .Y(exu_n29389));
AND2X1 exu_U8832(.A(exu_n3554), .B(exu_n16036), .Y(exu_n29390));
AND2X1 exu_U8833(.A(exu_n3555), .B(exu_n16036), .Y(exu_n29391));
AND2X1 exu_U8834(.A(exu_n3556), .B(exu_n16035), .Y(exu_n29392));
AND2X1 exu_U8835(.A(exu_n3557), .B(exu_n16035), .Y(exu_n29393));
AND2X1 exu_U8836(.A(exu_n3558), .B(exu_n16035), .Y(exu_n29394));
AND2X1 exu_U8837(.A(exu_n3559), .B(exu_n16035), .Y(exu_n29395));
AND2X1 exu_U8838(.A(exu_n3561), .B(exu_n16035), .Y(exu_n29396));
AND2X1 exu_U8839(.A(exu_n3562), .B(exu_n16035), .Y(exu_n29397));
AND2X1 exu_U8840(.A(exu_n3563), .B(exu_n16035), .Y(exu_n29398));
AND2X1 exu_U8841(.A(exu_n3564), .B(exu_n16035), .Y(exu_n29400));
AND2X1 exu_U8842(.A(exu_n3565), .B(exu_n16035), .Y(exu_n29401));
AND2X1 exu_U8843(.A(exu_n3566), .B(exu_n16035), .Y(exu_n29402));
AND2X1 exu_U8844(.A(exu_n3567), .B(exu_n16035), .Y(exu_n29403));
AND2X1 exu_U8845(.A(exu_n3568), .B(exu_n16035), .Y(exu_n29404));
AND2X1 exu_U8846(.A(exu_n3569), .B(exu_n16034), .Y(exu_n29405));
AND2X1 exu_U8847(.A(exu_n3570), .B(exu_n16034), .Y(exu_n29406));
AND2X1 exu_U8848(.A(exu_n3572), .B(exu_n16034), .Y(exu_n29407));
AND2X1 exu_U8849(.A(exu_n3573), .B(exu_n16034), .Y(exu_n29408));
AND2X1 exu_U8850(.A(exu_n3574), .B(exu_n16034), .Y(exu_n29409));
AND2X1 exu_U8851(.A(exu_n3575), .B(exu_n16034), .Y(exu_n29411));
AND2X1 exu_U8852(.A(exu_n3576), .B(exu_n16034), .Y(exu_n29412));
AND2X1 exu_U8853(.A(exu_n3577), .B(exu_n16034), .Y(exu_n29413));
AND2X1 exu_U8854(.A(exu_n3578), .B(exu_n16034), .Y(exu_n29414));
AND2X1 exu_U8855(.A(exu_n3579), .B(exu_n16034), .Y(exu_n29415));
AND2X1 exu_U8856(.A(exu_n3580), .B(exu_n16034), .Y(exu_n29416));
AND2X1 exu_U8857(.A(exu_n3581), .B(exu_n16034), .Y(exu_n29417));
AND2X1 exu_U8858(.A(exu_n3583), .B(exu_n16033), .Y(exu_n29418));
AND2X1 exu_U8859(.A(exu_n3584), .B(exu_n16033), .Y(exu_n29419));
AND2X1 exu_U8860(.A(exu_n3585), .B(exu_n16033), .Y(exu_n29420));
AND2X1 exu_U8861(.A(exu_n3586), .B(exu_n16033), .Y(exu_n29421));
AND2X1 exu_U8862(.A(exu_n3587), .B(exu_n16033), .Y(exu_n29422));
AND2X1 exu_U8863(.A(exu_n3588), .B(exu_n16033), .Y(exu_n29423));
AND2X1 exu_U8864(.A(exu_n3589), .B(exu_n16033), .Y(exu_n29424));
AND2X1 exu_U8865(.A(exu_n3590), .B(exu_n16033), .Y(exu_n29425));
AND2X1 exu_U8866(.A(exu_n3591), .B(exu_n16033), .Y(exu_n29426));
AND2X1 exu_U8867(.A(exu_n3592), .B(exu_n16033), .Y(exu_n29427));
AND2X1 exu_U8868(.A(exu_n3530), .B(exu_n16033), .Y(exu_n29428));
AND2X1 exu_U8869(.A(exu_n3531), .B(exu_n16033), .Y(exu_n29429));
AND2X1 exu_U8870(.A(exu_n3532), .B(exu_n16033), .Y(exu_n29430));
AND2X1 exu_U8871(.A(exu_n3533), .B(exu_n16037), .Y(exu_n29367));
AND2X1 exu_U8872(.A(exu_n3538), .B(exu_n16037), .Y(exu_n29368));
AND2X1 exu_U8873(.A(exu_n3549), .B(exu_n16037), .Y(exu_n29369));
AND2X1 exu_U8874(.A(exu_n3560), .B(exu_n16037), .Y(exu_n29377));
AND2X1 exu_U8875(.A(exu_n3571), .B(exu_n16036), .Y(exu_n29388));
AND2X1 exu_U8876(.A(exu_n3582), .B(exu_n16035), .Y(exu_n29399));
AND2X1 exu_U8877(.A(exu_n3593), .B(exu_n16034), .Y(exu_n29410));
AND2X1 exu_U8878(.A(exu_n3903), .B(exu_n16114), .Y(exu_n30084));
AND2X1 exu_U8879(.A(exu_n3904), .B(exu_n16114), .Y(exu_n30085));
AND2X1 exu_U8880(.A(exu_n3905), .B(exu_n16114), .Y(exu_n30086));
AND2X1 exu_U8881(.A(exu_n3906), .B(exu_n16114), .Y(exu_n30087));
AND2X1 exu_U8882(.A(exu_n3908), .B(exu_n16114), .Y(exu_n30088));
AND2X1 exu_U8883(.A(exu_n3909), .B(exu_n16114), .Y(exu_n30089));
AND2X1 exu_U8884(.A(exu_n3910), .B(exu_n16114), .Y(exu_n30090));
AND2X1 exu_U8885(.A(exu_n3911), .B(exu_n16114), .Y(exu_n30092));
AND2X1 exu_U8886(.A(exu_n3912), .B(exu_n16113), .Y(exu_n30093));
AND2X1 exu_U8887(.A(exu_n3913), .B(exu_n16113), .Y(exu_n30094));
AND2X1 exu_U8888(.A(exu_n3914), .B(exu_n16113), .Y(exu_n30095));
AND2X1 exu_U8889(.A(exu_n3915), .B(exu_n16113), .Y(exu_n30096));
AND2X1 exu_U8890(.A(exu_n3916), .B(exu_n16113), .Y(exu_n30097));
AND2X1 exu_U8891(.A(exu_n3917), .B(exu_n16113), .Y(exu_n30098));
AND2X1 exu_U8892(.A(exu_n3919), .B(exu_n16113), .Y(exu_n30099));
AND2X1 exu_U8893(.A(exu_n3920), .B(exu_n16113), .Y(exu_n30100));
AND2X1 exu_U8894(.A(exu_n3921), .B(exu_n16113), .Y(exu_n30101));
AND2X1 exu_U8895(.A(exu_n3922), .B(exu_n16113), .Y(exu_n30103));
AND2X1 exu_U8896(.A(exu_n3923), .B(exu_n16113), .Y(exu_n30104));
AND2X1 exu_U8897(.A(exu_n3924), .B(exu_n16113), .Y(exu_n30105));
AND2X1 exu_U8898(.A(exu_n3925), .B(exu_n16112), .Y(exu_n30106));
AND2X1 exu_U8899(.A(exu_n3926), .B(exu_n16112), .Y(exu_n30107));
AND2X1 exu_U8900(.A(exu_n3927), .B(exu_n16112), .Y(exu_n30108));
AND2X1 exu_U8901(.A(exu_n3928), .B(exu_n16112), .Y(exu_n30109));
AND2X1 exu_U8902(.A(exu_n3930), .B(exu_n16112), .Y(exu_n30110));
AND2X1 exu_U8903(.A(exu_n3931), .B(exu_n16112), .Y(exu_n30111));
AND2X1 exu_U8904(.A(exu_n3932), .B(exu_n16112), .Y(exu_n30112));
AND2X1 exu_U8905(.A(exu_n3933), .B(exu_n16112), .Y(exu_n30114));
AND2X1 exu_U8906(.A(exu_n3934), .B(exu_n16112), .Y(exu_n30115));
AND2X1 exu_U8907(.A(exu_n3935), .B(exu_n16112), .Y(exu_n30116));
AND2X1 exu_U8908(.A(exu_n3936), .B(exu_n16112), .Y(exu_n30117));
AND2X1 exu_U8909(.A(exu_n3937), .B(exu_n16112), .Y(exu_n30118));
AND2X1 exu_U8910(.A(exu_n3938), .B(exu_n16111), .Y(exu_n30119));
AND2X1 exu_U8911(.A(exu_n3939), .B(exu_n16111), .Y(exu_n30120));
AND2X1 exu_U8912(.A(exu_n3941), .B(exu_n16111), .Y(exu_n30121));
AND2X1 exu_U8913(.A(exu_n3942), .B(exu_n16111), .Y(exu_n30122));
AND2X1 exu_U8914(.A(exu_n3943), .B(exu_n16111), .Y(exu_n30123));
AND2X1 exu_U8915(.A(exu_n3944), .B(exu_n16111), .Y(exu_n30125));
AND2X1 exu_U8916(.A(exu_n3945), .B(exu_n16111), .Y(exu_n30126));
AND2X1 exu_U8917(.A(exu_n3946), .B(exu_n16111), .Y(exu_n30127));
AND2X1 exu_U8918(.A(exu_n3947), .B(exu_n16111), .Y(exu_n30128));
AND2X1 exu_U8919(.A(exu_n3948), .B(exu_n16111), .Y(exu_n30129));
AND2X1 exu_U8920(.A(exu_n3949), .B(exu_n16111), .Y(exu_n30130));
AND2X1 exu_U8921(.A(exu_n3950), .B(exu_n16111), .Y(exu_n30131));
AND2X1 exu_U8922(.A(exu_n3952), .B(exu_n16110), .Y(exu_n30132));
AND2X1 exu_U8923(.A(exu_n3953), .B(exu_n16110), .Y(exu_n30133));
AND2X1 exu_U8924(.A(exu_n3954), .B(exu_n16110), .Y(exu_n30134));
AND2X1 exu_U8925(.A(exu_n3955), .B(exu_n16110), .Y(exu_n30135));
AND2X1 exu_U8926(.A(exu_n3956), .B(exu_n16110), .Y(exu_n30136));
AND2X1 exu_U8927(.A(exu_n3957), .B(exu_n16110), .Y(exu_n30137));
AND2X1 exu_U8928(.A(exu_n3958), .B(exu_n16110), .Y(exu_n30138));
AND2X1 exu_U8929(.A(exu_n3959), .B(exu_n16110), .Y(exu_n30139));
AND2X1 exu_U8930(.A(exu_n3960), .B(exu_n16110), .Y(exu_n30140));
AND2X1 exu_U8931(.A(exu_n3961), .B(exu_n16110), .Y(exu_n30141));
AND2X1 exu_U8932(.A(exu_n3899), .B(exu_n16110), .Y(exu_n30142));
AND2X1 exu_U8933(.A(exu_n3900), .B(exu_n16110), .Y(exu_n30143));
AND2X1 exu_U8934(.A(exu_n3901), .B(exu_n16110), .Y(exu_n30144));
AND2X1 exu_U8935(.A(exu_n3902), .B(exu_n16114), .Y(exu_n30081));
AND2X1 exu_U8936(.A(exu_n3907), .B(exu_n16114), .Y(exu_n30082));
AND2X1 exu_U8937(.A(exu_n3918), .B(exu_n16114), .Y(exu_n30083));
AND2X1 exu_U8938(.A(exu_n3929), .B(exu_n16114), .Y(exu_n30091));
AND2X1 exu_U8939(.A(exu_n3940), .B(exu_n16113), .Y(exu_n30102));
AND2X1 exu_U8940(.A(exu_n3951), .B(exu_n16112), .Y(exu_n30113));
AND2X1 exu_U8941(.A(exu_n3962), .B(exu_n16111), .Y(exu_n30124));
AND2X1 exu_U8942(.A(exu_n4049), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n7));
AND2X1 exu_U8943(.A(exu_n4050), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n9));
AND2X1 exu_U8944(.A(exu_n4051), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n11));
AND2X1 exu_U8945(.A(exu_n4035), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n13));
AND2X1 exu_U8946(.A(exu_n4036), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n15));
AND2X1 exu_U8947(.A(exu_n4037), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n17));
AND2X1 exu_U8948(.A(exu_n4038), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n19));
AND2X1 exu_U8949(.A(exu_n4039), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n21));
AND2X1 exu_U8950(.A(exu_n4041), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n23));
AND2X1 exu_U8951(.A(exu_n4043), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n25));
AND2X1 exu_U8952(.A(exu_n4045), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n27));
AND2X1 exu_U8953(.A(exu_n4047), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n29));
AND2X1 exu_U8954(.A(exu_n4052), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n31));
AND2X1 exu_U8955(.A(exu_n4490), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n17));
AND2X1 exu_U8956(.A(exu_n4491), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n19));
AND2X1 exu_U8957(.A(exu_n4492), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n21));
AND2X1 exu_U8958(.A(exu_n4493), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n3));
AND2X1 exu_U8959(.A(exu_n4494), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n5));
AND2X1 exu_U8960(.A(exu_n4495), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n7));
AND2X1 exu_U8961(.A(exu_n4496), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n9));
AND2X1 exu_U8962(.A(exu_n4497), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n11));
AND2X1 exu_U8963(.A(exu_n4498), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n13));
AND2X1 exu_U8964(.A(exu_n4499), .B(ecl_mdqctl_mul_data_dff_n1), .Y(ecl_mdqctl_mul_data_dff_n15));
AND2X1 exu_U8965(.A(exu_n4065), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n2));
AND2X1 exu_U8966(.A(exu_n4064), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n5));
AND2X1 exu_U8967(.A(exu_n4062), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n9));
AND2X1 exu_U8968(.A(exu_n4061), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n11));
AND2X1 exu_U8969(.A(exu_n4060), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n13));
AND2X1 exu_U8970(.A(exu_n4059), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n15));
AND2X1 exu_U8971(.A(exu_n4058), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n17));
AND2X1 exu_U8972(.A(exu_n4057), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n19));
AND2X1 exu_U8973(.A(exu_n4056), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n21));
AND2X1 exu_U8974(.A(exu_n4055), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n23));
AND2X1 exu_U8975(.A(exu_n4054), .B(exu_n15947), .Y(ecl_mdqctl_div_data_dff_n25));
AND2X1 exu_U8976(.A(exu_n4502), .B(ecl_divcntl_divstate_dff_n1), .Y(ecl_divcntl_divstate_dff_n7));
AND2X1 exu_U8977(.A(exu_n4503), .B(ecl_divcntl_divstate_dff_n1), .Y(ecl_divcntl_divstate_dff_n9));
AND2X1 exu_U8978(.A(exu_n4504), .B(ecl_divcntl_divstate_dff_n1), .Y(ecl_divcntl_divstate_dff_n13));
AND2X1 exu_U8979(.A(exu_n15688), .B(ecl_writeback_valid_m), .Y(ecl_writeback_dff_wb_m2w_n2));
AND2X1 exu_U8980(.A(exu_n4891), .B(rml_oddwin_dff_n1), .Y(rml_oddwin_dff_n3));
AND2X1 exu_U8981(.A(exu_n4892), .B(rml_oddwin_dff_n1), .Y(rml_oddwin_dff_n5));
AND2X1 exu_U8982(.A(exu_n4893), .B(rml_oddwin_dff_n1), .Y(rml_oddwin_dff_n7));
AND2X1 exu_U8983(.A(exu_n4894), .B(rml_oddwin_dff_n1), .Y(rml_oddwin_dff_n9));
AND2X1 exu_U8984(.A(exu_n4353), .B(exu_n16119), .Y(div_d_dff_n189));
AND2X1 exu_U8985(.A(exu_n4355), .B(exu_n16119), .Y(div_d_dff_n193));
AND2X1 exu_U8986(.A(exu_n4357), .B(exu_n16119), .Y(div_d_dff_n195));
AND2X1 exu_U8987(.A(exu_n4359), .B(exu_n16119), .Y(div_d_dff_n197));
AND2X1 exu_U8988(.A(exu_n4361), .B(exu_n16119), .Y(div_d_dff_n199));
AND2X1 exu_U8989(.A(exu_n4363), .B(exu_n16119), .Y(div_d_dff_n201));
AND2X1 exu_U8990(.A(exu_n4365), .B(exu_n16119), .Y(div_d_dff_n203));
AND2X1 exu_U8991(.A(exu_n4367), .B(exu_n16119), .Y(div_d_dff_n205));
AND2X1 exu_U8992(.A(exu_n4371), .B(exu_n16118), .Y(div_d_dff_n207));
AND2X1 exu_U8993(.A(exu_n4373), .B(exu_n16118), .Y(div_d_dff_n209));
AND2X1 exu_U8994(.A(exu_n4375), .B(exu_n16118), .Y(div_d_dff_n211));
AND2X1 exu_U8995(.A(exu_n4377), .B(exu_n16118), .Y(div_d_dff_n215));
AND2X1 exu_U8996(.A(exu_n4379), .B(exu_n16118), .Y(div_d_dff_n217));
AND2X1 exu_U8997(.A(exu_n4381), .B(exu_n16118), .Y(div_d_dff_n219));
AND2X1 exu_U8998(.A(exu_n4383), .B(exu_n16118), .Y(div_d_dff_n221));
AND2X1 exu_U8999(.A(exu_n4385), .B(exu_n16118), .Y(div_d_dff_n223));
AND2X1 exu_U9000(.A(exu_n4387), .B(exu_n16118), .Y(div_d_dff_n225));
AND2X1 exu_U9001(.A(exu_n4389), .B(exu_n16118), .Y(div_d_dff_n227));
AND2X1 exu_U9002(.A(exu_n4393), .B(exu_n16118), .Y(div_d_dff_n229));
AND2X1 exu_U9003(.A(exu_n4395), .B(exu_n16118), .Y(div_d_dff_n231));
AND2X1 exu_U9004(.A(exu_n4397), .B(exu_n16117), .Y(div_d_dff_n233));
AND2X1 exu_U9005(.A(exu_n4399), .B(exu_n16117), .Y(div_d_dff_n237));
AND2X1 exu_U9006(.A(exu_n4401), .B(exu_n16117), .Y(div_d_dff_n239));
AND2X1 exu_U9007(.A(exu_n4403), .B(exu_n16117), .Y(div_d_dff_n241));
AND2X1 exu_U9008(.A(exu_n4405), .B(exu_n16117), .Y(div_d_dff_n243));
AND2X1 exu_U9009(.A(exu_n4407), .B(exu_n16117), .Y(div_d_dff_n245));
AND2X1 exu_U9010(.A(exu_n4409), .B(exu_n16117), .Y(div_d_dff_n247));
AND2X1 exu_U9011(.A(exu_n4411), .B(exu_n16117), .Y(div_d_dff_n249));
AND2X1 exu_U9012(.A(exu_n4161), .B(exu_n16117), .Y(div_d_dff_n251));
AND2X1 exu_U9013(.A(exu_n4163), .B(exu_n16117), .Y(div_d_dff_n253));
AND2X1 exu_U9014(.A(exu_n4165), .B(exu_n16117), .Y(div_d_dff_n255));
AND2X1 exu_U9015(.A(exu_n4167), .B(exu_n16126), .Y(div_d_dff_n3));
AND2X1 exu_U9016(.A(exu_n4169), .B(exu_n16126), .Y(div_d_dff_n5));
AND2X1 exu_U9017(.A(exu_n4171), .B(exu_n16126), .Y(div_d_dff_n7));
AND2X1 exu_U9018(.A(exu_n4173), .B(exu_n16126), .Y(div_d_dff_n9));
AND2X1 exu_U9019(.A(exu_n4175), .B(exu_n16126), .Y(div_d_dff_n11));
AND2X1 exu_U9020(.A(exu_n4177), .B(exu_n16126), .Y(div_d_dff_n13));
AND2X1 exu_U9021(.A(exu_n4179), .B(exu_n16126), .Y(div_d_dff_n15));
AND2X1 exu_U9022(.A(exu_n4183), .B(exu_n16126), .Y(div_d_dff_n17));
AND2X1 exu_U9023(.A(exu_n4185), .B(exu_n16126), .Y(div_d_dff_n19));
AND2X1 exu_U9024(.A(exu_n4187), .B(exu_n16126), .Y(div_d_dff_n21));
AND2X1 exu_U9025(.A(exu_n4189), .B(exu_n16125), .Y(div_d_dff_n25));
AND2X1 exu_U9026(.A(exu_n4191), .B(exu_n16125), .Y(div_d_dff_n27));
AND2X1 exu_U9027(.A(exu_n4193), .B(exu_n16125), .Y(div_d_dff_n29));
AND2X1 exu_U9028(.A(exu_n4195), .B(exu_n16125), .Y(div_d_dff_n31));
AND2X1 exu_U9029(.A(exu_n4197), .B(exu_n16125), .Y(div_d_dff_n33));
AND2X1 exu_U9030(.A(exu_n4199), .B(exu_n16125), .Y(div_d_dff_n35));
AND2X1 exu_U9031(.A(exu_n4201), .B(exu_n16125), .Y(div_d_dff_n37));
AND2X1 exu_U9032(.A(exu_n4205), .B(exu_n16125), .Y(div_d_dff_n39));
AND2X1 exu_U9033(.A(exu_n4207), .B(exu_n16125), .Y(div_d_dff_n41));
AND2X1 exu_U9034(.A(exu_n4209), .B(exu_n16125), .Y(div_d_dff_n43));
AND2X1 exu_U9035(.A(exu_n4211), .B(exu_n16125), .Y(div_d_dff_n47));
AND2X1 exu_U9036(.A(exu_n4213), .B(exu_n16125), .Y(div_d_dff_n49));
AND2X1 exu_U9037(.A(exu_n4215), .B(exu_n16124), .Y(div_d_dff_n51));
AND2X1 exu_U9038(.A(exu_n4217), .B(exu_n16124), .Y(div_d_dff_n53));
AND2X1 exu_U9039(.A(exu_n4219), .B(exu_n16124), .Y(div_d_dff_n55));
AND2X1 exu_U9040(.A(exu_n4221), .B(exu_n16124), .Y(div_d_dff_n57));
AND2X1 exu_U9041(.A(exu_n4223), .B(exu_n16124), .Y(div_d_dff_n59));
AND2X1 exu_U9042(.A(exu_n4227), .B(exu_n16124), .Y(div_d_dff_n61));
AND2X1 exu_U9043(.A(exu_n4229), .B(exu_n16124), .Y(div_d_dff_n63));
AND2X1 exu_U9044(.A(exu_n4231), .B(exu_n16124), .Y(div_d_dff_n65));
AND2X1 exu_U9045(.A(exu_n4233), .B(exu_n16124), .Y(div_d_dff_n69));
AND2X1 exu_U9046(.A(exu_n4235), .B(exu_n16124), .Y(div_d_dff_n71));
AND2X1 exu_U9047(.A(exu_n4237), .B(exu_n16124), .Y(div_d_dff_n73));
AND2X1 exu_U9048(.A(exu_n4239), .B(exu_n16124), .Y(div_d_dff_n75));
AND2X1 exu_U9049(.A(exu_n4241), .B(exu_n16123), .Y(div_d_dff_n77));
AND2X1 exu_U9050(.A(exu_n4243), .B(exu_n16123), .Y(div_d_dff_n79));
AND2X1 exu_U9051(.A(exu_n4245), .B(exu_n16123), .Y(div_d_dff_n81));
AND2X1 exu_U9052(.A(exu_n4249), .B(exu_n16123), .Y(div_d_dff_n83));
AND2X1 exu_U9053(.A(exu_n4251), .B(exu_n16123), .Y(div_d_dff_n85));
AND2X1 exu_U9054(.A(exu_n4253), .B(exu_n16123), .Y(div_d_dff_n87));
AND2X1 exu_U9055(.A(exu_n4255), .B(exu_n16123), .Y(div_d_dff_n91));
AND2X1 exu_U9056(.A(exu_n4257), .B(exu_n16123), .Y(div_d_dff_n93));
AND2X1 exu_U9057(.A(exu_n4259), .B(exu_n16123), .Y(div_d_dff_n95));
AND2X1 exu_U9058(.A(exu_n4261), .B(exu_n16123), .Y(div_d_dff_n97));
AND2X1 exu_U9059(.A(exu_n4263), .B(exu_n16123), .Y(div_d_dff_n99));
AND2X1 exu_U9060(.A(exu_n4265), .B(exu_n16123), .Y(div_d_dff_n101));
AND2X1 exu_U9061(.A(exu_n4267), .B(exu_n16122), .Y(div_d_dff_n103));
AND2X1 exu_U9062(.A(exu_n4271), .B(exu_n16122), .Y(div_d_dff_n105));
AND2X1 exu_U9063(.A(exu_n4273), .B(exu_n16122), .Y(div_d_dff_n107));
AND2X1 exu_U9064(.A(exu_n4275), .B(exu_n16122), .Y(div_d_dff_n109));
AND2X1 exu_U9065(.A(exu_n4277), .B(exu_n16122), .Y(div_d_dff_n113));
AND2X1 exu_U9066(.A(exu_n4279), .B(exu_n16122), .Y(div_d_dff_n115));
AND2X1 exu_U9067(.A(exu_n4281), .B(exu_n16122), .Y(div_d_dff_n117));
AND2X1 exu_U9068(.A(exu_n4283), .B(exu_n16122), .Y(div_d_dff_n119));
AND2X1 exu_U9069(.A(exu_n4285), .B(exu_n16122), .Y(div_d_dff_n121));
AND2X1 exu_U9070(.A(exu_n4287), .B(exu_n16122), .Y(div_d_dff_n123));
AND2X1 exu_U9071(.A(exu_n4289), .B(exu_n16122), .Y(div_d_dff_n125));
AND2X1 exu_U9072(.A(exu_n4293), .B(exu_n16122), .Y(div_d_dff_n127));
AND2X1 exu_U9073(.A(exu_n4295), .B(exu_n16121), .Y(div_d_dff_n129));
AND2X1 exu_U9074(.A(exu_n4297), .B(exu_n16121), .Y(div_d_dff_n131));
AND2X1 exu_U9075(.A(exu_n4299), .B(exu_n16121), .Y(div_d_dff_n135));
AND2X1 exu_U9076(.A(exu_n4301), .B(exu_n16121), .Y(div_d_dff_n137));
AND2X1 exu_U9077(.A(exu_n4303), .B(exu_n16121), .Y(div_d_dff_n139));
AND2X1 exu_U9078(.A(exu_n4305), .B(exu_n16121), .Y(div_d_dff_n141));
AND2X1 exu_U9079(.A(exu_n4307), .B(exu_n16121), .Y(div_d_dff_n143));
AND2X1 exu_U9080(.A(exu_n4309), .B(exu_n16121), .Y(div_d_dff_n145));
AND2X1 exu_U9081(.A(exu_n4311), .B(exu_n16121), .Y(div_d_dff_n147));
AND2X1 exu_U9082(.A(exu_n4315), .B(exu_n16121), .Y(div_d_dff_n149));
AND2X1 exu_U9083(.A(exu_n4317), .B(exu_n16121), .Y(div_d_dff_n151));
AND2X1 exu_U9084(.A(exu_n4319), .B(exu_n16121), .Y(div_d_dff_n153));
AND2X1 exu_U9085(.A(exu_n4321), .B(exu_n16120), .Y(div_d_dff_n157));
AND2X1 exu_U9086(.A(exu_n4323), .B(exu_n16120), .Y(div_d_dff_n159));
AND2X1 exu_U9087(.A(exu_n4325), .B(exu_n16120), .Y(div_d_dff_n161));
AND2X1 exu_U9088(.A(exu_n4327), .B(exu_n16120), .Y(div_d_dff_n163));
AND2X1 exu_U9089(.A(exu_n4329), .B(exu_n16120), .Y(div_d_dff_n165));
AND2X1 exu_U9090(.A(exu_n4331), .B(exu_n16120), .Y(div_d_dff_n167));
AND2X1 exu_U9091(.A(exu_n4333), .B(exu_n16120), .Y(div_d_dff_n169));
AND2X1 exu_U9092(.A(exu_n4337), .B(exu_n16120), .Y(div_d_dff_n171));
AND2X1 exu_U9093(.A(exu_n4339), .B(exu_n16120), .Y(div_d_dff_n173));
AND2X1 exu_U9094(.A(exu_n4341), .B(exu_n16120), .Y(div_d_dff_n175));
AND2X1 exu_U9095(.A(exu_n4343), .B(exu_n16120), .Y(div_d_dff_n177));
AND2X1 exu_U9096(.A(exu_n4345), .B(exu_n16120), .Y(div_d_dff_n179));
AND2X1 exu_U9097(.A(exu_n4347), .B(exu_n16119), .Y(div_d_dff_n181));
AND2X1 exu_U9098(.A(exu_n4349), .B(exu_n16119), .Y(div_d_dff_n183));
AND2X1 exu_U9099(.A(exu_n4351), .B(exu_n16119), .Y(div_d_dff_n185));
AND2X1 exu_U9100(.A(exu_n4369), .B(exu_n16119), .Y(div_d_dff_n187));
AND2X1 exu_U9101(.A(exu_n4391), .B(exu_n16119), .Y(div_d_dff_n191));
AND2X1 exu_U9102(.A(exu_n4159), .B(exu_n16118), .Y(div_d_dff_n213));
AND2X1 exu_U9103(.A(exu_n4181), .B(exu_n16117), .Y(div_d_dff_n235));
AND2X1 exu_U9104(.A(exu_n4203), .B(exu_n16117), .Y(div_d_dff_n257));
AND2X1 exu_U9105(.A(exu_n4225), .B(exu_n16126), .Y(div_d_dff_n23));
AND2X1 exu_U9106(.A(exu_n4247), .B(exu_n16125), .Y(div_d_dff_n45));
AND2X1 exu_U9107(.A(exu_n4269), .B(exu_n16124), .Y(div_d_dff_n67));
AND2X1 exu_U9108(.A(exu_n4291), .B(exu_n16123), .Y(div_d_dff_n89));
AND2X1 exu_U9109(.A(exu_n4313), .B(exu_n16122), .Y(div_d_dff_n111));
AND2X1 exu_U9110(.A(exu_n4335), .B(exu_n16121), .Y(div_d_dff_n133));
AND2X1 exu_U9111(.A(exu_n4413), .B(exu_n16120), .Y(div_d_dff_n155));
AND2X1 exu_U9112(.A(exu_n4569), .B(ecl_ttype_e2m_n1), .Y(ecl_ttype_e2m_n5));
AND2X1 exu_U9113(.A(exu_n4571), .B(ecl_ttype_e2m_n1), .Y(ecl_ttype_e2m_n7));
AND2X1 exu_U9114(.A(exu_n4574), .B(ecl_ttype_e2m_n1), .Y(ecl_ttype_e2m_n11));
AND2X1 exu_U9115(.A(exu_n4950), .B(exu_n15688), .Y(ecl_perr_dff_n2));
AND2X1 exu_U9116(.A(exu_n4951), .B(exu_n15688), .Y(ecl_perr_dff_n5));
AND2X1 exu_U9117(.A(exu_n4952), .B(exu_n15688), .Y(ecl_perr_dff_n7));
AND2X1 exu_U9118(.A(exu_n4953), .B(exu_n15688), .Y(ecl_perr_dff_n9));
AND2X1 exu_U9119(.A(exu_n4824), .B(exu_n16139), .Y(bypass_dfill_data_dff_n9));
AND2X1 exu_U9120(.A(exu_n4825), .B(exu_n16139), .Y(bypass_dfill_data_dff_n11));
AND2X1 exu_U9121(.A(exu_n4826), .B(exu_n16139), .Y(bypass_dfill_data_dff_n13));
AND2X1 exu_U9122(.A(exu_n4827), .B(exu_n16139), .Y(bypass_dfill_data_dff_n15));
AND2X1 exu_U9123(.A(exu_n4829), .B(exu_n16139), .Y(bypass_dfill_data_dff_n17));
AND2X1 exu_U9124(.A(exu_n4830), .B(exu_n16139), .Y(bypass_dfill_data_dff_n19));
AND2X1 exu_U9125(.A(exu_n4831), .B(exu_n16139), .Y(bypass_dfill_data_dff_n21));
AND2X1 exu_U9126(.A(exu_n4832), .B(exu_n16139), .Y(bypass_dfill_data_dff_n25));
AND2X1 exu_U9127(.A(exu_n4833), .B(exu_n16138), .Y(bypass_dfill_data_dff_n27));
AND2X1 exu_U9128(.A(exu_n4834), .B(exu_n16138), .Y(bypass_dfill_data_dff_n29));
AND2X1 exu_U9129(.A(exu_n4835), .B(exu_n16138), .Y(bypass_dfill_data_dff_n31));
AND2X1 exu_U9130(.A(exu_n4836), .B(exu_n16138), .Y(bypass_dfill_data_dff_n33));
AND2X1 exu_U9131(.A(exu_n4837), .B(exu_n16138), .Y(bypass_dfill_data_dff_n35));
AND2X1 exu_U9132(.A(exu_n4838), .B(exu_n16138), .Y(bypass_dfill_data_dff_n37));
AND2X1 exu_U9133(.A(exu_n4840), .B(exu_n16138), .Y(bypass_dfill_data_dff_n39));
AND2X1 exu_U9134(.A(exu_n4841), .B(exu_n16138), .Y(bypass_dfill_data_dff_n41));
AND2X1 exu_U9135(.A(exu_n4842), .B(exu_n16138), .Y(bypass_dfill_data_dff_n43));
AND2X1 exu_U9136(.A(exu_n4843), .B(exu_n16138), .Y(bypass_dfill_data_dff_n47));
AND2X1 exu_U9137(.A(exu_n4844), .B(exu_n16138), .Y(bypass_dfill_data_dff_n49));
AND2X1 exu_U9138(.A(exu_n4845), .B(exu_n16138), .Y(bypass_dfill_data_dff_n51));
AND2X1 exu_U9139(.A(exu_n4846), .B(exu_n16137), .Y(bypass_dfill_data_dff_n53));
AND2X1 exu_U9140(.A(exu_n4847), .B(exu_n16137), .Y(bypass_dfill_data_dff_n55));
AND2X1 exu_U9141(.A(exu_n4848), .B(exu_n16137), .Y(bypass_dfill_data_dff_n57));
AND2X1 exu_U9142(.A(exu_n4849), .B(exu_n16137), .Y(bypass_dfill_data_dff_n59));
AND2X1 exu_U9143(.A(exu_n4851), .B(exu_n16137), .Y(bypass_dfill_data_dff_n61));
AND2X1 exu_U9144(.A(exu_n4852), .B(exu_n16137), .Y(bypass_dfill_data_dff_n63));
AND2X1 exu_U9145(.A(exu_n4853), .B(exu_n16137), .Y(bypass_dfill_data_dff_n65));
AND2X1 exu_U9146(.A(exu_n4854), .B(exu_n16137), .Y(bypass_dfill_data_dff_n69));
AND2X1 exu_U9147(.A(exu_n4855), .B(exu_n16137), .Y(bypass_dfill_data_dff_n71));
AND2X1 exu_U9148(.A(exu_n4856), .B(exu_n16137), .Y(bypass_dfill_data_dff_n73));
AND2X1 exu_U9149(.A(exu_n4857), .B(exu_n16137), .Y(bypass_dfill_data_dff_n75));
AND2X1 exu_U9150(.A(exu_n4858), .B(exu_n16137), .Y(bypass_dfill_data_dff_n77));
AND2X1 exu_U9151(.A(exu_n4859), .B(exu_n16136), .Y(bypass_dfill_data_dff_n79));
AND2X1 exu_U9152(.A(exu_n4860), .B(exu_n16136), .Y(bypass_dfill_data_dff_n81));
AND2X1 exu_U9153(.A(exu_n4862), .B(exu_n16136), .Y(bypass_dfill_data_dff_n83));
AND2X1 exu_U9154(.A(exu_n4863), .B(exu_n16136), .Y(bypass_dfill_data_dff_n85));
AND2X1 exu_U9155(.A(exu_n4864), .B(exu_n16136), .Y(bypass_dfill_data_dff_n87));
AND2X1 exu_U9156(.A(exu_n4865), .B(exu_n16136), .Y(bypass_dfill_data_dff_n91));
AND2X1 exu_U9157(.A(exu_n4866), .B(exu_n16136), .Y(bypass_dfill_data_dff_n93));
AND2X1 exu_U9158(.A(exu_n4867), .B(exu_n16136), .Y(bypass_dfill_data_dff_n95));
AND2X1 exu_U9159(.A(exu_n4868), .B(exu_n16136), .Y(bypass_dfill_data_dff_n97));
AND2X1 exu_U9160(.A(exu_n4869), .B(exu_n16136), .Y(bypass_dfill_data_dff_n99));
AND2X1 exu_U9161(.A(exu_n4870), .B(exu_n16136), .Y(bypass_dfill_data_dff_n101));
AND2X1 exu_U9162(.A(exu_n4871), .B(exu_n16136), .Y(bypass_dfill_data_dff_n103));
AND2X1 exu_U9163(.A(exu_n4873), .B(exu_n16135), .Y(bypass_dfill_data_dff_n105));
AND2X1 exu_U9164(.A(exu_n4874), .B(exu_n16135), .Y(bypass_dfill_data_dff_n107));
AND2X1 exu_U9165(.A(exu_n4875), .B(exu_n16135), .Y(bypass_dfill_data_dff_n109));
AND2X1 exu_U9166(.A(exu_n4876), .B(exu_n16135), .Y(bypass_dfill_data_dff_n111));
AND2X1 exu_U9167(.A(exu_n4877), .B(exu_n16135), .Y(bypass_dfill_data_dff_n113));
AND2X1 exu_U9168(.A(exu_n4878), .B(exu_n16135), .Y(bypass_dfill_data_dff_n115));
AND2X1 exu_U9169(.A(exu_n4879), .B(exu_n16135), .Y(bypass_dfill_data_dff_n117));
AND2X1 exu_U9170(.A(exu_n4880), .B(exu_n16135), .Y(bypass_dfill_data_dff_n119));
AND2X1 exu_U9171(.A(exu_n4881), .B(exu_n16135), .Y(bypass_dfill_data_dff_n121));
AND2X1 exu_U9172(.A(exu_n4882), .B(exu_n16135), .Y(bypass_dfill_data_dff_n123));
AND2X1 exu_U9173(.A(exu_n4820), .B(exu_n16135), .Y(bypass_dfill_data_dff_n125));
AND2X1 exu_U9174(.A(exu_n4821), .B(exu_n16135), .Y(bypass_dfill_data_dff_n127));
AND2X1 exu_U9175(.A(exu_n4822), .B(exu_n16135), .Y(bypass_dfill_data_dff_n129));
AND2X1 exu_U9176(.A(exu_n4823), .B(exu_n16139), .Y(bypass_dfill_data_dff_n3));
AND2X1 exu_U9177(.A(exu_n4828), .B(exu_n16139), .Y(bypass_dfill_data_dff_n5));
AND2X1 exu_U9178(.A(exu_n4839), .B(exu_n16139), .Y(bypass_dfill_data_dff_n7));
AND2X1 exu_U9179(.A(exu_n4850), .B(exu_n16139), .Y(bypass_dfill_data_dff_n23));
AND2X1 exu_U9180(.A(exu_n4861), .B(exu_n16138), .Y(bypass_dfill_data_dff_n45));
AND2X1 exu_U9181(.A(exu_n4872), .B(exu_n16137), .Y(bypass_dfill_data_dff_n67));
AND2X1 exu_U9182(.A(exu_n4883), .B(exu_n16136), .Y(bypass_dfill_data_dff_n89));
INVX1 exu_U9183(.A(ecl_divcntl_subtract), .Y(exu_n16591));
INVX1 exu_U9184(.A(ecl_div_mul_wen), .Y(exu_n16186));
INVX1 exu_U9185(.A(ecl_shft_shift1_e[1]), .Y(exu_n16226));
INVX1 exu_U9186(.A(exu_n16147), .Y(exu_n16146));
AND2X1 exu_U9187(.A(exu_n19199), .B(exu_n5531), .Y(exu_n19187));
INVX1 exu_U9188(.A(ecl_byp_rs1_longmux_sel_g2), .Y(exu_n16284));
INVX1 exu_U9189(.A(ecl_byp_rs2_longmux_sel_g2), .Y(exu_n16281));
INVX1 exu_U9190(.A(ecl_byp_rs3_longmux_sel_g2), .Y(exu_n16278));
INVX1 exu_U9191(.A(ecl_byp_rs1_mux2_sel_ld), .Y(exu_n16313));
INVX1 exu_U9192(.A(ecl_byp_rcc_mux2_sel_ld), .Y(exu_n16304));
INVX1 exu_U9193(.A(ecl_byp_rs2_mux1_sel_w), .Y(exu_n16293));
INVX1 exu_U9194(.A(ecl_byp_rs2_mux2_sel_ld), .Y(exu_n16296));
INVX1 exu_U9195(.A(ecl_byp_rs3_mux1_sel_w), .Y(exu_n16289));
INVX1 exu_U9196(.A(ecl_byp_rs3_mux2_sel_ld), .Y(exu_n16291));
INVX1 exu_U9197(.A(ecl_alu_log_sel_move_e), .Y(exu_n16237));
INVX1 exu_U9198(.A(ecl_alu_log_sel_or_e), .Y(exu_n16239));
INVX1 exu_U9199(.A(ecl_byp_rs1_mux2_sel_usemux1), .Y(exu_n16312));
INVX1 exu_U9200(.A(ecl_byp_rcc_mux2_sel_usemux1), .Y(exu_n16303));
INVX1 exu_U9201(.A(ecl_byp_rs2_mux2_sel_e), .Y(exu_n16299));
INVX1 exu_U9202(.A(ecl_byp_rs2_mux2_sel_usemux1), .Y(exu_n16295));
INVX1 exu_U9203(.A(ecl_byp_rs3_mux2_sel_e), .Y(exu_n16292));
INVX1 exu_U9204(.A(ecl_alu_log_sel_xor_e), .Y(exu_n16238));
INVX1 exu_U9205(.A(ecl_alu_log_sel_and_e), .Y(exu_n16240));
INVX1 exu_U9206(.A(ecl_byp_sel_tlusr_m), .Y(exu_n16263));
AND2X1 exu_U9207(.A(exu_n774), .B(exu_n19222), .Y(exu_n19220));
INVX1 exu_U9208(.A(ecl_shft_shift4_e[1]), .Y(exu_n16231));
OR2X1 exu_U9209(.A(ecl_byp_restore_m), .B(se), .Y(ecl_writeback_restore_tid_dff_n6));
AND2X1 exu_U9210(.A(exu_n4905), .B(exu_n15821), .Y(rml_agp_wen_thr1_w));
AND2X1 exu_U9211(.A(exu_n4904), .B(exu_n15821), .Y(rml_agp_wen_thr2_w));
AND2X1 exu_U9212(.A(exu_n4903), .B(exu_n15821), .Y(rml_agp_wen_thr3_w));
AND2X1 exu_U9213(.A(exu_n4906), .B(exu_n15821), .Y(rml_agp_wen_thr0_w));
AND2X1 exu_U9214(.A(exu_n15238), .B(ecl_writeback_n54), .Y(ecl_writeback_n110));
AND2X1 exu_U9215(.A(exu_n15237), .B(exu_n16273), .Y(ecl_writeback_n198));
AND2X1 exu_U9216(.A(exu_n85), .B(exu_n5052), .Y(div_ecl_cout64));
AND2X1 exu_U9217(.A(ecl_wb_byplog_wen_g2), .B(exu_n15477), .Y(ecl_byp_sel_load_g));
AND2X1 exu_U9218(.A(ecl_tid_e[0]), .B(ecl_tid_e[1]), .Y(ecl_div_thr_e[3]));
INVX1 exu_U9219(.A(ecl_div_zero_rs2_e), .Y(exu_n16613));
INVX1 exu_U9220(.A(ecl_div_mul_get_32bit_data), .Y(exu_n16256));
AND2X1 exu_U9221(.A(ecl_mdqctl_mul_data[9]), .B(ecl_mdqctl_ismul_e), .Y(ecl_div_mul_get_new_data));
AND2X1 exu_U9222(.A(ecc_syn_mux_n21), .B(exu_n9370), .Y(ecc_err_m[1]));
AND2X1 exu_U9223(.A(exu_n15819), .B(exu_n15463), .Y(ecl_byp_rs3h_longmux_sel_w2));
INVX1 exu_U9224(.A(ecl_div_div64), .Y(exu_n16192));
AND2X1 exu_U9225(.A(ecc_syn_mux_n5), .B(exu_n9362), .Y(ecc_err_m[5]));
INVX1 exu_U9226(.A(ecl_tid_d[0]), .Y(exu_n15945));
INVX1 exu_U9227(.A(ecl_tid_d[1]), .Y(exu_n15944));
AND2X1 exu_U9228(.A(exu_n15348), .B(exu_n15420), .Y(ecl_byp_sel_yreg_e));
INVX1 exu_U9229(.A(ecl_sel_sum_e), .Y(exu_n16156));
INVX1 exu_U9230(.A(exu_n16155), .Y(exu_n16160));
AND2X1 exu_U9231(.A(exu_n4547), .B(ecl_mdqctl_wb_yreg_shift_g), .Y(ecl_writeback_n84));
AND2X1 exu_U9232(.A(exu_n4546), .B(ecl_mdqctl_wb_yreg_shift_g), .Y(ecl_writeback_n80));
AND2X1 exu_U9233(.A(exu_n4071), .B(ecl_divcntl_cntr[1]), .Y(ecl_divcntl_cnt6_n23));
AND2X1 exu_U9234(.A(exu_n15220), .B(exu_n9330), .Y(ecl_div_yreg_wen_l[0]));
AND2X1 exu_U9235(.A(exu_n15219), .B(ecl_writeback_n180), .Y(ecl_div_yreg_wen_w[1]));
AND2X1 exu_U9236(.A(exu_n15218), .B(ecl_writeback_n178), .Y(ecl_div_yreg_wen_w[2]));
AND2X1 exu_U9237(.A(exu_n15217), .B(ecl_writeback_n175), .Y(ecl_div_yreg_wen_w[3]));
AND2X1 exu_U9238(.A(exu_n4549), .B(ecl_writeback_n54), .Y(ecl_writeback_n129));
INVX1 exu_U9239(.A(exu_n16206), .Y(exu_n16203));
INVX1 exu_U9240(.A(ecl_div_ld_inputs), .Y(exu_n16206));
AND2X1 exu_U9241(.A(exu_n4548), .B(ecl_mdqctl_wb_yreg_shift_g), .Y(ecl_writeback_n191));
AND2X1 exu_U9242(.A(exu_n19235), .B(exu_n5536), .Y(exu_n19236));
AND2X1 exu_U9243(.A(exu_n15198), .B(exu_n9315), .Y(ecl_divcntl_n72));
AND2X1 exu_U9244(.A(exu_n4514), .B(ecl_ecl_div_signed_div), .Y(ecl_divcntl_n61));
INVX1 exu_U9245(.A(ecl_divcntl_N56), .Y(exu_n15979));
INVX1 exu_U9246(.A(ecl_mdqctl_ismul_e), .Y(exu_n15986));
INVX1 exu_U9247(.A(exu_n16194), .Y(exu_n16199));
INVX1 exu_U9248(.A(ecl_div_sel_div), .Y(exu_n16196));
INVX1 exu_U9249(.A(ecl_div_dividend_sign), .Y(exu_n16261));
INVX1 exu_U9250(.A(exu_n16261), .Y(exu_n16260));
AND2X1 exu_U9251(.A(alu_logic_rs1_data_bf1[31]), .B(ecl_mdqctl_mul_data[8]), .Y(ecl_div_mul_sext_rs1_e));
AND2X1 exu_U9252(.A(div_input_data_e[95]), .B(ecl_mdqctl_mul_data[8]), .Y(ecl_div_mul_sext_rs2_e));
AND2X1 exu_U9253(.A(div_input_data_e[95]), .B(ecl_ecl_div_signed_div), .Y(ecl_div_xinmask));
INVX1 exu_U9254(.A(sehold), .Y(ecl_writeback_n19));
INVX1 exu_U9255(.A(se), .Y(exu_n19277));
AND2X1 exu_U9256(.A(bypass_irf_write_clkbuf_tmb_l), .B(sehold), .Y(bypass_irf_write_clkbuf_N1));
INVX1 exu_U9257(.A(bypass_irf_write_clkbuf_N1), .Y(exu_n2));
INVX1 exu_U9258(.A(se), .Y(bypass_irf_write_clkbuf_tmb_l));
OR2X1 exu_U9259(.A(rml_tid_d[0]), .B(exu_n16574), .Y(exu_n15189));
INVX1 exu_U9260(.A(exu_n15189), .Y(exu_n3));
OR2X1 exu_U9261(.A(rml_tid_d[1]), .B(exu_n16573), .Y(exu_n15191));
OR2X1 exu_U9262(.A(rml_tid_d[1]), .B(rml_tid_d[0]), .Y(exu_n15193));
INVX1 exu_U9263(.A(exu_n15193), .Y(exu_n4));
INVX1 exu_U9264(.A(rml_tid_d[1]), .Y(exu_n16574));
INVX1 exu_U9265(.A(rml_tid_d[0]), .Y(exu_n16573));
AND2X1 exu_U9266(.A(exu_n16373), .B(exu_ifu_cc_d[7]), .Y(exu_n18011));
AND2X1 exu_U9267(.A(exu_ifu_cc_d[6]), .B(exu_n16373), .Y(exu_n18012));
AND2X1 exu_U9268(.A(shft_rshifterinput_b1[3]), .B(exu_n16148), .Y(exu_n27888));
INVX1 exu_U9269(.A(exu_n27888), .Y(exu_n5));
INVX1 exu_U9270(.A(exu_n16149), .Y(exu_n16148));
AND2X1 exu_U9271(.A(shft_rshifterinput_b1[2]), .B(shft_shift16_e[0]), .Y(exu_n27927));
INVX1 exu_U9272(.A(exu_n27927), .Y(exu_n6));
AND2X1 exu_U9273(.A(shft_rshifterinput_b1[1]), .B(exu_n16148), .Y(exu_n27958));
INVX1 exu_U9274(.A(exu_n27958), .Y(exu_n7));
AND2X1 exu_U9275(.A(shft_rshifterinput_b1[0]), .B(exu_n16148), .Y(exu_n27977));
INVX1 exu_U9276(.A(exu_n27977), .Y(exu_n8));
AND2X1 exu_U9277(.A(exu_n27977), .B(exu_n16230), .Y(exu_n28321));
OR2X1 exu_U9278(.A(exu_n16570), .B(rml_tid_e[1]), .Y(rml_n67));
INVX1 exu_U9279(.A(rml_n67), .Y(exu_n9));
AND2X1 exu_U9280(.A(exu_n10712), .B(exu_n9675), .Y(exu_n16634));
INVX1 exu_U9281(.A(exu_n16634), .Y(exu_n10));
AND2X1 exu_U9282(.A(exu_n10714), .B(exu_n9677), .Y(exu_n16648));
INVX1 exu_U9283(.A(exu_n16648), .Y(exu_n11));
AND2X1 exu_U9284(.A(exu_n10716), .B(exu_n9679), .Y(exu_n16662));
INVX1 exu_U9285(.A(exu_n16662), .Y(exu_n12));
OR2X1 exu_U9286(.A(exu_n11941), .B(exu_n14823), .Y(ecl_byplog_rs1_N1));
INVX1 exu_U9287(.A(ecl_byplog_rs1_N1), .Y(exu_n13));
AND2X1 exu_U9288(.A(exu_n10718), .B(exu_n9681), .Y(exu_n16676));
INVX1 exu_U9289(.A(exu_n16676), .Y(exu_n14));
OR2X1 exu_U9290(.A(exu_n11942), .B(exu_n14824), .Y(ecl_byplog_rs1_N0));
INVX1 exu_U9291(.A(ecl_byplog_rs1_N0), .Y(exu_n15));
AND2X1 exu_U9292(.A(exu_n10720), .B(exu_n9683), .Y(exu_n16690));
INVX1 exu_U9293(.A(exu_n16690), .Y(exu_n16));
AND2X1 exu_U9294(.A(exu_n10722), .B(exu_n9685), .Y(exu_n16704));
INVX1 exu_U9295(.A(exu_n16704), .Y(exu_n17));
AND2X1 exu_U9296(.A(exu_n10724), .B(exu_n9687), .Y(exu_n16718));
INVX1 exu_U9297(.A(exu_n16718), .Y(exu_n18));
OR2X1 exu_U9298(.A(exu_n11944), .B(exu_n14826), .Y(ecl_byplog_rs2_N1));
INVX1 exu_U9299(.A(ecl_byplog_rs2_N1), .Y(exu_n19));
AND2X1 exu_U9300(.A(exu_n10726), .B(exu_n9689), .Y(exu_n16732));
INVX1 exu_U9301(.A(exu_n16732), .Y(exu_n20));
OR2X1 exu_U9302(.A(exu_n11945), .B(exu_n14827), .Y(ecl_byplog_rs2_N0));
INVX1 exu_U9303(.A(ecl_byplog_rs2_N0), .Y(exu_n21));
AND2X1 exu_U9304(.A(div_adderin2[0]), .B(exu_n15859), .Y(exu_n16742));
INVX1 exu_U9305(.A(exu_n16742), .Y(exu_n22));
AND2X1 exu_U9306(.A(exu_n15910), .B(exu_n15559), .Y(exu_n16745));
INVX1 exu_U9307(.A(exu_n16745), .Y(exu_n23));
AND2X1 exu_U9308(.A(exu_n15899), .B(exu_n15560), .Y(exu_n16748));
INVX1 exu_U9309(.A(exu_n16748), .Y(exu_n24));
AND2X1 exu_U9310(.A(exu_n15889), .B(exu_n15561), .Y(exu_n16751));
INVX1 exu_U9311(.A(exu_n16751), .Y(exu_n25));
AND2X1 exu_U9312(.A(exu_n15878), .B(exu_n15562), .Y(exu_n16754));
INVX1 exu_U9313(.A(exu_n16754), .Y(exu_n26));
AND2X1 exu_U9314(.A(exu_n15867), .B(exu_n15563), .Y(exu_n16757));
INVX1 exu_U9315(.A(exu_n16757), .Y(exu_n27));
AND2X1 exu_U9316(.A(exu_n15863), .B(exu_n15564), .Y(exu_n16760));
INVX1 exu_U9317(.A(exu_n16760), .Y(exu_n28));
AND2X1 exu_U9318(.A(exu_n15862), .B(exu_n15565), .Y(exu_n16763));
INVX1 exu_U9319(.A(exu_n16763), .Y(exu_n29));
AND2X1 exu_U9320(.A(exu_n15861), .B(exu_n15566), .Y(exu_n16766));
INVX1 exu_U9321(.A(exu_n16766), .Y(exu_n30));
AND2X1 exu_U9322(.A(exu_n15860), .B(exu_n15567), .Y(exu_n16769));
INVX1 exu_U9323(.A(exu_n16769), .Y(exu_n31));
AND2X1 exu_U9324(.A(exu_n15920), .B(exu_n15595), .Y(exu_n16774));
INVX1 exu_U9325(.A(exu_n16774), .Y(exu_n32));
AND2X1 exu_U9326(.A(exu_n15919), .B(exu_n15596), .Y(exu_n16779));
INVX1 exu_U9327(.A(exu_n16779), .Y(exu_n33));
AND2X1 exu_U9328(.A(exu_n15918), .B(exu_n15597), .Y(exu_n16784));
INVX1 exu_U9329(.A(exu_n16784), .Y(exu_n34));
AND2X1 exu_U9330(.A(exu_n15917), .B(exu_n15598), .Y(exu_n16789));
INVX1 exu_U9331(.A(exu_n16789), .Y(exu_n35));
AND2X1 exu_U9332(.A(exu_n15916), .B(exu_n15599), .Y(exu_n16794));
INVX1 exu_U9333(.A(exu_n16794), .Y(exu_n36));
AND2X1 exu_U9334(.A(exu_n15915), .B(exu_n15600), .Y(exu_n16799));
INVX1 exu_U9335(.A(exu_n16799), .Y(exu_n37));
AND2X1 exu_U9336(.A(exu_n15914), .B(exu_n15601), .Y(exu_n16804));
INVX1 exu_U9337(.A(exu_n16804), .Y(exu_n38));
AND2X1 exu_U9338(.A(exu_n15913), .B(exu_n15602), .Y(exu_n16809));
INVX1 exu_U9339(.A(exu_n16809), .Y(exu_n39));
AND2X1 exu_U9340(.A(exu_n15912), .B(exu_n15603), .Y(exu_n16814));
INVX1 exu_U9341(.A(exu_n16814), .Y(exu_n40));
AND2X1 exu_U9342(.A(exu_n15911), .B(exu_n15604), .Y(exu_n16821));
INVX1 exu_U9343(.A(exu_n16821), .Y(exu_n41));
AND2X1 exu_U9344(.A(exu_n15909), .B(exu_n15605), .Y(exu_n16826));
INVX1 exu_U9345(.A(exu_n16826), .Y(exu_n42));
AND2X1 exu_U9346(.A(exu_n15908), .B(exu_n15606), .Y(exu_n16831));
INVX1 exu_U9347(.A(exu_n16831), .Y(exu_n43));
AND2X1 exu_U9348(.A(exu_n15907), .B(exu_n15607), .Y(exu_n16836));
INVX1 exu_U9349(.A(exu_n16836), .Y(exu_n44));
AND2X1 exu_U9350(.A(exu_n15906), .B(exu_n15608), .Y(exu_n16841));
INVX1 exu_U9351(.A(exu_n16841), .Y(exu_n45));
AND2X1 exu_U9352(.A(exu_n15905), .B(exu_n15609), .Y(exu_n16846));
INVX1 exu_U9353(.A(exu_n16846), .Y(exu_n46));
AND2X1 exu_U9354(.A(exu_n15904), .B(exu_n15610), .Y(exu_n16851));
INVX1 exu_U9355(.A(exu_n16851), .Y(exu_n47));
AND2X1 exu_U9356(.A(exu_n15903), .B(exu_n15611), .Y(exu_n16856));
INVX1 exu_U9357(.A(exu_n16856), .Y(exu_n48));
AND2X1 exu_U9358(.A(exu_n15902), .B(exu_n15612), .Y(exu_n16861));
INVX1 exu_U9359(.A(exu_n16861), .Y(exu_n49));
AND2X1 exu_U9360(.A(exu_n15901), .B(exu_n15613), .Y(exu_n16866));
INVX1 exu_U9361(.A(exu_n16866), .Y(exu_n50));
AND2X1 exu_U9362(.A(exu_n15900), .B(exu_n15614), .Y(exu_n16873));
INVX1 exu_U9363(.A(exu_n16873), .Y(exu_n51));
AND2X1 exu_U9364(.A(exu_n15898), .B(exu_n15615), .Y(exu_n16878));
INVX1 exu_U9365(.A(exu_n16878), .Y(exu_n52));
AND2X1 exu_U9366(.A(exu_n15897), .B(exu_n15616), .Y(exu_n16883));
INVX1 exu_U9367(.A(exu_n16883), .Y(exu_n53));
AND2X1 exu_U9368(.A(div_adderin2[32]), .B(exu_n15858), .Y(exu_n16901));
INVX1 exu_U9369(.A(exu_n16901), .Y(exu_n54));
AND2X1 exu_U9370(.A(exu_n15896), .B(exu_n15568), .Y(exu_n16904));
INVX1 exu_U9371(.A(exu_n16904), .Y(exu_n55));
AND2X1 exu_U9372(.A(exu_n15895), .B(exu_n15569), .Y(exu_n16907));
INVX1 exu_U9373(.A(exu_n16907), .Y(exu_n56));
AND2X1 exu_U9374(.A(exu_n15894), .B(exu_n15570), .Y(exu_n16910));
INVX1 exu_U9375(.A(exu_n16910), .Y(exu_n57));
AND2X1 exu_U9376(.A(exu_n15893), .B(exu_n15571), .Y(exu_n16913));
INVX1 exu_U9377(.A(exu_n16913), .Y(exu_n58));
AND2X1 exu_U9378(.A(exu_n15892), .B(exu_n15572), .Y(exu_n16916));
INVX1 exu_U9379(.A(exu_n16916), .Y(exu_n59));
AND2X1 exu_U9380(.A(exu_n15891), .B(exu_n15573), .Y(exu_n16919));
INVX1 exu_U9381(.A(exu_n16919), .Y(exu_n60));
AND2X1 exu_U9382(.A(exu_n15890), .B(exu_n15574), .Y(exu_n16922));
INVX1 exu_U9383(.A(exu_n16922), .Y(exu_n61));
AND2X1 exu_U9384(.A(exu_n15888), .B(exu_n15575), .Y(exu_n16925));
INVX1 exu_U9385(.A(exu_n16925), .Y(exu_n62));
AND2X1 exu_U9386(.A(exu_n15887), .B(exu_n15576), .Y(exu_n16928));
INVX1 exu_U9387(.A(exu_n16928), .Y(exu_n63));
AND2X1 exu_U9388(.A(exu_n15886), .B(exu_n15617), .Y(exu_n16933));
INVX1 exu_U9389(.A(exu_n16933), .Y(exu_n64));
AND2X1 exu_U9390(.A(exu_n15885), .B(exu_n15618), .Y(exu_n16938));
INVX1 exu_U9391(.A(exu_n16938), .Y(exu_n65));
AND2X1 exu_U9392(.A(exu_n15884), .B(exu_n15619), .Y(exu_n16943));
INVX1 exu_U9393(.A(exu_n16943), .Y(exu_n66));
AND2X1 exu_U9394(.A(exu_n15883), .B(exu_n15620), .Y(exu_n16948));
INVX1 exu_U9395(.A(exu_n16948), .Y(exu_n67));
AND2X1 exu_U9396(.A(exu_n15882), .B(exu_n15621), .Y(exu_n16953));
INVX1 exu_U9397(.A(exu_n16953), .Y(exu_n68));
AND2X1 exu_U9398(.A(exu_n15881), .B(exu_n15622), .Y(exu_n16958));
INVX1 exu_U9399(.A(exu_n16958), .Y(exu_n69));
AND2X1 exu_U9400(.A(exu_n15880), .B(exu_n15623), .Y(exu_n16963));
INVX1 exu_U9401(.A(exu_n16963), .Y(exu_n70));
AND2X1 exu_U9402(.A(exu_n15879), .B(exu_n15624), .Y(exu_n16968));
INVX1 exu_U9403(.A(exu_n16968), .Y(exu_n71));
AND2X1 exu_U9404(.A(exu_n15877), .B(exu_n15625), .Y(exu_n16973));
INVX1 exu_U9405(.A(exu_n16973), .Y(exu_n72));
AND2X1 exu_U9406(.A(exu_n15876), .B(exu_n15626), .Y(exu_n16980));
INVX1 exu_U9407(.A(exu_n16980), .Y(exu_n73));
AND2X1 exu_U9408(.A(exu_n15875), .B(exu_n15627), .Y(exu_n16985));
INVX1 exu_U9409(.A(exu_n16985), .Y(exu_n74));
AND2X1 exu_U9410(.A(exu_n15874), .B(exu_n15628), .Y(exu_n16990));
INVX1 exu_U9411(.A(exu_n16990), .Y(exu_n75));
AND2X1 exu_U9412(.A(exu_n15873), .B(exu_n15629), .Y(exu_n16995));
INVX1 exu_U9413(.A(exu_n16995), .Y(exu_n76));
AND2X1 exu_U9414(.A(exu_n15872), .B(exu_n15630), .Y(exu_n17000));
INVX1 exu_U9415(.A(exu_n17000), .Y(exu_n77));
AND2X1 exu_U9416(.A(exu_n15871), .B(exu_n15631), .Y(exu_n17005));
INVX1 exu_U9417(.A(exu_n17005), .Y(exu_n78));
AND2X1 exu_U9418(.A(exu_n15870), .B(exu_n15632), .Y(exu_n17010));
INVX1 exu_U9419(.A(exu_n17010), .Y(exu_n79));
AND2X1 exu_U9420(.A(exu_n15869), .B(exu_n15633), .Y(exu_n17015));
INVX1 exu_U9421(.A(exu_n17015), .Y(exu_n80));
AND2X1 exu_U9422(.A(exu_n15868), .B(exu_n15634), .Y(exu_n17020));
INVX1 exu_U9423(.A(exu_n17020), .Y(exu_n81));
AND2X1 exu_U9424(.A(exu_n15866), .B(exu_n15635), .Y(exu_n17025));
INVX1 exu_U9425(.A(exu_n17025), .Y(exu_n82));
AND2X1 exu_U9426(.A(exu_n15865), .B(exu_n15636), .Y(exu_n17032));
INVX1 exu_U9427(.A(exu_n17032), .Y(exu_n83));
AND2X1 exu_U9428(.A(exu_n15864), .B(exu_n15637), .Y(exu_n17037));
INVX1 exu_U9429(.A(exu_n17037), .Y(exu_n84));
AND2X1 exu_U9430(.A(exu_n15823), .B(exu_n15638), .Y(exu_n17042));
INVX1 exu_U9431(.A(exu_n17042), .Y(exu_n85));
AND2X1 exu_U9432(.A(alu_addsub_rs2_data_0), .B(alu_logic_rs1_data_bf1[0]), .Y(exu_n17060));
INVX1 exu_U9433(.A(exu_n17060), .Y(exu_n86));
AND2X1 exu_U9434(.A(alu_logic_rs1_data_bf1[1]), .B(exu_n15577), .Y(exu_n17063));
INVX1 exu_U9435(.A(exu_n17063), .Y(exu_n87));
AND2X1 exu_U9436(.A(alu_logic_rs1_data_bf1[2]), .B(exu_n15578), .Y(exu_n17066));
INVX1 exu_U9437(.A(exu_n17066), .Y(exu_n88));
AND2X1 exu_U9438(.A(alu_logic_rs1_data_bf1[3]), .B(exu_n15579), .Y(exu_n17069));
INVX1 exu_U9439(.A(exu_n17069), .Y(exu_n89));
AND2X1 exu_U9440(.A(alu_logic_rs1_data_bf1[4]), .B(exu_n15580), .Y(exu_n17072));
INVX1 exu_U9441(.A(exu_n17072), .Y(exu_n90));
AND2X1 exu_U9442(.A(alu_logic_rs1_data_bf1[5]), .B(exu_n15581), .Y(exu_n17075));
INVX1 exu_U9443(.A(exu_n17075), .Y(exu_n91));
AND2X1 exu_U9444(.A(alu_logic_rs1_data_bf1[6]), .B(exu_n15582), .Y(exu_n17078));
INVX1 exu_U9445(.A(exu_n17078), .Y(exu_n92));
AND2X1 exu_U9446(.A(alu_logic_rs1_data_bf1[7]), .B(exu_n15583), .Y(exu_n17081));
INVX1 exu_U9447(.A(exu_n17081), .Y(exu_n93));
AND2X1 exu_U9448(.A(alu_logic_rs1_data_bf1[8]), .B(exu_n15584), .Y(exu_n17084));
INVX1 exu_U9449(.A(exu_n17084), .Y(exu_n94));
AND2X1 exu_U9450(.A(alu_logic_rs1_data_bf1[9]), .B(exu_n15585), .Y(exu_n17087));
INVX1 exu_U9451(.A(exu_n17087), .Y(exu_n95));
AND2X1 exu_U9452(.A(alu_logic_rs1_data_bf1[10]), .B(exu_n15639), .Y(exu_n17092));
INVX1 exu_U9453(.A(exu_n17092), .Y(exu_n96));
AND2X1 exu_U9454(.A(alu_logic_rs1_data_bf1[11]), .B(exu_n15640), .Y(exu_n17097));
INVX1 exu_U9455(.A(exu_n17097), .Y(exu_n97));
AND2X1 exu_U9456(.A(alu_logic_rs1_data_bf1[12]), .B(exu_n15641), .Y(exu_n17102));
INVX1 exu_U9457(.A(exu_n17102), .Y(exu_n98));
AND2X1 exu_U9458(.A(alu_logic_rs1_data_bf1[13]), .B(exu_n15642), .Y(exu_n17107));
INVX1 exu_U9459(.A(exu_n17107), .Y(exu_n99));
AND2X1 exu_U9460(.A(alu_logic_rs1_data_bf1[14]), .B(exu_n15643), .Y(exu_n17112));
INVX1 exu_U9461(.A(exu_n17112), .Y(exu_n100));
AND2X1 exu_U9462(.A(alu_logic_rs1_data_bf1[15]), .B(exu_n15644), .Y(exu_n17117));
INVX1 exu_U9463(.A(exu_n17117), .Y(exu_n101));
AND2X1 exu_U9464(.A(alu_logic_rs1_data_bf1[16]), .B(exu_n15645), .Y(exu_n17122));
INVX1 exu_U9465(.A(exu_n17122), .Y(exu_n102));
AND2X1 exu_U9466(.A(alu_logic_rs1_data_bf1[17]), .B(exu_n15646), .Y(exu_n17127));
INVX1 exu_U9467(.A(exu_n17127), .Y(exu_n103));
AND2X1 exu_U9468(.A(alu_logic_rs1_data_bf1[18]), .B(exu_n15647), .Y(exu_n17132));
INVX1 exu_U9469(.A(exu_n17132), .Y(exu_n104));
AND2X1 exu_U9470(.A(alu_logic_rs1_data_bf1[19]), .B(exu_n15648), .Y(exu_n17139));
INVX1 exu_U9471(.A(exu_n17139), .Y(exu_n105));
AND2X1 exu_U9472(.A(alu_logic_rs1_data_bf1[20]), .B(exu_n15649), .Y(exu_n17144));
INVX1 exu_U9473(.A(exu_n17144), .Y(exu_n106));
AND2X1 exu_U9474(.A(alu_logic_rs1_data_bf1[21]), .B(exu_n15650), .Y(exu_n17149));
INVX1 exu_U9475(.A(exu_n17149), .Y(exu_n107));
AND2X1 exu_U9476(.A(alu_logic_rs1_data_bf1[22]), .B(exu_n15651), .Y(exu_n17154));
INVX1 exu_U9477(.A(exu_n17154), .Y(exu_n108));
AND2X1 exu_U9478(.A(alu_logic_rs1_data_bf1[23]), .B(exu_n15652), .Y(exu_n17159));
INVX1 exu_U9479(.A(exu_n17159), .Y(exu_n109));
AND2X1 exu_U9480(.A(alu_logic_rs1_data_bf1[24]), .B(exu_n15653), .Y(exu_n17164));
INVX1 exu_U9481(.A(exu_n17164), .Y(exu_n110));
AND2X1 exu_U9482(.A(alu_logic_rs1_data_bf1[25]), .B(exu_n15654), .Y(exu_n17169));
INVX1 exu_U9483(.A(exu_n17169), .Y(exu_n111));
AND2X1 exu_U9484(.A(alu_logic_rs1_data_bf1[26]), .B(exu_n15655), .Y(exu_n17174));
INVX1 exu_U9485(.A(exu_n17174), .Y(exu_n112));
AND2X1 exu_U9486(.A(alu_logic_rs1_data_bf1[27]), .B(exu_n15656), .Y(exu_n17179));
INVX1 exu_U9487(.A(exu_n17179), .Y(exu_n113));
AND2X1 exu_U9488(.A(alu_logic_rs1_data_bf1[28]), .B(exu_n15657), .Y(exu_n17184));
INVX1 exu_U9489(.A(exu_n17184), .Y(exu_n114));
AND2X1 exu_U9490(.A(alu_logic_rs1_data_bf1[29]), .B(exu_n15658), .Y(exu_n17191));
INVX1 exu_U9491(.A(exu_n17191), .Y(exu_n115));
AND2X1 exu_U9492(.A(alu_logic_rs1_data_bf1[30]), .B(exu_n15659), .Y(exu_n17196));
INVX1 exu_U9493(.A(exu_n17196), .Y(exu_n116));
AND2X1 exu_U9494(.A(alu_logic_rs1_data_bf1[31]), .B(exu_n15660), .Y(exu_n17201));
INVX1 exu_U9495(.A(exu_n17201), .Y(exu_n117));
AND2X1 exu_U9496(.A(alu_addsub_rs2_data[32]), .B(alu_logic_rs1_data_bf1[32]), .Y(exu_n17219));
INVX1 exu_U9497(.A(exu_n17219), .Y(exu_n118));
AND2X1 exu_U9498(.A(alu_logic_rs1_data_bf1[33]), .B(exu_n15586), .Y(exu_n17222));
INVX1 exu_U9499(.A(exu_n17222), .Y(exu_n119));
AND2X1 exu_U9500(.A(alu_logic_rs1_data_bf1[34]), .B(exu_n15587), .Y(exu_n17225));
INVX1 exu_U9501(.A(exu_n17225), .Y(exu_n120));
AND2X1 exu_U9502(.A(alu_logic_rs1_data_bf1[35]), .B(exu_n15588), .Y(exu_n17228));
INVX1 exu_U9503(.A(exu_n17228), .Y(exu_n121));
AND2X1 exu_U9504(.A(alu_logic_rs1_data_bf1[36]), .B(exu_n15589), .Y(exu_n17231));
INVX1 exu_U9505(.A(exu_n17231), .Y(exu_n122));
AND2X1 exu_U9506(.A(alu_logic_rs1_data_bf1[37]), .B(exu_n15590), .Y(exu_n17234));
INVX1 exu_U9507(.A(exu_n17234), .Y(exu_n123));
AND2X1 exu_U9508(.A(alu_logic_rs1_data_bf1[38]), .B(exu_n15591), .Y(exu_n17237));
INVX1 exu_U9509(.A(exu_n17237), .Y(exu_n124));
AND2X1 exu_U9510(.A(alu_logic_rs1_data_bf1[39]), .B(exu_n15592), .Y(exu_n17240));
INVX1 exu_U9511(.A(exu_n17240), .Y(exu_n125));
AND2X1 exu_U9512(.A(alu_logic_rs1_data_bf1[40]), .B(exu_n15593), .Y(exu_n17243));
INVX1 exu_U9513(.A(exu_n17243), .Y(exu_n126));
AND2X1 exu_U9514(.A(alu_logic_rs1_data_bf1[41]), .B(exu_n15594), .Y(exu_n17246));
INVX1 exu_U9515(.A(exu_n17246), .Y(exu_n127));
AND2X1 exu_U9516(.A(alu_logic_rs1_data_bf1[42]), .B(exu_n15661), .Y(exu_n17251));
INVX1 exu_U9517(.A(exu_n17251), .Y(exu_n128));
AND2X1 exu_U9518(.A(alu_logic_rs1_data_bf1[43]), .B(exu_n15662), .Y(exu_n17256));
INVX1 exu_U9519(.A(exu_n17256), .Y(exu_n129));
AND2X1 exu_U9520(.A(alu_logic_rs1_data_bf1[44]), .B(exu_n15663), .Y(exu_n17261));
INVX1 exu_U9521(.A(exu_n17261), .Y(exu_n130));
AND2X1 exu_U9522(.A(alu_logic_rs1_data_bf1[45]), .B(exu_n15664), .Y(exu_n17266));
INVX1 exu_U9523(.A(exu_n17266), .Y(exu_n131));
AND2X1 exu_U9524(.A(alu_logic_rs1_data_bf1[46]), .B(exu_n15665), .Y(exu_n17271));
INVX1 exu_U9525(.A(exu_n17271), .Y(exu_n132));
AND2X1 exu_U9526(.A(alu_logic_rs1_data_bf1[47]), .B(exu_n15666), .Y(exu_n17276));
INVX1 exu_U9527(.A(exu_n17276), .Y(exu_n133));
AND2X1 exu_U9528(.A(alu_logic_rs1_data_bf1[48]), .B(exu_n15667), .Y(exu_n17281));
INVX1 exu_U9529(.A(exu_n17281), .Y(exu_n134));
AND2X1 exu_U9530(.A(alu_logic_rs1_data_bf1[49]), .B(exu_n15668), .Y(exu_n17286));
INVX1 exu_U9531(.A(exu_n17286), .Y(exu_n135));
AND2X1 exu_U9532(.A(alu_logic_rs1_data_bf1[50]), .B(exu_n15669), .Y(exu_n17291));
INVX1 exu_U9533(.A(exu_n17291), .Y(exu_n136));
AND2X1 exu_U9534(.A(alu_logic_rs1_data_bf1[51]), .B(exu_n15670), .Y(exu_n17298));
INVX1 exu_U9535(.A(exu_n17298), .Y(exu_n137));
AND2X1 exu_U9536(.A(alu_logic_rs1_data_bf1[52]), .B(exu_n15671), .Y(exu_n17303));
INVX1 exu_U9537(.A(exu_n17303), .Y(exu_n138));
AND2X1 exu_U9538(.A(alu_logic_rs1_data_bf1[53]), .B(exu_n15672), .Y(exu_n17308));
INVX1 exu_U9539(.A(exu_n17308), .Y(exu_n139));
AND2X1 exu_U9540(.A(alu_logic_rs1_data_bf1[54]), .B(exu_n15673), .Y(exu_n17313));
INVX1 exu_U9541(.A(exu_n17313), .Y(exu_n140));
AND2X1 exu_U9542(.A(alu_logic_rs1_data_bf1[55]), .B(exu_n15674), .Y(exu_n17318));
INVX1 exu_U9543(.A(exu_n17318), .Y(exu_n141));
AND2X1 exu_U9544(.A(alu_logic_rs1_data_bf1[56]), .B(exu_n15675), .Y(exu_n17323));
INVX1 exu_U9545(.A(exu_n17323), .Y(exu_n142));
AND2X1 exu_U9546(.A(alu_logic_rs1_data_bf1[57]), .B(exu_n15676), .Y(exu_n17328));
INVX1 exu_U9547(.A(exu_n17328), .Y(exu_n143));
AND2X1 exu_U9548(.A(alu_logic_rs1_data_bf1[58]), .B(exu_n15677), .Y(exu_n17333));
INVX1 exu_U9549(.A(exu_n17333), .Y(exu_n144));
AND2X1 exu_U9550(.A(alu_logic_rs1_data_bf1[59]), .B(exu_n15678), .Y(exu_n17338));
INVX1 exu_U9551(.A(exu_n17338), .Y(exu_n145));
AND2X1 exu_U9552(.A(alu_logic_rs1_data_bf1[60]), .B(exu_n15679), .Y(exu_n17343));
INVX1 exu_U9553(.A(exu_n17343), .Y(exu_n146));
AND2X1 exu_U9554(.A(alu_logic_rs1_data_bf1[61]), .B(exu_n15680), .Y(exu_n17350));
INVX1 exu_U9555(.A(exu_n17350), .Y(exu_n147));
AND2X1 exu_U9556(.A(alu_logic_rs1_data_bf1[62]), .B(exu_n15681), .Y(exu_n17355));
INVX1 exu_U9557(.A(exu_n17355), .Y(exu_n148));
AND2X1 exu_U9558(.A(alu_logic_rs1_data_bf1[63]), .B(exu_n15682), .Y(exu_n17360));
INVX1 exu_U9559(.A(exu_n17360), .Y(exu_n149));
OR2X1 exu_U9560(.A(exu_n11947), .B(exu_n14829), .Y(ecl_byplog_rs3h_N1));
INVX1 exu_U9561(.A(ecl_byplog_rs3h_N1), .Y(exu_n150));
OR2X1 exu_U9562(.A(exu_n11948), .B(exu_n14830), .Y(ecl_byplog_rs3h_N0));
INVX1 exu_U9563(.A(ecl_byplog_rs3h_N0), .Y(exu_n151));
AND2X1 exu_U9564(.A(exu_n10728), .B(exu_n9691), .Y(exu_n17410));
INVX1 exu_U9565(.A(exu_n17410), .Y(exu_n152));
AND2X1 exu_U9566(.A(exu_n10730), .B(exu_n9693), .Y(exu_n17424));
INVX1 exu_U9567(.A(exu_n17424), .Y(exu_n153));
AND2X1 exu_U9568(.A(exu_n10732), .B(exu_n9695), .Y(exu_n17438));
INVX1 exu_U9569(.A(exu_n17438), .Y(exu_n154));
OR2X1 exu_U9570(.A(exu_n11950), .B(exu_n14832), .Y(ecl_byplog_rs3_N1));
INVX1 exu_U9571(.A(ecl_byplog_rs3_N1), .Y(exu_n155));
AND2X1 exu_U9572(.A(exu_n10734), .B(exu_n9697), .Y(exu_n17452));
INVX1 exu_U9573(.A(exu_n17452), .Y(exu_n156));
OR2X1 exu_U9574(.A(exu_n11951), .B(exu_n14833), .Y(ecl_byplog_rs3_N0));
INVX1 exu_U9575(.A(ecl_byplog_rs3_N0), .Y(exu_n157));
AND2X1 exu_U9576(.A(exu_n10736), .B(exu_n9699), .Y(rml_cwp_next_slot1_data[9]));
INVX1 exu_U9577(.A(rml_cwp_next_slot1_data[9]), .Y(exu_n158));
AND2X1 exu_U9578(.A(exu_n10737), .B(exu_n9700), .Y(rml_cwp_next_slot1_data[8]));
INVX1 exu_U9579(.A(rml_cwp_next_slot1_data[8]), .Y(exu_n159));
AND2X1 exu_U9580(.A(exu_n15488), .B(exu_n9701), .Y(rml_cwp_next_slot1_data[7]));
INVX1 exu_U9581(.A(rml_cwp_next_slot1_data[7]), .Y(exu_n160));
AND2X1 exu_U9582(.A(exu_n10738), .B(exu_n9702), .Y(rml_cwp_next_slot1_data[6]));
INVX1 exu_U9583(.A(rml_cwp_next_slot1_data[6]), .Y(exu_n161));
AND2X1 exu_U9584(.A(exu_n17513), .B(exu_n9703), .Y(rml_cwp_next_slot1_data[5]));
INVX1 exu_U9585(.A(rml_cwp_next_slot1_data[5]), .Y(exu_n162));
AND2X1 exu_U9586(.A(rml_cwp_tlu_exu_cwp_w[2]), .B(rml_cwp_n34), .Y(exu_n17515));
INVX1 exu_U9587(.A(exu_n17515), .Y(exu_n163));
AND2X1 exu_U9588(.A(exu_n17517), .B(exu_n9704), .Y(rml_cwp_next_slot1_data[4]));
INVX1 exu_U9589(.A(rml_cwp_next_slot1_data[4]), .Y(exu_n164));
AND2X1 exu_U9590(.A(rml_cwp_tlu_exu_cwp_w[1]), .B(rml_cwp_n34), .Y(exu_n17519));
INVX1 exu_U9591(.A(exu_n17519), .Y(exu_n165));
AND2X1 exu_U9592(.A(exu_n17521), .B(exu_n9705), .Y(rml_cwp_next_slot1_data[3]));
INVX1 exu_U9593(.A(rml_cwp_next_slot1_data[3]), .Y(exu_n166));
AND2X1 exu_U9594(.A(rml_cwp_tlu_exu_cwp_w[0]), .B(rml_cwp_n34), .Y(exu_n17523));
INVX1 exu_U9595(.A(exu_n17523), .Y(exu_n167));
AND2X1 exu_U9596(.A(exu_n17525), .B(exu_n9706), .Y(rml_cwp_next_slot1_data[2]));
INVX1 exu_U9597(.A(rml_cwp_next_slot1_data[2]), .Y(exu_n168));
AND2X1 exu_U9598(.A(rml_cwp_old_cwp_w[2]), .B(rml_cwp_n34), .Y(exu_n17527));
INVX1 exu_U9599(.A(exu_n17527), .Y(exu_n169));
AND2X1 exu_U9600(.A(exu_n17529), .B(exu_n9707), .Y(rml_cwp_next_slot1_data[1]));
INVX1 exu_U9601(.A(rml_cwp_next_slot1_data[1]), .Y(exu_n170));
AND2X1 exu_U9602(.A(rml_cwp_old_cwp_w[1]), .B(rml_cwp_n34), .Y(exu_n17531));
INVX1 exu_U9603(.A(exu_n17531), .Y(exu_n171));
AND2X1 exu_U9604(.A(exu_n10739), .B(exu_n9708), .Y(rml_cwp_next_slot1_data[12]));
INVX1 exu_U9605(.A(rml_cwp_next_slot1_data[12]), .Y(exu_n172));
AND2X1 exu_U9606(.A(exu_n10740), .B(exu_n9709), .Y(rml_cwp_next_slot1_data[11]));
INVX1 exu_U9607(.A(rml_cwp_next_slot1_data[11]), .Y(exu_n173));
AND2X1 exu_U9608(.A(exu_n10741), .B(exu_n9710), .Y(rml_cwp_next_slot1_data[10]));
INVX1 exu_U9609(.A(rml_cwp_next_slot1_data[10]), .Y(exu_n174));
AND2X1 exu_U9610(.A(exu_n17539), .B(exu_n9711), .Y(rml_cwp_next_slot1_data[0]));
INVX1 exu_U9611(.A(rml_cwp_next_slot1_data[0]), .Y(exu_n175));
AND2X1 exu_U9612(.A(rml_cwp_old_cwp_w[0]), .B(rml_cwp_n34), .Y(exu_n17541));
INVX1 exu_U9613(.A(exu_n17541), .Y(exu_n176));
AND2X1 exu_U9614(.A(exu_n10742), .B(exu_n9712), .Y(rml_cwp_next_slot2_data[9]));
INVX1 exu_U9615(.A(rml_cwp_next_slot2_data[9]), .Y(exu_n177));
AND2X1 exu_U9616(.A(exu_n10743), .B(exu_n9713), .Y(rml_cwp_next_slot2_data[8]));
INVX1 exu_U9617(.A(rml_cwp_next_slot2_data[8]), .Y(exu_n178));
AND2X1 exu_U9618(.A(exu_n15489), .B(exu_n9714), .Y(rml_cwp_next_slot2_data[7]));
INVX1 exu_U9619(.A(rml_cwp_next_slot2_data[7]), .Y(exu_n179));
AND2X1 exu_U9620(.A(exu_n10744), .B(exu_n9715), .Y(rml_cwp_next_slot2_data[6]));
INVX1 exu_U9621(.A(rml_cwp_next_slot2_data[6]), .Y(exu_n180));
AND2X1 exu_U9622(.A(exu_n17550), .B(exu_n9716), .Y(rml_cwp_next_slot2_data[5]));
INVX1 exu_U9623(.A(rml_cwp_next_slot2_data[5]), .Y(exu_n181));
AND2X1 exu_U9624(.A(rml_cwp_tlu_exu_cwp_w[2]), .B(rml_cwp_n33), .Y(exu_n17552));
INVX1 exu_U9625(.A(exu_n17552), .Y(exu_n182));
AND2X1 exu_U9626(.A(exu_n17554), .B(exu_n9717), .Y(rml_cwp_next_slot2_data[4]));
INVX1 exu_U9627(.A(rml_cwp_next_slot2_data[4]), .Y(exu_n183));
AND2X1 exu_U9628(.A(rml_cwp_tlu_exu_cwp_w[1]), .B(rml_cwp_n33), .Y(exu_n17556));
INVX1 exu_U9629(.A(exu_n17556), .Y(exu_n184));
AND2X1 exu_U9630(.A(exu_n17558), .B(exu_n9718), .Y(rml_cwp_next_slot2_data[3]));
INVX1 exu_U9631(.A(rml_cwp_next_slot2_data[3]), .Y(exu_n185));
AND2X1 exu_U9632(.A(rml_cwp_tlu_exu_cwp_w[0]), .B(rml_cwp_n33), .Y(exu_n17560));
INVX1 exu_U9633(.A(exu_n17560), .Y(exu_n186));
AND2X1 exu_U9634(.A(exu_n17562), .B(exu_n9719), .Y(rml_cwp_next_slot2_data[2]));
INVX1 exu_U9635(.A(rml_cwp_next_slot2_data[2]), .Y(exu_n187));
AND2X1 exu_U9636(.A(rml_cwp_old_cwp_w[2]), .B(rml_cwp_n33), .Y(exu_n17564));
INVX1 exu_U9637(.A(exu_n17564), .Y(exu_n188));
AND2X1 exu_U9638(.A(exu_n17566), .B(exu_n9720), .Y(rml_cwp_next_slot2_data[1]));
INVX1 exu_U9639(.A(rml_cwp_next_slot2_data[1]), .Y(exu_n189));
AND2X1 exu_U9640(.A(rml_cwp_old_cwp_w[1]), .B(rml_cwp_n33), .Y(exu_n17568));
INVX1 exu_U9641(.A(exu_n17568), .Y(exu_n190));
AND2X1 exu_U9642(.A(exu_n10745), .B(exu_n9721), .Y(rml_cwp_next_slot2_data[12]));
INVX1 exu_U9643(.A(rml_cwp_next_slot2_data[12]), .Y(exu_n191));
AND2X1 exu_U9644(.A(exu_n10746), .B(exu_n9722), .Y(rml_cwp_next_slot2_data[11]));
INVX1 exu_U9645(.A(rml_cwp_next_slot2_data[11]), .Y(exu_n192));
AND2X1 exu_U9646(.A(exu_n10747), .B(exu_n9723), .Y(rml_cwp_next_slot2_data[10]));
INVX1 exu_U9647(.A(rml_cwp_next_slot2_data[10]), .Y(exu_n193));
AND2X1 exu_U9648(.A(exu_n17576), .B(exu_n9724), .Y(rml_cwp_next_slot2_data[0]));
INVX1 exu_U9649(.A(rml_cwp_next_slot2_data[0]), .Y(exu_n194));
AND2X1 exu_U9650(.A(rml_cwp_old_cwp_w[0]), .B(rml_cwp_n33), .Y(exu_n17578));
INVX1 exu_U9651(.A(exu_n17578), .Y(exu_n195));
AND2X1 exu_U9652(.A(exu_n10748), .B(exu_n9725), .Y(rml_cwp_next_slot3_data[9]));
INVX1 exu_U9653(.A(rml_cwp_next_slot3_data[9]), .Y(exu_n196));
AND2X1 exu_U9654(.A(exu_n10749), .B(exu_n9726), .Y(rml_cwp_next_slot3_data[8]));
INVX1 exu_U9655(.A(rml_cwp_next_slot3_data[8]), .Y(exu_n197));
AND2X1 exu_U9656(.A(exu_n15490), .B(exu_n9727), .Y(rml_cwp_next_slot3_data[7]));
INVX1 exu_U9657(.A(rml_cwp_next_slot3_data[7]), .Y(exu_n198));
AND2X1 exu_U9658(.A(exu_n10750), .B(exu_n9728), .Y(rml_cwp_next_slot3_data[6]));
INVX1 exu_U9659(.A(rml_cwp_next_slot3_data[6]), .Y(exu_n199));
AND2X1 exu_U9660(.A(exu_n17587), .B(exu_n9729), .Y(rml_cwp_next_slot3_data[5]));
INVX1 exu_U9661(.A(rml_cwp_next_slot3_data[5]), .Y(exu_n200));
AND2X1 exu_U9662(.A(rml_cwp_tlu_exu_cwp_w[2]), .B(rml_cwp_n32), .Y(exu_n17589));
INVX1 exu_U9663(.A(exu_n17589), .Y(exu_n201));
AND2X1 exu_U9664(.A(exu_n17591), .B(exu_n9730), .Y(rml_cwp_next_slot3_data[4]));
INVX1 exu_U9665(.A(rml_cwp_next_slot3_data[4]), .Y(exu_n202));
AND2X1 exu_U9666(.A(rml_cwp_tlu_exu_cwp_w[1]), .B(rml_cwp_n32), .Y(exu_n17593));
INVX1 exu_U9667(.A(exu_n17593), .Y(exu_n203));
AND2X1 exu_U9668(.A(exu_n17595), .B(exu_n9731), .Y(rml_cwp_next_slot3_data[3]));
INVX1 exu_U9669(.A(rml_cwp_next_slot3_data[3]), .Y(exu_n204));
AND2X1 exu_U9670(.A(rml_cwp_tlu_exu_cwp_w[0]), .B(rml_cwp_n32), .Y(exu_n17597));
INVX1 exu_U9671(.A(exu_n17597), .Y(exu_n205));
AND2X1 exu_U9672(.A(exu_n17599), .B(exu_n9732), .Y(rml_cwp_next_slot3_data[2]));
INVX1 exu_U9673(.A(rml_cwp_next_slot3_data[2]), .Y(exu_n206));
AND2X1 exu_U9674(.A(rml_cwp_old_cwp_w[2]), .B(rml_cwp_n32), .Y(exu_n17601));
INVX1 exu_U9675(.A(exu_n17601), .Y(exu_n207));
AND2X1 exu_U9676(.A(exu_n17603), .B(exu_n9733), .Y(rml_cwp_next_slot3_data[1]));
INVX1 exu_U9677(.A(rml_cwp_next_slot3_data[1]), .Y(exu_n208));
AND2X1 exu_U9678(.A(rml_cwp_old_cwp_w[1]), .B(rml_cwp_n32), .Y(exu_n17605));
INVX1 exu_U9679(.A(exu_n17605), .Y(exu_n209));
AND2X1 exu_U9680(.A(exu_n10751), .B(exu_n9734), .Y(rml_cwp_next_slot3_data[12]));
INVX1 exu_U9681(.A(rml_cwp_next_slot3_data[12]), .Y(exu_n210));
AND2X1 exu_U9682(.A(exu_n10752), .B(exu_n9735), .Y(rml_cwp_next_slot3_data[11]));
INVX1 exu_U9683(.A(rml_cwp_next_slot3_data[11]), .Y(exu_n211));
AND2X1 exu_U9684(.A(exu_n10753), .B(exu_n9736), .Y(rml_cwp_next_slot3_data[10]));
INVX1 exu_U9685(.A(rml_cwp_next_slot3_data[10]), .Y(exu_n212));
AND2X1 exu_U9686(.A(exu_n17613), .B(exu_n9737), .Y(rml_cwp_next_slot3_data[0]));
INVX1 exu_U9687(.A(rml_cwp_next_slot3_data[0]), .Y(exu_n213));
AND2X1 exu_U9688(.A(rml_cwp_old_cwp_w[0]), .B(rml_cwp_n32), .Y(exu_n17615));
INVX1 exu_U9689(.A(exu_n17615), .Y(exu_n214));
AND2X1 exu_U9690(.A(exu_n10754), .B(exu_n9738), .Y(ecl_divcntl_sub_next));
INVX1 exu_U9691(.A(ecl_divcntl_sub_next), .Y(exu_n215));
OR2X1 exu_U9692(.A(exu_n17634), .B(exu_n14835), .Y(exu_n17626));
INVX1 exu_U9693(.A(exu_n17626), .Y(exu_n216));
OR2X1 exu_U9694(.A(exu_n17646), .B(exu_n14837), .Y(exu_n17638));
INVX1 exu_U9695(.A(exu_n17638), .Y(exu_n217));
OR2X1 exu_U9696(.A(exu_n17658), .B(exu_n14839), .Y(exu_n17650));
INVX1 exu_U9697(.A(exu_n17650), .Y(exu_n218));
OR2X1 exu_U9698(.A(exu_n17670), .B(exu_n14841), .Y(exu_n17662));
INVX1 exu_U9699(.A(exu_n17662), .Y(exu_n219));
OR2X1 exu_U9700(.A(exu_n17682), .B(exu_n14843), .Y(exu_n17674));
INVX1 exu_U9701(.A(exu_n17674), .Y(exu_n220));
OR2X1 exu_U9702(.A(exu_n17693), .B(exu_n14845), .Y(exu_n17686));
INVX1 exu_U9703(.A(exu_n17686), .Y(exu_n221));
OR2X1 exu_U9704(.A(exu_n17704), .B(exu_n14847), .Y(exu_n17697));
INVX1 exu_U9705(.A(exu_n17697), .Y(exu_n222));
AND2X1 exu_U9706(.A(ecl_ecc_log_rs2_m), .B(ecl_ifu_exu_rs2_m[4]), .Y(exu_n17710));
INVX1 exu_U9707(.A(exu_n17710), .Y(exu_n223));
AND2X1 exu_U9708(.A(ecl_ifu_exu_rs2_m[3]), .B(ecl_ecc_log_rs2_m), .Y(exu_n17714));
INVX1 exu_U9709(.A(exu_n17714), .Y(exu_n224));
AND2X1 exu_U9710(.A(ecl_ifu_exu_rs2_m[2]), .B(ecl_ecc_log_rs2_m), .Y(exu_n17718));
INVX1 exu_U9711(.A(exu_n17718), .Y(exu_n225));
AND2X1 exu_U9712(.A(ecl_ifu_exu_rs2_m[1]), .B(ecl_ecc_log_rs2_m), .Y(exu_n17722));
INVX1 exu_U9713(.A(exu_n17722), .Y(exu_n226));
AND2X1 exu_U9714(.A(ecl_ifu_exu_rs2_m[0]), .B(ecl_ecc_log_rs2_m), .Y(exu_n17726));
INVX1 exu_U9715(.A(exu_n17726), .Y(exu_n227));
AND2X1 exu_U9716(.A(ecl_rml_thr_w[3]), .B(exu_tlu_cwp3_w[2]), .Y(exu_n17730));
INVX1 exu_U9717(.A(exu_n17730), .Y(exu_n228));
AND2X1 exu_U9718(.A(exu_n15957), .B(exu_tlu_cwp1_w[2]), .Y(exu_n17732));
INVX1 exu_U9719(.A(exu_n17732), .Y(exu_n229));
AND2X1 exu_U9720(.A(exu_tlu_cwp3_w[1]), .B(ecl_rml_thr_w[3]), .Y(exu_n17736));
INVX1 exu_U9721(.A(exu_n17736), .Y(exu_n230));
AND2X1 exu_U9722(.A(exu_tlu_cwp1_w[1]), .B(exu_n15958), .Y(exu_n17738));
INVX1 exu_U9723(.A(exu_n17738), .Y(exu_n231));
AND2X1 exu_U9724(.A(exu_tlu_cwp3_w[0]), .B(ecl_rml_thr_w[3]), .Y(exu_n17742));
INVX1 exu_U9725(.A(exu_n17742), .Y(exu_n232));
AND2X1 exu_U9726(.A(exu_tlu_cwp1_w[0]), .B(exu_n15958), .Y(exu_n17744));
INVX1 exu_U9727(.A(exu_n17744), .Y(exu_n233));
AND2X1 exu_U9728(.A(rml_thr_d[3]), .B(exu_tlu_cwp3_w[2]), .Y(exu_n17748));
INVX1 exu_U9729(.A(exu_n17748), .Y(exu_n234));
AND2X1 exu_U9730(.A(exu_n15952), .B(exu_tlu_cwp1_w[2]), .Y(exu_n17750));
INVX1 exu_U9731(.A(exu_n17750), .Y(exu_n235));
AND2X1 exu_U9732(.A(exu_tlu_cwp3_w[1]), .B(exu_n15949), .Y(exu_n17754));
INVX1 exu_U9733(.A(exu_n17754), .Y(exu_n236));
AND2X1 exu_U9734(.A(exu_tlu_cwp1_w[1]), .B(exu_n15954), .Y(exu_n17756));
INVX1 exu_U9735(.A(exu_n17756), .Y(exu_n237));
AND2X1 exu_U9736(.A(exu_tlu_cwp3_w[0]), .B(exu_n15948), .Y(exu_n17760));
INVX1 exu_U9737(.A(exu_n17760), .Y(exu_n238));
AND2X1 exu_U9738(.A(exu_tlu_cwp1_w[0]), .B(exu_n15190), .Y(exu_n17762));
INVX1 exu_U9739(.A(exu_n17762), .Y(exu_n239));
AND2X1 exu_U9740(.A(rml_cwp_thr_e[3]), .B(exu_tlu_cwp3_w[2]), .Y(exu_n17766));
INVX1 exu_U9741(.A(exu_n17766), .Y(exu_n240));
AND2X1 exu_U9742(.A(exu_n9), .B(exu_tlu_cwp1_w[2]), .Y(exu_n17768));
INVX1 exu_U9743(.A(exu_n17768), .Y(exu_n241));
AND2X1 exu_U9744(.A(exu_tlu_cwp3_w[1]), .B(rml_cwp_thr_e[3]), .Y(exu_n17772));
INVX1 exu_U9745(.A(exu_n17772), .Y(exu_n242));
AND2X1 exu_U9746(.A(exu_tlu_cwp1_w[1]), .B(exu_n9), .Y(exu_n17774));
INVX1 exu_U9747(.A(exu_n17774), .Y(exu_n243));
AND2X1 exu_U9748(.A(exu_tlu_cwp3_w[0]), .B(rml_cwp_thr_e[3]), .Y(exu_n17778));
INVX1 exu_U9749(.A(exu_n17778), .Y(exu_n244));
AND2X1 exu_U9750(.A(exu_tlu_cwp1_w[0]), .B(exu_n9), .Y(exu_n17780));
INVX1 exu_U9751(.A(exu_n17780), .Y(exu_n245));
AND2X1 exu_U9752(.A(exu_n15921), .B(exu_tlu_cwp3_w[2]), .Y(exu_n17784));
INVX1 exu_U9753(.A(exu_n17784), .Y(exu_n246));
AND2X1 exu_U9754(.A(exu_n15923), .B(exu_tlu_cwp1_w[2]), .Y(exu_n17786));
INVX1 exu_U9755(.A(exu_n17786), .Y(exu_n247));
AND2X1 exu_U9756(.A(exu_tlu_cwp3_w[1]), .B(exu_n15921), .Y(exu_n17790));
INVX1 exu_U9757(.A(exu_n17790), .Y(exu_n248));
AND2X1 exu_U9758(.A(exu_tlu_cwp1_w[1]), .B(exu_n15923), .Y(exu_n17792));
INVX1 exu_U9759(.A(exu_n17792), .Y(exu_n249));
AND2X1 exu_U9760(.A(exu_tlu_cwp3_w[0]), .B(exu_n15921), .Y(exu_n17796));
INVX1 exu_U9761(.A(exu_n17796), .Y(exu_n250));
AND2X1 exu_U9762(.A(exu_tlu_cwp1_w[0]), .B(exu_n15923), .Y(exu_n17798));
INVX1 exu_U9763(.A(exu_n17798), .Y(exu_n251));
AND2X1 exu_U9764(.A(rml_cwp_n88), .B(rml_cwp_new_swap_cwp[2]), .Y(exu_n17802));
INVX1 exu_U9765(.A(exu_n17802), .Y(exu_n252));
AND2X1 exu_U9766(.A(rml_cwp_n89), .B(rml_next_cwp_noreset_w[2]), .Y(exu_n17804));
INVX1 exu_U9767(.A(exu_n17804), .Y(exu_n253));
AND2X1 exu_U9768(.A(rml_cwp_new_swap_cwp[1]), .B(rml_cwp_n88), .Y(exu_n17808));
INVX1 exu_U9769(.A(exu_n17808), .Y(exu_n254));
AND2X1 exu_U9770(.A(rml_next_cwp_noreset_w[1]), .B(rml_cwp_n89), .Y(exu_n17810));
INVX1 exu_U9771(.A(exu_n17810), .Y(exu_n255));
AND2X1 exu_U9772(.A(rml_cwp_new_swap_cwp[0]), .B(rml_cwp_n88), .Y(exu_n17814));
INVX1 exu_U9773(.A(exu_n17814), .Y(exu_n256));
AND2X1 exu_U9774(.A(rml_next_cwp_noreset_w[0]), .B(rml_cwp_n89), .Y(exu_n17816));
INVX1 exu_U9775(.A(exu_n17816), .Y(exu_n257));
AND2X1 exu_U9776(.A(rml_cwp_n85), .B(rml_cwp_new_swap_cwp[2]), .Y(exu_n17820));
INVX1 exu_U9777(.A(exu_n17820), .Y(exu_n258));
AND2X1 exu_U9778(.A(rml_cwp_n86), .B(rml_next_cwp_noreset_w[2]), .Y(exu_n17822));
INVX1 exu_U9779(.A(exu_n17822), .Y(exu_n259));
AND2X1 exu_U9780(.A(rml_cwp_new_swap_cwp[1]), .B(rml_cwp_n85), .Y(exu_n17826));
INVX1 exu_U9781(.A(exu_n17826), .Y(exu_n260));
AND2X1 exu_U9782(.A(rml_next_cwp_noreset_w[1]), .B(rml_cwp_n86), .Y(exu_n17828));
INVX1 exu_U9783(.A(exu_n17828), .Y(exu_n261));
AND2X1 exu_U9784(.A(rml_cwp_new_swap_cwp[0]), .B(rml_cwp_n85), .Y(exu_n17832));
INVX1 exu_U9785(.A(exu_n17832), .Y(exu_n262));
AND2X1 exu_U9786(.A(rml_next_cwp_noreset_w[0]), .B(rml_cwp_n86), .Y(exu_n17834));
INVX1 exu_U9787(.A(exu_n17834), .Y(exu_n263));
AND2X1 exu_U9788(.A(rml_cwp_n82), .B(rml_cwp_new_swap_cwp[2]), .Y(exu_n17838));
INVX1 exu_U9789(.A(exu_n17838), .Y(exu_n264));
AND2X1 exu_U9790(.A(rml_cwp_n83), .B(rml_next_cwp_noreset_w[2]), .Y(exu_n17840));
INVX1 exu_U9791(.A(exu_n17840), .Y(exu_n265));
AND2X1 exu_U9792(.A(rml_cwp_new_swap_cwp[1]), .B(rml_cwp_n82), .Y(exu_n17844));
INVX1 exu_U9793(.A(exu_n17844), .Y(exu_n266));
AND2X1 exu_U9794(.A(rml_next_cwp_noreset_w[1]), .B(rml_cwp_n83), .Y(exu_n17846));
INVX1 exu_U9795(.A(exu_n17846), .Y(exu_n267));
AND2X1 exu_U9796(.A(rml_cwp_new_swap_cwp[0]), .B(rml_cwp_n82), .Y(exu_n17850));
INVX1 exu_U9797(.A(exu_n17850), .Y(exu_n268));
AND2X1 exu_U9798(.A(rml_next_cwp_noreset_w[0]), .B(rml_cwp_n83), .Y(exu_n17852));
INVX1 exu_U9799(.A(exu_n17852), .Y(exu_n269));
AND2X1 exu_U9800(.A(rml_cwp_n79), .B(rml_cwp_new_swap_cwp[2]), .Y(exu_n17856));
INVX1 exu_U9801(.A(exu_n17856), .Y(exu_n270));
AND2X1 exu_U9802(.A(rml_cwp_n80), .B(rml_next_cwp_noreset_w[2]), .Y(exu_n17858));
INVX1 exu_U9803(.A(exu_n17858), .Y(exu_n271));
AND2X1 exu_U9804(.A(rml_cwp_new_swap_cwp[1]), .B(rml_cwp_n79), .Y(exu_n17862));
INVX1 exu_U9805(.A(exu_n17862), .Y(exu_n272));
AND2X1 exu_U9806(.A(rml_next_cwp_noreset_w[1]), .B(rml_cwp_n80), .Y(exu_n17864));
INVX1 exu_U9807(.A(exu_n17864), .Y(exu_n273));
AND2X1 exu_U9808(.A(rml_cwp_new_swap_cwp[0]), .B(rml_cwp_n79), .Y(exu_n17868));
INVX1 exu_U9809(.A(exu_n17868), .Y(exu_n274));
AND2X1 exu_U9810(.A(rml_next_cwp_noreset_w[0]), .B(rml_cwp_n80), .Y(exu_n17870));
INVX1 exu_U9811(.A(exu_n17870), .Y(exu_n275));
AND2X1 exu_U9812(.A(exu_n15948), .B(rml_cansave_reg_data_thr3[2]), .Y(exu_n17874));
INVX1 exu_U9813(.A(exu_n17874), .Y(exu_n276));
AND2X1 exu_U9814(.A(exu_n15953), .B(rml_cansave_reg_data_thr1[2]), .Y(exu_n17876));
INVX1 exu_U9815(.A(exu_n17876), .Y(exu_n277));
AND2X1 exu_U9816(.A(rml_cansave_reg_data_thr3[1]), .B(exu_n15948), .Y(exu_n17880));
INVX1 exu_U9817(.A(exu_n17880), .Y(exu_n278));
AND2X1 exu_U9818(.A(rml_cansave_reg_data_thr1[1]), .B(exu_n15954), .Y(exu_n17882));
INVX1 exu_U9819(.A(exu_n17882), .Y(exu_n279));
AND2X1 exu_U9820(.A(rml_cansave_reg_data_thr3[0]), .B(rml_thr_d[3]), .Y(exu_n17886));
INVX1 exu_U9821(.A(exu_n17886), .Y(exu_n280));
AND2X1 exu_U9822(.A(rml_cansave_reg_data_thr1[0]), .B(exu_n15952), .Y(exu_n17888));
INVX1 exu_U9823(.A(exu_n17888), .Y(exu_n281));
AND2X1 exu_U9824(.A(exu_n15949), .B(rml_canrestore_reg_data_thr3[2]), .Y(exu_n17892));
INVX1 exu_U9825(.A(exu_n17892), .Y(exu_n282));
AND2X1 exu_U9826(.A(exu_n15954), .B(rml_canrestore_reg_data_thr1[2]), .Y(exu_n17894));
INVX1 exu_U9827(.A(exu_n17894), .Y(exu_n283));
AND2X1 exu_U9828(.A(rml_canrestore_reg_data_thr3[1]), .B(rml_thr_d[3]), .Y(exu_n17898));
INVX1 exu_U9829(.A(exu_n17898), .Y(exu_n284));
AND2X1 exu_U9830(.A(rml_canrestore_reg_data_thr1[1]), .B(exu_n15953), .Y(exu_n17900));
INVX1 exu_U9831(.A(exu_n17900), .Y(exu_n285));
AND2X1 exu_U9832(.A(rml_canrestore_reg_data_thr3[0]), .B(exu_n15949), .Y(exu_n17904));
INVX1 exu_U9833(.A(exu_n17904), .Y(exu_n286));
AND2X1 exu_U9834(.A(rml_canrestore_reg_data_thr1[0]), .B(exu_n15954), .Y(exu_n17906));
INVX1 exu_U9835(.A(exu_n17906), .Y(exu_n287));
AND2X1 exu_U9836(.A(rml_thr_d[3]), .B(rml_otherwin_reg_data_thr3[2]), .Y(exu_n17910));
INVX1 exu_U9837(.A(exu_n17910), .Y(exu_n288));
AND2X1 exu_U9838(.A(exu_n15190), .B(rml_otherwin_reg_data_thr1[2]), .Y(exu_n17912));
INVX1 exu_U9839(.A(exu_n17912), .Y(exu_n289));
AND2X1 exu_U9840(.A(rml_otherwin_reg_data_thr3[1]), .B(exu_n15949), .Y(exu_n17916));
INVX1 exu_U9841(.A(exu_n17916), .Y(exu_n290));
AND2X1 exu_U9842(.A(rml_otherwin_reg_data_thr1[1]), .B(exu_n15952), .Y(exu_n17918));
INVX1 exu_U9843(.A(exu_n17918), .Y(exu_n291));
AND2X1 exu_U9844(.A(rml_otherwin_reg_data_thr3[0]), .B(exu_n15948), .Y(exu_n17922));
INVX1 exu_U9845(.A(exu_n17922), .Y(exu_n292));
AND2X1 exu_U9846(.A(rml_otherwin_reg_data_thr1[0]), .B(exu_n15953), .Y(exu_n17924));
INVX1 exu_U9847(.A(exu_n17924), .Y(exu_n293));
AND2X1 exu_U9848(.A(exu_n15948), .B(rml_cleanwin_reg_data_thr3[2]), .Y(exu_n17928));
INVX1 exu_U9849(.A(exu_n17928), .Y(exu_n294));
AND2X1 exu_U9850(.A(exu_n15190), .B(rml_cleanwin_reg_data_thr1[2]), .Y(exu_n17930));
INVX1 exu_U9851(.A(exu_n17930), .Y(exu_n295));
AND2X1 exu_U9852(.A(rml_cleanwin_reg_data_thr3[1]), .B(exu_n15948), .Y(exu_n17934));
INVX1 exu_U9853(.A(exu_n17934), .Y(exu_n296));
AND2X1 exu_U9854(.A(rml_cleanwin_reg_data_thr1[1]), .B(exu_n15190), .Y(exu_n17936));
INVX1 exu_U9855(.A(exu_n17936), .Y(exu_n297));
AND2X1 exu_U9856(.A(rml_cleanwin_reg_data_thr3[0]), .B(rml_thr_d[3]), .Y(exu_n17940));
INVX1 exu_U9857(.A(exu_n17940), .Y(exu_n298));
AND2X1 exu_U9858(.A(rml_cleanwin_reg_data_thr1[0]), .B(exu_n15952), .Y(exu_n17942));
INVX1 exu_U9859(.A(exu_n17942), .Y(exu_n299));
AND2X1 exu_U9860(.A(exu_n15949), .B(rml_hi_wstate_reg_data_thr3[2]), .Y(exu_n17946));
INVX1 exu_U9861(.A(exu_n17946), .Y(exu_n300));
AND2X1 exu_U9862(.A(exu_n15952), .B(rml_hi_wstate_reg_data_thr1[2]), .Y(exu_n17948));
INVX1 exu_U9863(.A(exu_n17948), .Y(exu_n301));
AND2X1 exu_U9864(.A(rml_hi_wstate_reg_data_thr3[1]), .B(rml_thr_d[3]), .Y(exu_n17952));
INVX1 exu_U9865(.A(exu_n17952), .Y(exu_n302));
AND2X1 exu_U9866(.A(rml_hi_wstate_reg_data_thr1[1]), .B(exu_n15953), .Y(exu_n17954));
INVX1 exu_U9867(.A(exu_n17954), .Y(exu_n303));
AND2X1 exu_U9868(.A(rml_hi_wstate_reg_data_thr3[0]), .B(exu_n15949), .Y(exu_n17958));
INVX1 exu_U9869(.A(exu_n17958), .Y(exu_n304));
AND2X1 exu_U9870(.A(rml_hi_wstate_reg_data_thr1[0]), .B(exu_n15954), .Y(exu_n17960));
INVX1 exu_U9871(.A(exu_n17960), .Y(exu_n305));
AND2X1 exu_U9872(.A(rml_thr_d[3]), .B(rml_lo_wstate_reg_data_thr3[2]), .Y(exu_n17964));
INVX1 exu_U9873(.A(exu_n17964), .Y(exu_n306));
AND2X1 exu_U9874(.A(exu_n15953), .B(rml_lo_wstate_reg_data_thr1[2]), .Y(exu_n17966));
INVX1 exu_U9875(.A(exu_n17966), .Y(exu_n307));
AND2X1 exu_U9876(.A(rml_lo_wstate_reg_data_thr3[1]), .B(exu_n15949), .Y(exu_n17970));
INVX1 exu_U9877(.A(exu_n17970), .Y(exu_n308));
AND2X1 exu_U9878(.A(rml_lo_wstate_reg_data_thr1[1]), .B(exu_n15190), .Y(exu_n17972));
INVX1 exu_U9879(.A(exu_n17972), .Y(exu_n309));
AND2X1 exu_U9880(.A(rml_lo_wstate_reg_data_thr3[0]), .B(exu_n15948), .Y(exu_n17976));
INVX1 exu_U9881(.A(exu_n17976), .Y(exu_n310));
AND2X1 exu_U9882(.A(rml_lo_wstate_reg_data_thr1[0]), .B(exu_n15953), .Y(exu_n17978));
INVX1 exu_U9883(.A(exu_n17978), .Y(exu_n311));
AND2X1 exu_U9884(.A(ecl_writeback_n130), .B(ecl_writeback_restore_rd[4]), .Y(exu_n17983));
INVX1 exu_U9885(.A(exu_n17983), .Y(exu_n312));
AND2X1 exu_U9886(.A(ecl_writeback_n167), .B(ecl_wb_byplog_rd_g2[4]), .Y(exu_n17985));
INVX1 exu_U9887(.A(exu_n17985), .Y(exu_n313));
AND2X1 exu_U9888(.A(ecl_writeback_restore_rd[3]), .B(ecl_writeback_n130), .Y(exu_n17989));
INVX1 exu_U9889(.A(exu_n17989), .Y(exu_n314));
AND2X1 exu_U9890(.A(ecl_wb_byplog_rd_g2[3]), .B(ecl_writeback_n167), .Y(exu_n17991));
INVX1 exu_U9891(.A(exu_n17991), .Y(exu_n315));
AND2X1 exu_U9892(.A(ecl_writeback_restore_rd[2]), .B(exu_n15989), .Y(exu_n17995));
INVX1 exu_U9893(.A(exu_n17995), .Y(exu_n316));
AND2X1 exu_U9894(.A(ecl_wb_byplog_rd_g2[2]), .B(exu_n15764), .Y(exu_n17997));
INVX1 exu_U9895(.A(exu_n17997), .Y(exu_n317));
AND2X1 exu_U9896(.A(ecl_writeback_restore_rd[1]), .B(ecl_writeback_n130), .Y(exu_n18001));
INVX1 exu_U9897(.A(exu_n18001), .Y(exu_n318));
AND2X1 exu_U9898(.A(ecl_wb_byplog_rd_g2[1]), .B(ecl_writeback_n167), .Y(exu_n18003));
INVX1 exu_U9899(.A(exu_n18003), .Y(exu_n319));
AND2X1 exu_U9900(.A(ecl_writeback_restore_rd[0]), .B(exu_n15989), .Y(exu_n18007));
INVX1 exu_U9901(.A(exu_n18007), .Y(exu_n320));
AND2X1 exu_U9902(.A(ecl_wb_byplog_rd_g2[0]), .B(ecl_writeback_n167), .Y(exu_n18009));
INVX1 exu_U9903(.A(exu_n18009), .Y(exu_n321));
AND2X1 exu_U9904(.A(ecl_writeback_rdpr_mux1_out[2]), .B(ecl_writeback_rdpr_mux2_sel3), .Y(exu_n18021));
INVX1 exu_U9905(.A(exu_n18021), .Y(exu_n322));
AND2X1 exu_U9906(.A(rml_ecl_cwp_d[2]), .B(exu_n15427), .Y(exu_n18023));
INVX1 exu_U9907(.A(exu_n18023), .Y(exu_n323));
AND2X1 exu_U9908(.A(ecl_writeback_rdpr_mux1_out[1]), .B(ecl_writeback_rdpr_mux2_sel3), .Y(exu_n18027));
INVX1 exu_U9909(.A(exu_n18027), .Y(exu_n324));
AND2X1 exu_U9910(.A(rml_ecl_cwp_d[1]), .B(exu_n15427), .Y(exu_n18029));
INVX1 exu_U9911(.A(exu_n18029), .Y(exu_n325));
AND2X1 exu_U9912(.A(ecl_writeback_rdpr_mux1_out[0]), .B(ecl_writeback_rdpr_mux2_sel3), .Y(exu_n18033));
INVX1 exu_U9913(.A(exu_n18033), .Y(exu_n326));
AND2X1 exu_U9914(.A(rml_ecl_cwp_d[0]), .B(exu_n15427), .Y(exu_n18035));
INVX1 exu_U9915(.A(exu_n18035), .Y(exu_n327));
AND2X1 exu_U9916(.A(exu_n18037), .B(exu_n9742), .Y(ecl_ccr_ccrin_thr1[7]));
INVX1 exu_U9917(.A(ecl_ccr_ccrin_thr1[7]), .Y(exu_n328));
AND2X1 exu_U9918(.A(ecl_ccr_n17), .B(ecl_divcntl_ccr_cc_w2[7]), .Y(exu_n18039));
INVX1 exu_U9919(.A(exu_n18039), .Y(exu_n329));
AND2X1 exu_U9920(.A(exu_n18041), .B(exu_n9743), .Y(ecl_ccr_ccrin_thr1[6]));
INVX1 exu_U9921(.A(ecl_ccr_ccrin_thr1[6]), .Y(exu_n330));
AND2X1 exu_U9922(.A(ecl_divcntl_ccr_cc_w2[6]), .B(ecl_ccr_n17), .Y(exu_n18043));
INVX1 exu_U9923(.A(exu_n18043), .Y(exu_n331));
AND2X1 exu_U9924(.A(exu_n10755), .B(exu_n9744), .Y(ecl_ccr_ccrin_thr1[5]));
INVX1 exu_U9925(.A(ecl_ccr_ccrin_thr1[5]), .Y(exu_n332));
AND2X1 exu_U9926(.A(exu_n10756), .B(exu_n9745), .Y(ecl_ccr_ccrin_thr1[4]));
INVX1 exu_U9927(.A(ecl_ccr_ccrin_thr1[4]), .Y(exu_n333));
AND2X1 exu_U9928(.A(exu_n18049), .B(exu_n9746), .Y(ecl_ccr_ccrin_thr1[3]));
INVX1 exu_U9929(.A(ecl_ccr_ccrin_thr1[3]), .Y(exu_n334));
AND2X1 exu_U9930(.A(exu_n15736), .B(ecl_ccr_n17), .Y(exu_n18051));
INVX1 exu_U9931(.A(exu_n18051), .Y(exu_n335));
AND2X1 exu_U9932(.A(exu_n18053), .B(exu_n9747), .Y(ecl_ccr_ccrin_thr1[2]));
INVX1 exu_U9933(.A(ecl_ccr_ccrin_thr1[2]), .Y(exu_n336));
AND2X1 exu_U9934(.A(exu_n15737), .B(ecl_ccr_n17), .Y(exu_n18055));
INVX1 exu_U9935(.A(exu_n18055), .Y(exu_n337));
AND2X1 exu_U9936(.A(exu_n18057), .B(exu_n9748), .Y(ecl_ccr_ccrin_thr1[1]));
INVX1 exu_U9937(.A(ecl_ccr_ccrin_thr1[1]), .Y(exu_n338));
AND2X1 exu_U9938(.A(exu_n15738), .B(ecl_ccr_n17), .Y(exu_n18059));
INVX1 exu_U9939(.A(exu_n18059), .Y(exu_n339));
AND2X1 exu_U9940(.A(exu_n18061), .B(exu_n9749), .Y(ecl_ccr_ccrin_thr1[0]));
INVX1 exu_U9941(.A(ecl_ccr_ccrin_thr1[0]), .Y(exu_n340));
AND2X1 exu_U9942(.A(ecl_divcntl_ccr_cc_w2[0]), .B(ecl_ccr_n17), .Y(exu_n18063));
INVX1 exu_U9943(.A(exu_n18063), .Y(exu_n341));
AND2X1 exu_U9944(.A(exu_n18065), .B(exu_n9750), .Y(ecl_ccr_ccrin_thr2[7]));
INVX1 exu_U9945(.A(ecl_ccr_ccrin_thr2[7]), .Y(exu_n342));
AND2X1 exu_U9946(.A(ecl_ccr_n15), .B(ecl_divcntl_ccr_cc_w2[7]), .Y(exu_n18067));
INVX1 exu_U9947(.A(exu_n18067), .Y(exu_n343));
AND2X1 exu_U9948(.A(exu_n18069), .B(exu_n9751), .Y(ecl_ccr_ccrin_thr2[6]));
INVX1 exu_U9949(.A(ecl_ccr_ccrin_thr2[6]), .Y(exu_n344));
AND2X1 exu_U9950(.A(ecl_divcntl_ccr_cc_w2[6]), .B(ecl_ccr_n15), .Y(exu_n18071));
INVX1 exu_U9951(.A(exu_n18071), .Y(exu_n345));
AND2X1 exu_U9952(.A(exu_n10757), .B(exu_n9752), .Y(ecl_ccr_ccrin_thr2[5]));
INVX1 exu_U9953(.A(ecl_ccr_ccrin_thr2[5]), .Y(exu_n346));
AND2X1 exu_U9954(.A(exu_n10758), .B(exu_n9753), .Y(ecl_ccr_ccrin_thr2[4]));
INVX1 exu_U9955(.A(ecl_ccr_ccrin_thr2[4]), .Y(exu_n347));
AND2X1 exu_U9956(.A(exu_n18077), .B(exu_n9754), .Y(ecl_ccr_ccrin_thr2[3]));
INVX1 exu_U9957(.A(ecl_ccr_ccrin_thr2[3]), .Y(exu_n348));
AND2X1 exu_U9958(.A(exu_n15736), .B(ecl_ccr_n15), .Y(exu_n18079));
INVX1 exu_U9959(.A(exu_n18079), .Y(exu_n349));
AND2X1 exu_U9960(.A(exu_n18081), .B(exu_n9755), .Y(ecl_ccr_ccrin_thr2[2]));
INVX1 exu_U9961(.A(ecl_ccr_ccrin_thr2[2]), .Y(exu_n350));
AND2X1 exu_U9962(.A(exu_n15737), .B(ecl_ccr_n15), .Y(exu_n18083));
INVX1 exu_U9963(.A(exu_n18083), .Y(exu_n351));
AND2X1 exu_U9964(.A(exu_n18085), .B(exu_n9756), .Y(ecl_ccr_ccrin_thr2[1]));
INVX1 exu_U9965(.A(ecl_ccr_ccrin_thr2[1]), .Y(exu_n352));
AND2X1 exu_U9966(.A(exu_n15738), .B(ecl_ccr_n15), .Y(exu_n18087));
INVX1 exu_U9967(.A(exu_n18087), .Y(exu_n353));
AND2X1 exu_U9968(.A(exu_n18089), .B(exu_n9757), .Y(ecl_ccr_ccrin_thr2[0]));
INVX1 exu_U9969(.A(ecl_ccr_ccrin_thr2[0]), .Y(exu_n354));
AND2X1 exu_U9970(.A(ecl_divcntl_ccr_cc_w2[0]), .B(ecl_ccr_n15), .Y(exu_n18091));
INVX1 exu_U9971(.A(exu_n18091), .Y(exu_n355));
AND2X1 exu_U9972(.A(exu_n18093), .B(exu_n9758), .Y(ecl_ccr_ccrin_thr3[7]));
INVX1 exu_U9973(.A(ecl_ccr_ccrin_thr3[7]), .Y(exu_n356));
AND2X1 exu_U9974(.A(ecl_ccr_n12), .B(ecl_divcntl_ccr_cc_w2[7]), .Y(exu_n18095));
INVX1 exu_U9975(.A(exu_n18095), .Y(exu_n357));
AND2X1 exu_U9976(.A(exu_n18097), .B(exu_n9759), .Y(ecl_ccr_ccrin_thr3[6]));
INVX1 exu_U9977(.A(ecl_ccr_ccrin_thr3[6]), .Y(exu_n358));
AND2X1 exu_U9978(.A(ecl_divcntl_ccr_cc_w2[6]), .B(ecl_ccr_n12), .Y(exu_n18099));
INVX1 exu_U9979(.A(exu_n18099), .Y(exu_n359));
AND2X1 exu_U9980(.A(exu_n10759), .B(exu_n9760), .Y(ecl_ccr_ccrin_thr3[5]));
INVX1 exu_U9981(.A(ecl_ccr_ccrin_thr3[5]), .Y(exu_n360));
AND2X1 exu_U9982(.A(exu_n10760), .B(exu_n9761), .Y(ecl_ccr_ccrin_thr3[4]));
INVX1 exu_U9983(.A(ecl_ccr_ccrin_thr3[4]), .Y(exu_n361));
AND2X1 exu_U9984(.A(exu_n18105), .B(exu_n9762), .Y(ecl_ccr_ccrin_thr3[3]));
INVX1 exu_U9985(.A(ecl_ccr_ccrin_thr3[3]), .Y(exu_n362));
AND2X1 exu_U9986(.A(exu_n15736), .B(ecl_ccr_n12), .Y(exu_n18107));
INVX1 exu_U9987(.A(exu_n18107), .Y(exu_n363));
AND2X1 exu_U9988(.A(exu_n18109), .B(exu_n9763), .Y(ecl_ccr_ccrin_thr3[2]));
INVX1 exu_U9989(.A(ecl_ccr_ccrin_thr3[2]), .Y(exu_n364));
AND2X1 exu_U9990(.A(exu_n15737), .B(ecl_ccr_n12), .Y(exu_n18111));
INVX1 exu_U9991(.A(exu_n18111), .Y(exu_n365));
AND2X1 exu_U9992(.A(exu_n18113), .B(exu_n9764), .Y(ecl_ccr_ccrin_thr3[1]));
INVX1 exu_U9993(.A(ecl_ccr_ccrin_thr3[1]), .Y(exu_n366));
AND2X1 exu_U9994(.A(exu_n15738), .B(ecl_ccr_n12), .Y(exu_n18115));
INVX1 exu_U9995(.A(exu_n18115), .Y(exu_n367));
AND2X1 exu_U9996(.A(exu_n18117), .B(exu_n9765), .Y(ecl_ccr_ccrin_thr3[0]));
INVX1 exu_U9997(.A(ecl_ccr_ccrin_thr3[0]), .Y(exu_n368));
AND2X1 exu_U9998(.A(ecl_divcntl_ccr_cc_w2[0]), .B(ecl_ccr_n12), .Y(exu_n18119));
INVX1 exu_U9999(.A(exu_n18119), .Y(exu_n369));
AND2X1 exu_U10000(.A(ecl_ccr_n24), .B(ecl_ccr_alu_cc_m[7]), .Y(exu_n18123));
INVX1 exu_U10001(.A(exu_n18123), .Y(exu_n370));
AND2X1 exu_U10002(.A(ecl_ccr_alu_cc_m[6]), .B(ecl_ccr_n24), .Y(exu_n18127));
INVX1 exu_U10003(.A(exu_n18127), .Y(exu_n371));
AND2X1 exu_U10004(.A(ecl_ccr_alu_cc_m[5]), .B(ecl_ccr_n24), .Y(exu_n18131));
INVX1 exu_U10005(.A(exu_n18131), .Y(exu_n372));
AND2X1 exu_U10006(.A(ecl_ccr_alu_cc_m[4]), .B(ecl_ccr_n24), .Y(exu_n18135));
INVX1 exu_U10007(.A(exu_n18135), .Y(exu_n373));
AND2X1 exu_U10008(.A(ecl_ccr_alu_cc_m[3]), .B(ecl_ccr_n24), .Y(exu_n18139));
INVX1 exu_U10009(.A(exu_n18139), .Y(exu_n374));
AND2X1 exu_U10010(.A(ecl_ccr_alu_cc_m[2]), .B(ecl_ccr_n24), .Y(exu_n18143));
INVX1 exu_U10011(.A(exu_n18143), .Y(exu_n375));
AND2X1 exu_U10012(.A(ecl_ccr_alu_cc_m[1]), .B(ecl_ccr_n24), .Y(exu_n18147));
INVX1 exu_U10013(.A(exu_n18147), .Y(exu_n376));
AND2X1 exu_U10014(.A(ecl_ccr_alu_cc_m[0]), .B(ecl_ccr_n24), .Y(exu_n18151));
INVX1 exu_U10015(.A(exu_n18151), .Y(exu_n377));
AND2X1 exu_U10016(.A(ecl_ccr_alu_cc_w[0]), .B(ecl_wb_ccr_wrccr_w), .Y(exu_n18153));
INVX1 exu_U10017(.A(exu_n18153), .Y(exu_n378));
AND2X1 exu_U10018(.A(ecl_ccr_alu_cc_w[1]), .B(ecl_wb_ccr_wrccr_w), .Y(exu_n18155));
INVX1 exu_U10019(.A(exu_n18155), .Y(exu_n379));
AND2X1 exu_U10020(.A(ecl_ccr_alu_cc_w[2]), .B(ecl_wb_ccr_wrccr_w), .Y(exu_n18157));
INVX1 exu_U10021(.A(exu_n18157), .Y(exu_n380));
AND2X1 exu_U10022(.A(ecl_ccr_alu_cc_w[3]), .B(ecl_wb_ccr_wrccr_w), .Y(exu_n18159));
INVX1 exu_U10023(.A(exu_n18159), .Y(exu_n381));
AND2X1 exu_U10024(.A(ecl_ccr_alu_cc_w[4]), .B(ecl_wb_ccr_wrccr_w), .Y(exu_n18161));
INVX1 exu_U10025(.A(exu_n18161), .Y(exu_n382));
AND2X1 exu_U10026(.A(ecl_ccr_alu_cc_w[5]), .B(ecl_wb_ccr_wrccr_w), .Y(exu_n18163));
INVX1 exu_U10027(.A(exu_n18163), .Y(exu_n383));
AND2X1 exu_U10028(.A(ecl_ccr_alu_cc_w[6]), .B(ecl_wb_ccr_wrccr_w), .Y(exu_n18165));
INVX1 exu_U10029(.A(exu_n18165), .Y(exu_n384));
AND2X1 exu_U10030(.A(ecl_ccr_alu_cc_w[7]), .B(ecl_wb_ccr_wrccr_w), .Y(exu_n18167));
INVX1 exu_U10031(.A(exu_n18167), .Y(exu_n385));
AND2X1 exu_U10032(.A(exu_n10769), .B(exu_n9766), .Y(rml_agp_thr1_next[0]));
INVX1 exu_U10033(.A(rml_agp_thr1_next[0]), .Y(exu_n386));
AND2X1 exu_U10034(.A(exu_n10770), .B(exu_n9767), .Y(rml_agp_thr1_next[1]));
INVX1 exu_U10035(.A(rml_agp_thr1_next[1]), .Y(exu_n387));
AND2X1 exu_U10036(.A(exu_n10771), .B(exu_n9768), .Y(rml_agp_thr2_next[0]));
INVX1 exu_U10037(.A(rml_agp_thr2_next[0]), .Y(exu_n388));
AND2X1 exu_U10038(.A(exu_n10772), .B(exu_n9769), .Y(rml_agp_thr2_next[1]));
INVX1 exu_U10039(.A(rml_agp_thr2_next[1]), .Y(exu_n389));
AND2X1 exu_U10040(.A(exu_n10773), .B(exu_n9770), .Y(rml_agp_thr3_next[0]));
INVX1 exu_U10041(.A(rml_agp_thr3_next[0]), .Y(exu_n390));
AND2X1 exu_U10042(.A(exu_n10774), .B(exu_n9771), .Y(rml_agp_thr3_next[1]));
INVX1 exu_U10043(.A(rml_agp_thr3_next[1]), .Y(exu_n391));
AND2X1 exu_U10044(.A(exu_n10784), .B(exu_n9776), .Y(rml_canrestore_reg_data_thr3_next[2]));
INVX1 exu_U10045(.A(rml_canrestore_reg_data_thr3_next[2]), .Y(exu_n392));
AND2X1 exu_U10046(.A(exu_n10785), .B(exu_n9777), .Y(rml_canrestore_reg_data_thr3_next[1]));
INVX1 exu_U10047(.A(rml_canrestore_reg_data_thr3_next[1]), .Y(exu_n393));
AND2X1 exu_U10048(.A(exu_n10786), .B(exu_n9778), .Y(rml_canrestore_reg_data_thr3_next[0]));
INVX1 exu_U10049(.A(rml_canrestore_reg_data_thr3_next[0]), .Y(exu_n394));
AND2X1 exu_U10050(.A(exu_n10787), .B(exu_n9779), .Y(rml_canrestore_reg_data_thr2_next[2]));
INVX1 exu_U10051(.A(rml_canrestore_reg_data_thr2_next[2]), .Y(exu_n395));
AND2X1 exu_U10052(.A(exu_n10788), .B(exu_n9780), .Y(rml_canrestore_reg_data_thr2_next[1]));
INVX1 exu_U10053(.A(rml_canrestore_reg_data_thr2_next[1]), .Y(exu_n396));
AND2X1 exu_U10054(.A(exu_n10789), .B(exu_n9781), .Y(rml_canrestore_reg_data_thr2_next[0]));
INVX1 exu_U10055(.A(rml_canrestore_reg_data_thr2_next[0]), .Y(exu_n397));
AND2X1 exu_U10056(.A(exu_n10790), .B(exu_n9782), .Y(rml_canrestore_reg_data_thr1_next[2]));
INVX1 exu_U10057(.A(rml_canrestore_reg_data_thr1_next[2]), .Y(exu_n398));
AND2X1 exu_U10058(.A(exu_n10791), .B(exu_n9783), .Y(rml_canrestore_reg_data_thr1_next[1]));
INVX1 exu_U10059(.A(rml_canrestore_reg_data_thr1_next[1]), .Y(exu_n399));
AND2X1 exu_U10060(.A(exu_n10792), .B(exu_n9784), .Y(rml_canrestore_reg_data_thr1_next[0]));
INVX1 exu_U10061(.A(rml_canrestore_reg_data_thr1_next[0]), .Y(exu_n400));
AND2X1 exu_U10062(.A(exu_n10793), .B(exu_n9785), .Y(rml_canrestore_reg_data_thr0_next[2]));
INVX1 exu_U10063(.A(rml_canrestore_reg_data_thr0_next[2]), .Y(exu_n401));
AND2X1 exu_U10064(.A(exu_n10794), .B(exu_n9786), .Y(rml_canrestore_reg_data_thr0_next[1]));
INVX1 exu_U10065(.A(rml_canrestore_reg_data_thr0_next[1]), .Y(exu_n402));
AND2X1 exu_U10066(.A(exu_n10795), .B(exu_n9787), .Y(rml_canrestore_reg_data_thr0_next[0]));
INVX1 exu_U10067(.A(rml_canrestore_reg_data_thr0_next[0]), .Y(exu_n403));
AND2X1 exu_U10068(.A(exu_n10796), .B(exu_n9788), .Y(rml_otherwin_reg_data_thr3_next[2]));
INVX1 exu_U10069(.A(rml_otherwin_reg_data_thr3_next[2]), .Y(exu_n404));
AND2X1 exu_U10070(.A(exu_n10797), .B(exu_n9789), .Y(rml_otherwin_reg_data_thr3_next[1]));
INVX1 exu_U10071(.A(rml_otherwin_reg_data_thr3_next[1]), .Y(exu_n405));
AND2X1 exu_U10072(.A(exu_n10798), .B(exu_n9790), .Y(rml_otherwin_reg_data_thr3_next[0]));
INVX1 exu_U10073(.A(rml_otherwin_reg_data_thr3_next[0]), .Y(exu_n406));
AND2X1 exu_U10074(.A(exu_n10799), .B(exu_n9791), .Y(rml_otherwin_reg_data_thr2_next[2]));
INVX1 exu_U10075(.A(rml_otherwin_reg_data_thr2_next[2]), .Y(exu_n407));
AND2X1 exu_U10076(.A(exu_n10800), .B(exu_n9792), .Y(rml_otherwin_reg_data_thr2_next[1]));
INVX1 exu_U10077(.A(rml_otherwin_reg_data_thr2_next[1]), .Y(exu_n408));
AND2X1 exu_U10078(.A(exu_n10801), .B(exu_n9793), .Y(rml_otherwin_reg_data_thr2_next[0]));
INVX1 exu_U10079(.A(rml_otherwin_reg_data_thr2_next[0]), .Y(exu_n409));
AND2X1 exu_U10080(.A(exu_n10802), .B(exu_n9794), .Y(rml_otherwin_reg_data_thr1_next[2]));
INVX1 exu_U10081(.A(rml_otherwin_reg_data_thr1_next[2]), .Y(exu_n410));
AND2X1 exu_U10082(.A(exu_n10803), .B(exu_n9795), .Y(rml_otherwin_reg_data_thr1_next[1]));
INVX1 exu_U10083(.A(rml_otherwin_reg_data_thr1_next[1]), .Y(exu_n411));
AND2X1 exu_U10084(.A(exu_n10804), .B(exu_n9796), .Y(rml_otherwin_reg_data_thr1_next[0]));
INVX1 exu_U10085(.A(rml_otherwin_reg_data_thr1_next[0]), .Y(exu_n412));
AND2X1 exu_U10086(.A(exu_n10805), .B(exu_n9797), .Y(rml_otherwin_reg_data_thr0_next[2]));
INVX1 exu_U10087(.A(rml_otherwin_reg_data_thr0_next[2]), .Y(exu_n413));
AND2X1 exu_U10088(.A(exu_n10806), .B(exu_n9798), .Y(rml_otherwin_reg_data_thr0_next[1]));
INVX1 exu_U10089(.A(rml_otherwin_reg_data_thr0_next[1]), .Y(exu_n414));
AND2X1 exu_U10090(.A(exu_n10807), .B(exu_n9799), .Y(rml_otherwin_reg_data_thr0_next[0]));
INVX1 exu_U10091(.A(rml_otherwin_reg_data_thr0_next[0]), .Y(exu_n415));
AND2X1 exu_U10092(.A(exu_n10808), .B(exu_n9800), .Y(rml_cleanwin_reg_data_thr3_next[2]));
INVX1 exu_U10093(.A(rml_cleanwin_reg_data_thr3_next[2]), .Y(exu_n416));
AND2X1 exu_U10094(.A(exu_n10809), .B(exu_n9801), .Y(rml_cleanwin_reg_data_thr3_next[1]));
INVX1 exu_U10095(.A(rml_cleanwin_reg_data_thr3_next[1]), .Y(exu_n417));
AND2X1 exu_U10096(.A(exu_n10810), .B(exu_n9802), .Y(rml_cleanwin_reg_data_thr3_next[0]));
INVX1 exu_U10097(.A(rml_cleanwin_reg_data_thr3_next[0]), .Y(exu_n418));
AND2X1 exu_U10098(.A(exu_n10811), .B(exu_n9803), .Y(rml_cleanwin_reg_data_thr2_next[2]));
INVX1 exu_U10099(.A(rml_cleanwin_reg_data_thr2_next[2]), .Y(exu_n419));
AND2X1 exu_U10100(.A(exu_n10812), .B(exu_n9804), .Y(rml_cleanwin_reg_data_thr2_next[1]));
INVX1 exu_U10101(.A(rml_cleanwin_reg_data_thr2_next[1]), .Y(exu_n420));
AND2X1 exu_U10102(.A(exu_n10813), .B(exu_n9805), .Y(rml_cleanwin_reg_data_thr2_next[0]));
INVX1 exu_U10103(.A(rml_cleanwin_reg_data_thr2_next[0]), .Y(exu_n421));
AND2X1 exu_U10104(.A(exu_n10814), .B(exu_n9806), .Y(rml_cleanwin_reg_data_thr1_next[2]));
INVX1 exu_U10105(.A(rml_cleanwin_reg_data_thr1_next[2]), .Y(exu_n422));
AND2X1 exu_U10106(.A(exu_n10815), .B(exu_n9807), .Y(rml_cleanwin_reg_data_thr1_next[1]));
INVX1 exu_U10107(.A(rml_cleanwin_reg_data_thr1_next[1]), .Y(exu_n423));
AND2X1 exu_U10108(.A(exu_n10816), .B(exu_n9808), .Y(rml_cleanwin_reg_data_thr1_next[0]));
INVX1 exu_U10109(.A(rml_cleanwin_reg_data_thr1_next[0]), .Y(exu_n424));
AND2X1 exu_U10110(.A(exu_n10817), .B(exu_n9809), .Y(rml_cleanwin_reg_data_thr0_next[2]));
INVX1 exu_U10111(.A(rml_cleanwin_reg_data_thr0_next[2]), .Y(exu_n425));
AND2X1 exu_U10112(.A(exu_n10818), .B(exu_n9810), .Y(rml_cleanwin_reg_data_thr0_next[1]));
INVX1 exu_U10113(.A(rml_cleanwin_reg_data_thr0_next[1]), .Y(exu_n426));
AND2X1 exu_U10114(.A(exu_n10819), .B(exu_n9811), .Y(rml_cleanwin_reg_data_thr0_next[0]));
INVX1 exu_U10115(.A(rml_cleanwin_reg_data_thr0_next[0]), .Y(exu_n427));
AND2X1 exu_U10116(.A(exu_n10820), .B(exu_n9812), .Y(rml_hi_wstate_reg_data_thr3_next[2]));
INVX1 exu_U10117(.A(rml_hi_wstate_reg_data_thr3_next[2]), .Y(exu_n428));
AND2X1 exu_U10118(.A(exu_n10821), .B(exu_n9813), .Y(rml_hi_wstate_reg_data_thr3_next[1]));
INVX1 exu_U10119(.A(rml_hi_wstate_reg_data_thr3_next[1]), .Y(exu_n429));
AND2X1 exu_U10120(.A(exu_n10822), .B(exu_n9814), .Y(rml_hi_wstate_reg_data_thr3_next[0]));
INVX1 exu_U10121(.A(rml_hi_wstate_reg_data_thr3_next[0]), .Y(exu_n430));
AND2X1 exu_U10122(.A(exu_n10823), .B(exu_n9815), .Y(rml_hi_wstate_reg_data_thr2_next[2]));
INVX1 exu_U10123(.A(rml_hi_wstate_reg_data_thr2_next[2]), .Y(exu_n431));
AND2X1 exu_U10124(.A(exu_n10824), .B(exu_n9816), .Y(rml_hi_wstate_reg_data_thr2_next[1]));
INVX1 exu_U10125(.A(rml_hi_wstate_reg_data_thr2_next[1]), .Y(exu_n432));
AND2X1 exu_U10126(.A(exu_n10825), .B(exu_n9817), .Y(rml_hi_wstate_reg_data_thr2_next[0]));
INVX1 exu_U10127(.A(rml_hi_wstate_reg_data_thr2_next[0]), .Y(exu_n433));
AND2X1 exu_U10128(.A(exu_n10826), .B(exu_n9818), .Y(rml_hi_wstate_reg_data_thr1_next[2]));
INVX1 exu_U10129(.A(rml_hi_wstate_reg_data_thr1_next[2]), .Y(exu_n434));
AND2X1 exu_U10130(.A(exu_n10827), .B(exu_n9819), .Y(rml_hi_wstate_reg_data_thr1_next[1]));
INVX1 exu_U10131(.A(rml_hi_wstate_reg_data_thr1_next[1]), .Y(exu_n435));
AND2X1 exu_U10132(.A(exu_n10828), .B(exu_n9820), .Y(rml_hi_wstate_reg_data_thr1_next[0]));
INVX1 exu_U10133(.A(rml_hi_wstate_reg_data_thr1_next[0]), .Y(exu_n436));
AND2X1 exu_U10134(.A(exu_n10829), .B(exu_n9821), .Y(rml_hi_wstate_reg_data_thr0_next[2]));
INVX1 exu_U10135(.A(rml_hi_wstate_reg_data_thr0_next[2]), .Y(exu_n437));
AND2X1 exu_U10136(.A(exu_n10830), .B(exu_n9822), .Y(rml_hi_wstate_reg_data_thr0_next[1]));
INVX1 exu_U10137(.A(rml_hi_wstate_reg_data_thr0_next[1]), .Y(exu_n438));
AND2X1 exu_U10138(.A(exu_n10831), .B(exu_n9823), .Y(rml_hi_wstate_reg_data_thr0_next[0]));
INVX1 exu_U10139(.A(rml_hi_wstate_reg_data_thr0_next[0]), .Y(exu_n439));
AND2X1 exu_U10140(.A(exu_n10832), .B(exu_n9824), .Y(rml_lo_wstate_reg_data_thr3_next[2]));
INVX1 exu_U10141(.A(rml_lo_wstate_reg_data_thr3_next[2]), .Y(exu_n440));
AND2X1 exu_U10142(.A(exu_n10833), .B(exu_n9825), .Y(rml_lo_wstate_reg_data_thr3_next[1]));
INVX1 exu_U10143(.A(rml_lo_wstate_reg_data_thr3_next[1]), .Y(exu_n441));
AND2X1 exu_U10144(.A(exu_n10834), .B(exu_n9826), .Y(rml_lo_wstate_reg_data_thr3_next[0]));
INVX1 exu_U10145(.A(rml_lo_wstate_reg_data_thr3_next[0]), .Y(exu_n442));
AND2X1 exu_U10146(.A(exu_n10835), .B(exu_n9827), .Y(rml_lo_wstate_reg_data_thr2_next[2]));
INVX1 exu_U10147(.A(rml_lo_wstate_reg_data_thr2_next[2]), .Y(exu_n443));
AND2X1 exu_U10148(.A(exu_n10836), .B(exu_n9828), .Y(rml_lo_wstate_reg_data_thr2_next[1]));
INVX1 exu_U10149(.A(rml_lo_wstate_reg_data_thr2_next[1]), .Y(exu_n444));
AND2X1 exu_U10150(.A(exu_n10837), .B(exu_n9829), .Y(rml_lo_wstate_reg_data_thr2_next[0]));
INVX1 exu_U10151(.A(rml_lo_wstate_reg_data_thr2_next[0]), .Y(exu_n445));
AND2X1 exu_U10152(.A(exu_n10838), .B(exu_n9830), .Y(rml_lo_wstate_reg_data_thr1_next[2]));
INVX1 exu_U10153(.A(rml_lo_wstate_reg_data_thr1_next[2]), .Y(exu_n446));
AND2X1 exu_U10154(.A(exu_n10839), .B(exu_n9831), .Y(rml_lo_wstate_reg_data_thr1_next[1]));
INVX1 exu_U10155(.A(rml_lo_wstate_reg_data_thr1_next[1]), .Y(exu_n447));
AND2X1 exu_U10156(.A(exu_n10840), .B(exu_n9832), .Y(rml_lo_wstate_reg_data_thr1_next[0]));
INVX1 exu_U10157(.A(rml_lo_wstate_reg_data_thr1_next[0]), .Y(exu_n448));
AND2X1 exu_U10158(.A(exu_n10841), .B(exu_n9833), .Y(rml_lo_wstate_reg_data_thr0_next[2]));
INVX1 exu_U10159(.A(rml_lo_wstate_reg_data_thr0_next[2]), .Y(exu_n449));
AND2X1 exu_U10160(.A(exu_n10842), .B(exu_n9834), .Y(rml_lo_wstate_reg_data_thr0_next[1]));
INVX1 exu_U10161(.A(rml_lo_wstate_reg_data_thr0_next[1]), .Y(exu_n450));
AND2X1 exu_U10162(.A(exu_n10843), .B(exu_n9835), .Y(rml_lo_wstate_reg_data_thr0_next[0]));
INVX1 exu_U10163(.A(rml_lo_wstate_reg_data_thr0_next[0]), .Y(exu_n451));
AND2X1 exu_U10164(.A(rml_rml_ecl_cansave_e[1]), .B(rml_rml_ecl_cansave_e[0]), .Y(exu_n18424));
INVX1 exu_U10165(.A(exu_n18424), .Y(exu_n452));
AND2X1 exu_U10166(.A(rml_rml_ecl_canrestore_e[1]), .B(rml_rml_ecl_canrestore_e[0]), .Y(exu_n18429));
INVX1 exu_U10167(.A(exu_n18429), .Y(exu_n453));
AND2X1 exu_U10168(.A(exu_n10844), .B(exu_n9836), .Y(rml_next_canrestore_e[0]));
INVX1 exu_U10169(.A(rml_next_canrestore_e[0]), .Y(exu_n454));
AND2X1 exu_U10170(.A(exu_n10845), .B(exu_n9837), .Y(rml_next_canrestore_e[1]));
INVX1 exu_U10171(.A(rml_next_canrestore_e[1]), .Y(exu_n455));
AND2X1 exu_U10172(.A(exu_n10846), .B(exu_n9838), .Y(rml_next_canrestore_e[2]));
INVX1 exu_U10173(.A(rml_next_canrestore_e[2]), .Y(exu_n456));
AND2X1 exu_U10174(.A(exu_n10847), .B(exu_n9839), .Y(rml_next_otherwin_e[0]));
INVX1 exu_U10175(.A(rml_next_otherwin_e[0]), .Y(exu_n457));
AND2X1 exu_U10176(.A(exu_n10848), .B(exu_n9840), .Y(rml_next_otherwin_e[1]));
INVX1 exu_U10177(.A(rml_next_otherwin_e[1]), .Y(exu_n458));
AND2X1 exu_U10178(.A(exu_n10849), .B(exu_n9841), .Y(rml_next_otherwin_e[2]));
INVX1 exu_U10179(.A(rml_next_otherwin_e[2]), .Y(exu_n459));
AND2X1 exu_U10180(.A(exu_n10850), .B(exu_n9842), .Y(rml_next_cleanwin_e[0]));
INVX1 exu_U10181(.A(rml_next_cleanwin_e[0]), .Y(exu_n460));
AND2X1 exu_U10182(.A(exu_n10851), .B(exu_n9843), .Y(rml_next_cleanwin_e[1]));
INVX1 exu_U10183(.A(rml_next_cleanwin_e[1]), .Y(exu_n461));
AND2X1 exu_U10184(.A(exu_n10852), .B(exu_n9844), .Y(rml_next_cleanwin_e[2]));
INVX1 exu_U10185(.A(rml_next_cleanwin_e[2]), .Y(exu_n462));
AND2X1 exu_U10186(.A(exu_n10853), .B(exu_n9845), .Y(rml_cansave_reg_data_thr0_next[0]));
INVX1 exu_U10187(.A(rml_cansave_reg_data_thr0_next[0]), .Y(exu_n463));
AND2X1 exu_U10188(.A(exu_n10854), .B(exu_n9846), .Y(rml_cansave_reg_data_thr0_next[1]));
INVX1 exu_U10189(.A(rml_cansave_reg_data_thr0_next[1]), .Y(exu_n464));
AND2X1 exu_U10190(.A(exu_n10855), .B(exu_n9847), .Y(rml_cansave_reg_data_thr0_next[2]));
INVX1 exu_U10191(.A(rml_cansave_reg_data_thr0_next[2]), .Y(exu_n465));
AND2X1 exu_U10192(.A(exu_n10856), .B(exu_n9848), .Y(rml_cansave_reg_data_thr1_next[0]));
INVX1 exu_U10193(.A(rml_cansave_reg_data_thr1_next[0]), .Y(exu_n466));
AND2X1 exu_U10194(.A(exu_n10857), .B(exu_n9849), .Y(rml_cansave_reg_data_thr1_next[1]));
INVX1 exu_U10195(.A(rml_cansave_reg_data_thr1_next[1]), .Y(exu_n467));
AND2X1 exu_U10196(.A(exu_n10858), .B(exu_n9850), .Y(rml_cansave_reg_data_thr1_next[2]));
INVX1 exu_U10197(.A(rml_cansave_reg_data_thr1_next[2]), .Y(exu_n468));
AND2X1 exu_U10198(.A(exu_n10859), .B(exu_n9851), .Y(rml_cansave_reg_data_thr2_next[0]));
INVX1 exu_U10199(.A(rml_cansave_reg_data_thr2_next[0]), .Y(exu_n469));
AND2X1 exu_U10200(.A(exu_n10860), .B(exu_n9852), .Y(rml_cansave_reg_data_thr2_next[1]));
INVX1 exu_U10201(.A(rml_cansave_reg_data_thr2_next[1]), .Y(exu_n470));
AND2X1 exu_U10202(.A(exu_n10861), .B(exu_n9853), .Y(rml_cansave_reg_data_thr2_next[2]));
INVX1 exu_U10203(.A(rml_cansave_reg_data_thr2_next[2]), .Y(exu_n471));
AND2X1 exu_U10204(.A(exu_n10862), .B(exu_n9854), .Y(rml_cansave_reg_data_thr3_next[0]));
INVX1 exu_U10205(.A(rml_cansave_reg_data_thr3_next[0]), .Y(exu_n472));
AND2X1 exu_U10206(.A(exu_n10863), .B(exu_n9855), .Y(rml_cansave_reg_data_thr3_next[1]));
INVX1 exu_U10207(.A(rml_cansave_reg_data_thr3_next[1]), .Y(exu_n473));
AND2X1 exu_U10208(.A(exu_n10864), .B(exu_n9856), .Y(rml_cansave_reg_data_thr3_next[2]));
INVX1 exu_U10209(.A(rml_cansave_reg_data_thr3_next[2]), .Y(exu_n474));
AND2X1 exu_U10210(.A(exu_n18603), .B(exu_n9857), .Y(div_next_mul_data[9]));
INVX1 exu_U10211(.A(div_next_mul_data[9]), .Y(exu_n475));
AND2X1 exu_U10212(.A(exu_n16256), .B(alu_logic_rs1_data_bf1[9]), .Y(exu_n18605));
INVX1 exu_U10213(.A(exu_n18605), .Y(exu_n476));
AND2X1 exu_U10214(.A(exu_n18607), .B(exu_n9858), .Y(div_next_mul_data[99]));
INVX1 exu_U10215(.A(div_next_mul_data[99]), .Y(exu_n477));
AND2X1 exu_U10216(.A(exu_n18610), .B(exu_n9859), .Y(div_next_mul_data[98]));
INVX1 exu_U10217(.A(div_next_mul_data[98]), .Y(exu_n478));
INVX1 exu_U10218(.A(exu_n483), .Y(exu_n479));
INVX1 exu_U10219(.A(exu_n479), .Y(exu_n480));
AND2X1 exu_U10220(.A(exu_n18613), .B(exu_n9860), .Y(div_next_mul_data[97]));
INVX1 exu_U10221(.A(div_next_mul_data[97]), .Y(exu_n481));
INVX1 exu_U10222(.A(exu_n486), .Y(exu_n482));
INVX1 exu_U10223(.A(exu_n482), .Y(exu_n483));
AND2X1 exu_U10224(.A(exu_n18616), .B(exu_n9861), .Y(div_next_mul_data[96]));
INVX1 exu_U10225(.A(div_next_mul_data[96]), .Y(exu_n484));
INVX1 exu_U10226(.A(exu_n678), .Y(exu_n485));
INVX1 exu_U10227(.A(exu_n485), .Y(exu_n486));
AND2X1 exu_U10228(.A(exu_n18619), .B(exu_n9862), .Y(div_next_mul_data[95]));
INVX1 exu_U10229(.A(div_next_mul_data[95]), .Y(exu_n487));
AND2X1 exu_U10230(.A(div_input_data_e[95]), .B(exu_n16256), .Y(exu_n18621));
INVX1 exu_U10231(.A(exu_n18621), .Y(exu_n488));
AND2X1 exu_U10232(.A(exu_n18623), .B(exu_n9863), .Y(div_next_mul_data[94]));
INVX1 exu_U10233(.A(div_next_mul_data[94]), .Y(exu_n489));
AND2X1 exu_U10234(.A(div_input_data_e[94]), .B(exu_n16256), .Y(exu_n18625));
INVX1 exu_U10235(.A(exu_n18625), .Y(exu_n490));
AND2X1 exu_U10236(.A(exu_n18627), .B(exu_n9864), .Y(div_next_mul_data[93]));
INVX1 exu_U10237(.A(div_next_mul_data[93]), .Y(exu_n491));
AND2X1 exu_U10238(.A(div_input_data_e[93]), .B(exu_n16256), .Y(exu_n18629));
INVX1 exu_U10239(.A(exu_n18629), .Y(exu_n492));
AND2X1 exu_U10240(.A(exu_n18631), .B(exu_n9865), .Y(div_next_mul_data[92]));
INVX1 exu_U10241(.A(div_next_mul_data[92]), .Y(exu_n493));
AND2X1 exu_U10242(.A(div_input_data_e[92]), .B(exu_n16256), .Y(exu_n18633));
INVX1 exu_U10243(.A(exu_n18633), .Y(exu_n494));
AND2X1 exu_U10244(.A(exu_n18635), .B(exu_n9866), .Y(div_next_mul_data[91]));
INVX1 exu_U10245(.A(div_next_mul_data[91]), .Y(exu_n495));
AND2X1 exu_U10246(.A(div_input_data_e[91]), .B(exu_n16256), .Y(exu_n18637));
INVX1 exu_U10247(.A(exu_n18637), .Y(exu_n496));
AND2X1 exu_U10248(.A(exu_n18639), .B(exu_n9867), .Y(div_next_mul_data[90]));
INVX1 exu_U10249(.A(div_next_mul_data[90]), .Y(exu_n497));
AND2X1 exu_U10250(.A(div_input_data_e[90]), .B(exu_n16256), .Y(exu_n18641));
INVX1 exu_U10251(.A(exu_n18641), .Y(exu_n498));
AND2X1 exu_U10252(.A(exu_n18643), .B(exu_n9868), .Y(div_next_mul_data[8]));
INVX1 exu_U10253(.A(div_next_mul_data[8]), .Y(exu_n499));
AND2X1 exu_U10254(.A(alu_logic_rs1_data_bf1[8]), .B(exu_n16256), .Y(exu_n18645));
INVX1 exu_U10255(.A(exu_n18645), .Y(exu_n500));
AND2X1 exu_U10256(.A(exu_n18647), .B(exu_n9869), .Y(div_next_mul_data[89]));
INVX1 exu_U10257(.A(div_next_mul_data[89]), .Y(exu_n501));
AND2X1 exu_U10258(.A(div_input_data_e[89]), .B(exu_n16256), .Y(exu_n18649));
INVX1 exu_U10259(.A(exu_n18649), .Y(exu_n502));
AND2X1 exu_U10260(.A(exu_n18651), .B(exu_n9870), .Y(div_next_mul_data[88]));
INVX1 exu_U10261(.A(div_next_mul_data[88]), .Y(exu_n503));
AND2X1 exu_U10262(.A(div_input_data_e[88]), .B(exu_n16256), .Y(exu_n18653));
INVX1 exu_U10263(.A(exu_n18653), .Y(exu_n504));
AND2X1 exu_U10264(.A(exu_n18655), .B(exu_n9871), .Y(div_next_mul_data[87]));
INVX1 exu_U10265(.A(div_next_mul_data[87]), .Y(exu_n505));
AND2X1 exu_U10266(.A(div_input_data_e[87]), .B(exu_n16256), .Y(exu_n18657));
INVX1 exu_U10267(.A(exu_n18657), .Y(exu_n506));
AND2X1 exu_U10268(.A(exu_n18659), .B(exu_n9872), .Y(div_next_mul_data[86]));
INVX1 exu_U10269(.A(div_next_mul_data[86]), .Y(exu_n507));
AND2X1 exu_U10270(.A(div_input_data_e[86]), .B(exu_n16256), .Y(exu_n18661));
INVX1 exu_U10271(.A(exu_n18661), .Y(exu_n508));
AND2X1 exu_U10272(.A(exu_n18663), .B(exu_n9873), .Y(div_next_mul_data[85]));
INVX1 exu_U10273(.A(div_next_mul_data[85]), .Y(exu_n509));
AND2X1 exu_U10274(.A(div_input_data_e[85]), .B(exu_n16256), .Y(exu_n18665));
INVX1 exu_U10275(.A(exu_n18665), .Y(exu_n510));
AND2X1 exu_U10276(.A(exu_n18667), .B(exu_n9874), .Y(div_next_mul_data[84]));
INVX1 exu_U10277(.A(div_next_mul_data[84]), .Y(exu_n511));
AND2X1 exu_U10278(.A(div_input_data_e[84]), .B(exu_n16256), .Y(exu_n18669));
INVX1 exu_U10279(.A(exu_n18669), .Y(exu_n512));
AND2X1 exu_U10280(.A(exu_n18671), .B(exu_n9875), .Y(div_next_mul_data[83]));
INVX1 exu_U10281(.A(div_next_mul_data[83]), .Y(exu_n513));
AND2X1 exu_U10282(.A(div_input_data_e[83]), .B(exu_n16256), .Y(exu_n18673));
INVX1 exu_U10283(.A(exu_n18673), .Y(exu_n514));
AND2X1 exu_U10284(.A(exu_n18675), .B(exu_n9876), .Y(div_next_mul_data[82]));
INVX1 exu_U10285(.A(div_next_mul_data[82]), .Y(exu_n515));
AND2X1 exu_U10286(.A(div_input_data_e[82]), .B(exu_n16256), .Y(exu_n18677));
INVX1 exu_U10287(.A(exu_n18677), .Y(exu_n516));
AND2X1 exu_U10288(.A(exu_n18679), .B(exu_n9877), .Y(div_next_mul_data[81]));
INVX1 exu_U10289(.A(div_next_mul_data[81]), .Y(exu_n517));
AND2X1 exu_U10290(.A(div_input_data_e[81]), .B(exu_n16256), .Y(exu_n18681));
INVX1 exu_U10291(.A(exu_n18681), .Y(exu_n518));
AND2X1 exu_U10292(.A(exu_n18683), .B(exu_n9878), .Y(div_next_mul_data[80]));
INVX1 exu_U10293(.A(div_next_mul_data[80]), .Y(exu_n519));
AND2X1 exu_U10294(.A(div_input_data_e[80]), .B(exu_n16256), .Y(exu_n18685));
INVX1 exu_U10295(.A(exu_n18685), .Y(exu_n520));
AND2X1 exu_U10296(.A(exu_n18687), .B(exu_n9879), .Y(div_next_mul_data[7]));
INVX1 exu_U10297(.A(div_next_mul_data[7]), .Y(exu_n521));
AND2X1 exu_U10298(.A(alu_logic_rs1_data_bf1[7]), .B(exu_n16256), .Y(exu_n18689));
INVX1 exu_U10299(.A(exu_n18689), .Y(exu_n522));
AND2X1 exu_U10300(.A(exu_n18691), .B(exu_n9880), .Y(div_next_mul_data[79]));
INVX1 exu_U10301(.A(div_next_mul_data[79]), .Y(exu_n523));
AND2X1 exu_U10302(.A(div_input_data_e[79]), .B(exu_n16256), .Y(exu_n18693));
INVX1 exu_U10303(.A(exu_n18693), .Y(exu_n524));
AND2X1 exu_U10304(.A(exu_n18695), .B(exu_n9881), .Y(div_next_mul_data[78]));
INVX1 exu_U10305(.A(div_next_mul_data[78]), .Y(exu_n525));
AND2X1 exu_U10306(.A(div_input_data_e[78]), .B(exu_n16256), .Y(exu_n18697));
INVX1 exu_U10307(.A(exu_n18697), .Y(exu_n526));
AND2X1 exu_U10308(.A(exu_n18699), .B(exu_n9882), .Y(div_next_mul_data[77]));
INVX1 exu_U10309(.A(div_next_mul_data[77]), .Y(exu_n527));
AND2X1 exu_U10310(.A(div_input_data_e[77]), .B(exu_n16256), .Y(exu_n18701));
INVX1 exu_U10311(.A(exu_n18701), .Y(exu_n528));
AND2X1 exu_U10312(.A(exu_n18703), .B(exu_n9883), .Y(div_next_mul_data[76]));
INVX1 exu_U10313(.A(div_next_mul_data[76]), .Y(exu_n529));
AND2X1 exu_U10314(.A(div_input_data_e[76]), .B(exu_n16256), .Y(exu_n18705));
INVX1 exu_U10315(.A(exu_n18705), .Y(exu_n530));
AND2X1 exu_U10316(.A(exu_n18707), .B(exu_n9884), .Y(div_next_mul_data[75]));
INVX1 exu_U10317(.A(div_next_mul_data[75]), .Y(exu_n531));
AND2X1 exu_U10318(.A(div_input_data_e[75]), .B(exu_n16256), .Y(exu_n18709));
INVX1 exu_U10319(.A(exu_n18709), .Y(exu_n532));
AND2X1 exu_U10320(.A(exu_n18711), .B(exu_n9885), .Y(div_next_mul_data[74]));
INVX1 exu_U10321(.A(div_next_mul_data[74]), .Y(exu_n533));
AND2X1 exu_U10322(.A(div_input_data_e[74]), .B(exu_n16256), .Y(exu_n18713));
INVX1 exu_U10323(.A(exu_n18713), .Y(exu_n534));
AND2X1 exu_U10324(.A(exu_n18715), .B(exu_n9886), .Y(div_next_mul_data[73]));
INVX1 exu_U10325(.A(div_next_mul_data[73]), .Y(exu_n535));
AND2X1 exu_U10326(.A(div_input_data_e[73]), .B(exu_n16256), .Y(exu_n18717));
INVX1 exu_U10327(.A(exu_n18717), .Y(exu_n536));
AND2X1 exu_U10328(.A(exu_n18719), .B(exu_n9887), .Y(div_next_mul_data[72]));
INVX1 exu_U10329(.A(div_next_mul_data[72]), .Y(exu_n537));
AND2X1 exu_U10330(.A(div_input_data_e[72]), .B(exu_n16256), .Y(exu_n18721));
INVX1 exu_U10331(.A(exu_n18721), .Y(exu_n538));
AND2X1 exu_U10332(.A(exu_n18723), .B(exu_n9888), .Y(div_next_mul_data[71]));
INVX1 exu_U10333(.A(div_next_mul_data[71]), .Y(exu_n539));
AND2X1 exu_U10334(.A(div_input_data_e[71]), .B(exu_n16256), .Y(exu_n18725));
INVX1 exu_U10335(.A(exu_n18725), .Y(exu_n540));
AND2X1 exu_U10336(.A(exu_n18727), .B(exu_n9889), .Y(div_next_mul_data[70]));
INVX1 exu_U10337(.A(div_next_mul_data[70]), .Y(exu_n541));
AND2X1 exu_U10338(.A(div_input_data_e[70]), .B(exu_n16256), .Y(exu_n18729));
INVX1 exu_U10339(.A(exu_n18729), .Y(exu_n542));
AND2X1 exu_U10340(.A(exu_n18731), .B(exu_n9890), .Y(div_next_mul_data[6]));
INVX1 exu_U10341(.A(div_next_mul_data[6]), .Y(exu_n543));
AND2X1 exu_U10342(.A(alu_logic_rs1_data_bf1[6]), .B(exu_n16256), .Y(exu_n18733));
INVX1 exu_U10343(.A(exu_n18733), .Y(exu_n544));
AND2X1 exu_U10344(.A(exu_n18735), .B(exu_n9891), .Y(div_next_mul_data[69]));
INVX1 exu_U10345(.A(div_next_mul_data[69]), .Y(exu_n545));
AND2X1 exu_U10346(.A(div_input_data_e[69]), .B(exu_n16256), .Y(exu_n18737));
INVX1 exu_U10347(.A(exu_n18737), .Y(exu_n546));
AND2X1 exu_U10348(.A(exu_n18739), .B(exu_n9892), .Y(div_next_mul_data[68]));
INVX1 exu_U10349(.A(div_next_mul_data[68]), .Y(exu_n547));
AND2X1 exu_U10350(.A(div_input_data_e[68]), .B(exu_n16256), .Y(exu_n18741));
INVX1 exu_U10351(.A(exu_n18741), .Y(exu_n548));
AND2X1 exu_U10352(.A(exu_n18743), .B(exu_n9893), .Y(div_next_mul_data[67]));
INVX1 exu_U10353(.A(div_next_mul_data[67]), .Y(exu_n549));
AND2X1 exu_U10354(.A(div_input_data_e[67]), .B(exu_n16256), .Y(exu_n18745));
INVX1 exu_U10355(.A(exu_n18745), .Y(exu_n550));
AND2X1 exu_U10356(.A(exu_n18747), .B(exu_n9894), .Y(div_next_mul_data[66]));
INVX1 exu_U10357(.A(div_next_mul_data[66]), .Y(exu_n551));
AND2X1 exu_U10358(.A(div_input_data_e[66]), .B(exu_n16256), .Y(exu_n18749));
INVX1 exu_U10359(.A(exu_n18749), .Y(exu_n552));
AND2X1 exu_U10360(.A(exu_n18751), .B(exu_n9895), .Y(div_next_mul_data[65]));
INVX1 exu_U10361(.A(div_next_mul_data[65]), .Y(exu_n553));
AND2X1 exu_U10362(.A(div_input_data_e[65]), .B(exu_n16256), .Y(exu_n18753));
INVX1 exu_U10363(.A(exu_n18753), .Y(exu_n554));
AND2X1 exu_U10364(.A(exu_n18755), .B(exu_n9896), .Y(div_next_mul_data[64]));
INVX1 exu_U10365(.A(div_next_mul_data[64]), .Y(exu_n555));
AND2X1 exu_U10366(.A(div_input_data_e[64]), .B(exu_n16256), .Y(exu_n18757));
INVX1 exu_U10367(.A(exu_n18757), .Y(exu_n556));
AND2X1 exu_U10368(.A(exu_n18759), .B(exu_n9897), .Y(div_next_mul_data[63]));
INVX1 exu_U10369(.A(div_next_mul_data[63]), .Y(exu_n557));
AND2X1 exu_U10370(.A(exu_n18762), .B(exu_n9898), .Y(div_next_mul_data[62]));
INVX1 exu_U10371(.A(div_next_mul_data[62]), .Y(exu_n558));
INVX1 exu_U10372(.A(exu_n563), .Y(exu_n559));
INVX1 exu_U10373(.A(exu_n559), .Y(exu_n560));
AND2X1 exu_U10374(.A(exu_n18765), .B(exu_n9899), .Y(div_next_mul_data[61]));
INVX1 exu_U10375(.A(div_next_mul_data[61]), .Y(exu_n561));
INVX1 exu_U10376(.A(exu_n566), .Y(exu_n562));
INVX1 exu_U10377(.A(exu_n562), .Y(exu_n563));
AND2X1 exu_U10378(.A(exu_n18768), .B(exu_n9900), .Y(div_next_mul_data[60]));
INVX1 exu_U10379(.A(div_next_mul_data[60]), .Y(exu_n564));
INVX1 exu_U10380(.A(exu_n571), .Y(exu_n565));
INVX1 exu_U10381(.A(exu_n565), .Y(exu_n566));
AND2X1 exu_U10382(.A(exu_n18771), .B(exu_n9901), .Y(div_next_mul_data[5]));
INVX1 exu_U10383(.A(div_next_mul_data[5]), .Y(exu_n567));
AND2X1 exu_U10384(.A(alu_logic_rs1_data_bf1[5]), .B(exu_n16256), .Y(exu_n18773));
INVX1 exu_U10385(.A(exu_n18773), .Y(exu_n568));
AND2X1 exu_U10386(.A(exu_n18775), .B(exu_n9902), .Y(div_next_mul_data[59]));
INVX1 exu_U10387(.A(div_next_mul_data[59]), .Y(exu_n569));
INVX1 exu_U10388(.A(exu_n574), .Y(exu_n570));
INVX1 exu_U10389(.A(exu_n570), .Y(exu_n571));
AND2X1 exu_U10390(.A(exu_n18778), .B(exu_n9903), .Y(div_next_mul_data[58]));
INVX1 exu_U10391(.A(div_next_mul_data[58]), .Y(exu_n572));
INVX1 exu_U10392(.A(exu_n577), .Y(exu_n573));
INVX1 exu_U10393(.A(exu_n573), .Y(exu_n574));
AND2X1 exu_U10394(.A(exu_n18781), .B(exu_n9904), .Y(div_next_mul_data[57]));
INVX1 exu_U10395(.A(div_next_mul_data[57]), .Y(exu_n575));
INVX1 exu_U10396(.A(exu_n580), .Y(exu_n576));
INVX1 exu_U10397(.A(exu_n576), .Y(exu_n577));
AND2X1 exu_U10398(.A(exu_n18784), .B(exu_n9905), .Y(div_next_mul_data[56]));
INVX1 exu_U10399(.A(div_next_mul_data[56]), .Y(exu_n578));
INVX1 exu_U10400(.A(exu_n583), .Y(exu_n579));
INVX1 exu_U10401(.A(exu_n579), .Y(exu_n580));
AND2X1 exu_U10402(.A(exu_n18787), .B(exu_n9906), .Y(div_next_mul_data[55]));
INVX1 exu_U10403(.A(div_next_mul_data[55]), .Y(exu_n581));
INVX1 exu_U10404(.A(exu_n586), .Y(exu_n582));
INVX1 exu_U10405(.A(exu_n582), .Y(exu_n583));
AND2X1 exu_U10406(.A(exu_n18790), .B(exu_n9907), .Y(div_next_mul_data[54]));
INVX1 exu_U10407(.A(div_next_mul_data[54]), .Y(exu_n584));
INVX1 exu_U10408(.A(exu_n589), .Y(exu_n585));
INVX1 exu_U10409(.A(exu_n585), .Y(exu_n586));
AND2X1 exu_U10410(.A(exu_n18793), .B(exu_n9908), .Y(div_next_mul_data[53]));
INVX1 exu_U10411(.A(div_next_mul_data[53]), .Y(exu_n587));
INVX1 exu_U10412(.A(exu_n592), .Y(exu_n588));
INVX1 exu_U10413(.A(exu_n588), .Y(exu_n589));
AND2X1 exu_U10414(.A(exu_n18796), .B(exu_n9909), .Y(div_next_mul_data[52]));
INVX1 exu_U10415(.A(div_next_mul_data[52]), .Y(exu_n590));
INVX1 exu_U10416(.A(exu_n595), .Y(exu_n591));
INVX1 exu_U10417(.A(exu_n591), .Y(exu_n592));
AND2X1 exu_U10418(.A(exu_n18799), .B(exu_n9910), .Y(div_next_mul_data[51]));
INVX1 exu_U10419(.A(div_next_mul_data[51]), .Y(exu_n593));
INVX1 exu_U10420(.A(exu_n598), .Y(exu_n594));
INVX1 exu_U10421(.A(exu_n594), .Y(exu_n595));
AND2X1 exu_U10422(.A(exu_n18802), .B(exu_n9911), .Y(div_next_mul_data[50]));
INVX1 exu_U10423(.A(div_next_mul_data[50]), .Y(exu_n596));
INVX1 exu_U10424(.A(exu_n603), .Y(exu_n597));
INVX1 exu_U10425(.A(exu_n597), .Y(exu_n598));
AND2X1 exu_U10426(.A(exu_n18805), .B(exu_n9912), .Y(div_next_mul_data[4]));
INVX1 exu_U10427(.A(div_next_mul_data[4]), .Y(exu_n599));
AND2X1 exu_U10428(.A(alu_logic_rs1_data_bf1[4]), .B(exu_n16256), .Y(exu_n18807));
INVX1 exu_U10429(.A(exu_n18807), .Y(exu_n600));
AND2X1 exu_U10430(.A(exu_n18809), .B(exu_n9913), .Y(div_next_mul_data[49]));
INVX1 exu_U10431(.A(div_next_mul_data[49]), .Y(exu_n601));
INVX1 exu_U10432(.A(exu_n606), .Y(exu_n602));
INVX1 exu_U10433(.A(exu_n602), .Y(exu_n603));
AND2X1 exu_U10434(.A(exu_n18812), .B(exu_n9914), .Y(div_next_mul_data[48]));
INVX1 exu_U10435(.A(div_next_mul_data[48]), .Y(exu_n604));
INVX1 exu_U10436(.A(exu_n609), .Y(exu_n605));
INVX1 exu_U10437(.A(exu_n605), .Y(exu_n606));
AND2X1 exu_U10438(.A(exu_n18815), .B(exu_n9915), .Y(div_next_mul_data[47]));
INVX1 exu_U10439(.A(div_next_mul_data[47]), .Y(exu_n607));
INVX1 exu_U10440(.A(exu_n612), .Y(exu_n608));
INVX1 exu_U10441(.A(exu_n608), .Y(exu_n609));
AND2X1 exu_U10442(.A(exu_n18818), .B(exu_n9916), .Y(div_next_mul_data[46]));
INVX1 exu_U10443(.A(div_next_mul_data[46]), .Y(exu_n610));
INVX1 exu_U10444(.A(exu_n615), .Y(exu_n611));
INVX1 exu_U10445(.A(exu_n611), .Y(exu_n612));
AND2X1 exu_U10446(.A(exu_n18821), .B(exu_n9917), .Y(div_next_mul_data[45]));
INVX1 exu_U10447(.A(div_next_mul_data[45]), .Y(exu_n613));
INVX1 exu_U10448(.A(exu_n631), .Y(exu_n614));
INVX1 exu_U10449(.A(exu_n614), .Y(exu_n615));
AND2X1 exu_U10450(.A(exu_n18824), .B(exu_n9918), .Y(div_next_mul_data[44]));
INVX1 exu_U10451(.A(div_next_mul_data[44]), .Y(exu_n616));
AND2X1 exu_U10452(.A(exu_n18827), .B(exu_n9919), .Y(div_next_mul_data[43]));
INVX1 exu_U10453(.A(div_next_mul_data[43]), .Y(exu_n617));
AND2X1 exu_U10454(.A(exu_n18830), .B(exu_n9920), .Y(div_next_mul_data[42]));
INVX1 exu_U10455(.A(div_next_mul_data[42]), .Y(exu_n618));
AND2X1 exu_U10456(.A(exu_n18833), .B(exu_n9921), .Y(div_next_mul_data[41]));
INVX1 exu_U10457(.A(div_next_mul_data[41]), .Y(exu_n619));
AND2X1 exu_U10458(.A(exu_n18836), .B(exu_n9922), .Y(div_next_mul_data[40]));
INVX1 exu_U10459(.A(div_next_mul_data[40]), .Y(exu_n620));
AND2X1 exu_U10460(.A(exu_n18839), .B(exu_n9923), .Y(div_next_mul_data[3]));
INVX1 exu_U10461(.A(div_next_mul_data[3]), .Y(exu_n621));
AND2X1 exu_U10462(.A(alu_logic_rs1_data_bf1[3]), .B(exu_n16256), .Y(exu_n18841));
INVX1 exu_U10463(.A(exu_n18841), .Y(exu_n622));
AND2X1 exu_U10464(.A(exu_n18843), .B(exu_n9924), .Y(div_next_mul_data[39]));
INVX1 exu_U10465(.A(div_next_mul_data[39]), .Y(exu_n623));
AND2X1 exu_U10466(.A(exu_n18846), .B(exu_n9925), .Y(div_next_mul_data[38]));
INVX1 exu_U10467(.A(div_next_mul_data[38]), .Y(exu_n624));
AND2X1 exu_U10468(.A(exu_n18849), .B(exu_n9926), .Y(div_next_mul_data[37]));
INVX1 exu_U10469(.A(div_next_mul_data[37]), .Y(exu_n625));
AND2X1 exu_U10470(.A(exu_n18852), .B(exu_n9927), .Y(div_next_mul_data[36]));
INVX1 exu_U10471(.A(div_next_mul_data[36]), .Y(exu_n626));
AND2X1 exu_U10472(.A(exu_n18855), .B(exu_n9928), .Y(div_next_mul_data[35]));
INVX1 exu_U10473(.A(div_next_mul_data[35]), .Y(exu_n627));
AND2X1 exu_U10474(.A(exu_n18858), .B(exu_n9929), .Y(div_next_mul_data[34]));
INVX1 exu_U10475(.A(div_next_mul_data[34]), .Y(exu_n628));
AND2X1 exu_U10476(.A(exu_n18861), .B(exu_n9930), .Y(div_next_mul_data[33]));
INVX1 exu_U10477(.A(div_next_mul_data[33]), .Y(exu_n629));
AND2X1 exu_U10478(.A(exu_n18864), .B(exu_n9931), .Y(div_next_mul_data[32]));
INVX1 exu_U10479(.A(div_next_mul_data[32]), .Y(exu_n630));
AND2X1 exu_U10480(.A(ecl_div_mul_sext_rs1_e), .B(exu_n16256), .Y(exu_n18866));
INVX1 exu_U10481(.A(exu_n18866), .Y(exu_n631));
AND2X1 exu_U10482(.A(exu_n18868), .B(exu_n9932), .Y(div_next_mul_data[31]));
INVX1 exu_U10483(.A(div_next_mul_data[31]), .Y(exu_n632));
AND2X1 exu_U10484(.A(alu_logic_rs1_data_bf1[31]), .B(exu_n16256), .Y(exu_n18870));
INVX1 exu_U10485(.A(exu_n18870), .Y(exu_n633));
AND2X1 exu_U10486(.A(exu_n18872), .B(exu_n9933), .Y(div_next_mul_data[30]));
INVX1 exu_U10487(.A(div_next_mul_data[30]), .Y(exu_n634));
AND2X1 exu_U10488(.A(alu_logic_rs1_data_bf1[30]), .B(exu_n16256), .Y(exu_n18874));
INVX1 exu_U10489(.A(exu_n18874), .Y(exu_n635));
AND2X1 exu_U10490(.A(exu_n18876), .B(exu_n9934), .Y(div_next_mul_data[2]));
INVX1 exu_U10491(.A(div_next_mul_data[2]), .Y(exu_n636));
AND2X1 exu_U10492(.A(alu_logic_rs1_data_bf1[2]), .B(exu_n16256), .Y(exu_n18878));
INVX1 exu_U10493(.A(exu_n18878), .Y(exu_n637));
AND2X1 exu_U10494(.A(exu_n18880), .B(exu_n9935), .Y(div_next_mul_data[29]));
INVX1 exu_U10495(.A(div_next_mul_data[29]), .Y(exu_n638));
AND2X1 exu_U10496(.A(alu_logic_rs1_data_bf1[29]), .B(exu_n16256), .Y(exu_n18882));
INVX1 exu_U10497(.A(exu_n18882), .Y(exu_n639));
AND2X1 exu_U10498(.A(exu_n18884), .B(exu_n9936), .Y(div_next_mul_data[28]));
INVX1 exu_U10499(.A(div_next_mul_data[28]), .Y(exu_n640));
AND2X1 exu_U10500(.A(alu_logic_rs1_data_bf1[28]), .B(exu_n16256), .Y(exu_n18886));
INVX1 exu_U10501(.A(exu_n18886), .Y(exu_n641));
AND2X1 exu_U10502(.A(exu_n18888), .B(exu_n9937), .Y(div_next_mul_data[27]));
INVX1 exu_U10503(.A(div_next_mul_data[27]), .Y(exu_n642));
AND2X1 exu_U10504(.A(alu_logic_rs1_data_bf1[27]), .B(exu_n16256), .Y(exu_n18890));
INVX1 exu_U10505(.A(exu_n18890), .Y(exu_n643));
AND2X1 exu_U10506(.A(exu_n18892), .B(exu_n9938), .Y(div_next_mul_data[26]));
INVX1 exu_U10507(.A(div_next_mul_data[26]), .Y(exu_n644));
AND2X1 exu_U10508(.A(alu_logic_rs1_data_bf1[26]), .B(exu_n16256), .Y(exu_n18894));
INVX1 exu_U10509(.A(exu_n18894), .Y(exu_n645));
AND2X1 exu_U10510(.A(exu_n18896), .B(exu_n9939), .Y(div_next_mul_data[25]));
INVX1 exu_U10511(.A(div_next_mul_data[25]), .Y(exu_n646));
AND2X1 exu_U10512(.A(alu_logic_rs1_data_bf1[25]), .B(exu_n16256), .Y(exu_n18898));
INVX1 exu_U10513(.A(exu_n18898), .Y(exu_n647));
AND2X1 exu_U10514(.A(exu_n18900), .B(exu_n9940), .Y(div_next_mul_data[24]));
INVX1 exu_U10515(.A(div_next_mul_data[24]), .Y(exu_n648));
AND2X1 exu_U10516(.A(alu_logic_rs1_data_bf1[24]), .B(exu_n16256), .Y(exu_n18902));
INVX1 exu_U10517(.A(exu_n18902), .Y(exu_n649));
AND2X1 exu_U10518(.A(exu_n18904), .B(exu_n9941), .Y(div_next_mul_data[23]));
INVX1 exu_U10519(.A(div_next_mul_data[23]), .Y(exu_n650));
AND2X1 exu_U10520(.A(alu_logic_rs1_data_bf1[23]), .B(exu_n16256), .Y(exu_n18906));
INVX1 exu_U10521(.A(exu_n18906), .Y(exu_n651));
AND2X1 exu_U10522(.A(exu_n18908), .B(exu_n9942), .Y(div_next_mul_data[22]));
INVX1 exu_U10523(.A(div_next_mul_data[22]), .Y(exu_n652));
AND2X1 exu_U10524(.A(alu_logic_rs1_data_bf1[22]), .B(exu_n16256), .Y(exu_n18910));
INVX1 exu_U10525(.A(exu_n18910), .Y(exu_n653));
AND2X1 exu_U10526(.A(exu_n18912), .B(exu_n9943), .Y(div_next_mul_data[21]));
INVX1 exu_U10527(.A(div_next_mul_data[21]), .Y(exu_n654));
AND2X1 exu_U10528(.A(alu_logic_rs1_data_bf1[21]), .B(exu_n16256), .Y(exu_n18914));
INVX1 exu_U10529(.A(exu_n18914), .Y(exu_n655));
AND2X1 exu_U10530(.A(exu_n18916), .B(exu_n9944), .Y(div_next_mul_data[20]));
INVX1 exu_U10531(.A(div_next_mul_data[20]), .Y(exu_n656));
AND2X1 exu_U10532(.A(alu_logic_rs1_data_bf1[20]), .B(exu_n16256), .Y(exu_n18918));
INVX1 exu_U10533(.A(exu_n18918), .Y(exu_n657));
AND2X1 exu_U10534(.A(exu_n18920), .B(exu_n9945), .Y(div_next_mul_data[1]));
INVX1 exu_U10535(.A(div_next_mul_data[1]), .Y(exu_n658));
AND2X1 exu_U10536(.A(alu_logic_rs1_data_bf1[1]), .B(exu_n16256), .Y(exu_n18922));
INVX1 exu_U10537(.A(exu_n18922), .Y(exu_n659));
AND2X1 exu_U10538(.A(exu_n18924), .B(exu_n9946), .Y(div_next_mul_data[19]));
INVX1 exu_U10539(.A(div_next_mul_data[19]), .Y(exu_n660));
AND2X1 exu_U10540(.A(alu_logic_rs1_data_bf1[19]), .B(exu_n16256), .Y(exu_n18926));
INVX1 exu_U10541(.A(exu_n18926), .Y(exu_n661));
AND2X1 exu_U10542(.A(exu_n18928), .B(exu_n9947), .Y(div_next_mul_data[18]));
INVX1 exu_U10543(.A(div_next_mul_data[18]), .Y(exu_n662));
AND2X1 exu_U10544(.A(alu_logic_rs1_data_bf1[18]), .B(exu_n16256), .Y(exu_n18930));
INVX1 exu_U10545(.A(exu_n18930), .Y(exu_n663));
AND2X1 exu_U10546(.A(exu_n18932), .B(exu_n9948), .Y(div_next_mul_data[17]));
INVX1 exu_U10547(.A(div_next_mul_data[17]), .Y(exu_n664));
AND2X1 exu_U10548(.A(alu_logic_rs1_data_bf1[17]), .B(exu_n16256), .Y(exu_n18934));
INVX1 exu_U10549(.A(exu_n18934), .Y(exu_n665));
AND2X1 exu_U10550(.A(exu_n18936), .B(exu_n9949), .Y(div_next_mul_data[16]));
INVX1 exu_U10551(.A(div_next_mul_data[16]), .Y(exu_n666));
AND2X1 exu_U10552(.A(alu_logic_rs1_data_bf1[16]), .B(exu_n16256), .Y(exu_n18938));
INVX1 exu_U10553(.A(exu_n18938), .Y(exu_n667));
AND2X1 exu_U10554(.A(exu_n18940), .B(exu_n9950), .Y(div_next_mul_data[15]));
INVX1 exu_U10555(.A(div_next_mul_data[15]), .Y(exu_n668));
AND2X1 exu_U10556(.A(alu_logic_rs1_data_bf1[15]), .B(exu_n16256), .Y(exu_n18942));
INVX1 exu_U10557(.A(exu_n18942), .Y(exu_n669));
AND2X1 exu_U10558(.A(exu_n18944), .B(exu_n9951), .Y(div_next_mul_data[14]));
INVX1 exu_U10559(.A(div_next_mul_data[14]), .Y(exu_n670));
AND2X1 exu_U10560(.A(alu_logic_rs1_data_bf1[14]), .B(exu_n16256), .Y(exu_n18946));
INVX1 exu_U10561(.A(exu_n18946), .Y(exu_n671));
AND2X1 exu_U10562(.A(exu_n18948), .B(exu_n9952), .Y(div_next_mul_data[13]));
INVX1 exu_U10563(.A(div_next_mul_data[13]), .Y(exu_n672));
AND2X1 exu_U10564(.A(alu_logic_rs1_data_bf1[13]), .B(exu_n16256), .Y(exu_n18950));
INVX1 exu_U10565(.A(exu_n18950), .Y(exu_n673));
AND2X1 exu_U10566(.A(exu_n18952), .B(exu_n9953), .Y(div_next_mul_data[12]));
INVX1 exu_U10567(.A(div_next_mul_data[12]), .Y(exu_n674));
AND2X1 exu_U10568(.A(alu_logic_rs1_data_bf1[12]), .B(exu_n16256), .Y(exu_n18954));
INVX1 exu_U10569(.A(exu_n18954), .Y(exu_n675));
AND2X1 exu_U10570(.A(exu_n18956), .B(exu_n9954), .Y(div_next_mul_data[127]));
INVX1 exu_U10571(.A(div_next_mul_data[127]), .Y(exu_n676));
INVX1 exu_U10572(.A(exu_n681), .Y(exu_n677));
INVX1 exu_U10573(.A(exu_n677), .Y(exu_n678));
AND2X1 exu_U10574(.A(exu_n18959), .B(exu_n9955), .Y(div_next_mul_data[126]));
INVX1 exu_U10575(.A(div_next_mul_data[126]), .Y(exu_n679));
INVX1 exu_U10576(.A(exu_n684), .Y(exu_n680));
INVX1 exu_U10577(.A(exu_n680), .Y(exu_n681));
AND2X1 exu_U10578(.A(exu_n18962), .B(exu_n9956), .Y(div_next_mul_data[125]));
INVX1 exu_U10579(.A(div_next_mul_data[125]), .Y(exu_n682));
INVX1 exu_U10580(.A(exu_n687), .Y(exu_n683));
INVX1 exu_U10581(.A(exu_n683), .Y(exu_n684));
AND2X1 exu_U10582(.A(exu_n18965), .B(exu_n9957), .Y(div_next_mul_data[124]));
INVX1 exu_U10583(.A(div_next_mul_data[124]), .Y(exu_n685));
INVX1 exu_U10584(.A(exu_n690), .Y(exu_n686));
INVX1 exu_U10585(.A(exu_n686), .Y(exu_n687));
AND2X1 exu_U10586(.A(exu_n18968), .B(exu_n9958), .Y(div_next_mul_data[123]));
INVX1 exu_U10587(.A(div_next_mul_data[123]), .Y(exu_n688));
INVX1 exu_U10588(.A(exu_n693), .Y(exu_n689));
INVX1 exu_U10589(.A(exu_n689), .Y(exu_n690));
AND2X1 exu_U10590(.A(exu_n18971), .B(exu_n9959), .Y(div_next_mul_data[122]));
INVX1 exu_U10591(.A(div_next_mul_data[122]), .Y(exu_n691));
INVX1 exu_U10592(.A(exu_n696), .Y(exu_n692));
INVX1 exu_U10593(.A(exu_n692), .Y(exu_n693));
AND2X1 exu_U10594(.A(exu_n18974), .B(exu_n9960), .Y(div_next_mul_data[121]));
INVX1 exu_U10595(.A(div_next_mul_data[121]), .Y(exu_n694));
INVX1 exu_U10596(.A(exu_n699), .Y(exu_n695));
INVX1 exu_U10597(.A(exu_n695), .Y(exu_n696));
AND2X1 exu_U10598(.A(exu_n18977), .B(exu_n9961), .Y(div_next_mul_data[120]));
INVX1 exu_U10599(.A(div_next_mul_data[120]), .Y(exu_n697));
INVX1 exu_U10600(.A(exu_n704), .Y(exu_n698));
INVX1 exu_U10601(.A(exu_n698), .Y(exu_n699));
AND2X1 exu_U10602(.A(exu_n18980), .B(exu_n9962), .Y(div_next_mul_data[11]));
INVX1 exu_U10603(.A(div_next_mul_data[11]), .Y(exu_n700));
AND2X1 exu_U10604(.A(alu_logic_rs1_data_bf1[11]), .B(exu_n16256), .Y(exu_n18982));
INVX1 exu_U10605(.A(exu_n18982), .Y(exu_n701));
AND2X1 exu_U10606(.A(exu_n18984), .B(exu_n9963), .Y(div_next_mul_data[119]));
INVX1 exu_U10607(.A(div_next_mul_data[119]), .Y(exu_n702));
INVX1 exu_U10608(.A(exu_n707), .Y(exu_n703));
INVX1 exu_U10609(.A(exu_n703), .Y(exu_n704));
AND2X1 exu_U10610(.A(exu_n18987), .B(exu_n9964), .Y(div_next_mul_data[118]));
INVX1 exu_U10611(.A(div_next_mul_data[118]), .Y(exu_n705));
INVX1 exu_U10612(.A(exu_n710), .Y(exu_n706));
INVX1 exu_U10613(.A(exu_n706), .Y(exu_n707));
AND2X1 exu_U10614(.A(exu_n18990), .B(exu_n9965), .Y(div_next_mul_data[117]));
INVX1 exu_U10615(.A(div_next_mul_data[117]), .Y(exu_n708));
INVX1 exu_U10616(.A(exu_n713), .Y(exu_n709));
INVX1 exu_U10617(.A(exu_n709), .Y(exu_n710));
AND2X1 exu_U10618(.A(exu_n18993), .B(exu_n9966), .Y(div_next_mul_data[116]));
INVX1 exu_U10619(.A(div_next_mul_data[116]), .Y(exu_n711));
INVX1 exu_U10620(.A(exu_n716), .Y(exu_n712));
INVX1 exu_U10621(.A(exu_n712), .Y(exu_n713));
AND2X1 exu_U10622(.A(exu_n18996), .B(exu_n9967), .Y(div_next_mul_data[115]));
INVX1 exu_U10623(.A(div_next_mul_data[115]), .Y(exu_n714));
INVX1 exu_U10624(.A(exu_n719), .Y(exu_n715));
INVX1 exu_U10625(.A(exu_n715), .Y(exu_n716));
AND2X1 exu_U10626(.A(exu_n18999), .B(exu_n9968), .Y(div_next_mul_data[114]));
INVX1 exu_U10627(.A(div_next_mul_data[114]), .Y(exu_n717));
INVX1 exu_U10628(.A(exu_n736), .Y(exu_n718));
INVX1 exu_U10629(.A(exu_n718), .Y(exu_n719));
AND2X1 exu_U10630(.A(exu_n19002), .B(exu_n9969), .Y(div_next_mul_data[113]));
INVX1 exu_U10631(.A(div_next_mul_data[113]), .Y(exu_n720));
AND2X1 exu_U10632(.A(exu_n19005), .B(exu_n9970), .Y(div_next_mul_data[112]));
INVX1 exu_U10633(.A(div_next_mul_data[112]), .Y(exu_n721));
AND2X1 exu_U10634(.A(exu_n19008), .B(exu_n9971), .Y(div_next_mul_data[111]));
INVX1 exu_U10635(.A(div_next_mul_data[111]), .Y(exu_n722));
AND2X1 exu_U10636(.A(exu_n19011), .B(exu_n9972), .Y(div_next_mul_data[110]));
INVX1 exu_U10637(.A(div_next_mul_data[110]), .Y(exu_n723));
AND2X1 exu_U10638(.A(exu_n19014), .B(exu_n9973), .Y(div_next_mul_data[10]));
INVX1 exu_U10639(.A(div_next_mul_data[10]), .Y(exu_n724));
AND2X1 exu_U10640(.A(alu_logic_rs1_data_bf1[10]), .B(exu_n16256), .Y(exu_n19016));
INVX1 exu_U10641(.A(exu_n19016), .Y(exu_n725));
AND2X1 exu_U10642(.A(exu_n19018), .B(exu_n9974), .Y(div_next_mul_data[109]));
INVX1 exu_U10643(.A(div_next_mul_data[109]), .Y(exu_n726));
AND2X1 exu_U10644(.A(exu_n19021), .B(exu_n9975), .Y(div_next_mul_data[108]));
INVX1 exu_U10645(.A(div_next_mul_data[108]), .Y(exu_n727));
AND2X1 exu_U10646(.A(exu_n19024), .B(exu_n9976), .Y(div_next_mul_data[107]));
INVX1 exu_U10647(.A(div_next_mul_data[107]), .Y(exu_n728));
AND2X1 exu_U10648(.A(exu_n19027), .B(exu_n9977), .Y(div_next_mul_data[106]));
INVX1 exu_U10649(.A(div_next_mul_data[106]), .Y(exu_n729));
AND2X1 exu_U10650(.A(exu_n19030), .B(exu_n9978), .Y(div_next_mul_data[105]));
INVX1 exu_U10651(.A(div_next_mul_data[105]), .Y(exu_n730));
AND2X1 exu_U10652(.A(exu_n19033), .B(exu_n9979), .Y(div_next_mul_data[104]));
INVX1 exu_U10653(.A(div_next_mul_data[104]), .Y(exu_n731));
AND2X1 exu_U10654(.A(exu_n19036), .B(exu_n9980), .Y(div_next_mul_data[103]));
INVX1 exu_U10655(.A(div_next_mul_data[103]), .Y(exu_n732));
AND2X1 exu_U10656(.A(exu_n19039), .B(exu_n9981), .Y(div_next_mul_data[102]));
INVX1 exu_U10657(.A(div_next_mul_data[102]), .Y(exu_n733));
AND2X1 exu_U10658(.A(exu_n19042), .B(exu_n9982), .Y(div_next_mul_data[101]));
INVX1 exu_U10659(.A(div_next_mul_data[101]), .Y(exu_n734));
AND2X1 exu_U10660(.A(exu_n19045), .B(exu_n9983), .Y(div_next_mul_data[100]));
INVX1 exu_U10661(.A(div_next_mul_data[100]), .Y(exu_n735));
AND2X1 exu_U10662(.A(ecl_div_mul_sext_rs2_e), .B(exu_n16256), .Y(exu_n19047));
INVX1 exu_U10663(.A(exu_n19047), .Y(exu_n736));
AND2X1 exu_U10664(.A(exu_n19049), .B(exu_n9984), .Y(div_next_mul_data[0]));
INVX1 exu_U10665(.A(div_next_mul_data[0]), .Y(exu_n737));
AND2X1 exu_U10666(.A(alu_logic_rs1_data_bf1[0]), .B(exu_n16256), .Y(exu_n19051));
INVX1 exu_U10667(.A(exu_n19051), .Y(exu_n738));
AND2X1 exu_U10668(.A(alu_logic_rs1_data_bf1[63]), .B(ecl_div_div64), .Y(exu_n19067));
INVX1 exu_U10669(.A(exu_n19067), .Y(exu_n739));
AND2X1 exu_U10670(.A(ecl_div_div64), .B(div_input_data_e[105]), .Y(exu_n19151));
INVX1 exu_U10671(.A(exu_n19151), .Y(exu_n740));
AND2X1 exu_U10672(.A(div_input_data_e[104]), .B(ecl_div_div64), .Y(exu_n19152));
INVX1 exu_U10673(.A(exu_n19152), .Y(exu_n741));
AND2X1 exu_U10674(.A(div_input_data_e[103]), .B(ecl_div_div64), .Y(exu_n19153));
INVX1 exu_U10675(.A(exu_n19153), .Y(exu_n742));
AND2X1 exu_U10676(.A(div_input_data_e[102]), .B(ecl_div_div64), .Y(exu_n19154));
INVX1 exu_U10677(.A(exu_n19154), .Y(exu_n743));
AND2X1 exu_U10678(.A(div_input_data_e[101]), .B(ecl_div_div64), .Y(exu_n19155));
INVX1 exu_U10679(.A(exu_n19155), .Y(exu_n744));
AND2X1 exu_U10680(.A(div_input_data_e[100]), .B(ecl_div_div64), .Y(exu_n19156));
INVX1 exu_U10681(.A(exu_n19156), .Y(exu_n745));
AND2X1 exu_U10682(.A(div_input_data_e[99]), .B(ecl_div_div64), .Y(exu_n19157));
INVX1 exu_U10683(.A(exu_n19157), .Y(exu_n746));
AND2X1 exu_U10684(.A(div_input_data_e[127]), .B(ecl_div_div64), .Y(exu_n19158));
INVX1 exu_U10685(.A(exu_n19158), .Y(exu_n747));
AND2X1 exu_U10686(.A(div_input_data_e[126]), .B(ecl_div_div64), .Y(exu_n19159));
INVX1 exu_U10687(.A(exu_n19159), .Y(exu_n748));
AND2X1 exu_U10688(.A(div_input_data_e[98]), .B(ecl_div_div64), .Y(exu_n19160));
INVX1 exu_U10689(.A(exu_n19160), .Y(exu_n749));
AND2X1 exu_U10690(.A(div_input_data_e[125]), .B(ecl_div_div64), .Y(exu_n19161));
INVX1 exu_U10691(.A(exu_n19161), .Y(exu_n750));
AND2X1 exu_U10692(.A(div_input_data_e[124]), .B(ecl_div_div64), .Y(exu_n19162));
INVX1 exu_U10693(.A(exu_n19162), .Y(exu_n751));
AND2X1 exu_U10694(.A(div_input_data_e[123]), .B(ecl_div_div64), .Y(exu_n19163));
INVX1 exu_U10695(.A(exu_n19163), .Y(exu_n752));
AND2X1 exu_U10696(.A(div_input_data_e[122]), .B(ecl_div_div64), .Y(exu_n19164));
INVX1 exu_U10697(.A(exu_n19164), .Y(exu_n753));
AND2X1 exu_U10698(.A(div_input_data_e[121]), .B(ecl_div_div64), .Y(exu_n19165));
INVX1 exu_U10699(.A(exu_n19165), .Y(exu_n754));
AND2X1 exu_U10700(.A(div_input_data_e[120]), .B(ecl_div_div64), .Y(exu_n19166));
INVX1 exu_U10701(.A(exu_n19166), .Y(exu_n755));
AND2X1 exu_U10702(.A(div_input_data_e[119]), .B(ecl_div_div64), .Y(exu_n19167));
INVX1 exu_U10703(.A(exu_n19167), .Y(exu_n756));
AND2X1 exu_U10704(.A(div_input_data_e[118]), .B(ecl_div_div64), .Y(exu_n19168));
INVX1 exu_U10705(.A(exu_n19168), .Y(exu_n757));
AND2X1 exu_U10706(.A(div_input_data_e[117]), .B(ecl_div_div64), .Y(exu_n19169));
INVX1 exu_U10707(.A(exu_n19169), .Y(exu_n758));
AND2X1 exu_U10708(.A(div_input_data_e[116]), .B(ecl_div_div64), .Y(exu_n19170));
INVX1 exu_U10709(.A(exu_n19170), .Y(exu_n759));
AND2X1 exu_U10710(.A(div_input_data_e[97]), .B(ecl_div_div64), .Y(exu_n19171));
INVX1 exu_U10711(.A(exu_n19171), .Y(exu_n760));
AND2X1 exu_U10712(.A(div_input_data_e[115]), .B(ecl_div_div64), .Y(exu_n19172));
INVX1 exu_U10713(.A(exu_n19172), .Y(exu_n761));
AND2X1 exu_U10714(.A(div_input_data_e[114]), .B(ecl_div_div64), .Y(exu_n19173));
INVX1 exu_U10715(.A(exu_n19173), .Y(exu_n762));
AND2X1 exu_U10716(.A(div_input_data_e[113]), .B(ecl_div_div64), .Y(exu_n19174));
INVX1 exu_U10717(.A(exu_n19174), .Y(exu_n763));
AND2X1 exu_U10718(.A(div_input_data_e[112]), .B(ecl_div_div64), .Y(exu_n19175));
INVX1 exu_U10719(.A(exu_n19175), .Y(exu_n764));
AND2X1 exu_U10720(.A(div_input_data_e[111]), .B(ecl_div_div64), .Y(exu_n19176));
INVX1 exu_U10721(.A(exu_n19176), .Y(exu_n765));
AND2X1 exu_U10722(.A(div_input_data_e[110]), .B(ecl_div_div64), .Y(exu_n19177));
INVX1 exu_U10723(.A(exu_n19177), .Y(exu_n766));
AND2X1 exu_U10724(.A(div_input_data_e[109]), .B(ecl_div_div64), .Y(exu_n19178));
INVX1 exu_U10725(.A(exu_n19178), .Y(exu_n767));
AND2X1 exu_U10726(.A(div_input_data_e[108]), .B(ecl_div_div64), .Y(exu_n19179));
INVX1 exu_U10727(.A(exu_n19179), .Y(exu_n768));
AND2X1 exu_U10728(.A(div_input_data_e[107]), .B(ecl_div_div64), .Y(exu_n19180));
INVX1 exu_U10729(.A(exu_n19180), .Y(exu_n769));
AND2X1 exu_U10730(.A(div_input_data_e[106]), .B(ecl_div_div64), .Y(exu_n19181));
INVX1 exu_U10731(.A(exu_n19181), .Y(exu_n770));
AND2X1 exu_U10732(.A(div_input_data_e[96]), .B(ecl_div_div64), .Y(exu_n19182));
INVX1 exu_U10733(.A(exu_n19182), .Y(exu_n771));
AND2X1 exu_U10734(.A(exu_n15376), .B(exu_n9985), .Y(exu_n19185));
INVX1 exu_U10735(.A(exu_n19185), .Y(exu_n772));
OR2X1 U10736 ( .A(1'b0), .B(sehold), .Y(n19215) );
INVX1 exu_U10737(.A(exu_n19215), .Y(exu_n773));
AND2X1 exu_U10738(.A(exu_n15377), .B(exu_n9989), .Y(exu_n19221));
INVX1 exu_U10739(.A(exu_n19221), .Y(exu_n774));
AND2X1 exu_U10740(.A(ecl_ecc_log_rs2_m), .B(ecc_rs2_err_m[6]), .Y(exu_n19924));
INVX1 exu_U10741(.A(exu_n19924), .Y(exu_n775));
AND2X1 exu_U10742(.A(ecc_rs2_err_m[5]), .B(ecl_ecc_log_rs2_m), .Y(exu_n19928));
INVX1 exu_U10743(.A(exu_n19928), .Y(exu_n776));
AND2X1 exu_U10744(.A(ecc_rs2_err_m[4]), .B(ecl_ecc_log_rs2_m), .Y(exu_n19932));
INVX1 exu_U10745(.A(exu_n19932), .Y(exu_n777));
AND2X1 exu_U10746(.A(ecc_rs2_err_m[3]), .B(ecl_ecc_log_rs2_m), .Y(exu_n19936));
INVX1 exu_U10747(.A(exu_n19936), .Y(exu_n778));
AND2X1 exu_U10748(.A(ecc_rs2_err_m[2]), .B(ecl_ecc_log_rs2_m), .Y(exu_n19940));
INVX1 exu_U10749(.A(exu_n19940), .Y(exu_n779));
AND2X1 exu_U10750(.A(ecc_rs2_err_m[1]), .B(ecl_ecc_log_rs2_m), .Y(exu_n19944));
INVX1 exu_U10751(.A(exu_n19944), .Y(exu_n780));
AND2X1 exu_U10752(.A(ecc_rs2_err_m[0]), .B(ecl_ecc_log_rs2_m), .Y(exu_n19948));
INVX1 exu_U10753(.A(exu_n19948), .Y(exu_n781));
AND2X1 exu_U10754(.A(exu_n10992), .B(exu_n19999), .Y(exu_n19997));
INVX1 exu_U10755(.A(exu_n19997), .Y(exu_n782));
OR2X1 exu_U10756(.A(ecc_rs2_err_e[4]), .B(ecc_rs2_err_e[3]), .Y(exu_n20000));
INVX1 exu_U10757(.A(exu_n20000), .Y(exu_n783));
AND2X1 exu_U10758(.A(exu_n10993), .B(exu_n20135), .Y(exu_n20133));
INVX1 exu_U10759(.A(exu_n20133), .Y(exu_n784));
OR2X1 exu_U10760(.A(ecc_rs3_err_e[4]), .B(ecc_rs3_err_e[3]), .Y(exu_n20136));
INVX1 exu_U10761(.A(exu_n20136), .Y(exu_n785));
AND2X1 exu_U10762(.A(exu_n16287), .B(lsu_exu_dfill_data_g[9]), .Y(exu_n20478));
INVX1 exu_U10763(.A(exu_n20478), .Y(exu_n786));
AND2X1 exu_U10764(.A(exu_n16005), .B(bypass_mux_rs3h_data_2_in1[9]), .Y(exu_n20480));
INVX1 exu_U10765(.A(exu_n20480), .Y(exu_n787));
AND2X1 exu_U10766(.A(lsu_exu_dfill_data_g[8]), .B(exu_n16287), .Y(exu_n20484));
INVX1 exu_U10767(.A(exu_n20484), .Y(exu_n788));
AND2X1 exu_U10768(.A(bypass_mux_rs3h_data_2_in1[8]), .B(exu_n16005), .Y(exu_n20486));
INVX1 exu_U10769(.A(exu_n20486), .Y(exu_n789));
AND2X1 exu_U10770(.A(lsu_exu_dfill_data_g[7]), .B(exu_n16287), .Y(exu_n20490));
INVX1 exu_U10771(.A(exu_n20490), .Y(exu_n790));
AND2X1 exu_U10772(.A(bypass_mux_rs3h_data_2_in1[7]), .B(exu_n16005), .Y(exu_n20492));
INVX1 exu_U10773(.A(exu_n20492), .Y(exu_n791));
AND2X1 exu_U10774(.A(lsu_exu_dfill_data_g[6]), .B(exu_n16287), .Y(exu_n20496));
INVX1 exu_U10775(.A(exu_n20496), .Y(exu_n792));
AND2X1 exu_U10776(.A(bypass_mux_rs3h_data_2_in1[6]), .B(exu_n16005), .Y(exu_n20498));
INVX1 exu_U10777(.A(exu_n20498), .Y(exu_n793));
AND2X1 exu_U10778(.A(lsu_exu_dfill_data_g[5]), .B(exu_n16287), .Y(exu_n20502));
INVX1 exu_U10779(.A(exu_n20502), .Y(exu_n794));
AND2X1 exu_U10780(.A(bypass_mux_rs3h_data_2_in1[5]), .B(exu_n16005), .Y(exu_n20504));
INVX1 exu_U10781(.A(exu_n20504), .Y(exu_n795));
AND2X1 exu_U10782(.A(lsu_exu_dfill_data_g[4]), .B(exu_n16287), .Y(exu_n20508));
INVX1 exu_U10783(.A(exu_n20508), .Y(exu_n796));
AND2X1 exu_U10784(.A(bypass_mux_rs3h_data_2_in1[4]), .B(exu_n16005), .Y(exu_n20510));
INVX1 exu_U10785(.A(exu_n20510), .Y(exu_n797));
AND2X1 exu_U10786(.A(lsu_exu_dfill_data_g[3]), .B(exu_n16287), .Y(exu_n20514));
INVX1 exu_U10787(.A(exu_n20514), .Y(exu_n798));
AND2X1 exu_U10788(.A(bypass_mux_rs3h_data_2_in1[3]), .B(exu_n16005), .Y(exu_n20516));
INVX1 exu_U10789(.A(exu_n20516), .Y(exu_n799));
AND2X1 exu_U10790(.A(lsu_exu_dfill_data_g[31]), .B(exu_n16287), .Y(exu_n20520));
INVX1 exu_U10791(.A(exu_n20520), .Y(exu_n800));
AND2X1 exu_U10792(.A(bypass_mux_rs3h_data_2_in1[31]), .B(exu_n16005), .Y(exu_n20522));
INVX1 exu_U10793(.A(exu_n20522), .Y(exu_n801));
AND2X1 exu_U10794(.A(lsu_exu_dfill_data_g[30]), .B(exu_n16287), .Y(exu_n20526));
INVX1 exu_U10795(.A(exu_n20526), .Y(exu_n802));
AND2X1 exu_U10796(.A(bypass_mux_rs3h_data_2_in1[30]), .B(exu_n16005), .Y(exu_n20528));
INVX1 exu_U10797(.A(exu_n20528), .Y(exu_n803));
AND2X1 exu_U10798(.A(lsu_exu_dfill_data_g[2]), .B(exu_n16287), .Y(exu_n20532));
INVX1 exu_U10799(.A(exu_n20532), .Y(exu_n804));
AND2X1 exu_U10800(.A(bypass_mux_rs3h_data_2_in1[2]), .B(exu_n16005), .Y(exu_n20534));
INVX1 exu_U10801(.A(exu_n20534), .Y(exu_n805));
AND2X1 exu_U10802(.A(lsu_exu_dfill_data_g[29]), .B(exu_n16287), .Y(exu_n20538));
INVX1 exu_U10803(.A(exu_n20538), .Y(exu_n806));
AND2X1 exu_U10804(.A(bypass_mux_rs3h_data_2_in1[29]), .B(exu_n16005), .Y(exu_n20540));
INVX1 exu_U10805(.A(exu_n20540), .Y(exu_n807));
AND2X1 exu_U10806(.A(lsu_exu_dfill_data_g[28]), .B(exu_n16287), .Y(exu_n20544));
INVX1 exu_U10807(.A(exu_n20544), .Y(exu_n808));
AND2X1 exu_U10808(.A(bypass_mux_rs3h_data_2_in1[28]), .B(exu_n16005), .Y(exu_n20546));
INVX1 exu_U10809(.A(exu_n20546), .Y(exu_n809));
AND2X1 exu_U10810(.A(lsu_exu_dfill_data_g[27]), .B(exu_n16287), .Y(exu_n20550));
INVX1 exu_U10811(.A(exu_n20550), .Y(exu_n810));
AND2X1 exu_U10812(.A(bypass_mux_rs3h_data_2_in1[27]), .B(exu_n16005), .Y(exu_n20552));
INVX1 exu_U10813(.A(exu_n20552), .Y(exu_n811));
AND2X1 exu_U10814(.A(lsu_exu_dfill_data_g[26]), .B(exu_n16287), .Y(exu_n20556));
INVX1 exu_U10815(.A(exu_n20556), .Y(exu_n812));
AND2X1 exu_U10816(.A(bypass_mux_rs3h_data_2_in1[26]), .B(exu_n16005), .Y(exu_n20558));
INVX1 exu_U10817(.A(exu_n20558), .Y(exu_n813));
AND2X1 exu_U10818(.A(lsu_exu_dfill_data_g[25]), .B(exu_n16287), .Y(exu_n20562));
INVX1 exu_U10819(.A(exu_n20562), .Y(exu_n814));
AND2X1 exu_U10820(.A(bypass_mux_rs3h_data_2_in1[25]), .B(exu_n16005), .Y(exu_n20564));
INVX1 exu_U10821(.A(exu_n20564), .Y(exu_n815));
AND2X1 exu_U10822(.A(lsu_exu_dfill_data_g[24]), .B(exu_n16287), .Y(exu_n20568));
INVX1 exu_U10823(.A(exu_n20568), .Y(exu_n816));
AND2X1 exu_U10824(.A(bypass_mux_rs3h_data_2_in1[24]), .B(exu_n16005), .Y(exu_n20570));
INVX1 exu_U10825(.A(exu_n20570), .Y(exu_n817));
AND2X1 exu_U10826(.A(lsu_exu_dfill_data_g[23]), .B(exu_n16287), .Y(exu_n20574));
INVX1 exu_U10827(.A(exu_n20574), .Y(exu_n818));
AND2X1 exu_U10828(.A(bypass_mux_rs3h_data_2_in1[23]), .B(exu_n16005), .Y(exu_n20576));
INVX1 exu_U10829(.A(exu_n20576), .Y(exu_n819));
AND2X1 exu_U10830(.A(lsu_exu_dfill_data_g[22]), .B(exu_n16287), .Y(exu_n20580));
INVX1 exu_U10831(.A(exu_n20580), .Y(exu_n820));
AND2X1 exu_U10832(.A(bypass_mux_rs3h_data_2_in1[22]), .B(exu_n16005), .Y(exu_n20582));
INVX1 exu_U10833(.A(exu_n20582), .Y(exu_n821));
AND2X1 exu_U10834(.A(lsu_exu_dfill_data_g[21]), .B(exu_n16287), .Y(exu_n20586));
INVX1 exu_U10835(.A(exu_n20586), .Y(exu_n822));
AND2X1 exu_U10836(.A(bypass_mux_rs3h_data_2_in1[21]), .B(exu_n16005), .Y(exu_n20588));
INVX1 exu_U10837(.A(exu_n20588), .Y(exu_n823));
AND2X1 exu_U10838(.A(lsu_exu_dfill_data_g[20]), .B(exu_n16287), .Y(exu_n20592));
INVX1 exu_U10839(.A(exu_n20592), .Y(exu_n824));
AND2X1 exu_U10840(.A(bypass_mux_rs3h_data_2_in1[20]), .B(exu_n16005), .Y(exu_n20594));
INVX1 exu_U10841(.A(exu_n20594), .Y(exu_n825));
AND2X1 exu_U10842(.A(lsu_exu_dfill_data_g[1]), .B(exu_n16287), .Y(exu_n20598));
INVX1 exu_U10843(.A(exu_n20598), .Y(exu_n826));
AND2X1 exu_U10844(.A(bypass_mux_rs3h_data_2_in1[1]), .B(exu_n16005), .Y(exu_n20600));
INVX1 exu_U10845(.A(exu_n20600), .Y(exu_n827));
AND2X1 exu_U10846(.A(lsu_exu_dfill_data_g[19]), .B(exu_n16287), .Y(exu_n20604));
INVX1 exu_U10847(.A(exu_n20604), .Y(exu_n828));
AND2X1 exu_U10848(.A(bypass_mux_rs3h_data_2_in1[19]), .B(exu_n16005), .Y(exu_n20606));
INVX1 exu_U10849(.A(exu_n20606), .Y(exu_n829));
AND2X1 exu_U10850(.A(lsu_exu_dfill_data_g[18]), .B(exu_n16287), .Y(exu_n20610));
INVX1 exu_U10851(.A(exu_n20610), .Y(exu_n830));
AND2X1 exu_U10852(.A(bypass_mux_rs3h_data_2_in1[18]), .B(exu_n16005), .Y(exu_n20612));
INVX1 exu_U10853(.A(exu_n20612), .Y(exu_n831));
AND2X1 exu_U10854(.A(lsu_exu_dfill_data_g[17]), .B(exu_n16287), .Y(exu_n20616));
INVX1 exu_U10855(.A(exu_n20616), .Y(exu_n832));
AND2X1 exu_U10856(.A(bypass_mux_rs3h_data_2_in1[17]), .B(exu_n16005), .Y(exu_n20618));
INVX1 exu_U10857(.A(exu_n20618), .Y(exu_n833));
AND2X1 exu_U10858(.A(lsu_exu_dfill_data_g[16]), .B(exu_n16287), .Y(exu_n20622));
INVX1 exu_U10859(.A(exu_n20622), .Y(exu_n834));
AND2X1 exu_U10860(.A(bypass_mux_rs3h_data_2_in1[16]), .B(exu_n16005), .Y(exu_n20624));
INVX1 exu_U10861(.A(exu_n20624), .Y(exu_n835));
AND2X1 exu_U10862(.A(lsu_exu_dfill_data_g[15]), .B(exu_n16287), .Y(exu_n20628));
INVX1 exu_U10863(.A(exu_n20628), .Y(exu_n836));
AND2X1 exu_U10864(.A(bypass_mux_rs3h_data_2_in1[15]), .B(exu_n16005), .Y(exu_n20630));
INVX1 exu_U10865(.A(exu_n20630), .Y(exu_n837));
AND2X1 exu_U10866(.A(lsu_exu_dfill_data_g[14]), .B(exu_n16287), .Y(exu_n20634));
INVX1 exu_U10867(.A(exu_n20634), .Y(exu_n838));
AND2X1 exu_U10868(.A(bypass_mux_rs3h_data_2_in1[14]), .B(exu_n16005), .Y(exu_n20636));
INVX1 exu_U10869(.A(exu_n20636), .Y(exu_n839));
AND2X1 exu_U10870(.A(lsu_exu_dfill_data_g[13]), .B(exu_n16287), .Y(exu_n20640));
INVX1 exu_U10871(.A(exu_n20640), .Y(exu_n840));
AND2X1 exu_U10872(.A(bypass_mux_rs3h_data_2_in1[13]), .B(exu_n16005), .Y(exu_n20642));
INVX1 exu_U10873(.A(exu_n20642), .Y(exu_n841));
AND2X1 exu_U10874(.A(lsu_exu_dfill_data_g[12]), .B(exu_n16287), .Y(exu_n20646));
INVX1 exu_U10875(.A(exu_n20646), .Y(exu_n842));
AND2X1 exu_U10876(.A(bypass_mux_rs3h_data_2_in1[12]), .B(exu_n16005), .Y(exu_n20648));
INVX1 exu_U10877(.A(exu_n20648), .Y(exu_n843));
AND2X1 exu_U10878(.A(lsu_exu_dfill_data_g[11]), .B(exu_n16287), .Y(exu_n20652));
INVX1 exu_U10879(.A(exu_n20652), .Y(exu_n844));
AND2X1 exu_U10880(.A(bypass_mux_rs3h_data_2_in1[11]), .B(exu_n16005), .Y(exu_n20654));
INVX1 exu_U10881(.A(exu_n20654), .Y(exu_n845));
AND2X1 exu_U10882(.A(lsu_exu_dfill_data_g[10]), .B(exu_n16287), .Y(exu_n20658));
INVX1 exu_U10883(.A(exu_n20658), .Y(exu_n846));
AND2X1 exu_U10884(.A(bypass_mux_rs3h_data_2_in1[10]), .B(exu_n16005), .Y(exu_n20660));
INVX1 exu_U10885(.A(exu_n20660), .Y(exu_n847));
AND2X1 exu_U10886(.A(lsu_exu_dfill_data_g[0]), .B(exu_n16287), .Y(exu_n20664));
INVX1 exu_U10887(.A(exu_n20664), .Y(exu_n848));
AND2X1 exu_U10888(.A(bypass_mux_rs3h_data_2_in1[0]), .B(exu_n16005), .Y(exu_n20666));
INVX1 exu_U10889(.A(exu_n20666), .Y(exu_n849));
AND2X1 exu_U10890(.A(ecl_div_thr_e[3]), .B(div_yreg_yreg_thr3[9]), .Y(exu_n20670));
INVX1 exu_U10891(.A(exu_n20670), .Y(exu_n850));
AND2X1 exu_U10892(.A(exu_n16221), .B(div_yreg_yreg_thr1[9]), .Y(exu_n20672));
INVX1 exu_U10893(.A(exu_n20672), .Y(exu_n851));
AND2X1 exu_U10894(.A(div_yreg_yreg_thr3[8]), .B(ecl_div_thr_e[3]), .Y(exu_n20676));
INVX1 exu_U10895(.A(exu_n20676), .Y(exu_n852));
AND2X1 exu_U10896(.A(div_yreg_yreg_thr1[8]), .B(exu_n16221), .Y(exu_n20678));
INVX1 exu_U10897(.A(exu_n20678), .Y(exu_n853));
AND2X1 exu_U10898(.A(div_yreg_yreg_thr3[7]), .B(ecl_div_thr_e[3]), .Y(exu_n20682));
INVX1 exu_U10899(.A(exu_n20682), .Y(exu_n854));
AND2X1 exu_U10900(.A(div_yreg_yreg_thr1[7]), .B(exu_n16221), .Y(exu_n20684));
INVX1 exu_U10901(.A(exu_n20684), .Y(exu_n855));
AND2X1 exu_U10902(.A(div_yreg_yreg_thr3[6]), .B(ecl_div_thr_e[3]), .Y(exu_n20688));
INVX1 exu_U10903(.A(exu_n20688), .Y(exu_n856));
AND2X1 exu_U10904(.A(div_yreg_yreg_thr1[6]), .B(exu_n16221), .Y(exu_n20690));
INVX1 exu_U10905(.A(exu_n20690), .Y(exu_n857));
AND2X1 exu_U10906(.A(div_yreg_yreg_thr3[5]), .B(ecl_div_thr_e[3]), .Y(exu_n20694));
INVX1 exu_U10907(.A(exu_n20694), .Y(exu_n858));
AND2X1 exu_U10908(.A(div_yreg_yreg_thr1[5]), .B(exu_n16221), .Y(exu_n20696));
INVX1 exu_U10909(.A(exu_n20696), .Y(exu_n859));
AND2X1 exu_U10910(.A(div_yreg_yreg_thr3[4]), .B(ecl_div_thr_e[3]), .Y(exu_n20700));
INVX1 exu_U10911(.A(exu_n20700), .Y(exu_n860));
AND2X1 exu_U10912(.A(div_yreg_yreg_thr1[4]), .B(exu_n16221), .Y(exu_n20702));
INVX1 exu_U10913(.A(exu_n20702), .Y(exu_n861));
AND2X1 exu_U10914(.A(div_yreg_yreg_thr3[3]), .B(ecl_div_thr_e[3]), .Y(exu_n20706));
INVX1 exu_U10915(.A(exu_n20706), .Y(exu_n862));
AND2X1 exu_U10916(.A(div_yreg_yreg_thr1[3]), .B(exu_n16221), .Y(exu_n20708));
INVX1 exu_U10917(.A(exu_n20708), .Y(exu_n863));
AND2X1 exu_U10918(.A(div_yreg_yreg_thr3[31]), .B(ecl_div_thr_e[3]), .Y(exu_n20712));
INVX1 exu_U10919(.A(exu_n20712), .Y(exu_n864));
AND2X1 exu_U10920(.A(div_yreg_yreg_thr1[31]), .B(exu_n16221), .Y(exu_n20714));
INVX1 exu_U10921(.A(exu_n20714), .Y(exu_n865));
AND2X1 exu_U10922(.A(div_yreg_yreg_thr3[30]), .B(ecl_div_thr_e[3]), .Y(exu_n20718));
INVX1 exu_U10923(.A(exu_n20718), .Y(exu_n866));
AND2X1 exu_U10924(.A(div_yreg_yreg_thr1[30]), .B(exu_n16221), .Y(exu_n20720));
INVX1 exu_U10925(.A(exu_n20720), .Y(exu_n867));
AND2X1 exu_U10926(.A(div_yreg_yreg_thr3[2]), .B(ecl_div_thr_e[3]), .Y(exu_n20724));
INVX1 exu_U10927(.A(exu_n20724), .Y(exu_n868));
AND2X1 exu_U10928(.A(div_yreg_yreg_thr1[2]), .B(exu_n16221), .Y(exu_n20726));
INVX1 exu_U10929(.A(exu_n20726), .Y(exu_n869));
AND2X1 exu_U10930(.A(div_yreg_yreg_thr3[29]), .B(ecl_div_thr_e[3]), .Y(exu_n20730));
INVX1 exu_U10931(.A(exu_n20730), .Y(exu_n870));
AND2X1 exu_U10932(.A(div_yreg_yreg_thr1[29]), .B(exu_n16221), .Y(exu_n20732));
INVX1 exu_U10933(.A(exu_n20732), .Y(exu_n871));
AND2X1 exu_U10934(.A(div_yreg_yreg_thr3[28]), .B(ecl_div_thr_e[3]), .Y(exu_n20736));
INVX1 exu_U10935(.A(exu_n20736), .Y(exu_n872));
AND2X1 exu_U10936(.A(div_yreg_yreg_thr1[28]), .B(exu_n16221), .Y(exu_n20738));
INVX1 exu_U10937(.A(exu_n20738), .Y(exu_n873));
AND2X1 exu_U10938(.A(div_yreg_yreg_thr3[27]), .B(ecl_div_thr_e[3]), .Y(exu_n20742));
INVX1 exu_U10939(.A(exu_n20742), .Y(exu_n874));
AND2X1 exu_U10940(.A(div_yreg_yreg_thr1[27]), .B(exu_n16221), .Y(exu_n20744));
INVX1 exu_U10941(.A(exu_n20744), .Y(exu_n875));
AND2X1 exu_U10942(.A(div_yreg_yreg_thr3[26]), .B(ecl_div_thr_e[3]), .Y(exu_n20748));
INVX1 exu_U10943(.A(exu_n20748), .Y(exu_n876));
AND2X1 exu_U10944(.A(div_yreg_yreg_thr1[26]), .B(exu_n16221), .Y(exu_n20750));
INVX1 exu_U10945(.A(exu_n20750), .Y(exu_n877));
AND2X1 exu_U10946(.A(div_yreg_yreg_thr3[25]), .B(ecl_div_thr_e[3]), .Y(exu_n20754));
INVX1 exu_U10947(.A(exu_n20754), .Y(exu_n878));
AND2X1 exu_U10948(.A(div_yreg_yreg_thr1[25]), .B(exu_n16221), .Y(exu_n20756));
INVX1 exu_U10949(.A(exu_n20756), .Y(exu_n879));
AND2X1 exu_U10950(.A(div_yreg_yreg_thr3[24]), .B(ecl_div_thr_e[3]), .Y(exu_n20760));
INVX1 exu_U10951(.A(exu_n20760), .Y(exu_n880));
AND2X1 exu_U10952(.A(div_yreg_yreg_thr1[24]), .B(exu_n16221), .Y(exu_n20762));
INVX1 exu_U10953(.A(exu_n20762), .Y(exu_n881));
AND2X1 exu_U10954(.A(div_yreg_yreg_thr3[23]), .B(ecl_div_thr_e[3]), .Y(exu_n20766));
INVX1 exu_U10955(.A(exu_n20766), .Y(exu_n882));
AND2X1 exu_U10956(.A(div_yreg_yreg_thr1[23]), .B(exu_n16221), .Y(exu_n20768));
INVX1 exu_U10957(.A(exu_n20768), .Y(exu_n883));
AND2X1 exu_U10958(.A(div_yreg_yreg_thr3[22]), .B(ecl_div_thr_e[3]), .Y(exu_n20772));
INVX1 exu_U10959(.A(exu_n20772), .Y(exu_n884));
AND2X1 exu_U10960(.A(div_yreg_yreg_thr1[22]), .B(exu_n16221), .Y(exu_n20774));
INVX1 exu_U10961(.A(exu_n20774), .Y(exu_n885));
AND2X1 exu_U10962(.A(div_yreg_yreg_thr3[21]), .B(ecl_div_thr_e[3]), .Y(exu_n20778));
INVX1 exu_U10963(.A(exu_n20778), .Y(exu_n886));
AND2X1 exu_U10964(.A(div_yreg_yreg_thr1[21]), .B(exu_n16221), .Y(exu_n20780));
INVX1 exu_U10965(.A(exu_n20780), .Y(exu_n887));
AND2X1 exu_U10966(.A(div_yreg_yreg_thr3[20]), .B(ecl_div_thr_e[3]), .Y(exu_n20784));
INVX1 exu_U10967(.A(exu_n20784), .Y(exu_n888));
AND2X1 exu_U10968(.A(div_yreg_yreg_thr1[20]), .B(exu_n16221), .Y(exu_n20786));
INVX1 exu_U10969(.A(exu_n20786), .Y(exu_n889));
AND2X1 exu_U10970(.A(div_yreg_yreg_thr3[1]), .B(ecl_div_thr_e[3]), .Y(exu_n20790));
INVX1 exu_U10971(.A(exu_n20790), .Y(exu_n890));
AND2X1 exu_U10972(.A(div_yreg_yreg_thr1[1]), .B(exu_n16221), .Y(exu_n20792));
INVX1 exu_U10973(.A(exu_n20792), .Y(exu_n891));
AND2X1 exu_U10974(.A(div_yreg_yreg_thr3[19]), .B(ecl_div_thr_e[3]), .Y(exu_n20796));
INVX1 exu_U10975(.A(exu_n20796), .Y(exu_n892));
AND2X1 exu_U10976(.A(div_yreg_yreg_thr1[19]), .B(exu_n16221), .Y(exu_n20798));
INVX1 exu_U10977(.A(exu_n20798), .Y(exu_n893));
AND2X1 exu_U10978(.A(div_yreg_yreg_thr3[18]), .B(ecl_div_thr_e[3]), .Y(exu_n20802));
INVX1 exu_U10979(.A(exu_n20802), .Y(exu_n894));
AND2X1 exu_U10980(.A(div_yreg_yreg_thr1[18]), .B(exu_n16221), .Y(exu_n20804));
INVX1 exu_U10981(.A(exu_n20804), .Y(exu_n895));
AND2X1 exu_U10982(.A(div_yreg_yreg_thr3[17]), .B(ecl_div_thr_e[3]), .Y(exu_n20808));
INVX1 exu_U10983(.A(exu_n20808), .Y(exu_n896));
AND2X1 exu_U10984(.A(div_yreg_yreg_thr1[17]), .B(exu_n16221), .Y(exu_n20810));
INVX1 exu_U10985(.A(exu_n20810), .Y(exu_n897));
AND2X1 exu_U10986(.A(div_yreg_yreg_thr3[16]), .B(ecl_div_thr_e[3]), .Y(exu_n20814));
INVX1 exu_U10987(.A(exu_n20814), .Y(exu_n898));
AND2X1 exu_U10988(.A(div_yreg_yreg_thr1[16]), .B(exu_n16221), .Y(exu_n20816));
INVX1 exu_U10989(.A(exu_n20816), .Y(exu_n899));
AND2X1 exu_U10990(.A(div_yreg_yreg_thr3[15]), .B(ecl_div_thr_e[3]), .Y(exu_n20820));
INVX1 exu_U10991(.A(exu_n20820), .Y(exu_n900));
AND2X1 exu_U10992(.A(div_yreg_yreg_thr1[15]), .B(exu_n16221), .Y(exu_n20822));
INVX1 exu_U10993(.A(exu_n20822), .Y(exu_n901));
AND2X1 exu_U10994(.A(div_yreg_yreg_thr3[14]), .B(ecl_div_thr_e[3]), .Y(exu_n20826));
INVX1 exu_U10995(.A(exu_n20826), .Y(exu_n902));
AND2X1 exu_U10996(.A(div_yreg_yreg_thr1[14]), .B(exu_n16221), .Y(exu_n20828));
INVX1 exu_U10997(.A(exu_n20828), .Y(exu_n903));
AND2X1 exu_U10998(.A(div_yreg_yreg_thr3[13]), .B(ecl_div_thr_e[3]), .Y(exu_n20832));
INVX1 exu_U10999(.A(exu_n20832), .Y(exu_n904));
AND2X1 exu_U11000(.A(div_yreg_yreg_thr1[13]), .B(exu_n16221), .Y(exu_n20834));
INVX1 exu_U11001(.A(exu_n20834), .Y(exu_n905));
AND2X1 exu_U11002(.A(div_yreg_yreg_thr3[12]), .B(ecl_div_thr_e[3]), .Y(exu_n20838));
INVX1 exu_U11003(.A(exu_n20838), .Y(exu_n906));
AND2X1 exu_U11004(.A(div_yreg_yreg_thr1[12]), .B(exu_n16221), .Y(exu_n20840));
INVX1 exu_U11005(.A(exu_n20840), .Y(exu_n907));
AND2X1 exu_U11006(.A(div_yreg_yreg_thr3[11]), .B(ecl_div_thr_e[3]), .Y(exu_n20844));
INVX1 exu_U11007(.A(exu_n20844), .Y(exu_n908));
AND2X1 exu_U11008(.A(div_yreg_yreg_thr1[11]), .B(exu_n16221), .Y(exu_n20846));
INVX1 exu_U11009(.A(exu_n20846), .Y(exu_n909));
AND2X1 exu_U11010(.A(div_yreg_yreg_thr3[10]), .B(ecl_div_thr_e[3]), .Y(exu_n20850));
INVX1 exu_U11011(.A(exu_n20850), .Y(exu_n910));
AND2X1 exu_U11012(.A(div_yreg_yreg_thr1[10]), .B(exu_n16221), .Y(exu_n20852));
INVX1 exu_U11013(.A(exu_n20852), .Y(exu_n911));
AND2X1 exu_U11014(.A(div_yreg_div_ecl_yreg_0[3]), .B(ecl_div_thr_e[3]), .Y(exu_n20856));
INVX1 exu_U11015(.A(exu_n20856), .Y(exu_n912));
AND2X1 exu_U11016(.A(div_yreg_div_ecl_yreg_0[1]), .B(exu_n16221), .Y(exu_n20858));
INVX1 exu_U11017(.A(exu_n20858), .Y(exu_n913));
AND2X1 exu_U11018(.A(ecl_writeback_n191), .B(div_yreg_yreg_thr0[10]), .Y(exu_n20862));
INVX1 exu_U11019(.A(exu_n20862), .Y(exu_n914));
AND2X1 exu_U11020(.A(exu_n16245), .B(mul_data_out[41]), .Y(exu_n20864));
INVX1 exu_U11021(.A(exu_n20864), .Y(exu_n915));
AND2X1 exu_U11022(.A(div_yreg_yreg_thr0[9]), .B(ecl_writeback_n191), .Y(exu_n20868));
INVX1 exu_U11023(.A(exu_n20868), .Y(exu_n916));
AND2X1 exu_U11024(.A(mul_data_out[40]), .B(exu_n16245), .Y(exu_n20870));
INVX1 exu_U11025(.A(exu_n20870), .Y(exu_n917));
AND2X1 exu_U11026(.A(div_yreg_yreg_thr0[8]), .B(ecl_writeback_n191), .Y(exu_n20874));
INVX1 exu_U11027(.A(exu_n20874), .Y(exu_n918));
AND2X1 exu_U11028(.A(mul_data_out[39]), .B(exu_n16245), .Y(exu_n20876));
INVX1 exu_U11029(.A(exu_n20876), .Y(exu_n919));
AND2X1 exu_U11030(.A(div_yreg_yreg_thr0[7]), .B(ecl_writeback_n191), .Y(exu_n20880));
INVX1 exu_U11031(.A(exu_n20880), .Y(exu_n920));
AND2X1 exu_U11032(.A(mul_data_out[38]), .B(exu_n16245), .Y(exu_n20882));
INVX1 exu_U11033(.A(exu_n20882), .Y(exu_n921));
AND2X1 exu_U11034(.A(div_yreg_yreg_thr0[6]), .B(ecl_writeback_n191), .Y(exu_n20886));
INVX1 exu_U11035(.A(exu_n20886), .Y(exu_n922));
AND2X1 exu_U11036(.A(mul_data_out[37]), .B(exu_n16245), .Y(exu_n20888));
INVX1 exu_U11037(.A(exu_n20888), .Y(exu_n923));
AND2X1 exu_U11038(.A(div_yreg_yreg_thr0[5]), .B(ecl_writeback_n191), .Y(exu_n20892));
INVX1 exu_U11039(.A(exu_n20892), .Y(exu_n924));
AND2X1 exu_U11040(.A(mul_data_out[36]), .B(exu_n16245), .Y(exu_n20894));
INVX1 exu_U11041(.A(exu_n20894), .Y(exu_n925));
AND2X1 exu_U11042(.A(div_yreg_yreg_thr0[4]), .B(ecl_writeback_n191), .Y(exu_n20898));
INVX1 exu_U11043(.A(exu_n20898), .Y(exu_n926));
AND2X1 exu_U11044(.A(mul_data_out[35]), .B(exu_n16245), .Y(exu_n20900));
INVX1 exu_U11045(.A(exu_n20900), .Y(exu_n927));
AND2X1 exu_U11046(.A(ecl_div_yreg_data_31_g), .B(ecl_writeback_n191), .Y(exu_n20904));
INVX1 exu_U11047(.A(exu_n20904), .Y(exu_n928));
AND2X1 exu_U11048(.A(mul_data_out[63]), .B(exu_n16245), .Y(exu_n20906));
INVX1 exu_U11049(.A(exu_n20906), .Y(exu_n929));
AND2X1 exu_U11050(.A(div_yreg_yreg_thr0[31]), .B(ecl_writeback_n191), .Y(exu_n20910));
INVX1 exu_U11051(.A(exu_n20910), .Y(exu_n930));
AND2X1 exu_U11052(.A(mul_data_out[62]), .B(exu_n16245), .Y(exu_n20912));
INVX1 exu_U11053(.A(exu_n20912), .Y(exu_n931));
AND2X1 exu_U11054(.A(div_yreg_yreg_thr0[3]), .B(ecl_writeback_n191), .Y(exu_n20916));
INVX1 exu_U11055(.A(exu_n20916), .Y(exu_n932));
AND2X1 exu_U11056(.A(mul_data_out[34]), .B(exu_n16245), .Y(exu_n20918));
INVX1 exu_U11057(.A(exu_n20918), .Y(exu_n933));
AND2X1 exu_U11058(.A(div_yreg_yreg_thr0[30]), .B(ecl_writeback_n191), .Y(exu_n20922));
INVX1 exu_U11059(.A(exu_n20922), .Y(exu_n934));
AND2X1 exu_U11060(.A(mul_data_out[61]), .B(exu_n16245), .Y(exu_n20924));
INVX1 exu_U11061(.A(exu_n20924), .Y(exu_n935));
AND2X1 exu_U11062(.A(div_yreg_yreg_thr0[29]), .B(ecl_writeback_n191), .Y(exu_n20928));
INVX1 exu_U11063(.A(exu_n20928), .Y(exu_n936));
AND2X1 exu_U11064(.A(mul_data_out[60]), .B(exu_n16245), .Y(exu_n20930));
INVX1 exu_U11065(.A(exu_n20930), .Y(exu_n937));
AND2X1 exu_U11066(.A(div_yreg_yreg_thr0[28]), .B(ecl_writeback_n191), .Y(exu_n20934));
INVX1 exu_U11067(.A(exu_n20934), .Y(exu_n938));
AND2X1 exu_U11068(.A(mul_data_out[59]), .B(exu_n16245), .Y(exu_n20936));
INVX1 exu_U11069(.A(exu_n20936), .Y(exu_n939));
AND2X1 exu_U11070(.A(div_yreg_yreg_thr0[27]), .B(ecl_writeback_n191), .Y(exu_n20940));
INVX1 exu_U11071(.A(exu_n20940), .Y(exu_n940));
AND2X1 exu_U11072(.A(mul_data_out[58]), .B(exu_n16245), .Y(exu_n20942));
INVX1 exu_U11073(.A(exu_n20942), .Y(exu_n941));
AND2X1 exu_U11074(.A(div_yreg_yreg_thr0[26]), .B(ecl_writeback_n191), .Y(exu_n20946));
INVX1 exu_U11075(.A(exu_n20946), .Y(exu_n942));
AND2X1 exu_U11076(.A(mul_data_out[57]), .B(exu_n16245), .Y(exu_n20948));
INVX1 exu_U11077(.A(exu_n20948), .Y(exu_n943));
AND2X1 exu_U11078(.A(div_yreg_yreg_thr0[25]), .B(ecl_writeback_n191), .Y(exu_n20952));
INVX1 exu_U11079(.A(exu_n20952), .Y(exu_n944));
AND2X1 exu_U11080(.A(mul_data_out[56]), .B(exu_n16245), .Y(exu_n20954));
INVX1 exu_U11081(.A(exu_n20954), .Y(exu_n945));
AND2X1 exu_U11082(.A(div_yreg_yreg_thr0[24]), .B(ecl_writeback_n191), .Y(exu_n20958));
INVX1 exu_U11083(.A(exu_n20958), .Y(exu_n946));
AND2X1 exu_U11084(.A(mul_data_out[55]), .B(exu_n16245), .Y(exu_n20960));
INVX1 exu_U11085(.A(exu_n20960), .Y(exu_n947));
AND2X1 exu_U11086(.A(div_yreg_yreg_thr0[23]), .B(ecl_writeback_n191), .Y(exu_n20964));
INVX1 exu_U11087(.A(exu_n20964), .Y(exu_n948));
AND2X1 exu_U11088(.A(mul_data_out[54]), .B(exu_n16245), .Y(exu_n20966));
INVX1 exu_U11089(.A(exu_n20966), .Y(exu_n949));
AND2X1 exu_U11090(.A(div_yreg_yreg_thr0[22]), .B(ecl_writeback_n191), .Y(exu_n20970));
INVX1 exu_U11091(.A(exu_n20970), .Y(exu_n950));
AND2X1 exu_U11092(.A(mul_data_out[53]), .B(exu_n16245), .Y(exu_n20972));
INVX1 exu_U11093(.A(exu_n20972), .Y(exu_n951));
AND2X1 exu_U11094(.A(div_yreg_yreg_thr0[21]), .B(ecl_writeback_n191), .Y(exu_n20976));
INVX1 exu_U11095(.A(exu_n20976), .Y(exu_n952));
AND2X1 exu_U11096(.A(mul_data_out[52]), .B(exu_n16245), .Y(exu_n20978));
INVX1 exu_U11097(.A(exu_n20978), .Y(exu_n953));
AND2X1 exu_U11098(.A(div_yreg_yreg_thr0[2]), .B(ecl_writeback_n191), .Y(exu_n20982));
INVX1 exu_U11099(.A(exu_n20982), .Y(exu_n954));
AND2X1 exu_U11100(.A(mul_data_out[33]), .B(exu_n16245), .Y(exu_n20984));
INVX1 exu_U11101(.A(exu_n20984), .Y(exu_n955));
AND2X1 exu_U11102(.A(div_yreg_yreg_thr0[20]), .B(ecl_writeback_n191), .Y(exu_n20988));
INVX1 exu_U11103(.A(exu_n20988), .Y(exu_n956));
AND2X1 exu_U11104(.A(mul_data_out[51]), .B(exu_n16245), .Y(exu_n20990));
INVX1 exu_U11105(.A(exu_n20990), .Y(exu_n957));
AND2X1 exu_U11106(.A(div_yreg_yreg_thr0[19]), .B(ecl_writeback_n191), .Y(exu_n20994));
INVX1 exu_U11107(.A(exu_n20994), .Y(exu_n958));
AND2X1 exu_U11108(.A(mul_data_out[50]), .B(exu_n16245), .Y(exu_n20996));
INVX1 exu_U11109(.A(exu_n20996), .Y(exu_n959));
AND2X1 exu_U11110(.A(div_yreg_yreg_thr0[18]), .B(ecl_writeback_n191), .Y(exu_n21000));
INVX1 exu_U11111(.A(exu_n21000), .Y(exu_n960));
AND2X1 exu_U11112(.A(mul_data_out[49]), .B(exu_n16245), .Y(exu_n21002));
INVX1 exu_U11113(.A(exu_n21002), .Y(exu_n961));
AND2X1 exu_U11114(.A(div_yreg_yreg_thr0[17]), .B(ecl_writeback_n191), .Y(exu_n21006));
INVX1 exu_U11115(.A(exu_n21006), .Y(exu_n962));
AND2X1 exu_U11116(.A(mul_data_out[48]), .B(exu_n16245), .Y(exu_n21008));
INVX1 exu_U11117(.A(exu_n21008), .Y(exu_n963));
AND2X1 exu_U11118(.A(div_yreg_yreg_thr0[16]), .B(ecl_writeback_n191), .Y(exu_n21012));
INVX1 exu_U11119(.A(exu_n21012), .Y(exu_n964));
AND2X1 exu_U11120(.A(mul_data_out[47]), .B(exu_n16245), .Y(exu_n21014));
INVX1 exu_U11121(.A(exu_n21014), .Y(exu_n965));
AND2X1 exu_U11122(.A(div_yreg_yreg_thr0[15]), .B(ecl_writeback_n191), .Y(exu_n21018));
INVX1 exu_U11123(.A(exu_n21018), .Y(exu_n966));
AND2X1 exu_U11124(.A(mul_data_out[46]), .B(exu_n16245), .Y(exu_n21020));
INVX1 exu_U11125(.A(exu_n21020), .Y(exu_n967));
AND2X1 exu_U11126(.A(div_yreg_yreg_thr0[14]), .B(ecl_writeback_n191), .Y(exu_n21024));
INVX1 exu_U11127(.A(exu_n21024), .Y(exu_n968));
AND2X1 exu_U11128(.A(mul_data_out[45]), .B(exu_n16245), .Y(exu_n21026));
INVX1 exu_U11129(.A(exu_n21026), .Y(exu_n969));
AND2X1 exu_U11130(.A(div_yreg_yreg_thr0[13]), .B(ecl_writeback_n191), .Y(exu_n21030));
INVX1 exu_U11131(.A(exu_n21030), .Y(exu_n970));
AND2X1 exu_U11132(.A(mul_data_out[44]), .B(exu_n16245), .Y(exu_n21032));
INVX1 exu_U11133(.A(exu_n21032), .Y(exu_n971));
AND2X1 exu_U11134(.A(div_yreg_yreg_thr0[12]), .B(ecl_writeback_n191), .Y(exu_n21036));
INVX1 exu_U11135(.A(exu_n21036), .Y(exu_n972));
AND2X1 exu_U11136(.A(mul_data_out[43]), .B(exu_n16245), .Y(exu_n21038));
INVX1 exu_U11137(.A(exu_n21038), .Y(exu_n973));
AND2X1 exu_U11138(.A(div_yreg_yreg_thr0[11]), .B(ecl_writeback_n191), .Y(exu_n21042));
INVX1 exu_U11139(.A(exu_n21042), .Y(exu_n974));
AND2X1 exu_U11140(.A(mul_data_out[42]), .B(exu_n16245), .Y(exu_n21044));
INVX1 exu_U11141(.A(exu_n21044), .Y(exu_n975));
AND2X1 exu_U11142(.A(div_yreg_yreg_thr0[1]), .B(ecl_writeback_n191), .Y(exu_n21048));
INVX1 exu_U11143(.A(exu_n21048), .Y(exu_n976));
AND2X1 exu_U11144(.A(mul_data_out[32]), .B(exu_n16245), .Y(exu_n21050));
INVX1 exu_U11145(.A(exu_n21050), .Y(exu_n977));
AND2X1 exu_U11146(.A(ecl_writeback_n84), .B(div_yreg_yreg_thr1[10]), .Y(exu_n21054));
INVX1 exu_U11147(.A(exu_n21054), .Y(exu_n978));
AND2X1 exu_U11148(.A(exu_n15980), .B(mul_data_out[41]), .Y(exu_n21056));
INVX1 exu_U11149(.A(exu_n21056), .Y(exu_n979));
AND2X1 exu_U11150(.A(div_yreg_yreg_thr1[9]), .B(ecl_writeback_n84), .Y(exu_n21060));
INVX1 exu_U11151(.A(exu_n21060), .Y(exu_n980));
AND2X1 exu_U11152(.A(mul_data_out[40]), .B(exu_n15980), .Y(exu_n21062));
INVX1 exu_U11153(.A(exu_n21062), .Y(exu_n981));
AND2X1 exu_U11154(.A(div_yreg_yreg_thr1[8]), .B(ecl_writeback_n84), .Y(exu_n21066));
INVX1 exu_U11155(.A(exu_n21066), .Y(exu_n982));
AND2X1 exu_U11156(.A(mul_data_out[39]), .B(exu_n15980), .Y(exu_n21068));
INVX1 exu_U11157(.A(exu_n21068), .Y(exu_n983));
AND2X1 exu_U11158(.A(div_yreg_yreg_thr1[7]), .B(ecl_writeback_n84), .Y(exu_n21072));
INVX1 exu_U11159(.A(exu_n21072), .Y(exu_n984));
AND2X1 exu_U11160(.A(mul_data_out[38]), .B(exu_n15980), .Y(exu_n21074));
INVX1 exu_U11161(.A(exu_n21074), .Y(exu_n985));
AND2X1 exu_U11162(.A(div_yreg_yreg_thr1[6]), .B(ecl_writeback_n84), .Y(exu_n21078));
INVX1 exu_U11163(.A(exu_n21078), .Y(exu_n986));
AND2X1 exu_U11164(.A(mul_data_out[37]), .B(exu_n15980), .Y(exu_n21080));
INVX1 exu_U11165(.A(exu_n21080), .Y(exu_n987));
AND2X1 exu_U11166(.A(div_yreg_yreg_thr1[5]), .B(ecl_writeback_n84), .Y(exu_n21084));
INVX1 exu_U11167(.A(exu_n21084), .Y(exu_n988));
AND2X1 exu_U11168(.A(mul_data_out[36]), .B(exu_n15980), .Y(exu_n21086));
INVX1 exu_U11169(.A(exu_n21086), .Y(exu_n989));
AND2X1 exu_U11170(.A(div_yreg_yreg_thr1[4]), .B(ecl_writeback_n84), .Y(exu_n21090));
INVX1 exu_U11171(.A(exu_n21090), .Y(exu_n990));
AND2X1 exu_U11172(.A(mul_data_out[35]), .B(exu_n15980), .Y(exu_n21092));
INVX1 exu_U11173(.A(exu_n21092), .Y(exu_n991));
AND2X1 exu_U11174(.A(ecl_div_yreg_data_31_g), .B(ecl_writeback_n84), .Y(exu_n21096));
INVX1 exu_U11175(.A(exu_n21096), .Y(exu_n992));
AND2X1 exu_U11176(.A(mul_data_out[63]), .B(exu_n15980), .Y(exu_n21098));
INVX1 exu_U11177(.A(exu_n21098), .Y(exu_n993));
AND2X1 exu_U11178(.A(div_yreg_yreg_thr1[31]), .B(ecl_writeback_n84), .Y(exu_n21102));
INVX1 exu_U11179(.A(exu_n21102), .Y(exu_n994));
AND2X1 exu_U11180(.A(mul_data_out[62]), .B(exu_n15980), .Y(exu_n21104));
INVX1 exu_U11181(.A(exu_n21104), .Y(exu_n995));
AND2X1 exu_U11182(.A(div_yreg_yreg_thr1[3]), .B(ecl_writeback_n84), .Y(exu_n21108));
INVX1 exu_U11183(.A(exu_n21108), .Y(exu_n996));
AND2X1 exu_U11184(.A(mul_data_out[34]), .B(exu_n15980), .Y(exu_n21110));
INVX1 exu_U11185(.A(exu_n21110), .Y(exu_n997));
AND2X1 exu_U11186(.A(div_yreg_yreg_thr1[30]), .B(ecl_writeback_n84), .Y(exu_n21114));
INVX1 exu_U11187(.A(exu_n21114), .Y(exu_n998));
AND2X1 exu_U11188(.A(mul_data_out[61]), .B(exu_n15980), .Y(exu_n21116));
INVX1 exu_U11189(.A(exu_n21116), .Y(exu_n999));
AND2X1 exu_U11190(.A(div_yreg_yreg_thr1[29]), .B(ecl_writeback_n84), .Y(exu_n21120));
INVX1 exu_U11191(.A(exu_n21120), .Y(exu_n1000));
AND2X1 exu_U11192(.A(mul_data_out[60]), .B(exu_n15980), .Y(exu_n21122));
INVX1 exu_U11193(.A(exu_n21122), .Y(exu_n1001));
AND2X1 exu_U11194(.A(div_yreg_yreg_thr1[28]), .B(ecl_writeback_n84), .Y(exu_n21126));
INVX1 exu_U11195(.A(exu_n21126), .Y(exu_n1002));
AND2X1 exu_U11196(.A(mul_data_out[59]), .B(exu_n15980), .Y(exu_n21128));
INVX1 exu_U11197(.A(exu_n21128), .Y(exu_n1003));
AND2X1 exu_U11198(.A(div_yreg_yreg_thr1[27]), .B(ecl_writeback_n84), .Y(exu_n21132));
INVX1 exu_U11199(.A(exu_n21132), .Y(exu_n1004));
AND2X1 exu_U11200(.A(mul_data_out[58]), .B(exu_n15980), .Y(exu_n21134));
INVX1 exu_U11201(.A(exu_n21134), .Y(exu_n1005));
AND2X1 exu_U11202(.A(div_yreg_yreg_thr1[26]), .B(ecl_writeback_n84), .Y(exu_n21138));
INVX1 exu_U11203(.A(exu_n21138), .Y(exu_n1006));
AND2X1 exu_U11204(.A(mul_data_out[57]), .B(exu_n15980), .Y(exu_n21140));
INVX1 exu_U11205(.A(exu_n21140), .Y(exu_n1007));
AND2X1 exu_U11206(.A(div_yreg_yreg_thr1[25]), .B(ecl_writeback_n84), .Y(exu_n21144));
INVX1 exu_U11207(.A(exu_n21144), .Y(exu_n1008));
AND2X1 exu_U11208(.A(mul_data_out[56]), .B(exu_n15980), .Y(exu_n21146));
INVX1 exu_U11209(.A(exu_n21146), .Y(exu_n1009));
AND2X1 exu_U11210(.A(div_yreg_yreg_thr1[24]), .B(ecl_writeback_n84), .Y(exu_n21150));
INVX1 exu_U11211(.A(exu_n21150), .Y(exu_n1010));
AND2X1 exu_U11212(.A(mul_data_out[55]), .B(exu_n15980), .Y(exu_n21152));
INVX1 exu_U11213(.A(exu_n21152), .Y(exu_n1011));
AND2X1 exu_U11214(.A(div_yreg_yreg_thr1[23]), .B(ecl_writeback_n84), .Y(exu_n21156));
INVX1 exu_U11215(.A(exu_n21156), .Y(exu_n1012));
AND2X1 exu_U11216(.A(mul_data_out[54]), .B(exu_n15980), .Y(exu_n21158));
INVX1 exu_U11217(.A(exu_n21158), .Y(exu_n1013));
AND2X1 exu_U11218(.A(div_yreg_yreg_thr1[22]), .B(ecl_writeback_n84), .Y(exu_n21162));
INVX1 exu_U11219(.A(exu_n21162), .Y(exu_n1014));
AND2X1 exu_U11220(.A(mul_data_out[53]), .B(exu_n15980), .Y(exu_n21164));
INVX1 exu_U11221(.A(exu_n21164), .Y(exu_n1015));
AND2X1 exu_U11222(.A(div_yreg_yreg_thr1[21]), .B(ecl_writeback_n84), .Y(exu_n21168));
INVX1 exu_U11223(.A(exu_n21168), .Y(exu_n1016));
AND2X1 exu_U11224(.A(mul_data_out[52]), .B(exu_n15980), .Y(exu_n21170));
INVX1 exu_U11225(.A(exu_n21170), .Y(exu_n1017));
AND2X1 exu_U11226(.A(div_yreg_yreg_thr1[2]), .B(ecl_writeback_n84), .Y(exu_n21174));
INVX1 exu_U11227(.A(exu_n21174), .Y(exu_n1018));
AND2X1 exu_U11228(.A(mul_data_out[33]), .B(exu_n15980), .Y(exu_n21176));
INVX1 exu_U11229(.A(exu_n21176), .Y(exu_n1019));
AND2X1 exu_U11230(.A(div_yreg_yreg_thr1[20]), .B(ecl_writeback_n84), .Y(exu_n21180));
INVX1 exu_U11231(.A(exu_n21180), .Y(exu_n1020));
AND2X1 exu_U11232(.A(mul_data_out[51]), .B(exu_n15980), .Y(exu_n21182));
INVX1 exu_U11233(.A(exu_n21182), .Y(exu_n1021));
AND2X1 exu_U11234(.A(div_yreg_yreg_thr1[19]), .B(ecl_writeback_n84), .Y(exu_n21186));
INVX1 exu_U11235(.A(exu_n21186), .Y(exu_n1022));
AND2X1 exu_U11236(.A(mul_data_out[50]), .B(exu_n15980), .Y(exu_n21188));
INVX1 exu_U11237(.A(exu_n21188), .Y(exu_n1023));
AND2X1 exu_U11238(.A(div_yreg_yreg_thr1[18]), .B(ecl_writeback_n84), .Y(exu_n21192));
INVX1 exu_U11239(.A(exu_n21192), .Y(exu_n1024));
AND2X1 exu_U11240(.A(mul_data_out[49]), .B(exu_n15980), .Y(exu_n21194));
INVX1 exu_U11241(.A(exu_n21194), .Y(exu_n1025));
AND2X1 exu_U11242(.A(div_yreg_yreg_thr1[17]), .B(ecl_writeback_n84), .Y(exu_n21198));
INVX1 exu_U11243(.A(exu_n21198), .Y(exu_n1026));
AND2X1 exu_U11244(.A(mul_data_out[48]), .B(exu_n15980), .Y(exu_n21200));
INVX1 exu_U11245(.A(exu_n21200), .Y(exu_n1027));
AND2X1 exu_U11246(.A(div_yreg_yreg_thr1[16]), .B(ecl_writeback_n84), .Y(exu_n21204));
INVX1 exu_U11247(.A(exu_n21204), .Y(exu_n1028));
AND2X1 exu_U11248(.A(mul_data_out[47]), .B(exu_n15980), .Y(exu_n21206));
INVX1 exu_U11249(.A(exu_n21206), .Y(exu_n1029));
AND2X1 exu_U11250(.A(div_yreg_yreg_thr1[15]), .B(ecl_writeback_n84), .Y(exu_n21210));
INVX1 exu_U11251(.A(exu_n21210), .Y(exu_n1030));
AND2X1 exu_U11252(.A(mul_data_out[46]), .B(exu_n15980), .Y(exu_n21212));
INVX1 exu_U11253(.A(exu_n21212), .Y(exu_n1031));
AND2X1 exu_U11254(.A(div_yreg_yreg_thr1[14]), .B(ecl_writeback_n84), .Y(exu_n21216));
INVX1 exu_U11255(.A(exu_n21216), .Y(exu_n1032));
AND2X1 exu_U11256(.A(mul_data_out[45]), .B(exu_n15980), .Y(exu_n21218));
INVX1 exu_U11257(.A(exu_n21218), .Y(exu_n1033));
AND2X1 exu_U11258(.A(div_yreg_yreg_thr1[13]), .B(ecl_writeback_n84), .Y(exu_n21222));
INVX1 exu_U11259(.A(exu_n21222), .Y(exu_n1034));
AND2X1 exu_U11260(.A(mul_data_out[44]), .B(exu_n15980), .Y(exu_n21224));
INVX1 exu_U11261(.A(exu_n21224), .Y(exu_n1035));
AND2X1 exu_U11262(.A(div_yreg_yreg_thr1[12]), .B(ecl_writeback_n84), .Y(exu_n21228));
INVX1 exu_U11263(.A(exu_n21228), .Y(exu_n1036));
AND2X1 exu_U11264(.A(mul_data_out[43]), .B(exu_n15980), .Y(exu_n21230));
INVX1 exu_U11265(.A(exu_n21230), .Y(exu_n1037));
AND2X1 exu_U11266(.A(div_yreg_yreg_thr1[11]), .B(ecl_writeback_n84), .Y(exu_n21234));
INVX1 exu_U11267(.A(exu_n21234), .Y(exu_n1038));
AND2X1 exu_U11268(.A(mul_data_out[42]), .B(exu_n15980), .Y(exu_n21236));
INVX1 exu_U11269(.A(exu_n21236), .Y(exu_n1039));
AND2X1 exu_U11270(.A(div_yreg_yreg_thr1[1]), .B(ecl_writeback_n84), .Y(exu_n21240));
INVX1 exu_U11271(.A(exu_n21240), .Y(exu_n1040));
AND2X1 exu_U11272(.A(mul_data_out[32]), .B(exu_n15980), .Y(exu_n21242));
INVX1 exu_U11273(.A(exu_n21242), .Y(exu_n1041));
AND2X1 exu_U11274(.A(ecl_writeback_n80), .B(div_yreg_yreg_thr2[10]), .Y(exu_n21246));
INVX1 exu_U11275(.A(exu_n21246), .Y(exu_n1042));
AND2X1 exu_U11276(.A(exu_n15981), .B(mul_data_out[41]), .Y(exu_n21248));
INVX1 exu_U11277(.A(exu_n21248), .Y(exu_n1043));
AND2X1 exu_U11278(.A(div_yreg_yreg_thr2[9]), .B(ecl_writeback_n80), .Y(exu_n21252));
INVX1 exu_U11279(.A(exu_n21252), .Y(exu_n1044));
AND2X1 exu_U11280(.A(mul_data_out[40]), .B(exu_n15981), .Y(exu_n21254));
INVX1 exu_U11281(.A(exu_n21254), .Y(exu_n1045));
AND2X1 exu_U11282(.A(div_yreg_yreg_thr2[8]), .B(ecl_writeback_n80), .Y(exu_n21258));
INVX1 exu_U11283(.A(exu_n21258), .Y(exu_n1046));
AND2X1 exu_U11284(.A(mul_data_out[39]), .B(exu_n15981), .Y(exu_n21260));
INVX1 exu_U11285(.A(exu_n21260), .Y(exu_n1047));
AND2X1 exu_U11286(.A(div_yreg_yreg_thr2[7]), .B(ecl_writeback_n80), .Y(exu_n21264));
INVX1 exu_U11287(.A(exu_n21264), .Y(exu_n1048));
AND2X1 exu_U11288(.A(mul_data_out[38]), .B(exu_n15981), .Y(exu_n21266));
INVX1 exu_U11289(.A(exu_n21266), .Y(exu_n1049));
AND2X1 exu_U11290(.A(div_yreg_yreg_thr2[6]), .B(ecl_writeback_n80), .Y(exu_n21270));
INVX1 exu_U11291(.A(exu_n21270), .Y(exu_n1050));
AND2X1 exu_U11292(.A(mul_data_out[37]), .B(exu_n15981), .Y(exu_n21272));
INVX1 exu_U11293(.A(exu_n21272), .Y(exu_n1051));
AND2X1 exu_U11294(.A(div_yreg_yreg_thr2[5]), .B(ecl_writeback_n80), .Y(exu_n21276));
INVX1 exu_U11295(.A(exu_n21276), .Y(exu_n1052));
AND2X1 exu_U11296(.A(mul_data_out[36]), .B(exu_n15981), .Y(exu_n21278));
INVX1 exu_U11297(.A(exu_n21278), .Y(exu_n1053));
AND2X1 exu_U11298(.A(div_yreg_yreg_thr2[4]), .B(ecl_writeback_n80), .Y(exu_n21282));
INVX1 exu_U11299(.A(exu_n21282), .Y(exu_n1054));
AND2X1 exu_U11300(.A(mul_data_out[35]), .B(exu_n15981), .Y(exu_n21284));
INVX1 exu_U11301(.A(exu_n21284), .Y(exu_n1055));
AND2X1 exu_U11302(.A(ecl_div_yreg_data_31_g), .B(ecl_writeback_n80), .Y(exu_n21288));
INVX1 exu_U11303(.A(exu_n21288), .Y(exu_n1056));
AND2X1 exu_U11304(.A(mul_data_out[63]), .B(exu_n15981), .Y(exu_n21290));
INVX1 exu_U11305(.A(exu_n21290), .Y(exu_n1057));
AND2X1 exu_U11306(.A(div_yreg_yreg_thr2[31]), .B(ecl_writeback_n80), .Y(exu_n21294));
INVX1 exu_U11307(.A(exu_n21294), .Y(exu_n1058));
AND2X1 exu_U11308(.A(mul_data_out[62]), .B(exu_n15981), .Y(exu_n21296));
INVX1 exu_U11309(.A(exu_n21296), .Y(exu_n1059));
AND2X1 exu_U11310(.A(div_yreg_yreg_thr2[3]), .B(ecl_writeback_n80), .Y(exu_n21300));
INVX1 exu_U11311(.A(exu_n21300), .Y(exu_n1060));
AND2X1 exu_U11312(.A(mul_data_out[34]), .B(exu_n15981), .Y(exu_n21302));
INVX1 exu_U11313(.A(exu_n21302), .Y(exu_n1061));
AND2X1 exu_U11314(.A(div_yreg_yreg_thr2[30]), .B(ecl_writeback_n80), .Y(exu_n21306));
INVX1 exu_U11315(.A(exu_n21306), .Y(exu_n1062));
AND2X1 exu_U11316(.A(mul_data_out[61]), .B(exu_n15981), .Y(exu_n21308));
INVX1 exu_U11317(.A(exu_n21308), .Y(exu_n1063));
AND2X1 exu_U11318(.A(div_yreg_yreg_thr2[29]), .B(ecl_writeback_n80), .Y(exu_n21312));
INVX1 exu_U11319(.A(exu_n21312), .Y(exu_n1064));
AND2X1 exu_U11320(.A(mul_data_out[60]), .B(exu_n15981), .Y(exu_n21314));
INVX1 exu_U11321(.A(exu_n21314), .Y(exu_n1065));
AND2X1 exu_U11322(.A(div_yreg_yreg_thr2[28]), .B(ecl_writeback_n80), .Y(exu_n21318));
INVX1 exu_U11323(.A(exu_n21318), .Y(exu_n1066));
AND2X1 exu_U11324(.A(mul_data_out[59]), .B(exu_n15981), .Y(exu_n21320));
INVX1 exu_U11325(.A(exu_n21320), .Y(exu_n1067));
AND2X1 exu_U11326(.A(div_yreg_yreg_thr2[27]), .B(ecl_writeback_n80), .Y(exu_n21324));
INVX1 exu_U11327(.A(exu_n21324), .Y(exu_n1068));
AND2X1 exu_U11328(.A(mul_data_out[58]), .B(exu_n15981), .Y(exu_n21326));
INVX1 exu_U11329(.A(exu_n21326), .Y(exu_n1069));
AND2X1 exu_U11330(.A(div_yreg_yreg_thr2[26]), .B(ecl_writeback_n80), .Y(exu_n21330));
INVX1 exu_U11331(.A(exu_n21330), .Y(exu_n1070));
AND2X1 exu_U11332(.A(mul_data_out[57]), .B(exu_n15981), .Y(exu_n21332));
INVX1 exu_U11333(.A(exu_n21332), .Y(exu_n1071));
AND2X1 exu_U11334(.A(div_yreg_yreg_thr2[25]), .B(ecl_writeback_n80), .Y(exu_n21336));
INVX1 exu_U11335(.A(exu_n21336), .Y(exu_n1072));
AND2X1 exu_U11336(.A(mul_data_out[56]), .B(exu_n15981), .Y(exu_n21338));
INVX1 exu_U11337(.A(exu_n21338), .Y(exu_n1073));
AND2X1 exu_U11338(.A(div_yreg_yreg_thr2[24]), .B(ecl_writeback_n80), .Y(exu_n21342));
INVX1 exu_U11339(.A(exu_n21342), .Y(exu_n1074));
AND2X1 exu_U11340(.A(mul_data_out[55]), .B(exu_n15981), .Y(exu_n21344));
INVX1 exu_U11341(.A(exu_n21344), .Y(exu_n1075));
AND2X1 exu_U11342(.A(div_yreg_yreg_thr2[23]), .B(ecl_writeback_n80), .Y(exu_n21348));
INVX1 exu_U11343(.A(exu_n21348), .Y(exu_n1076));
AND2X1 exu_U11344(.A(mul_data_out[54]), .B(exu_n15981), .Y(exu_n21350));
INVX1 exu_U11345(.A(exu_n21350), .Y(exu_n1077));
AND2X1 exu_U11346(.A(div_yreg_yreg_thr2[22]), .B(ecl_writeback_n80), .Y(exu_n21354));
INVX1 exu_U11347(.A(exu_n21354), .Y(exu_n1078));
AND2X1 exu_U11348(.A(mul_data_out[53]), .B(exu_n15981), .Y(exu_n21356));
INVX1 exu_U11349(.A(exu_n21356), .Y(exu_n1079));
AND2X1 exu_U11350(.A(div_yreg_yreg_thr2[21]), .B(ecl_writeback_n80), .Y(exu_n21360));
INVX1 exu_U11351(.A(exu_n21360), .Y(exu_n1080));
AND2X1 exu_U11352(.A(mul_data_out[52]), .B(exu_n15981), .Y(exu_n21362));
INVX1 exu_U11353(.A(exu_n21362), .Y(exu_n1081));
AND2X1 exu_U11354(.A(div_yreg_yreg_thr2[2]), .B(ecl_writeback_n80), .Y(exu_n21366));
INVX1 exu_U11355(.A(exu_n21366), .Y(exu_n1082));
AND2X1 exu_U11356(.A(mul_data_out[33]), .B(exu_n15981), .Y(exu_n21368));
INVX1 exu_U11357(.A(exu_n21368), .Y(exu_n1083));
AND2X1 exu_U11358(.A(div_yreg_yreg_thr2[20]), .B(ecl_writeback_n80), .Y(exu_n21372));
INVX1 exu_U11359(.A(exu_n21372), .Y(exu_n1084));
AND2X1 exu_U11360(.A(mul_data_out[51]), .B(exu_n15981), .Y(exu_n21374));
INVX1 exu_U11361(.A(exu_n21374), .Y(exu_n1085));
AND2X1 exu_U11362(.A(div_yreg_yreg_thr2[19]), .B(ecl_writeback_n80), .Y(exu_n21378));
INVX1 exu_U11363(.A(exu_n21378), .Y(exu_n1086));
AND2X1 exu_U11364(.A(mul_data_out[50]), .B(exu_n15981), .Y(exu_n21380));
INVX1 exu_U11365(.A(exu_n21380), .Y(exu_n1087));
AND2X1 exu_U11366(.A(div_yreg_yreg_thr2[18]), .B(ecl_writeback_n80), .Y(exu_n21384));
INVX1 exu_U11367(.A(exu_n21384), .Y(exu_n1088));
AND2X1 exu_U11368(.A(mul_data_out[49]), .B(exu_n15981), .Y(exu_n21386));
INVX1 exu_U11369(.A(exu_n21386), .Y(exu_n1089));
AND2X1 exu_U11370(.A(div_yreg_yreg_thr2[17]), .B(ecl_writeback_n80), .Y(exu_n21390));
INVX1 exu_U11371(.A(exu_n21390), .Y(exu_n1090));
AND2X1 exu_U11372(.A(mul_data_out[48]), .B(exu_n15981), .Y(exu_n21392));
INVX1 exu_U11373(.A(exu_n21392), .Y(exu_n1091));
AND2X1 exu_U11374(.A(div_yreg_yreg_thr2[16]), .B(ecl_writeback_n80), .Y(exu_n21396));
INVX1 exu_U11375(.A(exu_n21396), .Y(exu_n1092));
AND2X1 exu_U11376(.A(mul_data_out[47]), .B(exu_n15981), .Y(exu_n21398));
INVX1 exu_U11377(.A(exu_n21398), .Y(exu_n1093));
AND2X1 exu_U11378(.A(div_yreg_yreg_thr2[15]), .B(ecl_writeback_n80), .Y(exu_n21402));
INVX1 exu_U11379(.A(exu_n21402), .Y(exu_n1094));
AND2X1 exu_U11380(.A(mul_data_out[46]), .B(exu_n15981), .Y(exu_n21404));
INVX1 exu_U11381(.A(exu_n21404), .Y(exu_n1095));
AND2X1 exu_U11382(.A(div_yreg_yreg_thr2[14]), .B(ecl_writeback_n80), .Y(exu_n21408));
INVX1 exu_U11383(.A(exu_n21408), .Y(exu_n1096));
AND2X1 exu_U11384(.A(mul_data_out[45]), .B(exu_n15981), .Y(exu_n21410));
INVX1 exu_U11385(.A(exu_n21410), .Y(exu_n1097));
AND2X1 exu_U11386(.A(div_yreg_yreg_thr2[13]), .B(ecl_writeback_n80), .Y(exu_n21414));
INVX1 exu_U11387(.A(exu_n21414), .Y(exu_n1098));
AND2X1 exu_U11388(.A(mul_data_out[44]), .B(exu_n15981), .Y(exu_n21416));
INVX1 exu_U11389(.A(exu_n21416), .Y(exu_n1099));
AND2X1 exu_U11390(.A(div_yreg_yreg_thr2[12]), .B(ecl_writeback_n80), .Y(exu_n21420));
INVX1 exu_U11391(.A(exu_n21420), .Y(exu_n1100));
AND2X1 exu_U11392(.A(mul_data_out[43]), .B(exu_n15981), .Y(exu_n21422));
INVX1 exu_U11393(.A(exu_n21422), .Y(exu_n1101));
AND2X1 exu_U11394(.A(div_yreg_yreg_thr2[11]), .B(ecl_writeback_n80), .Y(exu_n21426));
INVX1 exu_U11395(.A(exu_n21426), .Y(exu_n1102));
AND2X1 exu_U11396(.A(mul_data_out[42]), .B(exu_n15981), .Y(exu_n21428));
INVX1 exu_U11397(.A(exu_n21428), .Y(exu_n1103));
AND2X1 exu_U11398(.A(div_yreg_yreg_thr2[1]), .B(ecl_writeback_n80), .Y(exu_n21432));
INVX1 exu_U11399(.A(exu_n21432), .Y(exu_n1104));
AND2X1 exu_U11400(.A(mul_data_out[32]), .B(exu_n15981), .Y(exu_n21434));
INVX1 exu_U11401(.A(exu_n21434), .Y(exu_n1105));
AND2X1 exu_U11402(.A(ecl_writeback_n76), .B(div_yreg_yreg_thr3[10]), .Y(exu_n21438));
INVX1 exu_U11403(.A(exu_n21438), .Y(exu_n1106));
AND2X1 exu_U11404(.A(exu_n15982), .B(mul_data_out[41]), .Y(exu_n21440));
INVX1 exu_U11405(.A(exu_n21440), .Y(exu_n1107));
AND2X1 exu_U11406(.A(div_yreg_yreg_thr3[9]), .B(ecl_writeback_n76), .Y(exu_n21444));
INVX1 exu_U11407(.A(exu_n21444), .Y(exu_n1108));
AND2X1 exu_U11408(.A(mul_data_out[40]), .B(exu_n15982), .Y(exu_n21446));
INVX1 exu_U11409(.A(exu_n21446), .Y(exu_n1109));
AND2X1 exu_U11410(.A(div_yreg_yreg_thr3[8]), .B(ecl_writeback_n76), .Y(exu_n21450));
INVX1 exu_U11411(.A(exu_n21450), .Y(exu_n1110));
AND2X1 exu_U11412(.A(mul_data_out[39]), .B(exu_n15982), .Y(exu_n21452));
INVX1 exu_U11413(.A(exu_n21452), .Y(exu_n1111));
AND2X1 exu_U11414(.A(div_yreg_yreg_thr3[7]), .B(ecl_writeback_n76), .Y(exu_n21456));
INVX1 exu_U11415(.A(exu_n21456), .Y(exu_n1112));
AND2X1 exu_U11416(.A(mul_data_out[38]), .B(exu_n15982), .Y(exu_n21458));
INVX1 exu_U11417(.A(exu_n21458), .Y(exu_n1113));
AND2X1 exu_U11418(.A(div_yreg_yreg_thr3[6]), .B(ecl_writeback_n76), .Y(exu_n21462));
INVX1 exu_U11419(.A(exu_n21462), .Y(exu_n1114));
AND2X1 exu_U11420(.A(mul_data_out[37]), .B(exu_n15982), .Y(exu_n21464));
INVX1 exu_U11421(.A(exu_n21464), .Y(exu_n1115));
AND2X1 exu_U11422(.A(div_yreg_yreg_thr3[5]), .B(ecl_writeback_n76), .Y(exu_n21468));
INVX1 exu_U11423(.A(exu_n21468), .Y(exu_n1116));
AND2X1 exu_U11424(.A(mul_data_out[36]), .B(exu_n15982), .Y(exu_n21470));
INVX1 exu_U11425(.A(exu_n21470), .Y(exu_n1117));
AND2X1 exu_U11426(.A(div_yreg_yreg_thr3[4]), .B(ecl_writeback_n76), .Y(exu_n21474));
INVX1 exu_U11427(.A(exu_n21474), .Y(exu_n1118));
AND2X1 exu_U11428(.A(mul_data_out[35]), .B(exu_n15982), .Y(exu_n21476));
INVX1 exu_U11429(.A(exu_n21476), .Y(exu_n1119));
AND2X1 exu_U11430(.A(ecl_div_yreg_data_31_g), .B(ecl_writeback_n76), .Y(exu_n21480));
INVX1 exu_U11431(.A(exu_n21480), .Y(exu_n1120));
AND2X1 exu_U11432(.A(mul_data_out[63]), .B(exu_n15982), .Y(exu_n21482));
INVX1 exu_U11433(.A(exu_n21482), .Y(exu_n1121));
AND2X1 exu_U11434(.A(div_yreg_yreg_thr3[31]), .B(ecl_writeback_n76), .Y(exu_n21486));
INVX1 exu_U11435(.A(exu_n21486), .Y(exu_n1122));
AND2X1 exu_U11436(.A(mul_data_out[62]), .B(exu_n15982), .Y(exu_n21488));
INVX1 exu_U11437(.A(exu_n21488), .Y(exu_n1123));
AND2X1 exu_U11438(.A(div_yreg_yreg_thr3[3]), .B(ecl_writeback_n76), .Y(exu_n21492));
INVX1 exu_U11439(.A(exu_n21492), .Y(exu_n1124));
AND2X1 exu_U11440(.A(mul_data_out[34]), .B(exu_n15982), .Y(exu_n21494));
INVX1 exu_U11441(.A(exu_n21494), .Y(exu_n1125));
AND2X1 exu_U11442(.A(div_yreg_yreg_thr3[30]), .B(ecl_writeback_n76), .Y(exu_n21498));
INVX1 exu_U11443(.A(exu_n21498), .Y(exu_n1126));
AND2X1 exu_U11444(.A(mul_data_out[61]), .B(exu_n15982), .Y(exu_n21500));
INVX1 exu_U11445(.A(exu_n21500), .Y(exu_n1127));
AND2X1 exu_U11446(.A(div_yreg_yreg_thr3[29]), .B(ecl_writeback_n76), .Y(exu_n21504));
INVX1 exu_U11447(.A(exu_n21504), .Y(exu_n1128));
AND2X1 exu_U11448(.A(mul_data_out[60]), .B(exu_n15982), .Y(exu_n21506));
INVX1 exu_U11449(.A(exu_n21506), .Y(exu_n1129));
AND2X1 exu_U11450(.A(div_yreg_yreg_thr3[28]), .B(ecl_writeback_n76), .Y(exu_n21510));
INVX1 exu_U11451(.A(exu_n21510), .Y(exu_n1130));
AND2X1 exu_U11452(.A(mul_data_out[59]), .B(exu_n15982), .Y(exu_n21512));
INVX1 exu_U11453(.A(exu_n21512), .Y(exu_n1131));
AND2X1 exu_U11454(.A(div_yreg_yreg_thr3[27]), .B(ecl_writeback_n76), .Y(exu_n21516));
INVX1 exu_U11455(.A(exu_n21516), .Y(exu_n1132));
AND2X1 exu_U11456(.A(mul_data_out[58]), .B(exu_n15982), .Y(exu_n21518));
INVX1 exu_U11457(.A(exu_n21518), .Y(exu_n1133));
AND2X1 exu_U11458(.A(div_yreg_yreg_thr3[26]), .B(ecl_writeback_n76), .Y(exu_n21522));
INVX1 exu_U11459(.A(exu_n21522), .Y(exu_n1134));
AND2X1 exu_U11460(.A(mul_data_out[57]), .B(exu_n15982), .Y(exu_n21524));
INVX1 exu_U11461(.A(exu_n21524), .Y(exu_n1135));
AND2X1 exu_U11462(.A(div_yreg_yreg_thr3[25]), .B(ecl_writeback_n76), .Y(exu_n21528));
INVX1 exu_U11463(.A(exu_n21528), .Y(exu_n1136));
AND2X1 exu_U11464(.A(mul_data_out[56]), .B(exu_n15982), .Y(exu_n21530));
INVX1 exu_U11465(.A(exu_n21530), .Y(exu_n1137));
AND2X1 exu_U11466(.A(div_yreg_yreg_thr3[24]), .B(ecl_writeback_n76), .Y(exu_n21534));
INVX1 exu_U11467(.A(exu_n21534), .Y(exu_n1138));
AND2X1 exu_U11468(.A(mul_data_out[55]), .B(exu_n15982), .Y(exu_n21536));
INVX1 exu_U11469(.A(exu_n21536), .Y(exu_n1139));
AND2X1 exu_U11470(.A(div_yreg_yreg_thr3[23]), .B(ecl_writeback_n76), .Y(exu_n21540));
INVX1 exu_U11471(.A(exu_n21540), .Y(exu_n1140));
AND2X1 exu_U11472(.A(mul_data_out[54]), .B(exu_n15982), .Y(exu_n21542));
INVX1 exu_U11473(.A(exu_n21542), .Y(exu_n1141));
AND2X1 exu_U11474(.A(div_yreg_yreg_thr3[22]), .B(ecl_writeback_n76), .Y(exu_n21546));
INVX1 exu_U11475(.A(exu_n21546), .Y(exu_n1142));
AND2X1 exu_U11476(.A(mul_data_out[53]), .B(exu_n15982), .Y(exu_n21548));
INVX1 exu_U11477(.A(exu_n21548), .Y(exu_n1143));
AND2X1 exu_U11478(.A(div_yreg_yreg_thr3[21]), .B(ecl_writeback_n76), .Y(exu_n21552));
INVX1 exu_U11479(.A(exu_n21552), .Y(exu_n1144));
AND2X1 exu_U11480(.A(mul_data_out[52]), .B(exu_n15982), .Y(exu_n21554));
INVX1 exu_U11481(.A(exu_n21554), .Y(exu_n1145));
AND2X1 exu_U11482(.A(div_yreg_yreg_thr3[2]), .B(ecl_writeback_n76), .Y(exu_n21558));
INVX1 exu_U11483(.A(exu_n21558), .Y(exu_n1146));
AND2X1 exu_U11484(.A(mul_data_out[33]), .B(exu_n15982), .Y(exu_n21560));
INVX1 exu_U11485(.A(exu_n21560), .Y(exu_n1147));
AND2X1 exu_U11486(.A(div_yreg_yreg_thr3[20]), .B(ecl_writeback_n76), .Y(exu_n21564));
INVX1 exu_U11487(.A(exu_n21564), .Y(exu_n1148));
AND2X1 exu_U11488(.A(mul_data_out[51]), .B(exu_n15982), .Y(exu_n21566));
INVX1 exu_U11489(.A(exu_n21566), .Y(exu_n1149));
AND2X1 exu_U11490(.A(div_yreg_yreg_thr3[19]), .B(ecl_writeback_n76), .Y(exu_n21570));
INVX1 exu_U11491(.A(exu_n21570), .Y(exu_n1150));
AND2X1 exu_U11492(.A(mul_data_out[50]), .B(exu_n15982), .Y(exu_n21572));
INVX1 exu_U11493(.A(exu_n21572), .Y(exu_n1151));
AND2X1 exu_U11494(.A(div_yreg_yreg_thr3[18]), .B(ecl_writeback_n76), .Y(exu_n21576));
INVX1 exu_U11495(.A(exu_n21576), .Y(exu_n1152));
AND2X1 exu_U11496(.A(mul_data_out[49]), .B(exu_n15982), .Y(exu_n21578));
INVX1 exu_U11497(.A(exu_n21578), .Y(exu_n1153));
AND2X1 exu_U11498(.A(div_yreg_yreg_thr3[17]), .B(ecl_writeback_n76), .Y(exu_n21582));
INVX1 exu_U11499(.A(exu_n21582), .Y(exu_n1154));
AND2X1 exu_U11500(.A(mul_data_out[48]), .B(exu_n15982), .Y(exu_n21584));
INVX1 exu_U11501(.A(exu_n21584), .Y(exu_n1155));
AND2X1 exu_U11502(.A(div_yreg_yreg_thr3[16]), .B(ecl_writeback_n76), .Y(exu_n21588));
INVX1 exu_U11503(.A(exu_n21588), .Y(exu_n1156));
AND2X1 exu_U11504(.A(mul_data_out[47]), .B(exu_n15982), .Y(exu_n21590));
INVX1 exu_U11505(.A(exu_n21590), .Y(exu_n1157));
AND2X1 exu_U11506(.A(div_yreg_yreg_thr3[15]), .B(ecl_writeback_n76), .Y(exu_n21594));
INVX1 exu_U11507(.A(exu_n21594), .Y(exu_n1158));
AND2X1 exu_U11508(.A(mul_data_out[46]), .B(exu_n15982), .Y(exu_n21596));
INVX1 exu_U11509(.A(exu_n21596), .Y(exu_n1159));
AND2X1 exu_U11510(.A(div_yreg_yreg_thr3[14]), .B(ecl_writeback_n76), .Y(exu_n21600));
INVX1 exu_U11511(.A(exu_n21600), .Y(exu_n1160));
AND2X1 exu_U11512(.A(mul_data_out[45]), .B(exu_n15982), .Y(exu_n21602));
INVX1 exu_U11513(.A(exu_n21602), .Y(exu_n1161));
AND2X1 exu_U11514(.A(div_yreg_yreg_thr3[13]), .B(ecl_writeback_n76), .Y(exu_n21606));
INVX1 exu_U11515(.A(exu_n21606), .Y(exu_n1162));
AND2X1 exu_U11516(.A(mul_data_out[44]), .B(exu_n15982), .Y(exu_n21608));
INVX1 exu_U11517(.A(exu_n21608), .Y(exu_n1163));
AND2X1 exu_U11518(.A(div_yreg_yreg_thr3[12]), .B(ecl_writeback_n76), .Y(exu_n21612));
INVX1 exu_U11519(.A(exu_n21612), .Y(exu_n1164));
AND2X1 exu_U11520(.A(mul_data_out[43]), .B(exu_n15982), .Y(exu_n21614));
INVX1 exu_U11521(.A(exu_n21614), .Y(exu_n1165));
AND2X1 exu_U11522(.A(div_yreg_yreg_thr3[11]), .B(ecl_writeback_n76), .Y(exu_n21618));
INVX1 exu_U11523(.A(exu_n21618), .Y(exu_n1166));
AND2X1 exu_U11524(.A(mul_data_out[42]), .B(exu_n15982), .Y(exu_n21620));
INVX1 exu_U11525(.A(exu_n21620), .Y(exu_n1167));
AND2X1 exu_U11526(.A(div_yreg_yreg_thr3[1]), .B(ecl_writeback_n76), .Y(exu_n21624));
INVX1 exu_U11527(.A(exu_n21624), .Y(exu_n1168));
AND2X1 exu_U11528(.A(mul_data_out[32]), .B(exu_n15982), .Y(exu_n21626));
INVX1 exu_U11529(.A(exu_n21626), .Y(exu_n1169));
AND2X1 exu_U11530(.A(exu_n16284), .B(bypass_dfill_data_g2[9]), .Y(exu_n21795));
INVX1 exu_U11531(.A(exu_n21795), .Y(exu_n1170));
AND2X1 exu_U11532(.A(bypass_dfill_data_g2[8]), .B(exu_n16284), .Y(exu_n21799));
INVX1 exu_U11533(.A(exu_n21799), .Y(exu_n1171));
AND2X1 exu_U11534(.A(bypass_dfill_data_g2[7]), .B(exu_n16284), .Y(exu_n21803));
INVX1 exu_U11535(.A(exu_n21803), .Y(exu_n1172));
AND2X1 exu_U11536(.A(bypass_dfill_data_g2[6]), .B(exu_n16284), .Y(exu_n21807));
INVX1 exu_U11537(.A(exu_n21807), .Y(exu_n1173));
AND2X1 exu_U11538(.A(bypass_dfill_data_g2[63]), .B(exu_n16284), .Y(exu_n21811));
INVX1 exu_U11539(.A(exu_n21811), .Y(exu_n1174));
AND2X1 exu_U11540(.A(bypass_dfill_data_g2[62]), .B(exu_n16284), .Y(exu_n21815));
INVX1 exu_U11541(.A(exu_n21815), .Y(exu_n1175));
AND2X1 exu_U11542(.A(bypass_dfill_data_g2[61]), .B(exu_n16284), .Y(exu_n21819));
INVX1 exu_U11543(.A(exu_n21819), .Y(exu_n1176));
AND2X1 exu_U11544(.A(bypass_dfill_data_g2[60]), .B(exu_n16284), .Y(exu_n21823));
INVX1 exu_U11545(.A(exu_n21823), .Y(exu_n1177));
AND2X1 exu_U11546(.A(bypass_dfill_data_g2[5]), .B(exu_n16284), .Y(exu_n21827));
INVX1 exu_U11547(.A(exu_n21827), .Y(exu_n1178));
AND2X1 exu_U11548(.A(bypass_dfill_data_g2[59]), .B(exu_n16284), .Y(exu_n21831));
INVX1 exu_U11549(.A(exu_n21831), .Y(exu_n1179));
AND2X1 exu_U11550(.A(bypass_dfill_data_g2[58]), .B(exu_n16284), .Y(exu_n21835));
INVX1 exu_U11551(.A(exu_n21835), .Y(exu_n1180));
AND2X1 exu_U11552(.A(bypass_dfill_data_g2[57]), .B(exu_n16284), .Y(exu_n21839));
INVX1 exu_U11553(.A(exu_n21839), .Y(exu_n1181));
AND2X1 exu_U11554(.A(bypass_dfill_data_g2[56]), .B(exu_n16284), .Y(exu_n21843));
INVX1 exu_U11555(.A(exu_n21843), .Y(exu_n1182));
AND2X1 exu_U11556(.A(bypass_dfill_data_g2[55]), .B(exu_n16284), .Y(exu_n21847));
INVX1 exu_U11557(.A(exu_n21847), .Y(exu_n1183));
AND2X1 exu_U11558(.A(bypass_dfill_data_g2[54]), .B(exu_n16284), .Y(exu_n21851));
INVX1 exu_U11559(.A(exu_n21851), .Y(exu_n1184));
AND2X1 exu_U11560(.A(bypass_dfill_data_g2[53]), .B(exu_n16284), .Y(exu_n21855));
INVX1 exu_U11561(.A(exu_n21855), .Y(exu_n1185));
AND2X1 exu_U11562(.A(bypass_dfill_data_g2[52]), .B(exu_n16284), .Y(exu_n21859));
INVX1 exu_U11563(.A(exu_n21859), .Y(exu_n1186));
AND2X1 exu_U11564(.A(bypass_dfill_data_g2[51]), .B(exu_n16284), .Y(exu_n21863));
INVX1 exu_U11565(.A(exu_n21863), .Y(exu_n1187));
AND2X1 exu_U11566(.A(bypass_dfill_data_g2[50]), .B(exu_n16284), .Y(exu_n21867));
INVX1 exu_U11567(.A(exu_n21867), .Y(exu_n1188));
AND2X1 exu_U11568(.A(bypass_dfill_data_g2[4]), .B(exu_n16284), .Y(exu_n21871));
INVX1 exu_U11569(.A(exu_n21871), .Y(exu_n1189));
AND2X1 exu_U11570(.A(bypass_dfill_data_g2[49]), .B(exu_n16284), .Y(exu_n21875));
INVX1 exu_U11571(.A(exu_n21875), .Y(exu_n1190));
AND2X1 exu_U11572(.A(bypass_dfill_data_g2[48]), .B(exu_n16284), .Y(exu_n21879));
INVX1 exu_U11573(.A(exu_n21879), .Y(exu_n1191));
AND2X1 exu_U11574(.A(bypass_dfill_data_g2[47]), .B(exu_n16284), .Y(exu_n21883));
INVX1 exu_U11575(.A(exu_n21883), .Y(exu_n1192));
AND2X1 exu_U11576(.A(bypass_dfill_data_g2[46]), .B(exu_n16284), .Y(exu_n21887));
INVX1 exu_U11577(.A(exu_n21887), .Y(exu_n1193));
AND2X1 exu_U11578(.A(bypass_dfill_data_g2[45]), .B(exu_n16284), .Y(exu_n21891));
INVX1 exu_U11579(.A(exu_n21891), .Y(exu_n1194));
AND2X1 exu_U11580(.A(bypass_dfill_data_g2[44]), .B(exu_n16284), .Y(exu_n21895));
INVX1 exu_U11581(.A(exu_n21895), .Y(exu_n1195));
AND2X1 exu_U11582(.A(bypass_dfill_data_g2[43]), .B(exu_n16284), .Y(exu_n21899));
INVX1 exu_U11583(.A(exu_n21899), .Y(exu_n1196));
AND2X1 exu_U11584(.A(bypass_dfill_data_g2[42]), .B(exu_n16284), .Y(exu_n21903));
INVX1 exu_U11585(.A(exu_n21903), .Y(exu_n1197));
AND2X1 exu_U11586(.A(bypass_dfill_data_g2[41]), .B(exu_n16284), .Y(exu_n21907));
INVX1 exu_U11587(.A(exu_n21907), .Y(exu_n1198));
AND2X1 exu_U11588(.A(bypass_dfill_data_g2[40]), .B(exu_n16284), .Y(exu_n21911));
INVX1 exu_U11589(.A(exu_n21911), .Y(exu_n1199));
AND2X1 exu_U11590(.A(bypass_dfill_data_g2[3]), .B(exu_n16284), .Y(exu_n21915));
INVX1 exu_U11591(.A(exu_n21915), .Y(exu_n1200));
AND2X1 exu_U11592(.A(bypass_dfill_data_g2[39]), .B(exu_n16284), .Y(exu_n21919));
INVX1 exu_U11593(.A(exu_n21919), .Y(exu_n1201));
AND2X1 exu_U11594(.A(bypass_dfill_data_g2[38]), .B(exu_n16284), .Y(exu_n21923));
INVX1 exu_U11595(.A(exu_n21923), .Y(exu_n1202));
AND2X1 exu_U11596(.A(bypass_dfill_data_g2[37]), .B(exu_n16284), .Y(exu_n21927));
INVX1 exu_U11597(.A(exu_n21927), .Y(exu_n1203));
AND2X1 exu_U11598(.A(bypass_dfill_data_g2[36]), .B(exu_n16284), .Y(exu_n21931));
INVX1 exu_U11599(.A(exu_n21931), .Y(exu_n1204));
AND2X1 exu_U11600(.A(bypass_dfill_data_g2[35]), .B(exu_n16284), .Y(exu_n21935));
INVX1 exu_U11601(.A(exu_n21935), .Y(exu_n1205));
AND2X1 exu_U11602(.A(bypass_dfill_data_g2[34]), .B(exu_n16284), .Y(exu_n21939));
INVX1 exu_U11603(.A(exu_n21939), .Y(exu_n1206));
AND2X1 exu_U11604(.A(bypass_dfill_data_g2[33]), .B(exu_n16284), .Y(exu_n21943));
INVX1 exu_U11605(.A(exu_n21943), .Y(exu_n1207));
AND2X1 exu_U11606(.A(bypass_dfill_data_g2[32]), .B(exu_n16284), .Y(exu_n21947));
INVX1 exu_U11607(.A(exu_n21947), .Y(exu_n1208));
AND2X1 exu_U11608(.A(bypass_dfill_data_g2[31]), .B(exu_n16284), .Y(exu_n21951));
INVX1 exu_U11609(.A(exu_n21951), .Y(exu_n1209));
AND2X1 exu_U11610(.A(bypass_dfill_data_g2[30]), .B(exu_n16284), .Y(exu_n21955));
INVX1 exu_U11611(.A(exu_n21955), .Y(exu_n1210));
AND2X1 exu_U11612(.A(bypass_dfill_data_g2[2]), .B(exu_n16284), .Y(exu_n21959));
INVX1 exu_U11613(.A(exu_n21959), .Y(exu_n1211));
AND2X1 exu_U11614(.A(bypass_dfill_data_g2[29]), .B(exu_n16284), .Y(exu_n21963));
INVX1 exu_U11615(.A(exu_n21963), .Y(exu_n1212));
AND2X1 exu_U11616(.A(bypass_dfill_data_g2[28]), .B(exu_n16284), .Y(exu_n21967));
INVX1 exu_U11617(.A(exu_n21967), .Y(exu_n1213));
AND2X1 exu_U11618(.A(bypass_dfill_data_g2[27]), .B(exu_n16284), .Y(exu_n21971));
INVX1 exu_U11619(.A(exu_n21971), .Y(exu_n1214));
AND2X1 exu_U11620(.A(bypass_dfill_data_g2[26]), .B(exu_n16284), .Y(exu_n21975));
INVX1 exu_U11621(.A(exu_n21975), .Y(exu_n1215));
AND2X1 exu_U11622(.A(bypass_dfill_data_g2[25]), .B(exu_n16284), .Y(exu_n21979));
INVX1 exu_U11623(.A(exu_n21979), .Y(exu_n1216));
AND2X1 exu_U11624(.A(bypass_dfill_data_g2[24]), .B(exu_n16284), .Y(exu_n21983));
INVX1 exu_U11625(.A(exu_n21983), .Y(exu_n1217));
AND2X1 exu_U11626(.A(bypass_dfill_data_g2[23]), .B(exu_n16284), .Y(exu_n21987));
INVX1 exu_U11627(.A(exu_n21987), .Y(exu_n1218));
AND2X1 exu_U11628(.A(bypass_dfill_data_g2[22]), .B(exu_n16284), .Y(exu_n21991));
INVX1 exu_U11629(.A(exu_n21991), .Y(exu_n1219));
AND2X1 exu_U11630(.A(bypass_dfill_data_g2[21]), .B(exu_n16284), .Y(exu_n21995));
INVX1 exu_U11631(.A(exu_n21995), .Y(exu_n1220));
AND2X1 exu_U11632(.A(bypass_dfill_data_g2[20]), .B(exu_n16284), .Y(exu_n21999));
INVX1 exu_U11633(.A(exu_n21999), .Y(exu_n1221));
AND2X1 exu_U11634(.A(bypass_dfill_data_g2[1]), .B(exu_n16284), .Y(exu_n22003));
INVX1 exu_U11635(.A(exu_n22003), .Y(exu_n1222));
AND2X1 exu_U11636(.A(bypass_dfill_data_g2[19]), .B(exu_n16284), .Y(exu_n22007));
INVX1 exu_U11637(.A(exu_n22007), .Y(exu_n1223));
AND2X1 exu_U11638(.A(bypass_dfill_data_g2[18]), .B(exu_n16284), .Y(exu_n22011));
INVX1 exu_U11639(.A(exu_n22011), .Y(exu_n1224));
AND2X1 exu_U11640(.A(bypass_dfill_data_g2[17]), .B(exu_n16284), .Y(exu_n22015));
INVX1 exu_U11641(.A(exu_n22015), .Y(exu_n1225));
AND2X1 exu_U11642(.A(bypass_dfill_data_g2[16]), .B(exu_n16284), .Y(exu_n22019));
INVX1 exu_U11643(.A(exu_n22019), .Y(exu_n1226));
AND2X1 exu_U11644(.A(bypass_dfill_data_g2[15]), .B(exu_n16284), .Y(exu_n22023));
INVX1 exu_U11645(.A(exu_n22023), .Y(exu_n1227));
AND2X1 exu_U11646(.A(bypass_dfill_data_g2[14]), .B(exu_n16284), .Y(exu_n22027));
INVX1 exu_U11647(.A(exu_n22027), .Y(exu_n1228));
AND2X1 exu_U11648(.A(bypass_dfill_data_g2[13]), .B(exu_n16284), .Y(exu_n22031));
INVX1 exu_U11649(.A(exu_n22031), .Y(exu_n1229));
AND2X1 exu_U11650(.A(bypass_dfill_data_g2[12]), .B(exu_n16284), .Y(exu_n22035));
INVX1 exu_U11651(.A(exu_n22035), .Y(exu_n1230));
AND2X1 exu_U11652(.A(bypass_dfill_data_g2[11]), .B(exu_n16284), .Y(exu_n22039));
INVX1 exu_U11653(.A(exu_n22039), .Y(exu_n1231));
AND2X1 exu_U11654(.A(bypass_dfill_data_g2[10]), .B(exu_n16284), .Y(exu_n22043));
INVX1 exu_U11655(.A(exu_n22043), .Y(exu_n1232));
AND2X1 exu_U11656(.A(bypass_dfill_data_g2[0]), .B(exu_n16284), .Y(exu_n22047));
INVX1 exu_U11657(.A(exu_n22047), .Y(exu_n1233));
AND2X1 exu_U11658(.A(exu_n16281), .B(bypass_dfill_data_g2[9]), .Y(exu_n22051));
INVX1 exu_U11659(.A(exu_n22051), .Y(exu_n1234));
AND2X1 exu_U11660(.A(bypass_dfill_data_g2[8]), .B(exu_n16281), .Y(exu_n22055));
INVX1 exu_U11661(.A(exu_n22055), .Y(exu_n1235));
AND2X1 exu_U11662(.A(bypass_dfill_data_g2[7]), .B(exu_n16281), .Y(exu_n22059));
INVX1 exu_U11663(.A(exu_n22059), .Y(exu_n1236));
AND2X1 exu_U11664(.A(bypass_dfill_data_g2[6]), .B(exu_n16281), .Y(exu_n22063));
INVX1 exu_U11665(.A(exu_n22063), .Y(exu_n1237));
AND2X1 exu_U11666(.A(bypass_dfill_data_g2[63]), .B(exu_n16281), .Y(exu_n22067));
INVX1 exu_U11667(.A(exu_n22067), .Y(exu_n1238));
AND2X1 exu_U11668(.A(bypass_dfill_data_g2[62]), .B(exu_n16281), .Y(exu_n22071));
INVX1 exu_U11669(.A(exu_n22071), .Y(exu_n1239));
AND2X1 exu_U11670(.A(bypass_dfill_data_g2[61]), .B(exu_n16281), .Y(exu_n22075));
INVX1 exu_U11671(.A(exu_n22075), .Y(exu_n1240));
AND2X1 exu_U11672(.A(bypass_dfill_data_g2[60]), .B(exu_n16281), .Y(exu_n22079));
INVX1 exu_U11673(.A(exu_n22079), .Y(exu_n1241));
AND2X1 exu_U11674(.A(bypass_dfill_data_g2[5]), .B(exu_n16281), .Y(exu_n22083));
INVX1 exu_U11675(.A(exu_n22083), .Y(exu_n1242));
AND2X1 exu_U11676(.A(bypass_dfill_data_g2[59]), .B(exu_n16281), .Y(exu_n22087));
INVX1 exu_U11677(.A(exu_n22087), .Y(exu_n1243));
AND2X1 exu_U11678(.A(bypass_dfill_data_g2[58]), .B(exu_n16281), .Y(exu_n22091));
INVX1 exu_U11679(.A(exu_n22091), .Y(exu_n1244));
AND2X1 exu_U11680(.A(bypass_dfill_data_g2[57]), .B(exu_n16281), .Y(exu_n22095));
INVX1 exu_U11681(.A(exu_n22095), .Y(exu_n1245));
AND2X1 exu_U11682(.A(bypass_dfill_data_g2[56]), .B(exu_n16281), .Y(exu_n22099));
INVX1 exu_U11683(.A(exu_n22099), .Y(exu_n1246));
AND2X1 exu_U11684(.A(bypass_dfill_data_g2[55]), .B(exu_n16281), .Y(exu_n22103));
INVX1 exu_U11685(.A(exu_n22103), .Y(exu_n1247));
AND2X1 exu_U11686(.A(bypass_dfill_data_g2[54]), .B(exu_n16281), .Y(exu_n22107));
INVX1 exu_U11687(.A(exu_n22107), .Y(exu_n1248));
AND2X1 exu_U11688(.A(bypass_dfill_data_g2[53]), .B(exu_n16281), .Y(exu_n22111));
INVX1 exu_U11689(.A(exu_n22111), .Y(exu_n1249));
AND2X1 exu_U11690(.A(bypass_dfill_data_g2[52]), .B(exu_n16281), .Y(exu_n22115));
INVX1 exu_U11691(.A(exu_n22115), .Y(exu_n1250));
AND2X1 exu_U11692(.A(bypass_dfill_data_g2[51]), .B(exu_n16281), .Y(exu_n22119));
INVX1 exu_U11693(.A(exu_n22119), .Y(exu_n1251));
AND2X1 exu_U11694(.A(bypass_dfill_data_g2[50]), .B(exu_n16281), .Y(exu_n22123));
INVX1 exu_U11695(.A(exu_n22123), .Y(exu_n1252));
AND2X1 exu_U11696(.A(bypass_dfill_data_g2[4]), .B(exu_n16281), .Y(exu_n22127));
INVX1 exu_U11697(.A(exu_n22127), .Y(exu_n1253));
AND2X1 exu_U11698(.A(bypass_dfill_data_g2[49]), .B(exu_n16281), .Y(exu_n22131));
INVX1 exu_U11699(.A(exu_n22131), .Y(exu_n1254));
AND2X1 exu_U11700(.A(bypass_dfill_data_g2[48]), .B(exu_n16281), .Y(exu_n22135));
INVX1 exu_U11701(.A(exu_n22135), .Y(exu_n1255));
AND2X1 exu_U11702(.A(bypass_dfill_data_g2[47]), .B(exu_n16281), .Y(exu_n22139));
INVX1 exu_U11703(.A(exu_n22139), .Y(exu_n1256));
AND2X1 exu_U11704(.A(bypass_dfill_data_g2[46]), .B(exu_n16281), .Y(exu_n22143));
INVX1 exu_U11705(.A(exu_n22143), .Y(exu_n1257));
AND2X1 exu_U11706(.A(bypass_dfill_data_g2[45]), .B(exu_n16281), .Y(exu_n22147));
INVX1 exu_U11707(.A(exu_n22147), .Y(exu_n1258));
AND2X1 exu_U11708(.A(bypass_dfill_data_g2[44]), .B(exu_n16281), .Y(exu_n22151));
INVX1 exu_U11709(.A(exu_n22151), .Y(exu_n1259));
AND2X1 exu_U11710(.A(bypass_dfill_data_g2[43]), .B(exu_n16281), .Y(exu_n22155));
INVX1 exu_U11711(.A(exu_n22155), .Y(exu_n1260));
AND2X1 exu_U11712(.A(bypass_dfill_data_g2[42]), .B(exu_n16281), .Y(exu_n22159));
INVX1 exu_U11713(.A(exu_n22159), .Y(exu_n1261));
AND2X1 exu_U11714(.A(bypass_dfill_data_g2[41]), .B(exu_n16281), .Y(exu_n22163));
INVX1 exu_U11715(.A(exu_n22163), .Y(exu_n1262));
AND2X1 exu_U11716(.A(bypass_dfill_data_g2[40]), .B(exu_n16281), .Y(exu_n22167));
INVX1 exu_U11717(.A(exu_n22167), .Y(exu_n1263));
AND2X1 exu_U11718(.A(bypass_dfill_data_g2[3]), .B(exu_n16281), .Y(exu_n22171));
INVX1 exu_U11719(.A(exu_n22171), .Y(exu_n1264));
AND2X1 exu_U11720(.A(bypass_dfill_data_g2[39]), .B(exu_n16281), .Y(exu_n22175));
INVX1 exu_U11721(.A(exu_n22175), .Y(exu_n1265));
AND2X1 exu_U11722(.A(bypass_dfill_data_g2[38]), .B(exu_n16281), .Y(exu_n22179));
INVX1 exu_U11723(.A(exu_n22179), .Y(exu_n1266));
AND2X1 exu_U11724(.A(bypass_dfill_data_g2[37]), .B(exu_n16281), .Y(exu_n22183));
INVX1 exu_U11725(.A(exu_n22183), .Y(exu_n1267));
AND2X1 exu_U11726(.A(bypass_dfill_data_g2[36]), .B(exu_n16281), .Y(exu_n22187));
INVX1 exu_U11727(.A(exu_n22187), .Y(exu_n1268));
AND2X1 exu_U11728(.A(bypass_dfill_data_g2[35]), .B(exu_n16281), .Y(exu_n22191));
INVX1 exu_U11729(.A(exu_n22191), .Y(exu_n1269));
AND2X1 exu_U11730(.A(bypass_dfill_data_g2[34]), .B(exu_n16281), .Y(exu_n22195));
INVX1 exu_U11731(.A(exu_n22195), .Y(exu_n1270));
AND2X1 exu_U11732(.A(bypass_dfill_data_g2[33]), .B(exu_n16281), .Y(exu_n22199));
INVX1 exu_U11733(.A(exu_n22199), .Y(exu_n1271));
AND2X1 exu_U11734(.A(bypass_dfill_data_g2[32]), .B(exu_n16281), .Y(exu_n22203));
INVX1 exu_U11735(.A(exu_n22203), .Y(exu_n1272));
AND2X1 exu_U11736(.A(bypass_dfill_data_g2[31]), .B(exu_n16281), .Y(exu_n22207));
INVX1 exu_U11737(.A(exu_n22207), .Y(exu_n1273));
AND2X1 exu_U11738(.A(bypass_dfill_data_g2[30]), .B(exu_n16281), .Y(exu_n22211));
INVX1 exu_U11739(.A(exu_n22211), .Y(exu_n1274));
AND2X1 exu_U11740(.A(bypass_dfill_data_g2[2]), .B(exu_n16281), .Y(exu_n22215));
INVX1 exu_U11741(.A(exu_n22215), .Y(exu_n1275));
AND2X1 exu_U11742(.A(bypass_dfill_data_g2[29]), .B(exu_n16281), .Y(exu_n22219));
INVX1 exu_U11743(.A(exu_n22219), .Y(exu_n1276));
AND2X1 exu_U11744(.A(bypass_dfill_data_g2[28]), .B(exu_n16281), .Y(exu_n22223));
INVX1 exu_U11745(.A(exu_n22223), .Y(exu_n1277));
AND2X1 exu_U11746(.A(bypass_dfill_data_g2[27]), .B(exu_n16281), .Y(exu_n22227));
INVX1 exu_U11747(.A(exu_n22227), .Y(exu_n1278));
AND2X1 exu_U11748(.A(bypass_dfill_data_g2[26]), .B(exu_n16281), .Y(exu_n22231));
INVX1 exu_U11749(.A(exu_n22231), .Y(exu_n1279));
AND2X1 exu_U11750(.A(bypass_dfill_data_g2[25]), .B(exu_n16281), .Y(exu_n22235));
INVX1 exu_U11751(.A(exu_n22235), .Y(exu_n1280));
AND2X1 exu_U11752(.A(bypass_dfill_data_g2[24]), .B(exu_n16281), .Y(exu_n22239));
INVX1 exu_U11753(.A(exu_n22239), .Y(exu_n1281));
AND2X1 exu_U11754(.A(bypass_dfill_data_g2[23]), .B(exu_n16281), .Y(exu_n22243));
INVX1 exu_U11755(.A(exu_n22243), .Y(exu_n1282));
AND2X1 exu_U11756(.A(bypass_dfill_data_g2[22]), .B(exu_n16281), .Y(exu_n22247));
INVX1 exu_U11757(.A(exu_n22247), .Y(exu_n1283));
AND2X1 exu_U11758(.A(bypass_dfill_data_g2[21]), .B(exu_n16281), .Y(exu_n22251));
INVX1 exu_U11759(.A(exu_n22251), .Y(exu_n1284));
AND2X1 exu_U11760(.A(bypass_dfill_data_g2[20]), .B(exu_n16281), .Y(exu_n22255));
INVX1 exu_U11761(.A(exu_n22255), .Y(exu_n1285));
AND2X1 exu_U11762(.A(bypass_dfill_data_g2[1]), .B(exu_n16281), .Y(exu_n22259));
INVX1 exu_U11763(.A(exu_n22259), .Y(exu_n1286));
AND2X1 exu_U11764(.A(bypass_dfill_data_g2[19]), .B(exu_n16281), .Y(exu_n22263));
INVX1 exu_U11765(.A(exu_n22263), .Y(exu_n1287));
AND2X1 exu_U11766(.A(bypass_dfill_data_g2[18]), .B(exu_n16281), .Y(exu_n22267));
INVX1 exu_U11767(.A(exu_n22267), .Y(exu_n1288));
AND2X1 exu_U11768(.A(bypass_dfill_data_g2[17]), .B(exu_n16281), .Y(exu_n22271));
INVX1 exu_U11769(.A(exu_n22271), .Y(exu_n1289));
AND2X1 exu_U11770(.A(bypass_dfill_data_g2[16]), .B(exu_n16281), .Y(exu_n22275));
INVX1 exu_U11771(.A(exu_n22275), .Y(exu_n1290));
AND2X1 exu_U11772(.A(bypass_dfill_data_g2[15]), .B(exu_n16281), .Y(exu_n22279));
INVX1 exu_U11773(.A(exu_n22279), .Y(exu_n1291));
AND2X1 exu_U11774(.A(bypass_dfill_data_g2[14]), .B(exu_n16281), .Y(exu_n22283));
INVX1 exu_U11775(.A(exu_n22283), .Y(exu_n1292));
AND2X1 exu_U11776(.A(bypass_dfill_data_g2[13]), .B(exu_n16281), .Y(exu_n22287));
INVX1 exu_U11777(.A(exu_n22287), .Y(exu_n1293));
AND2X1 exu_U11778(.A(bypass_dfill_data_g2[12]), .B(exu_n16281), .Y(exu_n22291));
INVX1 exu_U11779(.A(exu_n22291), .Y(exu_n1294));
AND2X1 exu_U11780(.A(bypass_dfill_data_g2[11]), .B(exu_n16281), .Y(exu_n22295));
INVX1 exu_U11781(.A(exu_n22295), .Y(exu_n1295));
AND2X1 exu_U11782(.A(bypass_dfill_data_g2[10]), .B(exu_n16281), .Y(exu_n22299));
INVX1 exu_U11783(.A(exu_n22299), .Y(exu_n1296));
AND2X1 exu_U11784(.A(bypass_dfill_data_g2[0]), .B(exu_n16281), .Y(exu_n22303));
INVX1 exu_U11785(.A(exu_n22303), .Y(exu_n1297));
AND2X1 exu_U11786(.A(exu_n16278), .B(bypass_dfill_data_g2[9]), .Y(exu_n22307));
INVX1 exu_U11787(.A(exu_n22307), .Y(exu_n1298));
AND2X1 exu_U11788(.A(exu_n22309), .B(exu_n10002), .Y(bypass_rs3_data_w2[8]));
INVX1 exu_U11789(.A(bypass_rs3_data_w2[8]), .Y(exu_n1299));
AND2X1 exu_U11790(.A(bypass_dfill_data_g2[8]), .B(exu_n16278), .Y(exu_n22311));
INVX1 exu_U11791(.A(exu_n22311), .Y(exu_n1300));
AND2X1 exu_U11792(.A(exu_n22313), .B(exu_n10003), .Y(bypass_rs3_data_w2[7]));
INVX1 exu_U11793(.A(bypass_rs3_data_w2[7]), .Y(exu_n1301));
AND2X1 exu_U11794(.A(bypass_dfill_data_g2[7]), .B(exu_n16278), .Y(exu_n22315));
INVX1 exu_U11795(.A(exu_n22315), .Y(exu_n1302));
AND2X1 exu_U11796(.A(exu_n22317), .B(exu_n10004), .Y(bypass_rs3_data_w2[6]));
INVX1 exu_U11797(.A(bypass_rs3_data_w2[6]), .Y(exu_n1303));
AND2X1 exu_U11798(.A(bypass_dfill_data_g2[6]), .B(exu_n16278), .Y(exu_n22319));
INVX1 exu_U11799(.A(exu_n22319), .Y(exu_n1304));
AND2X1 exu_U11800(.A(exu_n22321), .B(exu_n10005), .Y(bypass_rs3_data_w2[63]));
INVX1 exu_U11801(.A(bypass_rs3_data_w2[63]), .Y(exu_n1305));
AND2X1 exu_U11802(.A(bypass_dfill_data_g2[63]), .B(exu_n16278), .Y(exu_n22323));
INVX1 exu_U11803(.A(exu_n22323), .Y(exu_n1306));
AND2X1 exu_U11804(.A(exu_n22325), .B(exu_n10006), .Y(bypass_rs3_data_w2[62]));
INVX1 exu_U11805(.A(bypass_rs3_data_w2[62]), .Y(exu_n1307));
AND2X1 exu_U11806(.A(bypass_dfill_data_g2[62]), .B(exu_n16278), .Y(exu_n22327));
INVX1 exu_U11807(.A(exu_n22327), .Y(exu_n1308));
AND2X1 exu_U11808(.A(exu_n22329), .B(exu_n10007), .Y(bypass_rs3_data_w2[61]));
INVX1 exu_U11809(.A(bypass_rs3_data_w2[61]), .Y(exu_n1309));
AND2X1 exu_U11810(.A(bypass_dfill_data_g2[61]), .B(exu_n16278), .Y(exu_n22331));
INVX1 exu_U11811(.A(exu_n22331), .Y(exu_n1310));
AND2X1 exu_U11812(.A(exu_n22333), .B(exu_n10008), .Y(bypass_rs3_data_w2[60]));
INVX1 exu_U11813(.A(bypass_rs3_data_w2[60]), .Y(exu_n1311));
AND2X1 exu_U11814(.A(bypass_dfill_data_g2[60]), .B(exu_n16278), .Y(exu_n22335));
INVX1 exu_U11815(.A(exu_n22335), .Y(exu_n1312));
AND2X1 exu_U11816(.A(exu_n22337), .B(exu_n10009), .Y(bypass_rs3_data_w2[5]));
INVX1 exu_U11817(.A(bypass_rs3_data_w2[5]), .Y(exu_n1313));
AND2X1 exu_U11818(.A(bypass_dfill_data_g2[5]), .B(exu_n16278), .Y(exu_n22339));
INVX1 exu_U11819(.A(exu_n22339), .Y(exu_n1314));
AND2X1 exu_U11820(.A(exu_n22341), .B(exu_n10010), .Y(bypass_rs3_data_w2[59]));
INVX1 exu_U11821(.A(bypass_rs3_data_w2[59]), .Y(exu_n1315));
AND2X1 exu_U11822(.A(bypass_dfill_data_g2[59]), .B(exu_n16278), .Y(exu_n22343));
INVX1 exu_U11823(.A(exu_n22343), .Y(exu_n1316));
AND2X1 exu_U11824(.A(exu_n22345), .B(exu_n10011), .Y(bypass_rs3_data_w2[58]));
INVX1 exu_U11825(.A(bypass_rs3_data_w2[58]), .Y(exu_n1317));
AND2X1 exu_U11826(.A(bypass_dfill_data_g2[58]), .B(exu_n16278), .Y(exu_n22347));
INVX1 exu_U11827(.A(exu_n22347), .Y(exu_n1318));
AND2X1 exu_U11828(.A(exu_n22349), .B(exu_n10012), .Y(bypass_rs3_data_w2[57]));
INVX1 exu_U11829(.A(bypass_rs3_data_w2[57]), .Y(exu_n1319));
AND2X1 exu_U11830(.A(bypass_dfill_data_g2[57]), .B(exu_n16278), .Y(exu_n22351));
INVX1 exu_U11831(.A(exu_n22351), .Y(exu_n1320));
AND2X1 exu_U11832(.A(exu_n22353), .B(exu_n10013), .Y(bypass_rs3_data_w2[56]));
INVX1 exu_U11833(.A(bypass_rs3_data_w2[56]), .Y(exu_n1321));
AND2X1 exu_U11834(.A(bypass_dfill_data_g2[56]), .B(exu_n16278), .Y(exu_n22355));
INVX1 exu_U11835(.A(exu_n22355), .Y(exu_n1322));
AND2X1 exu_U11836(.A(exu_n22357), .B(exu_n10014), .Y(bypass_rs3_data_w2[55]));
INVX1 exu_U11837(.A(bypass_rs3_data_w2[55]), .Y(exu_n1323));
AND2X1 exu_U11838(.A(bypass_dfill_data_g2[55]), .B(exu_n16278), .Y(exu_n22359));
INVX1 exu_U11839(.A(exu_n22359), .Y(exu_n1324));
AND2X1 exu_U11840(.A(exu_n22361), .B(exu_n10015), .Y(bypass_rs3_data_w2[54]));
INVX1 exu_U11841(.A(bypass_rs3_data_w2[54]), .Y(exu_n1325));
AND2X1 exu_U11842(.A(bypass_dfill_data_g2[54]), .B(exu_n16278), .Y(exu_n22363));
INVX1 exu_U11843(.A(exu_n22363), .Y(exu_n1326));
AND2X1 exu_U11844(.A(exu_n22365), .B(exu_n10016), .Y(bypass_rs3_data_w2[53]));
INVX1 exu_U11845(.A(bypass_rs3_data_w2[53]), .Y(exu_n1327));
AND2X1 exu_U11846(.A(bypass_dfill_data_g2[53]), .B(exu_n16278), .Y(exu_n22367));
INVX1 exu_U11847(.A(exu_n22367), .Y(exu_n1328));
AND2X1 exu_U11848(.A(exu_n22369), .B(exu_n10017), .Y(bypass_rs3_data_w2[52]));
INVX1 exu_U11849(.A(bypass_rs3_data_w2[52]), .Y(exu_n1329));
AND2X1 exu_U11850(.A(bypass_dfill_data_g2[52]), .B(exu_n16278), .Y(exu_n22371));
INVX1 exu_U11851(.A(exu_n22371), .Y(exu_n1330));
AND2X1 exu_U11852(.A(exu_n22373), .B(exu_n10018), .Y(bypass_rs3_data_w2[51]));
INVX1 exu_U11853(.A(bypass_rs3_data_w2[51]), .Y(exu_n1331));
AND2X1 exu_U11854(.A(bypass_dfill_data_g2[51]), .B(exu_n16278), .Y(exu_n22375));
INVX1 exu_U11855(.A(exu_n22375), .Y(exu_n1332));
AND2X1 exu_U11856(.A(exu_n22377), .B(exu_n10019), .Y(bypass_rs3_data_w2[50]));
INVX1 exu_U11857(.A(bypass_rs3_data_w2[50]), .Y(exu_n1333));
AND2X1 exu_U11858(.A(bypass_dfill_data_g2[50]), .B(exu_n16278), .Y(exu_n22379));
INVX1 exu_U11859(.A(exu_n22379), .Y(exu_n1334));
AND2X1 exu_U11860(.A(exu_n22381), .B(exu_n10020), .Y(bypass_rs3_data_w2[4]));
INVX1 exu_U11861(.A(bypass_rs3_data_w2[4]), .Y(exu_n1335));
AND2X1 exu_U11862(.A(bypass_dfill_data_g2[4]), .B(exu_n16278), .Y(exu_n22383));
INVX1 exu_U11863(.A(exu_n22383), .Y(exu_n1336));
AND2X1 exu_U11864(.A(exu_n22385), .B(exu_n10021), .Y(bypass_rs3_data_w2[49]));
INVX1 exu_U11865(.A(bypass_rs3_data_w2[49]), .Y(exu_n1337));
AND2X1 exu_U11866(.A(bypass_dfill_data_g2[49]), .B(exu_n16278), .Y(exu_n22387));
INVX1 exu_U11867(.A(exu_n22387), .Y(exu_n1338));
AND2X1 exu_U11868(.A(exu_n22389), .B(exu_n10022), .Y(bypass_rs3_data_w2[48]));
INVX1 exu_U11869(.A(bypass_rs3_data_w2[48]), .Y(exu_n1339));
AND2X1 exu_U11870(.A(bypass_dfill_data_g2[48]), .B(exu_n16278), .Y(exu_n22391));
INVX1 exu_U11871(.A(exu_n22391), .Y(exu_n1340));
AND2X1 exu_U11872(.A(exu_n22393), .B(exu_n10023), .Y(bypass_rs3_data_w2[47]));
INVX1 exu_U11873(.A(bypass_rs3_data_w2[47]), .Y(exu_n1341));
AND2X1 exu_U11874(.A(bypass_dfill_data_g2[47]), .B(exu_n16278), .Y(exu_n22395));
INVX1 exu_U11875(.A(exu_n22395), .Y(exu_n1342));
AND2X1 exu_U11876(.A(exu_n22397), .B(exu_n10024), .Y(bypass_rs3_data_w2[46]));
INVX1 exu_U11877(.A(bypass_rs3_data_w2[46]), .Y(exu_n1343));
AND2X1 exu_U11878(.A(bypass_dfill_data_g2[46]), .B(exu_n16278), .Y(exu_n22399));
INVX1 exu_U11879(.A(exu_n22399), .Y(exu_n1344));
AND2X1 exu_U11880(.A(exu_n22401), .B(exu_n10025), .Y(bypass_rs3_data_w2[45]));
INVX1 exu_U11881(.A(bypass_rs3_data_w2[45]), .Y(exu_n1345));
AND2X1 exu_U11882(.A(bypass_dfill_data_g2[45]), .B(exu_n16278), .Y(exu_n22403));
INVX1 exu_U11883(.A(exu_n22403), .Y(exu_n1346));
AND2X1 exu_U11884(.A(exu_n22405), .B(exu_n10026), .Y(bypass_rs3_data_w2[44]));
INVX1 exu_U11885(.A(bypass_rs3_data_w2[44]), .Y(exu_n1347));
AND2X1 exu_U11886(.A(bypass_dfill_data_g2[44]), .B(exu_n16278), .Y(exu_n22407));
INVX1 exu_U11887(.A(exu_n22407), .Y(exu_n1348));
AND2X1 exu_U11888(.A(exu_n22409), .B(exu_n10027), .Y(bypass_rs3_data_w2[43]));
INVX1 exu_U11889(.A(bypass_rs3_data_w2[43]), .Y(exu_n1349));
AND2X1 exu_U11890(.A(bypass_dfill_data_g2[43]), .B(exu_n16278), .Y(exu_n22411));
INVX1 exu_U11891(.A(exu_n22411), .Y(exu_n1350));
AND2X1 exu_U11892(.A(exu_n22413), .B(exu_n10028), .Y(bypass_rs3_data_w2[42]));
INVX1 exu_U11893(.A(bypass_rs3_data_w2[42]), .Y(exu_n1351));
AND2X1 exu_U11894(.A(bypass_dfill_data_g2[42]), .B(exu_n16278), .Y(exu_n22415));
INVX1 exu_U11895(.A(exu_n22415), .Y(exu_n1352));
AND2X1 exu_U11896(.A(exu_n22417), .B(exu_n10029), .Y(bypass_rs3_data_w2[41]));
INVX1 exu_U11897(.A(bypass_rs3_data_w2[41]), .Y(exu_n1353));
AND2X1 exu_U11898(.A(bypass_dfill_data_g2[41]), .B(exu_n16278), .Y(exu_n22419));
INVX1 exu_U11899(.A(exu_n22419), .Y(exu_n1354));
AND2X1 exu_U11900(.A(exu_n22421), .B(exu_n10030), .Y(bypass_rs3_data_w2[40]));
INVX1 exu_U11901(.A(bypass_rs3_data_w2[40]), .Y(exu_n1355));
AND2X1 exu_U11902(.A(bypass_dfill_data_g2[40]), .B(exu_n16278), .Y(exu_n22423));
INVX1 exu_U11903(.A(exu_n22423), .Y(exu_n1356));
AND2X1 exu_U11904(.A(exu_n22425), .B(exu_n10031), .Y(bypass_rs3_data_w2[3]));
INVX1 exu_U11905(.A(bypass_rs3_data_w2[3]), .Y(exu_n1357));
AND2X1 exu_U11906(.A(bypass_dfill_data_g2[3]), .B(exu_n16278), .Y(exu_n22427));
INVX1 exu_U11907(.A(exu_n22427), .Y(exu_n1358));
AND2X1 exu_U11908(.A(exu_n22429), .B(exu_n10032), .Y(bypass_rs3_data_w2[39]));
INVX1 exu_U11909(.A(bypass_rs3_data_w2[39]), .Y(exu_n1359));
AND2X1 exu_U11910(.A(bypass_dfill_data_g2[39]), .B(exu_n16278), .Y(exu_n22431));
INVX1 exu_U11911(.A(exu_n22431), .Y(exu_n1360));
AND2X1 exu_U11912(.A(exu_n22433), .B(exu_n10033), .Y(bypass_rs3_data_w2[38]));
INVX1 exu_U11913(.A(bypass_rs3_data_w2[38]), .Y(exu_n1361));
AND2X1 exu_U11914(.A(bypass_dfill_data_g2[38]), .B(exu_n16278), .Y(exu_n22435));
INVX1 exu_U11915(.A(exu_n22435), .Y(exu_n1362));
AND2X1 exu_U11916(.A(exu_n22437), .B(exu_n10034), .Y(bypass_rs3_data_w2[37]));
INVX1 exu_U11917(.A(bypass_rs3_data_w2[37]), .Y(exu_n1363));
AND2X1 exu_U11918(.A(bypass_dfill_data_g2[37]), .B(exu_n16278), .Y(exu_n22439));
INVX1 exu_U11919(.A(exu_n22439), .Y(exu_n1364));
AND2X1 exu_U11920(.A(exu_n22441), .B(exu_n10035), .Y(bypass_rs3_data_w2[36]));
INVX1 exu_U11921(.A(bypass_rs3_data_w2[36]), .Y(exu_n1365));
AND2X1 exu_U11922(.A(bypass_dfill_data_g2[36]), .B(exu_n16278), .Y(exu_n22443));
INVX1 exu_U11923(.A(exu_n22443), .Y(exu_n1366));
AND2X1 exu_U11924(.A(exu_n22445), .B(exu_n10036), .Y(bypass_rs3_data_w2[35]));
INVX1 exu_U11925(.A(bypass_rs3_data_w2[35]), .Y(exu_n1367));
AND2X1 exu_U11926(.A(bypass_dfill_data_g2[35]), .B(exu_n16278), .Y(exu_n22447));
INVX1 exu_U11927(.A(exu_n22447), .Y(exu_n1368));
AND2X1 exu_U11928(.A(exu_n22449), .B(exu_n10037), .Y(bypass_rs3_data_w2[34]));
INVX1 exu_U11929(.A(bypass_rs3_data_w2[34]), .Y(exu_n1369));
AND2X1 exu_U11930(.A(bypass_dfill_data_g2[34]), .B(exu_n16278), .Y(exu_n22451));
INVX1 exu_U11931(.A(exu_n22451), .Y(exu_n1370));
AND2X1 exu_U11932(.A(exu_n22453), .B(exu_n10038), .Y(bypass_rs3_data_w2[33]));
INVX1 exu_U11933(.A(bypass_rs3_data_w2[33]), .Y(exu_n1371));
AND2X1 exu_U11934(.A(bypass_dfill_data_g2[33]), .B(exu_n16278), .Y(exu_n22455));
INVX1 exu_U11935(.A(exu_n22455), .Y(exu_n1372));
AND2X1 exu_U11936(.A(exu_n22457), .B(exu_n10039), .Y(bypass_rs3_data_w2[32]));
INVX1 exu_U11937(.A(bypass_rs3_data_w2[32]), .Y(exu_n1373));
AND2X1 exu_U11938(.A(bypass_dfill_data_g2[32]), .B(exu_n16278), .Y(exu_n22459));
INVX1 exu_U11939(.A(exu_n22459), .Y(exu_n1374));
AND2X1 exu_U11940(.A(exu_n22461), .B(exu_n10040), .Y(bypass_rs3_data_w2[31]));
INVX1 exu_U11941(.A(bypass_rs3_data_w2[31]), .Y(exu_n1375));
AND2X1 exu_U11942(.A(bypass_dfill_data_g2[31]), .B(exu_n16278), .Y(exu_n22463));
INVX1 exu_U11943(.A(exu_n22463), .Y(exu_n1376));
AND2X1 exu_U11944(.A(exu_n22465), .B(exu_n10041), .Y(bypass_rs3_data_w2[30]));
INVX1 exu_U11945(.A(bypass_rs3_data_w2[30]), .Y(exu_n1377));
AND2X1 exu_U11946(.A(bypass_dfill_data_g2[30]), .B(exu_n16278), .Y(exu_n22467));
INVX1 exu_U11947(.A(exu_n22467), .Y(exu_n1378));
AND2X1 exu_U11948(.A(exu_n22469), .B(exu_n10042), .Y(bypass_rs3_data_w2[2]));
INVX1 exu_U11949(.A(bypass_rs3_data_w2[2]), .Y(exu_n1379));
AND2X1 exu_U11950(.A(bypass_dfill_data_g2[2]), .B(exu_n16278), .Y(exu_n22471));
INVX1 exu_U11951(.A(exu_n22471), .Y(exu_n1380));
AND2X1 exu_U11952(.A(exu_n22473), .B(exu_n10043), .Y(bypass_rs3_data_w2[29]));
INVX1 exu_U11953(.A(bypass_rs3_data_w2[29]), .Y(exu_n1381));
AND2X1 exu_U11954(.A(bypass_dfill_data_g2[29]), .B(exu_n16278), .Y(exu_n22475));
INVX1 exu_U11955(.A(exu_n22475), .Y(exu_n1382));
AND2X1 exu_U11956(.A(exu_n22477), .B(exu_n10044), .Y(bypass_rs3_data_w2[28]));
INVX1 exu_U11957(.A(bypass_rs3_data_w2[28]), .Y(exu_n1383));
AND2X1 exu_U11958(.A(bypass_dfill_data_g2[28]), .B(exu_n16278), .Y(exu_n22479));
INVX1 exu_U11959(.A(exu_n22479), .Y(exu_n1384));
AND2X1 exu_U11960(.A(exu_n22481), .B(exu_n10045), .Y(bypass_rs3_data_w2[27]));
INVX1 exu_U11961(.A(bypass_rs3_data_w2[27]), .Y(exu_n1385));
AND2X1 exu_U11962(.A(bypass_dfill_data_g2[27]), .B(exu_n16278), .Y(exu_n22483));
INVX1 exu_U11963(.A(exu_n22483), .Y(exu_n1386));
AND2X1 exu_U11964(.A(exu_n22485), .B(exu_n10046), .Y(bypass_rs3_data_w2[26]));
INVX1 exu_U11965(.A(bypass_rs3_data_w2[26]), .Y(exu_n1387));
AND2X1 exu_U11966(.A(bypass_dfill_data_g2[26]), .B(exu_n16278), .Y(exu_n22487));
INVX1 exu_U11967(.A(exu_n22487), .Y(exu_n1388));
AND2X1 exu_U11968(.A(exu_n22489), .B(exu_n10047), .Y(bypass_rs3_data_w2[25]));
INVX1 exu_U11969(.A(bypass_rs3_data_w2[25]), .Y(exu_n1389));
AND2X1 exu_U11970(.A(bypass_dfill_data_g2[25]), .B(exu_n16278), .Y(exu_n22491));
INVX1 exu_U11971(.A(exu_n22491), .Y(exu_n1390));
AND2X1 exu_U11972(.A(exu_n22493), .B(exu_n10048), .Y(bypass_rs3_data_w2[24]));
INVX1 exu_U11973(.A(bypass_rs3_data_w2[24]), .Y(exu_n1391));
AND2X1 exu_U11974(.A(bypass_dfill_data_g2[24]), .B(exu_n16278), .Y(exu_n22495));
INVX1 exu_U11975(.A(exu_n22495), .Y(exu_n1392));
AND2X1 exu_U11976(.A(exu_n22497), .B(exu_n10049), .Y(bypass_rs3_data_w2[23]));
INVX1 exu_U11977(.A(bypass_rs3_data_w2[23]), .Y(exu_n1393));
AND2X1 exu_U11978(.A(bypass_dfill_data_g2[23]), .B(exu_n16278), .Y(exu_n22499));
INVX1 exu_U11979(.A(exu_n22499), .Y(exu_n1394));
AND2X1 exu_U11980(.A(exu_n22501), .B(exu_n10050), .Y(bypass_rs3_data_w2[22]));
INVX1 exu_U11981(.A(bypass_rs3_data_w2[22]), .Y(exu_n1395));
AND2X1 exu_U11982(.A(bypass_dfill_data_g2[22]), .B(exu_n16278), .Y(exu_n22503));
INVX1 exu_U11983(.A(exu_n22503), .Y(exu_n1396));
AND2X1 exu_U11984(.A(exu_n22505), .B(exu_n10051), .Y(bypass_rs3_data_w2[21]));
INVX1 exu_U11985(.A(bypass_rs3_data_w2[21]), .Y(exu_n1397));
AND2X1 exu_U11986(.A(bypass_dfill_data_g2[21]), .B(exu_n16278), .Y(exu_n22507));
INVX1 exu_U11987(.A(exu_n22507), .Y(exu_n1398));
AND2X1 exu_U11988(.A(exu_n22509), .B(exu_n10052), .Y(bypass_rs3_data_w2[20]));
INVX1 exu_U11989(.A(bypass_rs3_data_w2[20]), .Y(exu_n1399));
AND2X1 exu_U11990(.A(bypass_dfill_data_g2[20]), .B(exu_n16278), .Y(exu_n22511));
INVX1 exu_U11991(.A(exu_n22511), .Y(exu_n1400));
AND2X1 exu_U11992(.A(exu_n22513), .B(exu_n10053), .Y(bypass_rs3_data_w2[1]));
INVX1 exu_U11993(.A(bypass_rs3_data_w2[1]), .Y(exu_n1401));
AND2X1 exu_U11994(.A(bypass_dfill_data_g2[1]), .B(exu_n16278), .Y(exu_n22515));
INVX1 exu_U11995(.A(exu_n22515), .Y(exu_n1402));
AND2X1 exu_U11996(.A(exu_n22517), .B(exu_n10054), .Y(bypass_rs3_data_w2[19]));
INVX1 exu_U11997(.A(bypass_rs3_data_w2[19]), .Y(exu_n1403));
AND2X1 exu_U11998(.A(bypass_dfill_data_g2[19]), .B(exu_n16278), .Y(exu_n22519));
INVX1 exu_U11999(.A(exu_n22519), .Y(exu_n1404));
AND2X1 exu_U12000(.A(exu_n22521), .B(exu_n10055), .Y(bypass_rs3_data_w2[18]));
INVX1 exu_U12001(.A(bypass_rs3_data_w2[18]), .Y(exu_n1405));
AND2X1 exu_U12002(.A(bypass_dfill_data_g2[18]), .B(exu_n16278), .Y(exu_n22523));
INVX1 exu_U12003(.A(exu_n22523), .Y(exu_n1406));
AND2X1 exu_U12004(.A(exu_n22525), .B(exu_n10056), .Y(bypass_rs3_data_w2[17]));
INVX1 exu_U12005(.A(bypass_rs3_data_w2[17]), .Y(exu_n1407));
AND2X1 exu_U12006(.A(bypass_dfill_data_g2[17]), .B(exu_n16278), .Y(exu_n22527));
INVX1 exu_U12007(.A(exu_n22527), .Y(exu_n1408));
AND2X1 exu_U12008(.A(exu_n22529), .B(exu_n10057), .Y(bypass_rs3_data_w2[16]));
INVX1 exu_U12009(.A(bypass_rs3_data_w2[16]), .Y(exu_n1409));
AND2X1 exu_U12010(.A(bypass_dfill_data_g2[16]), .B(exu_n16278), .Y(exu_n22531));
INVX1 exu_U12011(.A(exu_n22531), .Y(exu_n1410));
AND2X1 exu_U12012(.A(exu_n22533), .B(exu_n10058), .Y(bypass_rs3_data_w2[15]));
INVX1 exu_U12013(.A(bypass_rs3_data_w2[15]), .Y(exu_n1411));
AND2X1 exu_U12014(.A(bypass_dfill_data_g2[15]), .B(exu_n16278), .Y(exu_n22535));
INVX1 exu_U12015(.A(exu_n22535), .Y(exu_n1412));
AND2X1 exu_U12016(.A(exu_n22537), .B(exu_n10059), .Y(bypass_rs3_data_w2[14]));
INVX1 exu_U12017(.A(bypass_rs3_data_w2[14]), .Y(exu_n1413));
AND2X1 exu_U12018(.A(bypass_dfill_data_g2[14]), .B(exu_n16278), .Y(exu_n22539));
INVX1 exu_U12019(.A(exu_n22539), .Y(exu_n1414));
AND2X1 exu_U12020(.A(exu_n22541), .B(exu_n10060), .Y(bypass_rs3_data_w2[13]));
INVX1 exu_U12021(.A(bypass_rs3_data_w2[13]), .Y(exu_n1415));
AND2X1 exu_U12022(.A(bypass_dfill_data_g2[13]), .B(exu_n16278), .Y(exu_n22543));
INVX1 exu_U12023(.A(exu_n22543), .Y(exu_n1416));
AND2X1 exu_U12024(.A(exu_n22545), .B(exu_n10061), .Y(bypass_rs3_data_w2[12]));
INVX1 exu_U12025(.A(bypass_rs3_data_w2[12]), .Y(exu_n1417));
AND2X1 exu_U12026(.A(bypass_dfill_data_g2[12]), .B(exu_n16278), .Y(exu_n22547));
INVX1 exu_U12027(.A(exu_n22547), .Y(exu_n1418));
AND2X1 exu_U12028(.A(exu_n22549), .B(exu_n10062), .Y(bypass_rs3_data_w2[11]));
INVX1 exu_U12029(.A(bypass_rs3_data_w2[11]), .Y(exu_n1419));
AND2X1 exu_U12030(.A(bypass_dfill_data_g2[11]), .B(exu_n16278), .Y(exu_n22551));
INVX1 exu_U12031(.A(exu_n22551), .Y(exu_n1420));
AND2X1 exu_U12032(.A(exu_n22553), .B(exu_n10063), .Y(bypass_rs3_data_w2[10]));
INVX1 exu_U12033(.A(bypass_rs3_data_w2[10]), .Y(exu_n1421));
AND2X1 exu_U12034(.A(bypass_dfill_data_g2[10]), .B(exu_n16278), .Y(exu_n22555));
INVX1 exu_U12035(.A(exu_n22555), .Y(exu_n1422));
AND2X1 exu_U12036(.A(exu_n22557), .B(exu_n10064), .Y(bypass_rs3_data_w2[0]));
INVX1 exu_U12037(.A(bypass_rs3_data_w2[0]), .Y(exu_n1423));
AND2X1 exu_U12038(.A(bypass_dfill_data_g2[0]), .B(exu_n16278), .Y(exu_n22559));
INVX1 exu_U12039(.A(exu_n22559), .Y(exu_n1424));
AND2X1 exu_U12040(.A(ecl_byp_sel_load_g), .B(bypass_dfill_data_g2[9]), .Y(exu_n22563));
INVX1 exu_U12041(.A(exu_n22563), .Y(exu_n1425));
AND2X1 exu_U12042(.A(bypass_dfill_data_g2[8]), .B(exu_n16271), .Y(exu_n22567));
INVX1 exu_U12043(.A(exu_n22567), .Y(exu_n1426));
AND2X1 exu_U12044(.A(bypass_dfill_data_g2[7]), .B(exu_n16271), .Y(exu_n22571));
INVX1 exu_U12045(.A(exu_n22571), .Y(exu_n1427));
AND2X1 exu_U12046(.A(bypass_dfill_data_g2[6]), .B(exu_n16271), .Y(exu_n22575));
INVX1 exu_U12047(.A(exu_n22575), .Y(exu_n1428));
AND2X1 exu_U12048(.A(bypass_dfill_data_g2[63]), .B(exu_n16271), .Y(exu_n22579));
INVX1 exu_U12049(.A(exu_n22579), .Y(exu_n1429));
AND2X1 exu_U12050(.A(bypass_dfill_data_g2[62]), .B(exu_n16271), .Y(exu_n22583));
INVX1 exu_U12051(.A(exu_n22583), .Y(exu_n1430));
AND2X1 exu_U12052(.A(bypass_dfill_data_g2[61]), .B(exu_n16271), .Y(exu_n22587));
INVX1 exu_U12053(.A(exu_n22587), .Y(exu_n1431));
AND2X1 exu_U12054(.A(bypass_dfill_data_g2[60]), .B(exu_n16271), .Y(exu_n22591));
INVX1 exu_U12055(.A(exu_n22591), .Y(exu_n1432));
AND2X1 exu_U12056(.A(bypass_dfill_data_g2[5]), .B(exu_n16271), .Y(exu_n22595));
INVX1 exu_U12057(.A(exu_n22595), .Y(exu_n1433));
AND2X1 exu_U12058(.A(bypass_dfill_data_g2[59]), .B(exu_n16271), .Y(exu_n22599));
INVX1 exu_U12059(.A(exu_n22599), .Y(exu_n1434));
AND2X1 exu_U12060(.A(bypass_dfill_data_g2[58]), .B(exu_n16271), .Y(exu_n22603));
INVX1 exu_U12061(.A(exu_n22603), .Y(exu_n1435));
AND2X1 exu_U12062(.A(bypass_dfill_data_g2[57]), .B(exu_n16271), .Y(exu_n22607));
INVX1 exu_U12063(.A(exu_n22607), .Y(exu_n1436));
AND2X1 exu_U12064(.A(bypass_dfill_data_g2[56]), .B(exu_n16271), .Y(exu_n22611));
INVX1 exu_U12065(.A(exu_n22611), .Y(exu_n1437));
AND2X1 exu_U12066(.A(bypass_dfill_data_g2[55]), .B(exu_n16271), .Y(exu_n22615));
INVX1 exu_U12067(.A(exu_n22615), .Y(exu_n1438));
AND2X1 exu_U12068(.A(bypass_dfill_data_g2[54]), .B(ecl_byp_sel_load_g), .Y(exu_n22619));
INVX1 exu_U12069(.A(exu_n22619), .Y(exu_n1439));
AND2X1 exu_U12070(.A(bypass_dfill_data_g2[53]), .B(exu_n16271), .Y(exu_n22623));
INVX1 exu_U12071(.A(exu_n22623), .Y(exu_n1440));
AND2X1 exu_U12072(.A(bypass_dfill_data_g2[52]), .B(ecl_byp_sel_load_g), .Y(exu_n22627));
INVX1 exu_U12073(.A(exu_n22627), .Y(exu_n1441));
AND2X1 exu_U12074(.A(bypass_dfill_data_g2[51]), .B(exu_n16271), .Y(exu_n22631));
INVX1 exu_U12075(.A(exu_n22631), .Y(exu_n1442));
AND2X1 exu_U12076(.A(bypass_dfill_data_g2[50]), .B(ecl_byp_sel_load_g), .Y(exu_n22635));
INVX1 exu_U12077(.A(exu_n22635), .Y(exu_n1443));
AND2X1 exu_U12078(.A(bypass_dfill_data_g2[4]), .B(exu_n16271), .Y(exu_n22639));
INVX1 exu_U12079(.A(exu_n22639), .Y(exu_n1444));
AND2X1 exu_U12080(.A(bypass_dfill_data_g2[49]), .B(ecl_byp_sel_load_g), .Y(exu_n22643));
INVX1 exu_U12081(.A(exu_n22643), .Y(exu_n1445));
AND2X1 exu_U12082(.A(bypass_dfill_data_g2[48]), .B(exu_n16271), .Y(exu_n22647));
INVX1 exu_U12083(.A(exu_n22647), .Y(exu_n1446));
AND2X1 exu_U12084(.A(bypass_dfill_data_g2[47]), .B(ecl_byp_sel_load_g), .Y(exu_n22651));
INVX1 exu_U12085(.A(exu_n22651), .Y(exu_n1447));
AND2X1 exu_U12086(.A(bypass_dfill_data_g2[46]), .B(exu_n16271), .Y(exu_n22655));
INVX1 exu_U12087(.A(exu_n22655), .Y(exu_n1448));
AND2X1 exu_U12088(.A(bypass_dfill_data_g2[45]), .B(ecl_byp_sel_load_g), .Y(exu_n22659));
INVX1 exu_U12089(.A(exu_n22659), .Y(exu_n1449));
AND2X1 exu_U12090(.A(bypass_dfill_data_g2[44]), .B(exu_n16271), .Y(exu_n22663));
INVX1 exu_U12091(.A(exu_n22663), .Y(exu_n1450));
AND2X1 exu_U12092(.A(bypass_dfill_data_g2[43]), .B(ecl_byp_sel_load_g), .Y(exu_n22667));
INVX1 exu_U12093(.A(exu_n22667), .Y(exu_n1451));
AND2X1 exu_U12094(.A(bypass_dfill_data_g2[42]), .B(exu_n16271), .Y(exu_n22671));
INVX1 exu_U12095(.A(exu_n22671), .Y(exu_n1452));
AND2X1 exu_U12096(.A(bypass_dfill_data_g2[41]), .B(ecl_byp_sel_load_g), .Y(exu_n22675));
INVX1 exu_U12097(.A(exu_n22675), .Y(exu_n1453));
AND2X1 exu_U12098(.A(bypass_dfill_data_g2[40]), .B(ecl_byp_sel_load_g), .Y(exu_n22679));
INVX1 exu_U12099(.A(exu_n22679), .Y(exu_n1454));
AND2X1 exu_U12100(.A(bypass_dfill_data_g2[3]), .B(ecl_byp_sel_load_g), .Y(exu_n22683));
INVX1 exu_U12101(.A(exu_n22683), .Y(exu_n1455));
AND2X1 exu_U12102(.A(bypass_dfill_data_g2[39]), .B(ecl_byp_sel_load_g), .Y(exu_n22687));
INVX1 exu_U12103(.A(exu_n22687), .Y(exu_n1456));
AND2X1 exu_U12104(.A(bypass_dfill_data_g2[38]), .B(ecl_byp_sel_load_g), .Y(exu_n22691));
INVX1 exu_U12105(.A(exu_n22691), .Y(exu_n1457));
AND2X1 exu_U12106(.A(bypass_dfill_data_g2[37]), .B(ecl_byp_sel_load_g), .Y(exu_n22695));
INVX1 exu_U12107(.A(exu_n22695), .Y(exu_n1458));
AND2X1 exu_U12108(.A(bypass_dfill_data_g2[36]), .B(exu_n16271), .Y(exu_n22699));
INVX1 exu_U12109(.A(exu_n22699), .Y(exu_n1459));
AND2X1 exu_U12110(.A(bypass_dfill_data_g2[35]), .B(ecl_byp_sel_load_g), .Y(exu_n22703));
INVX1 exu_U12111(.A(exu_n22703), .Y(exu_n1460));
AND2X1 exu_U12112(.A(bypass_dfill_data_g2[34]), .B(ecl_byp_sel_load_g), .Y(exu_n22707));
INVX1 exu_U12113(.A(exu_n22707), .Y(exu_n1461));
AND2X1 exu_U12114(.A(bypass_dfill_data_g2[33]), .B(exu_n16271), .Y(exu_n22711));
INVX1 exu_U12115(.A(exu_n22711), .Y(exu_n1462));
AND2X1 exu_U12116(.A(bypass_dfill_data_g2[32]), .B(ecl_byp_sel_load_g), .Y(exu_n22715));
INVX1 exu_U12117(.A(exu_n22715), .Y(exu_n1463));
AND2X1 exu_U12118(.A(bypass_dfill_data_g2[31]), .B(ecl_byp_sel_load_g), .Y(exu_n22719));
INVX1 exu_U12119(.A(exu_n22719), .Y(exu_n1464));
AND2X1 exu_U12120(.A(bypass_dfill_data_g2[30]), .B(ecl_byp_sel_load_g), .Y(exu_n22723));
INVX1 exu_U12121(.A(exu_n22723), .Y(exu_n1465));
AND2X1 exu_U12122(.A(bypass_dfill_data_g2[2]), .B(ecl_byp_sel_load_g), .Y(exu_n22727));
INVX1 exu_U12123(.A(exu_n22727), .Y(exu_n1466));
AND2X1 exu_U12124(.A(bypass_dfill_data_g2[29]), .B(ecl_byp_sel_load_g), .Y(exu_n22731));
INVX1 exu_U12125(.A(exu_n22731), .Y(exu_n1467));
AND2X1 exu_U12126(.A(bypass_dfill_data_g2[28]), .B(ecl_byp_sel_load_g), .Y(exu_n22735));
INVX1 exu_U12127(.A(exu_n22735), .Y(exu_n1468));
AND2X1 exu_U12128(.A(bypass_dfill_data_g2[27]), .B(exu_n16271), .Y(exu_n22739));
INVX1 exu_U12129(.A(exu_n22739), .Y(exu_n1469));
AND2X1 exu_U12130(.A(bypass_dfill_data_g2[26]), .B(ecl_byp_sel_load_g), .Y(exu_n22743));
INVX1 exu_U12131(.A(exu_n22743), .Y(exu_n1470));
AND2X1 exu_U12132(.A(bypass_dfill_data_g2[25]), .B(exu_n16271), .Y(exu_n22747));
INVX1 exu_U12133(.A(exu_n22747), .Y(exu_n1471));
AND2X1 exu_U12134(.A(bypass_dfill_data_g2[24]), .B(exu_n16271), .Y(exu_n22751));
INVX1 exu_U12135(.A(exu_n22751), .Y(exu_n1472));
AND2X1 exu_U12136(.A(bypass_dfill_data_g2[23]), .B(ecl_byp_sel_load_g), .Y(exu_n22755));
INVX1 exu_U12137(.A(exu_n22755), .Y(exu_n1473));
AND2X1 exu_U12138(.A(bypass_dfill_data_g2[22]), .B(ecl_byp_sel_load_g), .Y(exu_n22759));
INVX1 exu_U12139(.A(exu_n22759), .Y(exu_n1474));
AND2X1 exu_U12140(.A(bypass_dfill_data_g2[21]), .B(ecl_byp_sel_load_g), .Y(exu_n22763));
INVX1 exu_U12141(.A(exu_n22763), .Y(exu_n1475));
AND2X1 exu_U12142(.A(bypass_dfill_data_g2[20]), .B(exu_n16271), .Y(exu_n22767));
INVX1 exu_U12143(.A(exu_n22767), .Y(exu_n1476));
AND2X1 exu_U12144(.A(bypass_dfill_data_g2[1]), .B(exu_n16271), .Y(exu_n22771));
INVX1 exu_U12145(.A(exu_n22771), .Y(exu_n1477));
AND2X1 exu_U12146(.A(bypass_dfill_data_g2[19]), .B(ecl_byp_sel_load_g), .Y(exu_n22775));
INVX1 exu_U12147(.A(exu_n22775), .Y(exu_n1478));
AND2X1 exu_U12148(.A(bypass_dfill_data_g2[18]), .B(ecl_byp_sel_load_g), .Y(exu_n22779));
INVX1 exu_U12149(.A(exu_n22779), .Y(exu_n1479));
AND2X1 exu_U12150(.A(bypass_dfill_data_g2[17]), .B(exu_n16271), .Y(exu_n22783));
INVX1 exu_U12151(.A(exu_n22783), .Y(exu_n1480));
AND2X1 exu_U12152(.A(bypass_dfill_data_g2[16]), .B(exu_n16271), .Y(exu_n22787));
INVX1 exu_U12153(.A(exu_n22787), .Y(exu_n1481));
AND2X1 exu_U12154(.A(bypass_dfill_data_g2[15]), .B(ecl_byp_sel_load_g), .Y(exu_n22791));
INVX1 exu_U12155(.A(exu_n22791), .Y(exu_n1482));
AND2X1 exu_U12156(.A(bypass_dfill_data_g2[14]), .B(ecl_byp_sel_load_g), .Y(exu_n22795));
INVX1 exu_U12157(.A(exu_n22795), .Y(exu_n1483));
AND2X1 exu_U12158(.A(bypass_dfill_data_g2[13]), .B(exu_n16271), .Y(exu_n22799));
INVX1 exu_U12159(.A(exu_n22799), .Y(exu_n1484));
AND2X1 exu_U12160(.A(bypass_dfill_data_g2[12]), .B(ecl_byp_sel_load_g), .Y(exu_n22803));
INVX1 exu_U12161(.A(exu_n22803), .Y(exu_n1485));
AND2X1 exu_U12162(.A(bypass_dfill_data_g2[11]), .B(exu_n16271), .Y(exu_n22807));
INVX1 exu_U12163(.A(exu_n22807), .Y(exu_n1486));
AND2X1 exu_U12164(.A(bypass_dfill_data_g2[10]), .B(exu_n16271), .Y(exu_n22811));
INVX1 exu_U12165(.A(exu_n22811), .Y(exu_n1487));
AND2X1 exu_U12166(.A(bypass_dfill_data_g2[0]), .B(exu_n16271), .Y(exu_n22815));
INVX1 exu_U12167(.A(exu_n22815), .Y(exu_n1488));
AND2X1 exu_U12168(.A(ecl_ecc_sel_rs2_m_l), .B(ecc_byp_alu_rs2_data_m[9]), .Y(exu_n22819));
INVX1 exu_U12169(.A(exu_n22819), .Y(exu_n1489));
AND2X1 exu_U12170(.A(ecc_byp_alu_rs2_data_m[8]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22823));
INVX1 exu_U12171(.A(exu_n22823), .Y(exu_n1490));
AND2X1 exu_U12172(.A(ecc_byp_alu_rs2_data_m[7]), .B(exu_n15974), .Y(exu_n22827));
INVX1 exu_U12173(.A(exu_n22827), .Y(exu_n1491));
AND2X1 exu_U12174(.A(ecc_byp_alu_rs2_data_m[6]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22831));
INVX1 exu_U12175(.A(exu_n22831), .Y(exu_n1492));
AND2X1 exu_U12176(.A(ecc_byp_alu_rs2_data_m[63]), .B(exu_n15974), .Y(exu_n22835));
INVX1 exu_U12177(.A(exu_n22835), .Y(exu_n1493));
AND2X1 exu_U12178(.A(ecc_byp_alu_rs2_data_m[62]), .B(exu_n15974), .Y(exu_n22839));
INVX1 exu_U12179(.A(exu_n22839), .Y(exu_n1494));
AND2X1 exu_U12180(.A(ecc_byp_alu_rs2_data_m[61]), .B(exu_n15974), .Y(exu_n22843));
INVX1 exu_U12181(.A(exu_n22843), .Y(exu_n1495));
AND2X1 exu_U12182(.A(ecc_byp_alu_rs2_data_m[60]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22847));
INVX1 exu_U12183(.A(exu_n22847), .Y(exu_n1496));
AND2X1 exu_U12184(.A(ecc_byp_alu_rs2_data_m[5]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22851));
INVX1 exu_U12185(.A(exu_n22851), .Y(exu_n1497));
AND2X1 exu_U12186(.A(ecc_byp_alu_rs2_data_m[59]), .B(exu_n15974), .Y(exu_n22855));
INVX1 exu_U12187(.A(exu_n22855), .Y(exu_n1498));
AND2X1 exu_U12188(.A(ecc_byp_alu_rs2_data_m[58]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22859));
INVX1 exu_U12189(.A(exu_n22859), .Y(exu_n1499));
AND2X1 exu_U12190(.A(ecc_byp_alu_rs2_data_m[57]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22863));
INVX1 exu_U12191(.A(exu_n22863), .Y(exu_n1500));
AND2X1 exu_U12192(.A(ecc_byp_alu_rs2_data_m[56]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22867));
INVX1 exu_U12193(.A(exu_n22867), .Y(exu_n1501));
AND2X1 exu_U12194(.A(ecc_byp_alu_rs2_data_m[55]), .B(exu_n15974), .Y(exu_n22871));
INVX1 exu_U12195(.A(exu_n22871), .Y(exu_n1502));
AND2X1 exu_U12196(.A(ecc_byp_alu_rs2_data_m[54]), .B(exu_n15974), .Y(exu_n22875));
INVX1 exu_U12197(.A(exu_n22875), .Y(exu_n1503));
AND2X1 exu_U12198(.A(ecc_byp_alu_rs2_data_m[53]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22879));
INVX1 exu_U12199(.A(exu_n22879), .Y(exu_n1504));
AND2X1 exu_U12200(.A(ecc_byp_alu_rs2_data_m[52]), .B(exu_n15974), .Y(exu_n22883));
INVX1 exu_U12201(.A(exu_n22883), .Y(exu_n1505));
AND2X1 exu_U12202(.A(ecc_byp_alu_rs2_data_m[51]), .B(exu_n15974), .Y(exu_n22887));
INVX1 exu_U12203(.A(exu_n22887), .Y(exu_n1506));
AND2X1 exu_U12204(.A(ecc_byp_alu_rs2_data_m[50]), .B(exu_n15974), .Y(exu_n22891));
INVX1 exu_U12205(.A(exu_n22891), .Y(exu_n1507));
AND2X1 exu_U12206(.A(ecc_byp_alu_rs2_data_m[4]), .B(exu_n15974), .Y(exu_n22895));
INVX1 exu_U12207(.A(exu_n22895), .Y(exu_n1508));
AND2X1 exu_U12208(.A(ecc_byp_alu_rs2_data_m[49]), .B(exu_n15974), .Y(exu_n22899));
INVX1 exu_U12209(.A(exu_n22899), .Y(exu_n1509));
AND2X1 exu_U12210(.A(ecc_byp_alu_rs2_data_m[48]), .B(exu_n15974), .Y(exu_n22903));
INVX1 exu_U12211(.A(exu_n22903), .Y(exu_n1510));
AND2X1 exu_U12212(.A(ecc_byp_alu_rs2_data_m[47]), .B(exu_n15974), .Y(exu_n22907));
INVX1 exu_U12213(.A(exu_n22907), .Y(exu_n1511));
AND2X1 exu_U12214(.A(ecc_byp_alu_rs2_data_m[46]), .B(exu_n15974), .Y(exu_n22911));
INVX1 exu_U12215(.A(exu_n22911), .Y(exu_n1512));
AND2X1 exu_U12216(.A(ecc_byp_alu_rs2_data_m[45]), .B(exu_n15974), .Y(exu_n22915));
INVX1 exu_U12217(.A(exu_n22915), .Y(exu_n1513));
AND2X1 exu_U12218(.A(ecc_byp_alu_rs2_data_m[44]), .B(exu_n15974), .Y(exu_n22919));
INVX1 exu_U12219(.A(exu_n22919), .Y(exu_n1514));
AND2X1 exu_U12220(.A(ecc_byp_alu_rs2_data_m[43]), .B(exu_n15974), .Y(exu_n22923));
INVX1 exu_U12221(.A(exu_n22923), .Y(exu_n1515));
AND2X1 exu_U12222(.A(ecc_byp_alu_rs2_data_m[42]), .B(exu_n15974), .Y(exu_n22927));
INVX1 exu_U12223(.A(exu_n22927), .Y(exu_n1516));
AND2X1 exu_U12224(.A(ecc_byp_alu_rs2_data_m[41]), .B(exu_n15974), .Y(exu_n22931));
INVX1 exu_U12225(.A(exu_n22931), .Y(exu_n1517));
AND2X1 exu_U12226(.A(ecc_byp_alu_rs2_data_m[40]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22935));
INVX1 exu_U12227(.A(exu_n22935), .Y(exu_n1518));
AND2X1 exu_U12228(.A(ecc_byp_alu_rs2_data_m[3]), .B(exu_n15974), .Y(exu_n22939));
INVX1 exu_U12229(.A(exu_n22939), .Y(exu_n1519));
AND2X1 exu_U12230(.A(ecc_byp_alu_rs2_data_m[39]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22943));
INVX1 exu_U12231(.A(exu_n22943), .Y(exu_n1520));
AND2X1 exu_U12232(.A(ecc_byp_alu_rs2_data_m[38]), .B(exu_n15974), .Y(exu_n22947));
INVX1 exu_U12233(.A(exu_n22947), .Y(exu_n1521));
AND2X1 exu_U12234(.A(ecc_byp_alu_rs2_data_m[37]), .B(exu_n15974), .Y(exu_n22951));
INVX1 exu_U12235(.A(exu_n22951), .Y(exu_n1522));
AND2X1 exu_U12236(.A(ecc_byp_alu_rs2_data_m[36]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22955));
INVX1 exu_U12237(.A(exu_n22955), .Y(exu_n1523));
AND2X1 exu_U12238(.A(ecc_byp_alu_rs2_data_m[35]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22959));
INVX1 exu_U12239(.A(exu_n22959), .Y(exu_n1524));
AND2X1 exu_U12240(.A(ecc_byp_alu_rs2_data_m[34]), .B(exu_n15974), .Y(exu_n22963));
INVX1 exu_U12241(.A(exu_n22963), .Y(exu_n1525));
AND2X1 exu_U12242(.A(ecc_byp_alu_rs2_data_m[33]), .B(exu_n15974), .Y(exu_n22967));
INVX1 exu_U12243(.A(exu_n22967), .Y(exu_n1526));
AND2X1 exu_U12244(.A(ecc_byp_alu_rs2_data_m[32]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22971));
INVX1 exu_U12245(.A(exu_n22971), .Y(exu_n1527));
AND2X1 exu_U12246(.A(ecc_byp_alu_rs2_data_m[31]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22975));
INVX1 exu_U12247(.A(exu_n22975), .Y(exu_n1528));
AND2X1 exu_U12248(.A(ecc_byp_alu_rs2_data_m[30]), .B(exu_n15974), .Y(exu_n22979));
INVX1 exu_U12249(.A(exu_n22979), .Y(exu_n1529));
AND2X1 exu_U12250(.A(ecc_byp_alu_rs2_data_m[2]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22983));
INVX1 exu_U12251(.A(exu_n22983), .Y(exu_n1530));
AND2X1 exu_U12252(.A(ecc_byp_alu_rs2_data_m[29]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22987));
INVX1 exu_U12253(.A(exu_n22987), .Y(exu_n1531));
AND2X1 exu_U12254(.A(ecc_byp_alu_rs2_data_m[28]), .B(exu_n15974), .Y(exu_n22991));
INVX1 exu_U12255(.A(exu_n22991), .Y(exu_n1532));
AND2X1 exu_U12256(.A(ecc_byp_alu_rs2_data_m[27]), .B(exu_n15974), .Y(exu_n22995));
INVX1 exu_U12257(.A(exu_n22995), .Y(exu_n1533));
AND2X1 exu_U12258(.A(ecc_byp_alu_rs2_data_m[26]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n22999));
INVX1 exu_U12259(.A(exu_n22999), .Y(exu_n1534));
AND2X1 exu_U12260(.A(ecc_byp_alu_rs2_data_m[25]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23003));
INVX1 exu_U12261(.A(exu_n23003), .Y(exu_n1535));
AND2X1 exu_U12262(.A(ecc_byp_alu_rs2_data_m[24]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23007));
INVX1 exu_U12263(.A(exu_n23007), .Y(exu_n1536));
AND2X1 exu_U12264(.A(ecc_byp_alu_rs2_data_m[23]), .B(exu_n15974), .Y(exu_n23011));
INVX1 exu_U12265(.A(exu_n23011), .Y(exu_n1537));
AND2X1 exu_U12266(.A(ecc_byp_alu_rs2_data_m[22]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23015));
INVX1 exu_U12267(.A(exu_n23015), .Y(exu_n1538));
AND2X1 exu_U12268(.A(ecc_byp_alu_rs2_data_m[21]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23019));
INVX1 exu_U12269(.A(exu_n23019), .Y(exu_n1539));
AND2X1 exu_U12270(.A(ecc_byp_alu_rs2_data_m[20]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23023));
INVX1 exu_U12271(.A(exu_n23023), .Y(exu_n1540));
AND2X1 exu_U12272(.A(ecc_byp_alu_rs2_data_m[1]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23027));
INVX1 exu_U12273(.A(exu_n23027), .Y(exu_n1541));
AND2X1 exu_U12274(.A(ecc_byp_alu_rs2_data_m[19]), .B(exu_n15974), .Y(exu_n23031));
INVX1 exu_U12275(.A(exu_n23031), .Y(exu_n1542));
AND2X1 exu_U12276(.A(ecc_byp_alu_rs2_data_m[18]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23035));
INVX1 exu_U12277(.A(exu_n23035), .Y(exu_n1543));
AND2X1 exu_U12278(.A(ecc_byp_alu_rs2_data_m[17]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23039));
INVX1 exu_U12279(.A(exu_n23039), .Y(exu_n1544));
AND2X1 exu_U12280(.A(ecc_byp_alu_rs2_data_m[16]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23043));
INVX1 exu_U12281(.A(exu_n23043), .Y(exu_n1545));
AND2X1 exu_U12282(.A(ecc_byp_alu_rs2_data_m[15]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23047));
INVX1 exu_U12283(.A(exu_n23047), .Y(exu_n1546));
AND2X1 exu_U12284(.A(ecc_byp_alu_rs2_data_m[14]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23051));
INVX1 exu_U12285(.A(exu_n23051), .Y(exu_n1547));
AND2X1 exu_U12286(.A(ecc_byp_alu_rs2_data_m[13]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23055));
INVX1 exu_U12287(.A(exu_n23055), .Y(exu_n1548));
AND2X1 exu_U12288(.A(ecc_byp_alu_rs2_data_m[12]), .B(exu_n15974), .Y(exu_n23059));
INVX1 exu_U12289(.A(exu_n23059), .Y(exu_n1549));
AND2X1 exu_U12290(.A(ecc_byp_alu_rs2_data_m[11]), .B(ecl_ecc_sel_rs2_m_l), .Y(exu_n23063));
INVX1 exu_U12291(.A(exu_n23063), .Y(exu_n1550));
AND2X1 exu_U12292(.A(ecc_byp_alu_rs2_data_m[10]), .B(exu_n15974), .Y(exu_n23067));
INVX1 exu_U12293(.A(exu_n23067), .Y(exu_n1551));
AND2X1 exu_U12294(.A(ecc_byp_alu_rs2_data_m[0]), .B(exu_n15974), .Y(exu_n23071));
INVX1 exu_U12295(.A(exu_n23071), .Y(exu_n1552));
AND2X1 exu_U12296(.A(ecl_writeback_n130), .B(bypass_restore_rd_data[9]), .Y(exu_n23203));
INVX1 exu_U12297(.A(exu_n23203), .Y(exu_n1553));
AND2X1 exu_U12298(.A(ecl_writeback_n167), .B(bypass_dfill_data_g2[9]), .Y(exu_n23205));
INVX1 exu_U12299(.A(exu_n23205), .Y(exu_n1554));
AND2X1 exu_U12300(.A(bypass_restore_rd_data[8]), .B(ecl_writeback_n130), .Y(exu_n23209));
INVX1 exu_U12301(.A(exu_n23209), .Y(exu_n1555));
AND2X1 exu_U12302(.A(bypass_dfill_data_g2[8]), .B(ecl_writeback_n167), .Y(exu_n23211));
INVX1 exu_U12303(.A(exu_n23211), .Y(exu_n1556));
AND2X1 exu_U12304(.A(bypass_restore_rd_data[7]), .B(ecl_writeback_n130), .Y(exu_n23215));
INVX1 exu_U12305(.A(exu_n23215), .Y(exu_n1557));
AND2X1 exu_U12306(.A(bypass_dfill_data_g2[7]), .B(exu_n15764), .Y(exu_n23217));
INVX1 exu_U12307(.A(exu_n23217), .Y(exu_n1558));
AND2X1 exu_U12308(.A(bypass_restore_rd_data[6]), .B(exu_n15989), .Y(exu_n23221));
INVX1 exu_U12309(.A(exu_n23221), .Y(exu_n1559));
AND2X1 exu_U12310(.A(bypass_dfill_data_g2[6]), .B(ecl_writeback_n167), .Y(exu_n23223));
INVX1 exu_U12311(.A(exu_n23223), .Y(exu_n1560));
AND2X1 exu_U12312(.A(bypass_restore_rd_data[63]), .B(ecl_writeback_n130), .Y(exu_n23227));
INVX1 exu_U12313(.A(exu_n23227), .Y(exu_n1561));
AND2X1 exu_U12314(.A(bypass_dfill_data_g2[63]), .B(exu_n15764), .Y(exu_n23229));
INVX1 exu_U12315(.A(exu_n23229), .Y(exu_n1562));
AND2X1 exu_U12316(.A(bypass_restore_rd_data[62]), .B(ecl_writeback_n130), .Y(exu_n23233));
INVX1 exu_U12317(.A(exu_n23233), .Y(exu_n1563));
AND2X1 exu_U12318(.A(bypass_dfill_data_g2[62]), .B(ecl_writeback_n167), .Y(exu_n23235));
INVX1 exu_U12319(.A(exu_n23235), .Y(exu_n1564));
AND2X1 exu_U12320(.A(bypass_restore_rd_data[61]), .B(ecl_writeback_n130), .Y(exu_n23239));
INVX1 exu_U12321(.A(exu_n23239), .Y(exu_n1565));
AND2X1 exu_U12322(.A(bypass_dfill_data_g2[61]), .B(exu_n15764), .Y(exu_n23241));
INVX1 exu_U12323(.A(exu_n23241), .Y(exu_n1566));
AND2X1 exu_U12324(.A(bypass_restore_rd_data[60]), .B(ecl_writeback_n130), .Y(exu_n23245));
INVX1 exu_U12325(.A(exu_n23245), .Y(exu_n1567));
AND2X1 exu_U12326(.A(bypass_dfill_data_g2[60]), .B(ecl_writeback_n167), .Y(exu_n23247));
INVX1 exu_U12327(.A(exu_n23247), .Y(exu_n1568));
AND2X1 exu_U12328(.A(bypass_restore_rd_data[5]), .B(ecl_writeback_n130), .Y(exu_n23251));
INVX1 exu_U12329(.A(exu_n23251), .Y(exu_n1569));
AND2X1 exu_U12330(.A(bypass_dfill_data_g2[5]), .B(exu_n15764), .Y(exu_n23253));
INVX1 exu_U12331(.A(exu_n23253), .Y(exu_n1570));
AND2X1 exu_U12332(.A(bypass_restore_rd_data[59]), .B(exu_n15989), .Y(exu_n23257));
INVX1 exu_U12333(.A(exu_n23257), .Y(exu_n1571));
AND2X1 exu_U12334(.A(bypass_dfill_data_g2[59]), .B(ecl_writeback_n167), .Y(exu_n23259));
INVX1 exu_U12335(.A(exu_n23259), .Y(exu_n1572));
AND2X1 exu_U12336(.A(bypass_restore_rd_data[58]), .B(exu_n15989), .Y(exu_n23263));
INVX1 exu_U12337(.A(exu_n23263), .Y(exu_n1573));
AND2X1 exu_U12338(.A(bypass_dfill_data_g2[58]), .B(exu_n15764), .Y(exu_n23265));
INVX1 exu_U12339(.A(exu_n23265), .Y(exu_n1574));
AND2X1 exu_U12340(.A(bypass_restore_rd_data[57]), .B(ecl_writeback_n130), .Y(exu_n23269));
INVX1 exu_U12341(.A(exu_n23269), .Y(exu_n1575));
AND2X1 exu_U12342(.A(bypass_dfill_data_g2[57]), .B(ecl_writeback_n167), .Y(exu_n23271));
INVX1 exu_U12343(.A(exu_n23271), .Y(exu_n1576));
AND2X1 exu_U12344(.A(bypass_restore_rd_data[56]), .B(exu_n15989), .Y(exu_n23275));
INVX1 exu_U12345(.A(exu_n23275), .Y(exu_n1577));
AND2X1 exu_U12346(.A(bypass_dfill_data_g2[56]), .B(exu_n15764), .Y(exu_n23277));
INVX1 exu_U12347(.A(exu_n23277), .Y(exu_n1578));
AND2X1 exu_U12348(.A(bypass_restore_rd_data[55]), .B(exu_n15989), .Y(exu_n23281));
INVX1 exu_U12349(.A(exu_n23281), .Y(exu_n1579));
AND2X1 exu_U12350(.A(bypass_dfill_data_g2[55]), .B(ecl_writeback_n167), .Y(exu_n23283));
INVX1 exu_U12351(.A(exu_n23283), .Y(exu_n1580));
AND2X1 exu_U12352(.A(bypass_restore_rd_data[54]), .B(ecl_writeback_n130), .Y(exu_n23287));
INVX1 exu_U12353(.A(exu_n23287), .Y(exu_n1581));
AND2X1 exu_U12354(.A(bypass_dfill_data_g2[54]), .B(exu_n15764), .Y(exu_n23289));
INVX1 exu_U12355(.A(exu_n23289), .Y(exu_n1582));
AND2X1 exu_U12356(.A(bypass_restore_rd_data[53]), .B(ecl_writeback_n130), .Y(exu_n23293));
INVX1 exu_U12357(.A(exu_n23293), .Y(exu_n1583));
AND2X1 exu_U12358(.A(bypass_dfill_data_g2[53]), .B(exu_n15764), .Y(exu_n23295));
INVX1 exu_U12359(.A(exu_n23295), .Y(exu_n1584));
AND2X1 exu_U12360(.A(bypass_restore_rd_data[52]), .B(ecl_writeback_n130), .Y(exu_n23299));
INVX1 exu_U12361(.A(exu_n23299), .Y(exu_n1585));
AND2X1 exu_U12362(.A(bypass_dfill_data_g2[52]), .B(ecl_writeback_n167), .Y(exu_n23301));
INVX1 exu_U12363(.A(exu_n23301), .Y(exu_n1586));
AND2X1 exu_U12364(.A(bypass_restore_rd_data[51]), .B(exu_n15989), .Y(exu_n23305));
INVX1 exu_U12365(.A(exu_n23305), .Y(exu_n1587));
AND2X1 exu_U12366(.A(bypass_dfill_data_g2[51]), .B(ecl_writeback_n167), .Y(exu_n23307));
INVX1 exu_U12367(.A(exu_n23307), .Y(exu_n1588));
AND2X1 exu_U12368(.A(bypass_restore_rd_data[50]), .B(ecl_writeback_n130), .Y(exu_n23311));
INVX1 exu_U12369(.A(exu_n23311), .Y(exu_n1589));
AND2X1 exu_U12370(.A(bypass_dfill_data_g2[50]), .B(exu_n15764), .Y(exu_n23313));
INVX1 exu_U12371(.A(exu_n23313), .Y(exu_n1590));
AND2X1 exu_U12372(.A(bypass_restore_rd_data[4]), .B(ecl_writeback_n130), .Y(exu_n23317));
INVX1 exu_U12373(.A(exu_n23317), .Y(exu_n1591));
AND2X1 exu_U12374(.A(bypass_dfill_data_g2[4]), .B(ecl_writeback_n167), .Y(exu_n23319));
INVX1 exu_U12375(.A(exu_n23319), .Y(exu_n1592));
AND2X1 exu_U12376(.A(bypass_restore_rd_data[49]), .B(exu_n15989), .Y(exu_n23323));
INVX1 exu_U12377(.A(exu_n23323), .Y(exu_n1593));
AND2X1 exu_U12378(.A(bypass_dfill_data_g2[49]), .B(exu_n15764), .Y(exu_n23325));
INVX1 exu_U12379(.A(exu_n23325), .Y(exu_n1594));
AND2X1 exu_U12380(.A(bypass_restore_rd_data[48]), .B(exu_n15989), .Y(exu_n23329));
INVX1 exu_U12381(.A(exu_n23329), .Y(exu_n1595));
AND2X1 exu_U12382(.A(bypass_dfill_data_g2[48]), .B(ecl_writeback_n167), .Y(exu_n23331));
INVX1 exu_U12383(.A(exu_n23331), .Y(exu_n1596));
AND2X1 exu_U12384(.A(bypass_restore_rd_data[47]), .B(exu_n15989), .Y(exu_n23335));
INVX1 exu_U12385(.A(exu_n23335), .Y(exu_n1597));
AND2X1 exu_U12386(.A(bypass_dfill_data_g2[47]), .B(exu_n15764), .Y(exu_n23337));
INVX1 exu_U12387(.A(exu_n23337), .Y(exu_n1598));
AND2X1 exu_U12388(.A(bypass_restore_rd_data[46]), .B(exu_n15989), .Y(exu_n23341));
INVX1 exu_U12389(.A(exu_n23341), .Y(exu_n1599));
AND2X1 exu_U12390(.A(bypass_dfill_data_g2[46]), .B(ecl_writeback_n167), .Y(exu_n23343));
INVX1 exu_U12391(.A(exu_n23343), .Y(exu_n1600));
AND2X1 exu_U12392(.A(bypass_restore_rd_data[45]), .B(exu_n15989), .Y(exu_n23347));
INVX1 exu_U12393(.A(exu_n23347), .Y(exu_n1601));
AND2X1 exu_U12394(.A(bypass_dfill_data_g2[45]), .B(exu_n15764), .Y(exu_n23349));
INVX1 exu_U12395(.A(exu_n23349), .Y(exu_n1602));
AND2X1 exu_U12396(.A(bypass_restore_rd_data[44]), .B(exu_n15989), .Y(exu_n23353));
INVX1 exu_U12397(.A(exu_n23353), .Y(exu_n1603));
AND2X1 exu_U12398(.A(bypass_dfill_data_g2[44]), .B(ecl_writeback_n167), .Y(exu_n23355));
INVX1 exu_U12399(.A(exu_n23355), .Y(exu_n1604));
AND2X1 exu_U12400(.A(bypass_restore_rd_data[43]), .B(exu_n15989), .Y(exu_n23359));
INVX1 exu_U12401(.A(exu_n23359), .Y(exu_n1605));
AND2X1 exu_U12402(.A(bypass_dfill_data_g2[43]), .B(exu_n15764), .Y(exu_n23361));
INVX1 exu_U12403(.A(exu_n23361), .Y(exu_n1606));
AND2X1 exu_U12404(.A(bypass_restore_rd_data[42]), .B(exu_n15989), .Y(exu_n23365));
INVX1 exu_U12405(.A(exu_n23365), .Y(exu_n1607));
AND2X1 exu_U12406(.A(bypass_dfill_data_g2[42]), .B(ecl_writeback_n167), .Y(exu_n23367));
INVX1 exu_U12407(.A(exu_n23367), .Y(exu_n1608));
AND2X1 exu_U12408(.A(bypass_restore_rd_data[41]), .B(exu_n15989), .Y(exu_n23371));
INVX1 exu_U12409(.A(exu_n23371), .Y(exu_n1609));
AND2X1 exu_U12410(.A(bypass_dfill_data_g2[41]), .B(exu_n15764), .Y(exu_n23373));
INVX1 exu_U12411(.A(exu_n23373), .Y(exu_n1610));
AND2X1 exu_U12412(.A(bypass_restore_rd_data[40]), .B(exu_n15989), .Y(exu_n23377));
INVX1 exu_U12413(.A(exu_n23377), .Y(exu_n1611));
AND2X1 exu_U12414(.A(bypass_dfill_data_g2[40]), .B(ecl_writeback_n167), .Y(exu_n23379));
INVX1 exu_U12415(.A(exu_n23379), .Y(exu_n1612));
AND2X1 exu_U12416(.A(bypass_restore_rd_data[3]), .B(exu_n15989), .Y(exu_n23383));
INVX1 exu_U12417(.A(exu_n23383), .Y(exu_n1613));
AND2X1 exu_U12418(.A(bypass_dfill_data_g2[3]), .B(exu_n15764), .Y(exu_n23385));
INVX1 exu_U12419(.A(exu_n23385), .Y(exu_n1614));
AND2X1 exu_U12420(.A(bypass_restore_rd_data[39]), .B(exu_n15989), .Y(exu_n23389));
INVX1 exu_U12421(.A(exu_n23389), .Y(exu_n1615));
AND2X1 exu_U12422(.A(bypass_dfill_data_g2[39]), .B(ecl_writeback_n167), .Y(exu_n23391));
INVX1 exu_U12423(.A(exu_n23391), .Y(exu_n1616));
AND2X1 exu_U12424(.A(bypass_restore_rd_data[38]), .B(exu_n15989), .Y(exu_n23395));
INVX1 exu_U12425(.A(exu_n23395), .Y(exu_n1617));
AND2X1 exu_U12426(.A(bypass_dfill_data_g2[38]), .B(exu_n15764), .Y(exu_n23397));
INVX1 exu_U12427(.A(exu_n23397), .Y(exu_n1618));
AND2X1 exu_U12428(.A(bypass_restore_rd_data[37]), .B(exu_n15989), .Y(exu_n23401));
INVX1 exu_U12429(.A(exu_n23401), .Y(exu_n1619));
AND2X1 exu_U12430(.A(bypass_dfill_data_g2[37]), .B(ecl_writeback_n167), .Y(exu_n23403));
INVX1 exu_U12431(.A(exu_n23403), .Y(exu_n1620));
AND2X1 exu_U12432(.A(bypass_restore_rd_data[36]), .B(ecl_writeback_n130), .Y(exu_n23407));
INVX1 exu_U12433(.A(exu_n23407), .Y(exu_n1621));
AND2X1 exu_U12434(.A(bypass_dfill_data_g2[36]), .B(exu_n15764), .Y(exu_n23409));
INVX1 exu_U12435(.A(exu_n23409), .Y(exu_n1622));
AND2X1 exu_U12436(.A(bypass_restore_rd_data[35]), .B(ecl_writeback_n130), .Y(exu_n23413));
INVX1 exu_U12437(.A(exu_n23413), .Y(exu_n1623));
AND2X1 exu_U12438(.A(bypass_dfill_data_g2[35]), .B(ecl_writeback_n167), .Y(exu_n23415));
INVX1 exu_U12439(.A(exu_n23415), .Y(exu_n1624));
AND2X1 exu_U12440(.A(bypass_restore_rd_data[34]), .B(ecl_writeback_n130), .Y(exu_n23419));
INVX1 exu_U12441(.A(exu_n23419), .Y(exu_n1625));
AND2X1 exu_U12442(.A(bypass_dfill_data_g2[34]), .B(ecl_writeback_n167), .Y(exu_n23421));
INVX1 exu_U12443(.A(exu_n23421), .Y(exu_n1626));
AND2X1 exu_U12444(.A(bypass_restore_rd_data[33]), .B(ecl_writeback_n130), .Y(exu_n23425));
INVX1 exu_U12445(.A(exu_n23425), .Y(exu_n1627));
AND2X1 exu_U12446(.A(bypass_dfill_data_g2[33]), .B(exu_n15764), .Y(exu_n23427));
INVX1 exu_U12447(.A(exu_n23427), .Y(exu_n1628));
AND2X1 exu_U12448(.A(bypass_restore_rd_data[32]), .B(exu_n15989), .Y(exu_n23431));
INVX1 exu_U12449(.A(exu_n23431), .Y(exu_n1629));
AND2X1 exu_U12450(.A(bypass_dfill_data_g2[32]), .B(exu_n15764), .Y(exu_n23433));
INVX1 exu_U12451(.A(exu_n23433), .Y(exu_n1630));
AND2X1 exu_U12452(.A(bypass_restore_rd_data[31]), .B(exu_n15989), .Y(exu_n23437));
INVX1 exu_U12453(.A(exu_n23437), .Y(exu_n1631));
AND2X1 exu_U12454(.A(bypass_dfill_data_g2[31]), .B(ecl_writeback_n167), .Y(exu_n23439));
INVX1 exu_U12455(.A(exu_n23439), .Y(exu_n1632));
AND2X1 exu_U12456(.A(bypass_restore_rd_data[30]), .B(exu_n15989), .Y(exu_n23443));
INVX1 exu_U12457(.A(exu_n23443), .Y(exu_n1633));
AND2X1 exu_U12458(.A(bypass_dfill_data_g2[30]), .B(exu_n15764), .Y(exu_n23445));
INVX1 exu_U12459(.A(exu_n23445), .Y(exu_n1634));
AND2X1 exu_U12460(.A(bypass_restore_rd_data[2]), .B(exu_n15989), .Y(exu_n23449));
INVX1 exu_U12461(.A(exu_n23449), .Y(exu_n1635));
AND2X1 exu_U12462(.A(bypass_dfill_data_g2[2]), .B(exu_n15764), .Y(exu_n23451));
INVX1 exu_U12463(.A(exu_n23451), .Y(exu_n1636));
AND2X1 exu_U12464(.A(bypass_restore_rd_data[29]), .B(ecl_writeback_n130), .Y(exu_n23455));
INVX1 exu_U12465(.A(exu_n23455), .Y(exu_n1637));
AND2X1 exu_U12466(.A(bypass_dfill_data_g2[29]), .B(exu_n15764), .Y(exu_n23457));
INVX1 exu_U12467(.A(exu_n23457), .Y(exu_n1638));
AND2X1 exu_U12468(.A(bypass_restore_rd_data[28]), .B(exu_n15989), .Y(exu_n23461));
INVX1 exu_U12469(.A(exu_n23461), .Y(exu_n1639));
AND2X1 exu_U12470(.A(bypass_dfill_data_g2[28]), .B(exu_n15764), .Y(exu_n23463));
INVX1 exu_U12471(.A(exu_n23463), .Y(exu_n1640));
AND2X1 exu_U12472(.A(bypass_restore_rd_data[27]), .B(exu_n15989), .Y(exu_n23467));
INVX1 exu_U12473(.A(exu_n23467), .Y(exu_n1641));
AND2X1 exu_U12474(.A(bypass_dfill_data_g2[27]), .B(ecl_writeback_n167), .Y(exu_n23469));
INVX1 exu_U12475(.A(exu_n23469), .Y(exu_n1642));
AND2X1 exu_U12476(.A(bypass_restore_rd_data[26]), .B(exu_n15989), .Y(exu_n23473));
INVX1 exu_U12477(.A(exu_n23473), .Y(exu_n1643));
AND2X1 exu_U12478(.A(bypass_dfill_data_g2[26]), .B(exu_n15764), .Y(exu_n23475));
INVX1 exu_U12479(.A(exu_n23475), .Y(exu_n1644));
AND2X1 exu_U12480(.A(bypass_restore_rd_data[25]), .B(ecl_writeback_n130), .Y(exu_n23479));
INVX1 exu_U12481(.A(exu_n23479), .Y(exu_n1645));
AND2X1 exu_U12482(.A(bypass_dfill_data_g2[25]), .B(ecl_writeback_n167), .Y(exu_n23481));
INVX1 exu_U12483(.A(exu_n23481), .Y(exu_n1646));
AND2X1 exu_U12484(.A(bypass_restore_rd_data[24]), .B(ecl_writeback_n130), .Y(exu_n23485));
INVX1 exu_U12485(.A(exu_n23485), .Y(exu_n1647));
AND2X1 exu_U12486(.A(bypass_dfill_data_g2[24]), .B(ecl_writeback_n167), .Y(exu_n23487));
INVX1 exu_U12487(.A(exu_n23487), .Y(exu_n1648));
AND2X1 exu_U12488(.A(bypass_restore_rd_data[23]), .B(exu_n15989), .Y(exu_n23491));
INVX1 exu_U12489(.A(exu_n23491), .Y(exu_n1649));
AND2X1 exu_U12490(.A(bypass_dfill_data_g2[23]), .B(exu_n15764), .Y(exu_n23493));
INVX1 exu_U12491(.A(exu_n23493), .Y(exu_n1650));
AND2X1 exu_U12492(.A(bypass_restore_rd_data[22]), .B(ecl_writeback_n130), .Y(exu_n23497));
INVX1 exu_U12493(.A(exu_n23497), .Y(exu_n1651));
AND2X1 exu_U12494(.A(bypass_dfill_data_g2[22]), .B(ecl_writeback_n167), .Y(exu_n23499));
INVX1 exu_U12495(.A(exu_n23499), .Y(exu_n1652));
AND2X1 exu_U12496(.A(bypass_restore_rd_data[21]), .B(ecl_writeback_n130), .Y(exu_n23503));
INVX1 exu_U12497(.A(exu_n23503), .Y(exu_n1653));
AND2X1 exu_U12498(.A(bypass_dfill_data_g2[21]), .B(exu_n15764), .Y(exu_n23505));
INVX1 exu_U12499(.A(exu_n23505), .Y(exu_n1654));
AND2X1 exu_U12500(.A(bypass_restore_rd_data[20]), .B(ecl_writeback_n130), .Y(exu_n23509));
INVX1 exu_U12501(.A(exu_n23509), .Y(exu_n1655));
AND2X1 exu_U12502(.A(bypass_dfill_data_g2[20]), .B(ecl_writeback_n167), .Y(exu_n23511));
INVX1 exu_U12503(.A(exu_n23511), .Y(exu_n1656));
AND2X1 exu_U12504(.A(bypass_restore_rd_data[1]), .B(exu_n15989), .Y(exu_n23515));
INVX1 exu_U12505(.A(exu_n23515), .Y(exu_n1657));
AND2X1 exu_U12506(.A(bypass_dfill_data_g2[1]), .B(ecl_writeback_n167), .Y(exu_n23517));
INVX1 exu_U12507(.A(exu_n23517), .Y(exu_n1658));
AND2X1 exu_U12508(.A(bypass_restore_rd_data[19]), .B(ecl_writeback_n130), .Y(exu_n23521));
INVX1 exu_U12509(.A(exu_n23521), .Y(exu_n1659));
AND2X1 exu_U12510(.A(bypass_dfill_data_g2[19]), .B(exu_n15764), .Y(exu_n23523));
INVX1 exu_U12511(.A(exu_n23523), .Y(exu_n1660));
AND2X1 exu_U12512(.A(bypass_restore_rd_data[18]), .B(exu_n15989), .Y(exu_n23527));
INVX1 exu_U12513(.A(exu_n23527), .Y(exu_n1661));
AND2X1 exu_U12514(.A(bypass_dfill_data_g2[18]), .B(exu_n15764), .Y(exu_n23529));
INVX1 exu_U12515(.A(exu_n23529), .Y(exu_n1662));
AND2X1 exu_U12516(.A(bypass_restore_rd_data[17]), .B(ecl_writeback_n130), .Y(exu_n23533));
INVX1 exu_U12517(.A(exu_n23533), .Y(exu_n1663));
AND2X1 exu_U12518(.A(bypass_dfill_data_g2[17]), .B(ecl_writeback_n167), .Y(exu_n23535));
INVX1 exu_U12519(.A(exu_n23535), .Y(exu_n1664));
AND2X1 exu_U12520(.A(bypass_restore_rd_data[16]), .B(ecl_writeback_n130), .Y(exu_n23539));
INVX1 exu_U12521(.A(exu_n23539), .Y(exu_n1665));
AND2X1 exu_U12522(.A(bypass_dfill_data_g2[16]), .B(exu_n15764), .Y(exu_n23541));
INVX1 exu_U12523(.A(exu_n23541), .Y(exu_n1666));
AND2X1 exu_U12524(.A(bypass_restore_rd_data[15]), .B(exu_n15989), .Y(exu_n23545));
INVX1 exu_U12525(.A(exu_n23545), .Y(exu_n1667));
AND2X1 exu_U12526(.A(bypass_dfill_data_g2[15]), .B(exu_n15764), .Y(exu_n23547));
INVX1 exu_U12527(.A(exu_n23547), .Y(exu_n1668));
AND2X1 exu_U12528(.A(bypass_restore_rd_data[14]), .B(ecl_writeback_n130), .Y(exu_n23551));
INVX1 exu_U12529(.A(exu_n23551), .Y(exu_n1669));
AND2X1 exu_U12530(.A(bypass_dfill_data_g2[14]), .B(ecl_writeback_n167), .Y(exu_n23553));
INVX1 exu_U12531(.A(exu_n23553), .Y(exu_n1670));
AND2X1 exu_U12532(.A(bypass_restore_rd_data[13]), .B(ecl_writeback_n130), .Y(exu_n23557));
INVX1 exu_U12533(.A(exu_n23557), .Y(exu_n1671));
AND2X1 exu_U12534(.A(bypass_dfill_data_g2[13]), .B(exu_n15764), .Y(exu_n23559));
INVX1 exu_U12535(.A(exu_n23559), .Y(exu_n1672));
AND2X1 exu_U12536(.A(bypass_restore_rd_data[12]), .B(ecl_writeback_n130), .Y(exu_n23563));
INVX1 exu_U12537(.A(exu_n23563), .Y(exu_n1673));
AND2X1 exu_U12538(.A(bypass_dfill_data_g2[12]), .B(exu_n15764), .Y(exu_n23565));
INVX1 exu_U12539(.A(exu_n23565), .Y(exu_n1674));
AND2X1 exu_U12540(.A(bypass_restore_rd_data[11]), .B(ecl_writeback_n130), .Y(exu_n23569));
INVX1 exu_U12541(.A(exu_n23569), .Y(exu_n1675));
AND2X1 exu_U12542(.A(bypass_dfill_data_g2[11]), .B(ecl_writeback_n167), .Y(exu_n23571));
INVX1 exu_U12543(.A(exu_n23571), .Y(exu_n1676));
AND2X1 exu_U12544(.A(bypass_restore_rd_data[10]), .B(exu_n15989), .Y(exu_n23575));
INVX1 exu_U12545(.A(exu_n23575), .Y(exu_n1677));
AND2X1 exu_U12546(.A(bypass_dfill_data_g2[10]), .B(exu_n15764), .Y(exu_n23577));
INVX1 exu_U12547(.A(exu_n23577), .Y(exu_n1678));
AND2X1 exu_U12548(.A(bypass_restore_rd_data[0]), .B(ecl_writeback_n130), .Y(exu_n23581));
INVX1 exu_U12549(.A(exu_n23581), .Y(exu_n1679));
AND2X1 exu_U12550(.A(bypass_dfill_data_g2[0]), .B(exu_n15764), .Y(exu_n23583));
INVX1 exu_U12551(.A(exu_n23583), .Y(exu_n1680));
AND2X1 exu_U12552(.A(exu_n15397), .B(ifu_exu_pc_d[9]), .Y(exu_n23587));
INVX1 exu_U12553(.A(exu_n23587), .Y(exu_n1681));
AND2X1 exu_U12554(.A(exu_n16308), .B(byp_irf_rd_data_w[9]), .Y(exu_n23589));
INVX1 exu_U12555(.A(exu_n23589), .Y(exu_n1682));
AND2X1 exu_U12556(.A(ifu_exu_pc_d[8]), .B(exu_n15397), .Y(exu_n23593));
INVX1 exu_U12557(.A(exu_n23593), .Y(exu_n1683));
AND2X1 exu_U12558(.A(byp_irf_rd_data_w[8]), .B(exu_n16308), .Y(exu_n23595));
INVX1 exu_U12559(.A(exu_n23595), .Y(exu_n1684));
AND2X1 exu_U12560(.A(ifu_exu_pc_d[7]), .B(exu_n15397), .Y(exu_n23599));
INVX1 exu_U12561(.A(exu_n23599), .Y(exu_n1685));
AND2X1 exu_U12562(.A(byp_irf_rd_data_w[7]), .B(exu_n16308), .Y(exu_n23601));
INVX1 exu_U12563(.A(exu_n23601), .Y(exu_n1686));
AND2X1 exu_U12564(.A(ifu_exu_pc_d[6]), .B(exu_n15397), .Y(exu_n23605));
INVX1 exu_U12565(.A(exu_n23605), .Y(exu_n1687));
AND2X1 exu_U12566(.A(byp_irf_rd_data_w[6]), .B(exu_n16308), .Y(exu_n23607));
INVX1 exu_U12567(.A(exu_n23607), .Y(exu_n1688));
AND2X1 exu_U12568(.A(byp_irf_rd_data_w[63]), .B(exu_n16308), .Y(exu_n23612));
INVX1 exu_U12569(.A(exu_n23612), .Y(exu_n1689));
INVX1 exu_U12570(.A(exu_n1694), .Y(exu_n1690));
INVX1 exu_U12571(.A(exu_n1690), .Y(exu_n1691));
AND2X1 exu_U12572(.A(byp_irf_rd_data_w[62]), .B(exu_n16308), .Y(exu_n23617));
INVX1 exu_U12573(.A(exu_n23617), .Y(exu_n1692));
INVX1 exu_U12574(.A(exu_n1713), .Y(exu_n1693));
INVX1 exu_U12575(.A(exu_n1693), .Y(exu_n1694));
AND2X1 exu_U12576(.A(byp_irf_rd_data_w[61]), .B(exu_n16308), .Y(exu_n23622));
INVX1 exu_U12577(.A(exu_n23622), .Y(exu_n1695));
AND2X1 exu_U12578(.A(byp_irf_rd_data_w[60]), .B(exu_n16308), .Y(exu_n23627));
INVX1 exu_U12579(.A(exu_n23627), .Y(exu_n1696));
AND2X1 exu_U12580(.A(ifu_exu_pc_d[5]), .B(exu_n15397), .Y(exu_n23631));
INVX1 exu_U12581(.A(exu_n23631), .Y(exu_n1697));
AND2X1 exu_U12582(.A(byp_irf_rd_data_w[5]), .B(exu_n16308), .Y(exu_n23633));
INVX1 exu_U12583(.A(exu_n23633), .Y(exu_n1698));
AND2X1 exu_U12584(.A(byp_irf_rd_data_w[59]), .B(exu_n16308), .Y(exu_n23638));
INVX1 exu_U12585(.A(exu_n23638), .Y(exu_n1699));
AND2X1 exu_U12586(.A(byp_irf_rd_data_w[58]), .B(exu_n16308), .Y(exu_n23643));
INVX1 exu_U12587(.A(exu_n23643), .Y(exu_n1700));
AND2X1 exu_U12588(.A(byp_irf_rd_data_w[57]), .B(exu_n16308), .Y(exu_n23648));
INVX1 exu_U12589(.A(exu_n23648), .Y(exu_n1701));
AND2X1 exu_U12590(.A(byp_irf_rd_data_w[56]), .B(exu_n16308), .Y(exu_n23653));
INVX1 exu_U12591(.A(exu_n23653), .Y(exu_n1702));
AND2X1 exu_U12592(.A(byp_irf_rd_data_w[55]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23658));
INVX1 exu_U12593(.A(exu_n23658), .Y(exu_n1703));
AND2X1 exu_U12594(.A(byp_irf_rd_data_w[54]), .B(exu_n16308), .Y(exu_n23663));
INVX1 exu_U12595(.A(exu_n23663), .Y(exu_n1704));
AND2X1 exu_U12596(.A(byp_irf_rd_data_w[53]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23668));
INVX1 exu_U12597(.A(exu_n23668), .Y(exu_n1705));
AND2X1 exu_U12598(.A(byp_irf_rd_data_w[52]), .B(exu_n16308), .Y(exu_n23673));
INVX1 exu_U12599(.A(exu_n23673), .Y(exu_n1706));
AND2X1 exu_U12600(.A(byp_irf_rd_data_w[51]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23678));
INVX1 exu_U12601(.A(exu_n23678), .Y(exu_n1707));
AND2X1 exu_U12602(.A(byp_irf_rd_data_w[50]), .B(exu_n16308), .Y(exu_n23683));
INVX1 exu_U12603(.A(exu_n23683), .Y(exu_n1708));
AND2X1 exu_U12604(.A(ifu_exu_pc_d[4]), .B(exu_n15397), .Y(exu_n23687));
INVX1 exu_U12605(.A(exu_n23687), .Y(exu_n1709));
AND2X1 exu_U12606(.A(byp_irf_rd_data_w[4]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23689));
INVX1 exu_U12607(.A(exu_n23689), .Y(exu_n1710));
AND2X1 exu_U12608(.A(byp_irf_rd_data_w[49]), .B(exu_n16308), .Y(exu_n23694));
INVX1 exu_U12609(.A(exu_n23694), .Y(exu_n1711));
AND2X1 exu_U12610(.A(byp_irf_rd_data_w[48]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23699));
INVX1 exu_U12611(.A(exu_n23699), .Y(exu_n1712));
AND2X1 exu_U12612(.A(ifu_exu_pc_d[47]), .B(exu_n15397), .Y(exu_n23703));
INVX1 exu_U12613(.A(exu_n23703), .Y(exu_n1713));
AND2X1 exu_U12614(.A(byp_irf_rd_data_w[47]), .B(exu_n16308), .Y(exu_n23705));
INVX1 exu_U12615(.A(exu_n23705), .Y(exu_n1714));
AND2X1 exu_U12616(.A(ifu_exu_pc_d[46]), .B(exu_n15397), .Y(exu_n23709));
INVX1 exu_U12617(.A(exu_n23709), .Y(exu_n1715));
AND2X1 exu_U12618(.A(byp_irf_rd_data_w[46]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23711));
INVX1 exu_U12619(.A(exu_n23711), .Y(exu_n1716));
AND2X1 exu_U12620(.A(ifu_exu_pc_d[45]), .B(exu_n15397), .Y(exu_n23715));
INVX1 exu_U12621(.A(exu_n23715), .Y(exu_n1717));
AND2X1 exu_U12622(.A(byp_irf_rd_data_w[45]), .B(exu_n16308), .Y(exu_n23717));
INVX1 exu_U12623(.A(exu_n23717), .Y(exu_n1718));
AND2X1 exu_U12624(.A(ifu_exu_pc_d[44]), .B(exu_n15397), .Y(exu_n23721));
INVX1 exu_U12625(.A(exu_n23721), .Y(exu_n1719));
AND2X1 exu_U12626(.A(byp_irf_rd_data_w[44]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23723));
INVX1 exu_U12627(.A(exu_n23723), .Y(exu_n1720));
AND2X1 exu_U12628(.A(ifu_exu_pc_d[43]), .B(exu_n15397), .Y(exu_n23727));
INVX1 exu_U12629(.A(exu_n23727), .Y(exu_n1721));
AND2X1 exu_U12630(.A(byp_irf_rd_data_w[43]), .B(exu_n16308), .Y(exu_n23729));
INVX1 exu_U12631(.A(exu_n23729), .Y(exu_n1722));
AND2X1 exu_U12632(.A(ifu_exu_pc_d[42]), .B(exu_n15397), .Y(exu_n23733));
INVX1 exu_U12633(.A(exu_n23733), .Y(exu_n1723));
AND2X1 exu_U12634(.A(byp_irf_rd_data_w[42]), .B(exu_n16308), .Y(exu_n23735));
INVX1 exu_U12635(.A(exu_n23735), .Y(exu_n1724));
AND2X1 exu_U12636(.A(ifu_exu_pc_d[41]), .B(exu_n15397), .Y(exu_n23739));
INVX1 exu_U12637(.A(exu_n23739), .Y(exu_n1725));
AND2X1 exu_U12638(.A(byp_irf_rd_data_w[41]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23741));
INVX1 exu_U12639(.A(exu_n23741), .Y(exu_n1726));
AND2X1 exu_U12640(.A(ifu_exu_pc_d[40]), .B(exu_n15397), .Y(exu_n23745));
INVX1 exu_U12641(.A(exu_n23745), .Y(exu_n1727));
AND2X1 exu_U12642(.A(byp_irf_rd_data_w[40]), .B(exu_n16308), .Y(exu_n23747));
INVX1 exu_U12643(.A(exu_n23747), .Y(exu_n1728));
AND2X1 exu_U12644(.A(ifu_exu_pc_d[3]), .B(exu_n15397), .Y(exu_n23751));
INVX1 exu_U12645(.A(exu_n23751), .Y(exu_n1729));
AND2X1 exu_U12646(.A(byp_irf_rd_data_w[3]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23753));
INVX1 exu_U12647(.A(exu_n23753), .Y(exu_n1730));
AND2X1 exu_U12648(.A(ifu_exu_pc_d[39]), .B(exu_n15397), .Y(exu_n23757));
INVX1 exu_U12649(.A(exu_n23757), .Y(exu_n1731));
AND2X1 exu_U12650(.A(byp_irf_rd_data_w[39]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23759));
INVX1 exu_U12651(.A(exu_n23759), .Y(exu_n1732));
AND2X1 exu_U12652(.A(ifu_exu_pc_d[38]), .B(exu_n15397), .Y(exu_n23763));
INVX1 exu_U12653(.A(exu_n23763), .Y(exu_n1733));
AND2X1 exu_U12654(.A(byp_irf_rd_data_w[38]), .B(exu_n16308), .Y(exu_n23765));
INVX1 exu_U12655(.A(exu_n23765), .Y(exu_n1734));
AND2X1 exu_U12656(.A(ifu_exu_pc_d[37]), .B(exu_n15397), .Y(exu_n23769));
INVX1 exu_U12657(.A(exu_n23769), .Y(exu_n1735));
AND2X1 exu_U12658(.A(byp_irf_rd_data_w[37]), .B(exu_n16308), .Y(exu_n23771));
INVX1 exu_U12659(.A(exu_n23771), .Y(exu_n1736));
AND2X1 exu_U12660(.A(ifu_exu_pc_d[36]), .B(exu_n15397), .Y(exu_n23775));
INVX1 exu_U12661(.A(exu_n23775), .Y(exu_n1737));
AND2X1 exu_U12662(.A(byp_irf_rd_data_w[36]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23777));
INVX1 exu_U12663(.A(exu_n23777), .Y(exu_n1738));
AND2X1 exu_U12664(.A(ifu_exu_pc_d[35]), .B(exu_n15397), .Y(exu_n23781));
INVX1 exu_U12665(.A(exu_n23781), .Y(exu_n1739));
AND2X1 exu_U12666(.A(byp_irf_rd_data_w[35]), .B(exu_n16308), .Y(exu_n23783));
INVX1 exu_U12667(.A(exu_n23783), .Y(exu_n1740));
AND2X1 exu_U12668(.A(ifu_exu_pc_d[34]), .B(exu_n15397), .Y(exu_n23787));
INVX1 exu_U12669(.A(exu_n23787), .Y(exu_n1741));
AND2X1 exu_U12670(.A(byp_irf_rd_data_w[34]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23789));
INVX1 exu_U12671(.A(exu_n23789), .Y(exu_n1742));
AND2X1 exu_U12672(.A(ifu_exu_pc_d[33]), .B(exu_n15397), .Y(exu_n23793));
INVX1 exu_U12673(.A(exu_n23793), .Y(exu_n1743));
AND2X1 exu_U12674(.A(byp_irf_rd_data_w[33]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23795));
INVX1 exu_U12675(.A(exu_n23795), .Y(exu_n1744));
AND2X1 exu_U12676(.A(ifu_exu_pc_d[32]), .B(exu_n15397), .Y(exu_n23799));
INVX1 exu_U12677(.A(exu_n23799), .Y(exu_n1745));
AND2X1 exu_U12678(.A(byp_irf_rd_data_w[32]), .B(exu_n16308), .Y(exu_n23801));
INVX1 exu_U12679(.A(exu_n23801), .Y(exu_n1746));
AND2X1 exu_U12680(.A(ifu_exu_pc_d[31]), .B(exu_n15397), .Y(exu_n23805));
INVX1 exu_U12681(.A(exu_n23805), .Y(exu_n1747));
AND2X1 exu_U12682(.A(byp_irf_rd_data_w[31]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23807));
INVX1 exu_U12683(.A(exu_n23807), .Y(exu_n1748));
AND2X1 exu_U12684(.A(ifu_exu_pc_d[30]), .B(exu_n15397), .Y(exu_n23811));
INVX1 exu_U12685(.A(exu_n23811), .Y(exu_n1749));
AND2X1 exu_U12686(.A(byp_irf_rd_data_w[30]), .B(exu_n16308), .Y(exu_n23813));
INVX1 exu_U12687(.A(exu_n23813), .Y(exu_n1750));
AND2X1 exu_U12688(.A(ifu_exu_pc_d[2]), .B(exu_n15397), .Y(exu_n23817));
INVX1 exu_U12689(.A(exu_n23817), .Y(exu_n1751));
AND2X1 exu_U12690(.A(byp_irf_rd_data_w[2]), .B(exu_n16308), .Y(exu_n23819));
INVX1 exu_U12691(.A(exu_n23819), .Y(exu_n1752));
AND2X1 exu_U12692(.A(ifu_exu_pc_d[29]), .B(exu_n15397), .Y(exu_n23823));
INVX1 exu_U12693(.A(exu_n23823), .Y(exu_n1753));
AND2X1 exu_U12694(.A(byp_irf_rd_data_w[29]), .B(exu_n16308), .Y(exu_n23825));
INVX1 exu_U12695(.A(exu_n23825), .Y(exu_n1754));
AND2X1 exu_U12696(.A(ifu_exu_pc_d[28]), .B(exu_n15397), .Y(exu_n23829));
INVX1 exu_U12697(.A(exu_n23829), .Y(exu_n1755));
AND2X1 exu_U12698(.A(byp_irf_rd_data_w[28]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23831));
INVX1 exu_U12699(.A(exu_n23831), .Y(exu_n1756));
AND2X1 exu_U12700(.A(ifu_exu_pc_d[27]), .B(exu_n15397), .Y(exu_n23835));
INVX1 exu_U12701(.A(exu_n23835), .Y(exu_n1757));
AND2X1 exu_U12702(.A(byp_irf_rd_data_w[27]), .B(exu_n16308), .Y(exu_n23837));
INVX1 exu_U12703(.A(exu_n23837), .Y(exu_n1758));
AND2X1 exu_U12704(.A(ifu_exu_pc_d[26]), .B(exu_n15397), .Y(exu_n23841));
INVX1 exu_U12705(.A(exu_n23841), .Y(exu_n1759));
AND2X1 exu_U12706(.A(byp_irf_rd_data_w[26]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23843));
INVX1 exu_U12707(.A(exu_n23843), .Y(exu_n1760));
AND2X1 exu_U12708(.A(ifu_exu_pc_d[25]), .B(exu_n15397), .Y(exu_n23847));
INVX1 exu_U12709(.A(exu_n23847), .Y(exu_n1761));
AND2X1 exu_U12710(.A(byp_irf_rd_data_w[25]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23849));
INVX1 exu_U12711(.A(exu_n23849), .Y(exu_n1762));
AND2X1 exu_U12712(.A(ifu_exu_pc_d[24]), .B(exu_n15397), .Y(exu_n23853));
INVX1 exu_U12713(.A(exu_n23853), .Y(exu_n1763));
AND2X1 exu_U12714(.A(byp_irf_rd_data_w[24]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23855));
INVX1 exu_U12715(.A(exu_n23855), .Y(exu_n1764));
AND2X1 exu_U12716(.A(ifu_exu_pc_d[23]), .B(exu_n15397), .Y(exu_n23859));
INVX1 exu_U12717(.A(exu_n23859), .Y(exu_n1765));
AND2X1 exu_U12718(.A(byp_irf_rd_data_w[23]), .B(exu_n16308), .Y(exu_n23861));
INVX1 exu_U12719(.A(exu_n23861), .Y(exu_n1766));
AND2X1 exu_U12720(.A(ifu_exu_pc_d[22]), .B(exu_n15397), .Y(exu_n23865));
INVX1 exu_U12721(.A(exu_n23865), .Y(exu_n1767));
AND2X1 exu_U12722(.A(byp_irf_rd_data_w[22]), .B(exu_n16308), .Y(exu_n23867));
INVX1 exu_U12723(.A(exu_n23867), .Y(exu_n1768));
AND2X1 exu_U12724(.A(ifu_exu_pc_d[21]), .B(exu_n15397), .Y(exu_n23871));
INVX1 exu_U12725(.A(exu_n23871), .Y(exu_n1769));
AND2X1 exu_U12726(.A(byp_irf_rd_data_w[21]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23873));
INVX1 exu_U12727(.A(exu_n23873), .Y(exu_n1770));
AND2X1 exu_U12728(.A(ifu_exu_pc_d[20]), .B(exu_n15397), .Y(exu_n23877));
INVX1 exu_U12729(.A(exu_n23877), .Y(exu_n1771));
AND2X1 exu_U12730(.A(byp_irf_rd_data_w[20]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23879));
INVX1 exu_U12731(.A(exu_n23879), .Y(exu_n1772));
AND2X1 exu_U12732(.A(ifu_exu_pc_d[1]), .B(exu_n15397), .Y(exu_n23883));
INVX1 exu_U12733(.A(exu_n23883), .Y(exu_n1773));
AND2X1 exu_U12734(.A(byp_irf_rd_data_w[1]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23885));
INVX1 exu_U12735(.A(exu_n23885), .Y(exu_n1774));
AND2X1 exu_U12736(.A(ifu_exu_pc_d[19]), .B(exu_n15397), .Y(exu_n23889));
INVX1 exu_U12737(.A(exu_n23889), .Y(exu_n1775));
AND2X1 exu_U12738(.A(byp_irf_rd_data_w[19]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23891));
INVX1 exu_U12739(.A(exu_n23891), .Y(exu_n1776));
AND2X1 exu_U12740(.A(ifu_exu_pc_d[18]), .B(exu_n15397), .Y(exu_n23895));
INVX1 exu_U12741(.A(exu_n23895), .Y(exu_n1777));
AND2X1 exu_U12742(.A(byp_irf_rd_data_w[18]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23897));
INVX1 exu_U12743(.A(exu_n23897), .Y(exu_n1778));
AND2X1 exu_U12744(.A(ifu_exu_pc_d[17]), .B(exu_n15397), .Y(exu_n23901));
INVX1 exu_U12745(.A(exu_n23901), .Y(exu_n1779));
AND2X1 exu_U12746(.A(byp_irf_rd_data_w[17]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23903));
INVX1 exu_U12747(.A(exu_n23903), .Y(exu_n1780));
AND2X1 exu_U12748(.A(ifu_exu_pc_d[16]), .B(exu_n15397), .Y(exu_n23907));
INVX1 exu_U12749(.A(exu_n23907), .Y(exu_n1781));
AND2X1 exu_U12750(.A(byp_irf_rd_data_w[16]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23909));
INVX1 exu_U12751(.A(exu_n23909), .Y(exu_n1782));
AND2X1 exu_U12752(.A(ifu_exu_pc_d[15]), .B(exu_n15397), .Y(exu_n23913));
INVX1 exu_U12753(.A(exu_n23913), .Y(exu_n1783));
AND2X1 exu_U12754(.A(byp_irf_rd_data_w[15]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23915));
INVX1 exu_U12755(.A(exu_n23915), .Y(exu_n1784));
AND2X1 exu_U12756(.A(ifu_exu_pc_d[14]), .B(exu_n15397), .Y(exu_n23919));
INVX1 exu_U12757(.A(exu_n23919), .Y(exu_n1785));
AND2X1 exu_U12758(.A(byp_irf_rd_data_w[14]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23921));
INVX1 exu_U12759(.A(exu_n23921), .Y(exu_n1786));
AND2X1 exu_U12760(.A(ifu_exu_pc_d[13]), .B(exu_n15397), .Y(exu_n23925));
INVX1 exu_U12761(.A(exu_n23925), .Y(exu_n1787));
AND2X1 exu_U12762(.A(byp_irf_rd_data_w[13]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23927));
INVX1 exu_U12763(.A(exu_n23927), .Y(exu_n1788));
AND2X1 exu_U12764(.A(ifu_exu_pc_d[12]), .B(exu_n15397), .Y(exu_n23931));
INVX1 exu_U12765(.A(exu_n23931), .Y(exu_n1789));
AND2X1 exu_U12766(.A(byp_irf_rd_data_w[12]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23933));
INVX1 exu_U12767(.A(exu_n23933), .Y(exu_n1790));
AND2X1 exu_U12768(.A(ifu_exu_pc_d[11]), .B(exu_n15397), .Y(exu_n23937));
INVX1 exu_U12769(.A(exu_n23937), .Y(exu_n1791));
AND2X1 exu_U12770(.A(byp_irf_rd_data_w[11]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23939));
INVX1 exu_U12771(.A(exu_n23939), .Y(exu_n1792));
AND2X1 exu_U12772(.A(ifu_exu_pc_d[10]), .B(exu_n15397), .Y(exu_n23943));
INVX1 exu_U12773(.A(exu_n23943), .Y(exu_n1793));
AND2X1 exu_U12774(.A(byp_irf_rd_data_w[10]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23945));
INVX1 exu_U12775(.A(exu_n23945), .Y(exu_n1794));
AND2X1 exu_U12776(.A(ifu_exu_pc_d[0]), .B(exu_n15397), .Y(exu_n23949));
INVX1 exu_U12777(.A(exu_n23949), .Y(exu_n1795));
AND2X1 exu_U12778(.A(byp_irf_rd_data_w[0]), .B(ecl_byp_rs1_mux1_sel_w), .Y(exu_n23951));
INVX1 exu_U12779(.A(exu_n23951), .Y(exu_n1796));
AND2X1 exu_U12780(.A(exu_n16313), .B(lsu_exu_dfill_data_g[9]), .Y(exu_n23955));
INVX1 exu_U12781(.A(exu_n23955), .Y(exu_n1797));
AND2X1 exu_U12782(.A(ecl_byp_rs1_mux2_sel_rf), .B(bypass_mux_rcc_data_2_in1[9]), .Y(exu_n23957));
INVX1 exu_U12783(.A(exu_n23957), .Y(exu_n1798));
AND2X1 exu_U12784(.A(lsu_exu_dfill_data_g[8]), .B(exu_n16313), .Y(exu_n23961));
INVX1 exu_U12785(.A(exu_n23961), .Y(exu_n1799));
AND2X1 exu_U12786(.A(bypass_mux_rcc_data_2_in1[8]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n23963));
INVX1 exu_U12787(.A(exu_n23963), .Y(exu_n1800));
AND2X1 exu_U12788(.A(lsu_exu_dfill_data_g[7]), .B(exu_n16313), .Y(exu_n23967));
INVX1 exu_U12789(.A(exu_n23967), .Y(exu_n1801));
AND2X1 exu_U12790(.A(bypass_mux_rcc_data_2_in1[7]), .B(exu_n16314), .Y(exu_n23969));
INVX1 exu_U12791(.A(exu_n23969), .Y(exu_n1802));
AND2X1 exu_U12792(.A(lsu_exu_dfill_data_g[6]), .B(exu_n16313), .Y(exu_n23973));
INVX1 exu_U12793(.A(exu_n23973), .Y(exu_n1803));
AND2X1 exu_U12794(.A(bypass_mux_rcc_data_2_in1[6]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n23975));
INVX1 exu_U12795(.A(exu_n23975), .Y(exu_n1804));
AND2X1 exu_U12796(.A(lsu_exu_dfill_data_g[63]), .B(exu_n16313), .Y(exu_n23979));
INVX1 exu_U12797(.A(exu_n23979), .Y(exu_n1805));
AND2X1 exu_U12798(.A(bypass_mux_rcc_data_2_in1[63]), .B(exu_n16314), .Y(exu_n23981));
INVX1 exu_U12799(.A(exu_n23981), .Y(exu_n1806));
AND2X1 exu_U12800(.A(lsu_exu_dfill_data_g[62]), .B(exu_n16313), .Y(exu_n23985));
INVX1 exu_U12801(.A(exu_n23985), .Y(exu_n1807));
AND2X1 exu_U12802(.A(bypass_mux_rcc_data_2_in1[62]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n23987));
INVX1 exu_U12803(.A(exu_n23987), .Y(exu_n1808));
AND2X1 exu_U12804(.A(lsu_exu_dfill_data_g[61]), .B(exu_n16313), .Y(exu_n23991));
INVX1 exu_U12805(.A(exu_n23991), .Y(exu_n1809));
AND2X1 exu_U12806(.A(bypass_mux_rcc_data_2_in1[61]), .B(exu_n16314), .Y(exu_n23993));
INVX1 exu_U12807(.A(exu_n23993), .Y(exu_n1810));
AND2X1 exu_U12808(.A(lsu_exu_dfill_data_g[60]), .B(exu_n16313), .Y(exu_n23997));
INVX1 exu_U12809(.A(exu_n23997), .Y(exu_n1811));
AND2X1 exu_U12810(.A(bypass_mux_rcc_data_2_in1[60]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n23999));
INVX1 exu_U12811(.A(exu_n23999), .Y(exu_n1812));
AND2X1 exu_U12812(.A(lsu_exu_dfill_data_g[5]), .B(exu_n16313), .Y(exu_n24003));
INVX1 exu_U12813(.A(exu_n24003), .Y(exu_n1813));
AND2X1 exu_U12814(.A(bypass_mux_rcc_data_2_in1[5]), .B(exu_n16314), .Y(exu_n24005));
INVX1 exu_U12815(.A(exu_n24005), .Y(exu_n1814));
AND2X1 exu_U12816(.A(lsu_exu_dfill_data_g[59]), .B(exu_n16313), .Y(exu_n24009));
INVX1 exu_U12817(.A(exu_n24009), .Y(exu_n1815));
AND2X1 exu_U12818(.A(bypass_mux_rcc_data_2_in1[59]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24011));
INVX1 exu_U12819(.A(exu_n24011), .Y(exu_n1816));
AND2X1 exu_U12820(.A(lsu_exu_dfill_data_g[58]), .B(exu_n16313), .Y(exu_n24015));
INVX1 exu_U12821(.A(exu_n24015), .Y(exu_n1817));
AND2X1 exu_U12822(.A(bypass_mux_rcc_data_2_in1[58]), .B(exu_n16314), .Y(exu_n24017));
INVX1 exu_U12823(.A(exu_n24017), .Y(exu_n1818));
AND2X1 exu_U12824(.A(lsu_exu_dfill_data_g[57]), .B(exu_n16313), .Y(exu_n24021));
INVX1 exu_U12825(.A(exu_n24021), .Y(exu_n1819));
AND2X1 exu_U12826(.A(bypass_mux_rcc_data_2_in1[57]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24023));
INVX1 exu_U12827(.A(exu_n24023), .Y(exu_n1820));
AND2X1 exu_U12828(.A(lsu_exu_dfill_data_g[56]), .B(exu_n16313), .Y(exu_n24027));
INVX1 exu_U12829(.A(exu_n24027), .Y(exu_n1821));
AND2X1 exu_U12830(.A(bypass_mux_rcc_data_2_in1[56]), .B(exu_n16314), .Y(exu_n24029));
INVX1 exu_U12831(.A(exu_n24029), .Y(exu_n1822));
AND2X1 exu_U12832(.A(lsu_exu_dfill_data_g[55]), .B(exu_n16313), .Y(exu_n24033));
INVX1 exu_U12833(.A(exu_n24033), .Y(exu_n1823));
AND2X1 exu_U12834(.A(bypass_mux_rcc_data_2_in1[55]), .B(exu_n16314), .Y(exu_n24035));
INVX1 exu_U12835(.A(exu_n24035), .Y(exu_n1824));
AND2X1 exu_U12836(.A(lsu_exu_dfill_data_g[54]), .B(exu_n16313), .Y(exu_n24039));
INVX1 exu_U12837(.A(exu_n24039), .Y(exu_n1825));
AND2X1 exu_U12838(.A(bypass_mux_rcc_data_2_in1[54]), .B(exu_n16314), .Y(exu_n24041));
INVX1 exu_U12839(.A(exu_n24041), .Y(exu_n1826));
AND2X1 exu_U12840(.A(lsu_exu_dfill_data_g[53]), .B(exu_n16313), .Y(exu_n24045));
INVX1 exu_U12841(.A(exu_n24045), .Y(exu_n1827));
AND2X1 exu_U12842(.A(bypass_mux_rcc_data_2_in1[53]), .B(exu_n16314), .Y(exu_n24047));
INVX1 exu_U12843(.A(exu_n24047), .Y(exu_n1828));
AND2X1 exu_U12844(.A(lsu_exu_dfill_data_g[52]), .B(exu_n16313), .Y(exu_n24051));
INVX1 exu_U12845(.A(exu_n24051), .Y(exu_n1829));
AND2X1 exu_U12846(.A(bypass_mux_rcc_data_2_in1[52]), .B(exu_n16314), .Y(exu_n24053));
INVX1 exu_U12847(.A(exu_n24053), .Y(exu_n1830));
AND2X1 exu_U12848(.A(lsu_exu_dfill_data_g[51]), .B(exu_n16313), .Y(exu_n24057));
INVX1 exu_U12849(.A(exu_n24057), .Y(exu_n1831));
AND2X1 exu_U12850(.A(bypass_mux_rcc_data_2_in1[51]), .B(exu_n16314), .Y(exu_n24059));
INVX1 exu_U12851(.A(exu_n24059), .Y(exu_n1832));
AND2X1 exu_U12852(.A(lsu_exu_dfill_data_g[50]), .B(exu_n16313), .Y(exu_n24063));
INVX1 exu_U12853(.A(exu_n24063), .Y(exu_n1833));
AND2X1 exu_U12854(.A(bypass_mux_rcc_data_2_in1[50]), .B(exu_n16314), .Y(exu_n24065));
INVX1 exu_U12855(.A(exu_n24065), .Y(exu_n1834));
AND2X1 exu_U12856(.A(lsu_exu_dfill_data_g[4]), .B(exu_n16313), .Y(exu_n24069));
INVX1 exu_U12857(.A(exu_n24069), .Y(exu_n1835));
AND2X1 exu_U12858(.A(bypass_mux_rcc_data_2_in1[4]), .B(exu_n16314), .Y(exu_n24071));
INVX1 exu_U12859(.A(exu_n24071), .Y(exu_n1836));
AND2X1 exu_U12860(.A(lsu_exu_dfill_data_g[49]), .B(exu_n16313), .Y(exu_n24075));
INVX1 exu_U12861(.A(exu_n24075), .Y(exu_n1837));
AND2X1 exu_U12862(.A(bypass_mux_rcc_data_2_in1[49]), .B(exu_n16314), .Y(exu_n24077));
INVX1 exu_U12863(.A(exu_n24077), .Y(exu_n1838));
AND2X1 exu_U12864(.A(lsu_exu_dfill_data_g[48]), .B(exu_n16313), .Y(exu_n24081));
INVX1 exu_U12865(.A(exu_n24081), .Y(exu_n1839));
AND2X1 exu_U12866(.A(bypass_mux_rcc_data_2_in1[48]), .B(exu_n16314), .Y(exu_n24083));
INVX1 exu_U12867(.A(exu_n24083), .Y(exu_n1840));
AND2X1 exu_U12868(.A(lsu_exu_dfill_data_g[47]), .B(exu_n16313), .Y(exu_n24087));
INVX1 exu_U12869(.A(exu_n24087), .Y(exu_n1841));
AND2X1 exu_U12870(.A(bypass_mux_rcc_data_2_in1[47]), .B(exu_n16314), .Y(exu_n24089));
INVX1 exu_U12871(.A(exu_n24089), .Y(exu_n1842));
AND2X1 exu_U12872(.A(lsu_exu_dfill_data_g[46]), .B(exu_n16313), .Y(exu_n24093));
INVX1 exu_U12873(.A(exu_n24093), .Y(exu_n1843));
AND2X1 exu_U12874(.A(bypass_mux_rcc_data_2_in1[46]), .B(exu_n16314), .Y(exu_n24095));
INVX1 exu_U12875(.A(exu_n24095), .Y(exu_n1844));
AND2X1 exu_U12876(.A(lsu_exu_dfill_data_g[45]), .B(exu_n16313), .Y(exu_n24099));
INVX1 exu_U12877(.A(exu_n24099), .Y(exu_n1845));
AND2X1 exu_U12878(.A(bypass_mux_rcc_data_2_in1[45]), .B(exu_n16314), .Y(exu_n24101));
INVX1 exu_U12879(.A(exu_n24101), .Y(exu_n1846));
AND2X1 exu_U12880(.A(lsu_exu_dfill_data_g[44]), .B(exu_n16313), .Y(exu_n24105));
INVX1 exu_U12881(.A(exu_n24105), .Y(exu_n1847));
AND2X1 exu_U12882(.A(bypass_mux_rcc_data_2_in1[44]), .B(exu_n16314), .Y(exu_n24107));
INVX1 exu_U12883(.A(exu_n24107), .Y(exu_n1848));
AND2X1 exu_U12884(.A(lsu_exu_dfill_data_g[43]), .B(exu_n16313), .Y(exu_n24111));
INVX1 exu_U12885(.A(exu_n24111), .Y(exu_n1849));
AND2X1 exu_U12886(.A(bypass_mux_rcc_data_2_in1[43]), .B(exu_n16314), .Y(exu_n24113));
INVX1 exu_U12887(.A(exu_n24113), .Y(exu_n1850));
AND2X1 exu_U12888(.A(lsu_exu_dfill_data_g[42]), .B(exu_n16313), .Y(exu_n24117));
INVX1 exu_U12889(.A(exu_n24117), .Y(exu_n1851));
AND2X1 exu_U12890(.A(bypass_mux_rcc_data_2_in1[42]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24119));
INVX1 exu_U12891(.A(exu_n24119), .Y(exu_n1852));
AND2X1 exu_U12892(.A(lsu_exu_dfill_data_g[41]), .B(exu_n16313), .Y(exu_n24123));
INVX1 exu_U12893(.A(exu_n24123), .Y(exu_n1853));
AND2X1 exu_U12894(.A(bypass_mux_rcc_data_2_in1[41]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24125));
INVX1 exu_U12895(.A(exu_n24125), .Y(exu_n1854));
AND2X1 exu_U12896(.A(lsu_exu_dfill_data_g[40]), .B(exu_n16313), .Y(exu_n24129));
INVX1 exu_U12897(.A(exu_n24129), .Y(exu_n1855));
AND2X1 exu_U12898(.A(bypass_mux_rcc_data_2_in1[40]), .B(exu_n16314), .Y(exu_n24131));
INVX1 exu_U12899(.A(exu_n24131), .Y(exu_n1856));
AND2X1 exu_U12900(.A(lsu_exu_dfill_data_g[3]), .B(exu_n16313), .Y(exu_n24135));
INVX1 exu_U12901(.A(exu_n24135), .Y(exu_n1857));
AND2X1 exu_U12902(.A(bypass_mux_rcc_data_2_in1[3]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24137));
INVX1 exu_U12903(.A(exu_n24137), .Y(exu_n1858));
AND2X1 exu_U12904(.A(lsu_exu_dfill_data_g[39]), .B(exu_n16313), .Y(exu_n24141));
INVX1 exu_U12905(.A(exu_n24141), .Y(exu_n1859));
AND2X1 exu_U12906(.A(bypass_mux_rcc_data_2_in1[39]), .B(exu_n16314), .Y(exu_n24143));
INVX1 exu_U12907(.A(exu_n24143), .Y(exu_n1860));
AND2X1 exu_U12908(.A(lsu_exu_dfill_data_g[38]), .B(exu_n16313), .Y(exu_n24147));
INVX1 exu_U12909(.A(exu_n24147), .Y(exu_n1861));
AND2X1 exu_U12910(.A(bypass_mux_rcc_data_2_in1[38]), .B(exu_n16314), .Y(exu_n24149));
INVX1 exu_U12911(.A(exu_n24149), .Y(exu_n1862));
AND2X1 exu_U12912(.A(lsu_exu_dfill_data_g[37]), .B(exu_n16313), .Y(exu_n24153));
INVX1 exu_U12913(.A(exu_n24153), .Y(exu_n1863));
AND2X1 exu_U12914(.A(bypass_mux_rcc_data_2_in1[37]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24155));
INVX1 exu_U12915(.A(exu_n24155), .Y(exu_n1864));
AND2X1 exu_U12916(.A(lsu_exu_dfill_data_g[36]), .B(exu_n16313), .Y(exu_n24159));
INVX1 exu_U12917(.A(exu_n24159), .Y(exu_n1865));
AND2X1 exu_U12918(.A(bypass_mux_rcc_data_2_in1[36]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24161));
INVX1 exu_U12919(.A(exu_n24161), .Y(exu_n1866));
AND2X1 exu_U12920(.A(lsu_exu_dfill_data_g[35]), .B(exu_n16313), .Y(exu_n24165));
INVX1 exu_U12921(.A(exu_n24165), .Y(exu_n1867));
AND2X1 exu_U12922(.A(bypass_mux_rcc_data_2_in1[35]), .B(exu_n16314), .Y(exu_n24167));
INVX1 exu_U12923(.A(exu_n24167), .Y(exu_n1868));
AND2X1 exu_U12924(.A(lsu_exu_dfill_data_g[34]), .B(exu_n16313), .Y(exu_n24171));
INVX1 exu_U12925(.A(exu_n24171), .Y(exu_n1869));
AND2X1 exu_U12926(.A(bypass_mux_rcc_data_2_in1[34]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24173));
INVX1 exu_U12927(.A(exu_n24173), .Y(exu_n1870));
AND2X1 exu_U12928(.A(lsu_exu_dfill_data_g[33]), .B(exu_n16313), .Y(exu_n24177));
INVX1 exu_U12929(.A(exu_n24177), .Y(exu_n1871));
AND2X1 exu_U12930(.A(bypass_mux_rcc_data_2_in1[33]), .B(exu_n16314), .Y(exu_n24179));
INVX1 exu_U12931(.A(exu_n24179), .Y(exu_n1872));
AND2X1 exu_U12932(.A(lsu_exu_dfill_data_g[32]), .B(exu_n16313), .Y(exu_n24183));
INVX1 exu_U12933(.A(exu_n24183), .Y(exu_n1873));
AND2X1 exu_U12934(.A(bypass_mux_rcc_data_2_in1[32]), .B(exu_n16314), .Y(exu_n24185));
INVX1 exu_U12935(.A(exu_n24185), .Y(exu_n1874));
AND2X1 exu_U12936(.A(lsu_exu_dfill_data_g[31]), .B(exu_n16313), .Y(exu_n24189));
INVX1 exu_U12937(.A(exu_n24189), .Y(exu_n1875));
AND2X1 exu_U12938(.A(bypass_mux_rcc_data_2_in1[31]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24191));
INVX1 exu_U12939(.A(exu_n24191), .Y(exu_n1876));
AND2X1 exu_U12940(.A(lsu_exu_dfill_data_g[30]), .B(exu_n16313), .Y(exu_n24195));
INVX1 exu_U12941(.A(exu_n24195), .Y(exu_n1877));
AND2X1 exu_U12942(.A(bypass_mux_rcc_data_2_in1[30]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24197));
INVX1 exu_U12943(.A(exu_n24197), .Y(exu_n1878));
AND2X1 exu_U12944(.A(lsu_exu_dfill_data_g[2]), .B(exu_n16313), .Y(exu_n24201));
INVX1 exu_U12945(.A(exu_n24201), .Y(exu_n1879));
AND2X1 exu_U12946(.A(bypass_mux_rcc_data_2_in1[2]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24203));
INVX1 exu_U12947(.A(exu_n24203), .Y(exu_n1880));
AND2X1 exu_U12948(.A(lsu_exu_dfill_data_g[29]), .B(exu_n16313), .Y(exu_n24207));
INVX1 exu_U12949(.A(exu_n24207), .Y(exu_n1881));
AND2X1 exu_U12950(.A(bypass_mux_rcc_data_2_in1[29]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24209));
INVX1 exu_U12951(.A(exu_n24209), .Y(exu_n1882));
AND2X1 exu_U12952(.A(lsu_exu_dfill_data_g[28]), .B(exu_n16313), .Y(exu_n24213));
INVX1 exu_U12953(.A(exu_n24213), .Y(exu_n1883));
AND2X1 exu_U12954(.A(bypass_mux_rcc_data_2_in1[28]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24215));
INVX1 exu_U12955(.A(exu_n24215), .Y(exu_n1884));
AND2X1 exu_U12956(.A(lsu_exu_dfill_data_g[27]), .B(exu_n16313), .Y(exu_n24219));
INVX1 exu_U12957(.A(exu_n24219), .Y(exu_n1885));
AND2X1 exu_U12958(.A(bypass_mux_rcc_data_2_in1[27]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24221));
INVX1 exu_U12959(.A(exu_n24221), .Y(exu_n1886));
AND2X1 exu_U12960(.A(lsu_exu_dfill_data_g[26]), .B(exu_n16313), .Y(exu_n24225));
INVX1 exu_U12961(.A(exu_n24225), .Y(exu_n1887));
AND2X1 exu_U12962(.A(bypass_mux_rcc_data_2_in1[26]), .B(exu_n16314), .Y(exu_n24227));
INVX1 exu_U12963(.A(exu_n24227), .Y(exu_n1888));
AND2X1 exu_U12964(.A(lsu_exu_dfill_data_g[25]), .B(exu_n16313), .Y(exu_n24231));
INVX1 exu_U12965(.A(exu_n24231), .Y(exu_n1889));
AND2X1 exu_U12966(.A(bypass_mux_rcc_data_2_in1[25]), .B(exu_n16314), .Y(exu_n24233));
INVX1 exu_U12967(.A(exu_n24233), .Y(exu_n1890));
AND2X1 exu_U12968(.A(lsu_exu_dfill_data_g[24]), .B(exu_n16313), .Y(exu_n24237));
INVX1 exu_U12969(.A(exu_n24237), .Y(exu_n1891));
AND2X1 exu_U12970(.A(bypass_mux_rcc_data_2_in1[24]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24239));
INVX1 exu_U12971(.A(exu_n24239), .Y(exu_n1892));
AND2X1 exu_U12972(.A(lsu_exu_dfill_data_g[23]), .B(exu_n16313), .Y(exu_n24243));
INVX1 exu_U12973(.A(exu_n24243), .Y(exu_n1893));
AND2X1 exu_U12974(.A(bypass_mux_rcc_data_2_in1[23]), .B(exu_n16314), .Y(exu_n24245));
INVX1 exu_U12975(.A(exu_n24245), .Y(exu_n1894));
AND2X1 exu_U12976(.A(lsu_exu_dfill_data_g[22]), .B(exu_n16313), .Y(exu_n24249));
INVX1 exu_U12977(.A(exu_n24249), .Y(exu_n1895));
AND2X1 exu_U12978(.A(bypass_mux_rcc_data_2_in1[22]), .B(exu_n16314), .Y(exu_n24251));
INVX1 exu_U12979(.A(exu_n24251), .Y(exu_n1896));
AND2X1 exu_U12980(.A(lsu_exu_dfill_data_g[21]), .B(exu_n16313), .Y(exu_n24255));
INVX1 exu_U12981(.A(exu_n24255), .Y(exu_n1897));
AND2X1 exu_U12982(.A(bypass_mux_rcc_data_2_in1[21]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24257));
INVX1 exu_U12983(.A(exu_n24257), .Y(exu_n1898));
AND2X1 exu_U12984(.A(lsu_exu_dfill_data_g[20]), .B(exu_n16313), .Y(exu_n24261));
INVX1 exu_U12985(.A(exu_n24261), .Y(exu_n1899));
AND2X1 exu_U12986(.A(bypass_mux_rcc_data_2_in1[20]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24263));
INVX1 exu_U12987(.A(exu_n24263), .Y(exu_n1900));
AND2X1 exu_U12988(.A(lsu_exu_dfill_data_g[1]), .B(exu_n16313), .Y(exu_n24267));
INVX1 exu_U12989(.A(exu_n24267), .Y(exu_n1901));
AND2X1 exu_U12990(.A(bypass_mux_rcc_data_2_in1[1]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24269));
INVX1 exu_U12991(.A(exu_n24269), .Y(exu_n1902));
AND2X1 exu_U12992(.A(lsu_exu_dfill_data_g[19]), .B(exu_n16313), .Y(exu_n24273));
INVX1 exu_U12993(.A(exu_n24273), .Y(exu_n1903));
AND2X1 exu_U12994(.A(bypass_mux_rcc_data_2_in1[19]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24275));
INVX1 exu_U12995(.A(exu_n24275), .Y(exu_n1904));
AND2X1 exu_U12996(.A(lsu_exu_dfill_data_g[18]), .B(exu_n16313), .Y(exu_n24279));
INVX1 exu_U12997(.A(exu_n24279), .Y(exu_n1905));
AND2X1 exu_U12998(.A(bypass_mux_rcc_data_2_in1[18]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24281));
INVX1 exu_U12999(.A(exu_n24281), .Y(exu_n1906));
AND2X1 exu_U13000(.A(lsu_exu_dfill_data_g[17]), .B(exu_n16313), .Y(exu_n24285));
INVX1 exu_U13001(.A(exu_n24285), .Y(exu_n1907));
AND2X1 exu_U13002(.A(bypass_mux_rcc_data_2_in1[17]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24287));
INVX1 exu_U13003(.A(exu_n24287), .Y(exu_n1908));
AND2X1 exu_U13004(.A(lsu_exu_dfill_data_g[16]), .B(exu_n16313), .Y(exu_n24291));
INVX1 exu_U13005(.A(exu_n24291), .Y(exu_n1909));
AND2X1 exu_U13006(.A(bypass_mux_rcc_data_2_in1[16]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24293));
INVX1 exu_U13007(.A(exu_n24293), .Y(exu_n1910));
AND2X1 exu_U13008(.A(lsu_exu_dfill_data_g[15]), .B(exu_n16313), .Y(exu_n24297));
INVX1 exu_U13009(.A(exu_n24297), .Y(exu_n1911));
AND2X1 exu_U13010(.A(bypass_mux_rcc_data_2_in1[15]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24299));
INVX1 exu_U13011(.A(exu_n24299), .Y(exu_n1912));
AND2X1 exu_U13012(.A(lsu_exu_dfill_data_g[14]), .B(exu_n16313), .Y(exu_n24303));
INVX1 exu_U13013(.A(exu_n24303), .Y(exu_n1913));
AND2X1 exu_U13014(.A(bypass_mux_rcc_data_2_in1[14]), .B(exu_n16314), .Y(exu_n24305));
INVX1 exu_U13015(.A(exu_n24305), .Y(exu_n1914));
AND2X1 exu_U13016(.A(lsu_exu_dfill_data_g[13]), .B(exu_n16313), .Y(exu_n24309));
INVX1 exu_U13017(.A(exu_n24309), .Y(exu_n1915));
AND2X1 exu_U13018(.A(bypass_mux_rcc_data_2_in1[13]), .B(exu_n16314), .Y(exu_n24311));
INVX1 exu_U13019(.A(exu_n24311), .Y(exu_n1916));
AND2X1 exu_U13020(.A(lsu_exu_dfill_data_g[12]), .B(exu_n16313), .Y(exu_n24315));
INVX1 exu_U13021(.A(exu_n24315), .Y(exu_n1917));
AND2X1 exu_U13022(.A(bypass_mux_rcc_data_2_in1[12]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24317));
INVX1 exu_U13023(.A(exu_n24317), .Y(exu_n1918));
AND2X1 exu_U13024(.A(lsu_exu_dfill_data_g[11]), .B(exu_n16313), .Y(exu_n24321));
INVX1 exu_U13025(.A(exu_n24321), .Y(exu_n1919));
AND2X1 exu_U13026(.A(bypass_mux_rcc_data_2_in1[11]), .B(ecl_byp_rs1_mux2_sel_rf), .Y(exu_n24323));
INVX1 exu_U13027(.A(exu_n24323), .Y(exu_n1920));
AND2X1 exu_U13028(.A(lsu_exu_dfill_data_g[10]), .B(exu_n16313), .Y(exu_n24327));
INVX1 exu_U13029(.A(exu_n24327), .Y(exu_n1921));
AND2X1 exu_U13030(.A(bypass_mux_rcc_data_2_in1[10]), .B(exu_n16314), .Y(exu_n24329));
INVX1 exu_U13031(.A(exu_n24329), .Y(exu_n1922));
AND2X1 exu_U13032(.A(lsu_exu_dfill_data_g[0]), .B(exu_n16313), .Y(exu_n24333));
INVX1 exu_U13033(.A(exu_n24333), .Y(exu_n1923));
AND2X1 exu_U13034(.A(bypass_mux_rcc_data_2_in1[0]), .B(exu_n16314), .Y(exu_n24335));
INVX1 exu_U13035(.A(exu_n24335), .Y(exu_n1924));
AND2X1 exu_U13036(.A(exu_n16301), .B(byp_irf_rd_data_w[9]), .Y(exu_n24339));
INVX1 exu_U13037(.A(exu_n24339), .Y(exu_n1925));
AND2X1 exu_U13038(.A(byp_irf_rd_data_w[8]), .B(exu_n16301), .Y(exu_n24343));
INVX1 exu_U13039(.A(exu_n24343), .Y(exu_n1926));
AND2X1 exu_U13040(.A(byp_irf_rd_data_w[7]), .B(exu_n16301), .Y(exu_n24347));
INVX1 exu_U13041(.A(exu_n24347), .Y(exu_n1927));
AND2X1 exu_U13042(.A(byp_irf_rd_data_w[6]), .B(exu_n16301), .Y(exu_n24351));
INVX1 exu_U13043(.A(exu_n24351), .Y(exu_n1928));
AND2X1 exu_U13044(.A(byp_irf_rd_data_w[63]), .B(exu_n16301), .Y(exu_n24355));
INVX1 exu_U13045(.A(exu_n24355), .Y(exu_n1929));
AND2X1 exu_U13046(.A(byp_irf_rd_data_w[62]), .B(exu_n16301), .Y(exu_n24359));
INVX1 exu_U13047(.A(exu_n24359), .Y(exu_n1930));
AND2X1 exu_U13048(.A(byp_irf_rd_data_w[61]), .B(exu_n16301), .Y(exu_n24363));
INVX1 exu_U13049(.A(exu_n24363), .Y(exu_n1931));
AND2X1 exu_U13050(.A(byp_irf_rd_data_w[60]), .B(exu_n16301), .Y(exu_n24367));
INVX1 exu_U13051(.A(exu_n24367), .Y(exu_n1932));
AND2X1 exu_U13052(.A(byp_irf_rd_data_w[5]), .B(exu_n16301), .Y(exu_n24371));
INVX1 exu_U13053(.A(exu_n24371), .Y(exu_n1933));
AND2X1 exu_U13054(.A(byp_irf_rd_data_w[59]), .B(exu_n16301), .Y(exu_n24375));
INVX1 exu_U13055(.A(exu_n24375), .Y(exu_n1934));
AND2X1 exu_U13056(.A(byp_irf_rd_data_w[58]), .B(exu_n16301), .Y(exu_n24379));
INVX1 exu_U13057(.A(exu_n24379), .Y(exu_n1935));
AND2X1 exu_U13058(.A(byp_irf_rd_data_w[57]), .B(exu_n16301), .Y(exu_n24383));
INVX1 exu_U13059(.A(exu_n24383), .Y(exu_n1936));
AND2X1 exu_U13060(.A(byp_irf_rd_data_w[56]), .B(exu_n16301), .Y(exu_n24387));
INVX1 exu_U13061(.A(exu_n24387), .Y(exu_n1937));
AND2X1 exu_U13062(.A(byp_irf_rd_data_w[55]), .B(exu_n16301), .Y(exu_n24391));
INVX1 exu_U13063(.A(exu_n24391), .Y(exu_n1938));
AND2X1 exu_U13064(.A(byp_irf_rd_data_w[54]), .B(exu_n16301), .Y(exu_n24395));
INVX1 exu_U13065(.A(exu_n24395), .Y(exu_n1939));
AND2X1 exu_U13066(.A(byp_irf_rd_data_w[53]), .B(exu_n16301), .Y(exu_n24399));
INVX1 exu_U13067(.A(exu_n24399), .Y(exu_n1940));
AND2X1 exu_U13068(.A(byp_irf_rd_data_w[52]), .B(exu_n16301), .Y(exu_n24403));
INVX1 exu_U13069(.A(exu_n24403), .Y(exu_n1941));
AND2X1 exu_U13070(.A(byp_irf_rd_data_w[51]), .B(exu_n16301), .Y(exu_n24407));
INVX1 exu_U13071(.A(exu_n24407), .Y(exu_n1942));
AND2X1 exu_U13072(.A(byp_irf_rd_data_w[50]), .B(exu_n16301), .Y(exu_n24411));
INVX1 exu_U13073(.A(exu_n24411), .Y(exu_n1943));
AND2X1 exu_U13074(.A(byp_irf_rd_data_w[4]), .B(exu_n16301), .Y(exu_n24415));
INVX1 exu_U13075(.A(exu_n24415), .Y(exu_n1944));
AND2X1 exu_U13076(.A(byp_irf_rd_data_w[49]), .B(exu_n16301), .Y(exu_n24419));
INVX1 exu_U13077(.A(exu_n24419), .Y(exu_n1945));
AND2X1 exu_U13078(.A(byp_irf_rd_data_w[48]), .B(exu_n16301), .Y(exu_n24423));
INVX1 exu_U13079(.A(exu_n24423), .Y(exu_n1946));
AND2X1 exu_U13080(.A(byp_irf_rd_data_w[47]), .B(exu_n16301), .Y(exu_n24427));
INVX1 exu_U13081(.A(exu_n24427), .Y(exu_n1947));
AND2X1 exu_U13082(.A(byp_irf_rd_data_w[46]), .B(exu_n16301), .Y(exu_n24431));
INVX1 exu_U13083(.A(exu_n24431), .Y(exu_n1948));
AND2X1 exu_U13084(.A(byp_irf_rd_data_w[45]), .B(exu_n16301), .Y(exu_n24435));
INVX1 exu_U13085(.A(exu_n24435), .Y(exu_n1949));
AND2X1 exu_U13086(.A(byp_irf_rd_data_w[44]), .B(exu_n16301), .Y(exu_n24439));
INVX1 exu_U13087(.A(exu_n24439), .Y(exu_n1950));
AND2X1 exu_U13088(.A(byp_irf_rd_data_w[43]), .B(exu_n16301), .Y(exu_n24443));
INVX1 exu_U13089(.A(exu_n24443), .Y(exu_n1951));
AND2X1 exu_U13090(.A(byp_irf_rd_data_w[42]), .B(exu_n16301), .Y(exu_n24447));
INVX1 exu_U13091(.A(exu_n24447), .Y(exu_n1952));
AND2X1 exu_U13092(.A(byp_irf_rd_data_w[41]), .B(exu_n16301), .Y(exu_n24451));
INVX1 exu_U13093(.A(exu_n24451), .Y(exu_n1953));
AND2X1 exu_U13094(.A(byp_irf_rd_data_w[40]), .B(exu_n16301), .Y(exu_n24455));
INVX1 exu_U13095(.A(exu_n24455), .Y(exu_n1954));
AND2X1 exu_U13096(.A(byp_irf_rd_data_w[3]), .B(exu_n16301), .Y(exu_n24459));
INVX1 exu_U13097(.A(exu_n24459), .Y(exu_n1955));
AND2X1 exu_U13098(.A(byp_irf_rd_data_w[39]), .B(exu_n16301), .Y(exu_n24463));
INVX1 exu_U13099(.A(exu_n24463), .Y(exu_n1956));
AND2X1 exu_U13100(.A(byp_irf_rd_data_w[38]), .B(exu_n16301), .Y(exu_n24467));
INVX1 exu_U13101(.A(exu_n24467), .Y(exu_n1957));
AND2X1 exu_U13102(.A(byp_irf_rd_data_w[37]), .B(exu_n16301), .Y(exu_n24471));
INVX1 exu_U13103(.A(exu_n24471), .Y(exu_n1958));
AND2X1 exu_U13104(.A(byp_irf_rd_data_w[36]), .B(exu_n16301), .Y(exu_n24475));
INVX1 exu_U13105(.A(exu_n24475), .Y(exu_n1959));
AND2X1 exu_U13106(.A(byp_irf_rd_data_w[35]), .B(exu_n16301), .Y(exu_n24479));
INVX1 exu_U13107(.A(exu_n24479), .Y(exu_n1960));
AND2X1 exu_U13108(.A(byp_irf_rd_data_w[34]), .B(exu_n16301), .Y(exu_n24483));
INVX1 exu_U13109(.A(exu_n24483), .Y(exu_n1961));
AND2X1 exu_U13110(.A(byp_irf_rd_data_w[33]), .B(exu_n16301), .Y(exu_n24487));
INVX1 exu_U13111(.A(exu_n24487), .Y(exu_n1962));
AND2X1 exu_U13112(.A(byp_irf_rd_data_w[32]), .B(exu_n16301), .Y(exu_n24491));
INVX1 exu_U13113(.A(exu_n24491), .Y(exu_n1963));
AND2X1 exu_U13114(.A(byp_irf_rd_data_w[31]), .B(exu_n16301), .Y(exu_n24495));
INVX1 exu_U13115(.A(exu_n24495), .Y(exu_n1964));
AND2X1 exu_U13116(.A(byp_irf_rd_data_w[30]), .B(exu_n16301), .Y(exu_n24499));
INVX1 exu_U13117(.A(exu_n24499), .Y(exu_n1965));
AND2X1 exu_U13118(.A(byp_irf_rd_data_w[2]), .B(exu_n16301), .Y(exu_n24503));
INVX1 exu_U13119(.A(exu_n24503), .Y(exu_n1966));
AND2X1 exu_U13120(.A(byp_irf_rd_data_w[29]), .B(exu_n16301), .Y(exu_n24507));
INVX1 exu_U13121(.A(exu_n24507), .Y(exu_n1967));
AND2X1 exu_U13122(.A(byp_irf_rd_data_w[28]), .B(exu_n16301), .Y(exu_n24511));
INVX1 exu_U13123(.A(exu_n24511), .Y(exu_n1968));
AND2X1 exu_U13124(.A(byp_irf_rd_data_w[27]), .B(exu_n16301), .Y(exu_n24515));
INVX1 exu_U13125(.A(exu_n24515), .Y(exu_n1969));
AND2X1 exu_U13126(.A(byp_irf_rd_data_w[26]), .B(exu_n16301), .Y(exu_n24519));
INVX1 exu_U13127(.A(exu_n24519), .Y(exu_n1970));
AND2X1 exu_U13128(.A(byp_irf_rd_data_w[25]), .B(exu_n16301), .Y(exu_n24523));
INVX1 exu_U13129(.A(exu_n24523), .Y(exu_n1971));
AND2X1 exu_U13130(.A(byp_irf_rd_data_w[24]), .B(exu_n16301), .Y(exu_n24527));
INVX1 exu_U13131(.A(exu_n24527), .Y(exu_n1972));
AND2X1 exu_U13132(.A(byp_irf_rd_data_w[23]), .B(exu_n16301), .Y(exu_n24531));
INVX1 exu_U13133(.A(exu_n24531), .Y(exu_n1973));
AND2X1 exu_U13134(.A(byp_irf_rd_data_w[22]), .B(exu_n16301), .Y(exu_n24535));
INVX1 exu_U13135(.A(exu_n24535), .Y(exu_n1974));
AND2X1 exu_U13136(.A(byp_irf_rd_data_w[21]), .B(exu_n16301), .Y(exu_n24539));
INVX1 exu_U13137(.A(exu_n24539), .Y(exu_n1975));
AND2X1 exu_U13138(.A(byp_irf_rd_data_w[20]), .B(exu_n16301), .Y(exu_n24543));
INVX1 exu_U13139(.A(exu_n24543), .Y(exu_n1976));
AND2X1 exu_U13140(.A(byp_irf_rd_data_w[1]), .B(exu_n16301), .Y(exu_n24547));
INVX1 exu_U13141(.A(exu_n24547), .Y(exu_n1977));
AND2X1 exu_U13142(.A(byp_irf_rd_data_w[19]), .B(exu_n16301), .Y(exu_n24551));
INVX1 exu_U13143(.A(exu_n24551), .Y(exu_n1978));
AND2X1 exu_U13144(.A(byp_irf_rd_data_w[18]), .B(exu_n16301), .Y(exu_n24555));
INVX1 exu_U13145(.A(exu_n24555), .Y(exu_n1979));
AND2X1 exu_U13146(.A(byp_irf_rd_data_w[17]), .B(exu_n16301), .Y(exu_n24559));
INVX1 exu_U13147(.A(exu_n24559), .Y(exu_n1980));
AND2X1 exu_U13148(.A(byp_irf_rd_data_w[16]), .B(exu_n16301), .Y(exu_n24563));
INVX1 exu_U13149(.A(exu_n24563), .Y(exu_n1981));
AND2X1 exu_U13150(.A(byp_irf_rd_data_w[15]), .B(exu_n16301), .Y(exu_n24567));
INVX1 exu_U13151(.A(exu_n24567), .Y(exu_n1982));
AND2X1 exu_U13152(.A(byp_irf_rd_data_w[14]), .B(exu_n16301), .Y(exu_n24571));
INVX1 exu_U13153(.A(exu_n24571), .Y(exu_n1983));
AND2X1 exu_U13154(.A(byp_irf_rd_data_w[13]), .B(exu_n16301), .Y(exu_n24575));
INVX1 exu_U13155(.A(exu_n24575), .Y(exu_n1984));
AND2X1 exu_U13156(.A(byp_irf_rd_data_w[12]), .B(exu_n16301), .Y(exu_n24579));
INVX1 exu_U13157(.A(exu_n24579), .Y(exu_n1985));
AND2X1 exu_U13158(.A(byp_irf_rd_data_w[11]), .B(exu_n16301), .Y(exu_n24583));
INVX1 exu_U13159(.A(exu_n24583), .Y(exu_n1986));
AND2X1 exu_U13160(.A(byp_irf_rd_data_w[10]), .B(exu_n16301), .Y(exu_n24587));
INVX1 exu_U13161(.A(exu_n24587), .Y(exu_n1987));
AND2X1 exu_U13162(.A(byp_irf_rd_data_w[0]), .B(exu_n16301), .Y(exu_n24591));
INVX1 exu_U13163(.A(exu_n24591), .Y(exu_n1988));
AND2X1 exu_U13164(.A(exu_n16304), .B(lsu_exu_dfill_data_g[9]), .Y(exu_n24595));
INVX1 exu_U13165(.A(exu_n24595), .Y(exu_n1989));
AND2X1 exu_U13166(.A(exu_n16305), .B(bypass_mux_rcc_data_2_in1[9]), .Y(exu_n24597));
INVX1 exu_U13167(.A(exu_n24597), .Y(exu_n1990));
AND2X1 exu_U13168(.A(lsu_exu_dfill_data_g[8]), .B(exu_n16304), .Y(exu_n24601));
INVX1 exu_U13169(.A(exu_n24601), .Y(exu_n1991));
AND2X1 exu_U13170(.A(bypass_mux_rcc_data_2_in1[8]), .B(exu_n16305), .Y(exu_n24603));
INVX1 exu_U13171(.A(exu_n24603), .Y(exu_n1992));
AND2X1 exu_U13172(.A(lsu_exu_dfill_data_g[7]), .B(exu_n16304), .Y(exu_n24607));
INVX1 exu_U13173(.A(exu_n24607), .Y(exu_n1993));
AND2X1 exu_U13174(.A(bypass_mux_rcc_data_2_in1[7]), .B(exu_n16305), .Y(exu_n24609));
INVX1 exu_U13175(.A(exu_n24609), .Y(exu_n1994));
AND2X1 exu_U13176(.A(lsu_exu_dfill_data_g[6]), .B(exu_n16304), .Y(exu_n24613));
INVX1 exu_U13177(.A(exu_n24613), .Y(exu_n1995));
AND2X1 exu_U13178(.A(bypass_mux_rcc_data_2_in1[6]), .B(exu_n16305), .Y(exu_n24615));
INVX1 exu_U13179(.A(exu_n24615), .Y(exu_n1996));
AND2X1 exu_U13180(.A(lsu_exu_dfill_data_g[63]), .B(exu_n16304), .Y(exu_n24619));
INVX1 exu_U13181(.A(exu_n24619), .Y(exu_n1997));
AND2X1 exu_U13182(.A(bypass_mux_rcc_data_2_in1[63]), .B(exu_n16305), .Y(exu_n24621));
INVX1 exu_U13183(.A(exu_n24621), .Y(exu_n1998));
AND2X1 exu_U13184(.A(lsu_exu_dfill_data_g[62]), .B(exu_n16304), .Y(exu_n24625));
INVX1 exu_U13185(.A(exu_n24625), .Y(exu_n1999));
AND2X1 exu_U13186(.A(bypass_mux_rcc_data_2_in1[62]), .B(exu_n16305), .Y(exu_n24627));
INVX1 exu_U13187(.A(exu_n24627), .Y(exu_n2000));
AND2X1 exu_U13188(.A(lsu_exu_dfill_data_g[61]), .B(exu_n16304), .Y(exu_n24631));
INVX1 exu_U13189(.A(exu_n24631), .Y(exu_n2001));
AND2X1 exu_U13190(.A(bypass_mux_rcc_data_2_in1[61]), .B(exu_n16305), .Y(exu_n24633));
INVX1 exu_U13191(.A(exu_n24633), .Y(exu_n2002));
AND2X1 exu_U13192(.A(lsu_exu_dfill_data_g[60]), .B(exu_n16304), .Y(exu_n24637));
INVX1 exu_U13193(.A(exu_n24637), .Y(exu_n2003));
AND2X1 exu_U13194(.A(bypass_mux_rcc_data_2_in1[60]), .B(exu_n16305), .Y(exu_n24639));
INVX1 exu_U13195(.A(exu_n24639), .Y(exu_n2004));
AND2X1 exu_U13196(.A(lsu_exu_dfill_data_g[5]), .B(exu_n16304), .Y(exu_n24643));
INVX1 exu_U13197(.A(exu_n24643), .Y(exu_n2005));
AND2X1 exu_U13198(.A(bypass_mux_rcc_data_2_in1[5]), .B(exu_n16305), .Y(exu_n24645));
INVX1 exu_U13199(.A(exu_n24645), .Y(exu_n2006));
AND2X1 exu_U13200(.A(lsu_exu_dfill_data_g[59]), .B(exu_n16304), .Y(exu_n24649));
INVX1 exu_U13201(.A(exu_n24649), .Y(exu_n2007));
AND2X1 exu_U13202(.A(bypass_mux_rcc_data_2_in1[59]), .B(exu_n16305), .Y(exu_n24651));
INVX1 exu_U13203(.A(exu_n24651), .Y(exu_n2008));
AND2X1 exu_U13204(.A(lsu_exu_dfill_data_g[58]), .B(exu_n16304), .Y(exu_n24655));
INVX1 exu_U13205(.A(exu_n24655), .Y(exu_n2009));
AND2X1 exu_U13206(.A(bypass_mux_rcc_data_2_in1[58]), .B(exu_n16305), .Y(exu_n24657));
INVX1 exu_U13207(.A(exu_n24657), .Y(exu_n2010));
AND2X1 exu_U13208(.A(lsu_exu_dfill_data_g[57]), .B(exu_n16304), .Y(exu_n24661));
INVX1 exu_U13209(.A(exu_n24661), .Y(exu_n2011));
AND2X1 exu_U13210(.A(bypass_mux_rcc_data_2_in1[57]), .B(exu_n16305), .Y(exu_n24663));
INVX1 exu_U13211(.A(exu_n24663), .Y(exu_n2012));
AND2X1 exu_U13212(.A(lsu_exu_dfill_data_g[56]), .B(exu_n16304), .Y(exu_n24667));
INVX1 exu_U13213(.A(exu_n24667), .Y(exu_n2013));
AND2X1 exu_U13214(.A(bypass_mux_rcc_data_2_in1[56]), .B(exu_n16305), .Y(exu_n24669));
INVX1 exu_U13215(.A(exu_n24669), .Y(exu_n2014));
AND2X1 exu_U13216(.A(lsu_exu_dfill_data_g[55]), .B(exu_n16304), .Y(exu_n24673));
INVX1 exu_U13217(.A(exu_n24673), .Y(exu_n2015));
AND2X1 exu_U13218(.A(bypass_mux_rcc_data_2_in1[55]), .B(exu_n16305), .Y(exu_n24675));
INVX1 exu_U13219(.A(exu_n24675), .Y(exu_n2016));
AND2X1 exu_U13220(.A(lsu_exu_dfill_data_g[54]), .B(exu_n16304), .Y(exu_n24679));
INVX1 exu_U13221(.A(exu_n24679), .Y(exu_n2017));
AND2X1 exu_U13222(.A(bypass_mux_rcc_data_2_in1[54]), .B(exu_n16305), .Y(exu_n24681));
INVX1 exu_U13223(.A(exu_n24681), .Y(exu_n2018));
AND2X1 exu_U13224(.A(lsu_exu_dfill_data_g[53]), .B(exu_n16304), .Y(exu_n24685));
INVX1 exu_U13225(.A(exu_n24685), .Y(exu_n2019));
AND2X1 exu_U13226(.A(bypass_mux_rcc_data_2_in1[53]), .B(exu_n16305), .Y(exu_n24687));
INVX1 exu_U13227(.A(exu_n24687), .Y(exu_n2020));
AND2X1 exu_U13228(.A(lsu_exu_dfill_data_g[52]), .B(exu_n16304), .Y(exu_n24691));
INVX1 exu_U13229(.A(exu_n24691), .Y(exu_n2021));
AND2X1 exu_U13230(.A(bypass_mux_rcc_data_2_in1[52]), .B(exu_n16305), .Y(exu_n24693));
INVX1 exu_U13231(.A(exu_n24693), .Y(exu_n2022));
AND2X1 exu_U13232(.A(lsu_exu_dfill_data_g[51]), .B(exu_n16304), .Y(exu_n24697));
INVX1 exu_U13233(.A(exu_n24697), .Y(exu_n2023));
AND2X1 exu_U13234(.A(bypass_mux_rcc_data_2_in1[51]), .B(exu_n16305), .Y(exu_n24699));
INVX1 exu_U13235(.A(exu_n24699), .Y(exu_n2024));
AND2X1 exu_U13236(.A(lsu_exu_dfill_data_g[50]), .B(exu_n16304), .Y(exu_n24703));
INVX1 exu_U13237(.A(exu_n24703), .Y(exu_n2025));
AND2X1 exu_U13238(.A(bypass_mux_rcc_data_2_in1[50]), .B(exu_n16305), .Y(exu_n24705));
INVX1 exu_U13239(.A(exu_n24705), .Y(exu_n2026));
AND2X1 exu_U13240(.A(lsu_exu_dfill_data_g[4]), .B(exu_n16304), .Y(exu_n24709));
INVX1 exu_U13241(.A(exu_n24709), .Y(exu_n2027));
AND2X1 exu_U13242(.A(bypass_mux_rcc_data_2_in1[4]), .B(exu_n16305), .Y(exu_n24711));
INVX1 exu_U13243(.A(exu_n24711), .Y(exu_n2028));
AND2X1 exu_U13244(.A(lsu_exu_dfill_data_g[49]), .B(exu_n16304), .Y(exu_n24715));
INVX1 exu_U13245(.A(exu_n24715), .Y(exu_n2029));
AND2X1 exu_U13246(.A(bypass_mux_rcc_data_2_in1[49]), .B(exu_n16305), .Y(exu_n24717));
INVX1 exu_U13247(.A(exu_n24717), .Y(exu_n2030));
AND2X1 exu_U13248(.A(lsu_exu_dfill_data_g[48]), .B(exu_n16304), .Y(exu_n24721));
INVX1 exu_U13249(.A(exu_n24721), .Y(exu_n2031));
AND2X1 exu_U13250(.A(bypass_mux_rcc_data_2_in1[48]), .B(exu_n16305), .Y(exu_n24723));
INVX1 exu_U13251(.A(exu_n24723), .Y(exu_n2032));
AND2X1 exu_U13252(.A(lsu_exu_dfill_data_g[47]), .B(exu_n16304), .Y(exu_n24727));
INVX1 exu_U13253(.A(exu_n24727), .Y(exu_n2033));
AND2X1 exu_U13254(.A(bypass_mux_rcc_data_2_in1[47]), .B(exu_n16305), .Y(exu_n24729));
INVX1 exu_U13255(.A(exu_n24729), .Y(exu_n2034));
AND2X1 exu_U13256(.A(lsu_exu_dfill_data_g[46]), .B(exu_n16304), .Y(exu_n24733));
INVX1 exu_U13257(.A(exu_n24733), .Y(exu_n2035));
AND2X1 exu_U13258(.A(bypass_mux_rcc_data_2_in1[46]), .B(exu_n16305), .Y(exu_n24735));
INVX1 exu_U13259(.A(exu_n24735), .Y(exu_n2036));
AND2X1 exu_U13260(.A(lsu_exu_dfill_data_g[45]), .B(exu_n16304), .Y(exu_n24739));
INVX1 exu_U13261(.A(exu_n24739), .Y(exu_n2037));
AND2X1 exu_U13262(.A(bypass_mux_rcc_data_2_in1[45]), .B(exu_n16305), .Y(exu_n24741));
INVX1 exu_U13263(.A(exu_n24741), .Y(exu_n2038));
AND2X1 exu_U13264(.A(lsu_exu_dfill_data_g[44]), .B(exu_n16304), .Y(exu_n24745));
INVX1 exu_U13265(.A(exu_n24745), .Y(exu_n2039));
AND2X1 exu_U13266(.A(bypass_mux_rcc_data_2_in1[44]), .B(exu_n16305), .Y(exu_n24747));
INVX1 exu_U13267(.A(exu_n24747), .Y(exu_n2040));
AND2X1 exu_U13268(.A(lsu_exu_dfill_data_g[43]), .B(exu_n16304), .Y(exu_n24751));
INVX1 exu_U13269(.A(exu_n24751), .Y(exu_n2041));
AND2X1 exu_U13270(.A(bypass_mux_rcc_data_2_in1[43]), .B(exu_n16305), .Y(exu_n24753));
INVX1 exu_U13271(.A(exu_n24753), .Y(exu_n2042));
AND2X1 exu_U13272(.A(lsu_exu_dfill_data_g[42]), .B(exu_n16304), .Y(exu_n24757));
INVX1 exu_U13273(.A(exu_n24757), .Y(exu_n2043));
AND2X1 exu_U13274(.A(bypass_mux_rcc_data_2_in1[42]), .B(exu_n16305), .Y(exu_n24759));
INVX1 exu_U13275(.A(exu_n24759), .Y(exu_n2044));
AND2X1 exu_U13276(.A(lsu_exu_dfill_data_g[41]), .B(exu_n16304), .Y(exu_n24763));
INVX1 exu_U13277(.A(exu_n24763), .Y(exu_n2045));
AND2X1 exu_U13278(.A(bypass_mux_rcc_data_2_in1[41]), .B(exu_n16305), .Y(exu_n24765));
INVX1 exu_U13279(.A(exu_n24765), .Y(exu_n2046));
AND2X1 exu_U13280(.A(lsu_exu_dfill_data_g[40]), .B(exu_n16304), .Y(exu_n24769));
INVX1 exu_U13281(.A(exu_n24769), .Y(exu_n2047));
AND2X1 exu_U13282(.A(bypass_mux_rcc_data_2_in1[40]), .B(exu_n16305), .Y(exu_n24771));
INVX1 exu_U13283(.A(exu_n24771), .Y(exu_n2048));
AND2X1 exu_U13284(.A(lsu_exu_dfill_data_g[3]), .B(exu_n16304), .Y(exu_n24775));
INVX1 exu_U13285(.A(exu_n24775), .Y(exu_n2049));
AND2X1 exu_U13286(.A(bypass_mux_rcc_data_2_in1[3]), .B(exu_n16305), .Y(exu_n24777));
INVX1 exu_U13287(.A(exu_n24777), .Y(exu_n2050));
AND2X1 exu_U13288(.A(lsu_exu_dfill_data_g[39]), .B(exu_n16304), .Y(exu_n24781));
INVX1 exu_U13289(.A(exu_n24781), .Y(exu_n2051));
AND2X1 exu_U13290(.A(bypass_mux_rcc_data_2_in1[39]), .B(exu_n16305), .Y(exu_n24783));
INVX1 exu_U13291(.A(exu_n24783), .Y(exu_n2052));
AND2X1 exu_U13292(.A(lsu_exu_dfill_data_g[38]), .B(exu_n16304), .Y(exu_n24787));
INVX1 exu_U13293(.A(exu_n24787), .Y(exu_n2053));
AND2X1 exu_U13294(.A(bypass_mux_rcc_data_2_in1[38]), .B(exu_n16305), .Y(exu_n24789));
INVX1 exu_U13295(.A(exu_n24789), .Y(exu_n2054));
AND2X1 exu_U13296(.A(lsu_exu_dfill_data_g[37]), .B(exu_n16304), .Y(exu_n24793));
INVX1 exu_U13297(.A(exu_n24793), .Y(exu_n2055));
AND2X1 exu_U13298(.A(bypass_mux_rcc_data_2_in1[37]), .B(exu_n16305), .Y(exu_n24795));
INVX1 exu_U13299(.A(exu_n24795), .Y(exu_n2056));
AND2X1 exu_U13300(.A(lsu_exu_dfill_data_g[36]), .B(exu_n16304), .Y(exu_n24799));
INVX1 exu_U13301(.A(exu_n24799), .Y(exu_n2057));
AND2X1 exu_U13302(.A(bypass_mux_rcc_data_2_in1[36]), .B(exu_n16305), .Y(exu_n24801));
INVX1 exu_U13303(.A(exu_n24801), .Y(exu_n2058));
AND2X1 exu_U13304(.A(lsu_exu_dfill_data_g[35]), .B(exu_n16304), .Y(exu_n24805));
INVX1 exu_U13305(.A(exu_n24805), .Y(exu_n2059));
AND2X1 exu_U13306(.A(bypass_mux_rcc_data_2_in1[35]), .B(exu_n16305), .Y(exu_n24807));
INVX1 exu_U13307(.A(exu_n24807), .Y(exu_n2060));
AND2X1 exu_U13308(.A(lsu_exu_dfill_data_g[34]), .B(exu_n16304), .Y(exu_n24811));
INVX1 exu_U13309(.A(exu_n24811), .Y(exu_n2061));
AND2X1 exu_U13310(.A(bypass_mux_rcc_data_2_in1[34]), .B(exu_n16305), .Y(exu_n24813));
INVX1 exu_U13311(.A(exu_n24813), .Y(exu_n2062));
AND2X1 exu_U13312(.A(lsu_exu_dfill_data_g[33]), .B(exu_n16304), .Y(exu_n24817));
INVX1 exu_U13313(.A(exu_n24817), .Y(exu_n2063));
AND2X1 exu_U13314(.A(bypass_mux_rcc_data_2_in1[33]), .B(exu_n16305), .Y(exu_n24819));
INVX1 exu_U13315(.A(exu_n24819), .Y(exu_n2064));
AND2X1 exu_U13316(.A(lsu_exu_dfill_data_g[32]), .B(exu_n16304), .Y(exu_n24823));
INVX1 exu_U13317(.A(exu_n24823), .Y(exu_n2065));
AND2X1 exu_U13318(.A(bypass_mux_rcc_data_2_in1[32]), .B(exu_n16305), .Y(exu_n24825));
INVX1 exu_U13319(.A(exu_n24825), .Y(exu_n2066));
AND2X1 exu_U13320(.A(lsu_exu_dfill_data_g[31]), .B(exu_n16304), .Y(exu_n24829));
INVX1 exu_U13321(.A(exu_n24829), .Y(exu_n2067));
AND2X1 exu_U13322(.A(bypass_mux_rcc_data_2_in1[31]), .B(exu_n16305), .Y(exu_n24831));
INVX1 exu_U13323(.A(exu_n24831), .Y(exu_n2068));
AND2X1 exu_U13324(.A(lsu_exu_dfill_data_g[30]), .B(exu_n16304), .Y(exu_n24835));
INVX1 exu_U13325(.A(exu_n24835), .Y(exu_n2069));
AND2X1 exu_U13326(.A(bypass_mux_rcc_data_2_in1[30]), .B(exu_n16305), .Y(exu_n24837));
INVX1 exu_U13327(.A(exu_n24837), .Y(exu_n2070));
AND2X1 exu_U13328(.A(lsu_exu_dfill_data_g[2]), .B(exu_n16304), .Y(exu_n24841));
INVX1 exu_U13329(.A(exu_n24841), .Y(exu_n2071));
AND2X1 exu_U13330(.A(bypass_mux_rcc_data_2_in1[2]), .B(exu_n16305), .Y(exu_n24843));
INVX1 exu_U13331(.A(exu_n24843), .Y(exu_n2072));
AND2X1 exu_U13332(.A(lsu_exu_dfill_data_g[29]), .B(exu_n16304), .Y(exu_n24847));
INVX1 exu_U13333(.A(exu_n24847), .Y(exu_n2073));
AND2X1 exu_U13334(.A(bypass_mux_rcc_data_2_in1[29]), .B(exu_n16305), .Y(exu_n24849));
INVX1 exu_U13335(.A(exu_n24849), .Y(exu_n2074));
AND2X1 exu_U13336(.A(lsu_exu_dfill_data_g[28]), .B(exu_n16304), .Y(exu_n24853));
INVX1 exu_U13337(.A(exu_n24853), .Y(exu_n2075));
AND2X1 exu_U13338(.A(bypass_mux_rcc_data_2_in1[28]), .B(exu_n16305), .Y(exu_n24855));
INVX1 exu_U13339(.A(exu_n24855), .Y(exu_n2076));
AND2X1 exu_U13340(.A(lsu_exu_dfill_data_g[27]), .B(exu_n16304), .Y(exu_n24859));
INVX1 exu_U13341(.A(exu_n24859), .Y(exu_n2077));
AND2X1 exu_U13342(.A(bypass_mux_rcc_data_2_in1[27]), .B(exu_n16305), .Y(exu_n24861));
INVX1 exu_U13343(.A(exu_n24861), .Y(exu_n2078));
AND2X1 exu_U13344(.A(lsu_exu_dfill_data_g[26]), .B(exu_n16304), .Y(exu_n24865));
INVX1 exu_U13345(.A(exu_n24865), .Y(exu_n2079));
AND2X1 exu_U13346(.A(bypass_mux_rcc_data_2_in1[26]), .B(exu_n16305), .Y(exu_n24867));
INVX1 exu_U13347(.A(exu_n24867), .Y(exu_n2080));
AND2X1 exu_U13348(.A(lsu_exu_dfill_data_g[25]), .B(exu_n16304), .Y(exu_n24871));
INVX1 exu_U13349(.A(exu_n24871), .Y(exu_n2081));
AND2X1 exu_U13350(.A(bypass_mux_rcc_data_2_in1[25]), .B(exu_n16305), .Y(exu_n24873));
INVX1 exu_U13351(.A(exu_n24873), .Y(exu_n2082));
AND2X1 exu_U13352(.A(lsu_exu_dfill_data_g[24]), .B(exu_n16304), .Y(exu_n24877));
INVX1 exu_U13353(.A(exu_n24877), .Y(exu_n2083));
AND2X1 exu_U13354(.A(bypass_mux_rcc_data_2_in1[24]), .B(exu_n16305), .Y(exu_n24879));
INVX1 exu_U13355(.A(exu_n24879), .Y(exu_n2084));
AND2X1 exu_U13356(.A(lsu_exu_dfill_data_g[23]), .B(exu_n16304), .Y(exu_n24883));
INVX1 exu_U13357(.A(exu_n24883), .Y(exu_n2085));
AND2X1 exu_U13358(.A(bypass_mux_rcc_data_2_in1[23]), .B(exu_n16305), .Y(exu_n24885));
INVX1 exu_U13359(.A(exu_n24885), .Y(exu_n2086));
AND2X1 exu_U13360(.A(lsu_exu_dfill_data_g[22]), .B(exu_n16304), .Y(exu_n24889));
INVX1 exu_U13361(.A(exu_n24889), .Y(exu_n2087));
AND2X1 exu_U13362(.A(bypass_mux_rcc_data_2_in1[22]), .B(exu_n16305), .Y(exu_n24891));
INVX1 exu_U13363(.A(exu_n24891), .Y(exu_n2088));
AND2X1 exu_U13364(.A(lsu_exu_dfill_data_g[21]), .B(exu_n16304), .Y(exu_n24895));
INVX1 exu_U13365(.A(exu_n24895), .Y(exu_n2089));
AND2X1 exu_U13366(.A(bypass_mux_rcc_data_2_in1[21]), .B(exu_n16305), .Y(exu_n24897));
INVX1 exu_U13367(.A(exu_n24897), .Y(exu_n2090));
AND2X1 exu_U13368(.A(lsu_exu_dfill_data_g[20]), .B(exu_n16304), .Y(exu_n24901));
INVX1 exu_U13369(.A(exu_n24901), .Y(exu_n2091));
AND2X1 exu_U13370(.A(bypass_mux_rcc_data_2_in1[20]), .B(exu_n16305), .Y(exu_n24903));
INVX1 exu_U13371(.A(exu_n24903), .Y(exu_n2092));
AND2X1 exu_U13372(.A(lsu_exu_dfill_data_g[1]), .B(exu_n16304), .Y(exu_n24907));
INVX1 exu_U13373(.A(exu_n24907), .Y(exu_n2093));
AND2X1 exu_U13374(.A(bypass_mux_rcc_data_2_in1[1]), .B(exu_n16305), .Y(exu_n24909));
INVX1 exu_U13375(.A(exu_n24909), .Y(exu_n2094));
AND2X1 exu_U13376(.A(lsu_exu_dfill_data_g[19]), .B(exu_n16304), .Y(exu_n24913));
INVX1 exu_U13377(.A(exu_n24913), .Y(exu_n2095));
AND2X1 exu_U13378(.A(bypass_mux_rcc_data_2_in1[19]), .B(exu_n16305), .Y(exu_n24915));
INVX1 exu_U13379(.A(exu_n24915), .Y(exu_n2096));
AND2X1 exu_U13380(.A(lsu_exu_dfill_data_g[18]), .B(exu_n16304), .Y(exu_n24919));
INVX1 exu_U13381(.A(exu_n24919), .Y(exu_n2097));
AND2X1 exu_U13382(.A(bypass_mux_rcc_data_2_in1[18]), .B(exu_n16305), .Y(exu_n24921));
INVX1 exu_U13383(.A(exu_n24921), .Y(exu_n2098));
AND2X1 exu_U13384(.A(lsu_exu_dfill_data_g[17]), .B(exu_n16304), .Y(exu_n24925));
INVX1 exu_U13385(.A(exu_n24925), .Y(exu_n2099));
AND2X1 exu_U13386(.A(bypass_mux_rcc_data_2_in1[17]), .B(exu_n16305), .Y(exu_n24927));
INVX1 exu_U13387(.A(exu_n24927), .Y(exu_n2100));
AND2X1 exu_U13388(.A(lsu_exu_dfill_data_g[16]), .B(exu_n16304), .Y(exu_n24931));
INVX1 exu_U13389(.A(exu_n24931), .Y(exu_n2101));
AND2X1 exu_U13390(.A(bypass_mux_rcc_data_2_in1[16]), .B(exu_n16305), .Y(exu_n24933));
INVX1 exu_U13391(.A(exu_n24933), .Y(exu_n2102));
AND2X1 exu_U13392(.A(lsu_exu_dfill_data_g[15]), .B(exu_n16304), .Y(exu_n24937));
INVX1 exu_U13393(.A(exu_n24937), .Y(exu_n2103));
AND2X1 exu_U13394(.A(bypass_mux_rcc_data_2_in1[15]), .B(exu_n16305), .Y(exu_n24939));
INVX1 exu_U13395(.A(exu_n24939), .Y(exu_n2104));
AND2X1 exu_U13396(.A(lsu_exu_dfill_data_g[14]), .B(exu_n16304), .Y(exu_n24943));
INVX1 exu_U13397(.A(exu_n24943), .Y(exu_n2105));
AND2X1 exu_U13398(.A(bypass_mux_rcc_data_2_in1[14]), .B(exu_n16305), .Y(exu_n24945));
INVX1 exu_U13399(.A(exu_n24945), .Y(exu_n2106));
AND2X1 exu_U13400(.A(lsu_exu_dfill_data_g[13]), .B(exu_n16304), .Y(exu_n24949));
INVX1 exu_U13401(.A(exu_n24949), .Y(exu_n2107));
AND2X1 exu_U13402(.A(bypass_mux_rcc_data_2_in1[13]), .B(exu_n16305), .Y(exu_n24951));
INVX1 exu_U13403(.A(exu_n24951), .Y(exu_n2108));
AND2X1 exu_U13404(.A(lsu_exu_dfill_data_g[12]), .B(exu_n16304), .Y(exu_n24955));
INVX1 exu_U13405(.A(exu_n24955), .Y(exu_n2109));
AND2X1 exu_U13406(.A(bypass_mux_rcc_data_2_in1[12]), .B(exu_n16305), .Y(exu_n24957));
INVX1 exu_U13407(.A(exu_n24957), .Y(exu_n2110));
AND2X1 exu_U13408(.A(lsu_exu_dfill_data_g[11]), .B(exu_n16304), .Y(exu_n24961));
INVX1 exu_U13409(.A(exu_n24961), .Y(exu_n2111));
AND2X1 exu_U13410(.A(bypass_mux_rcc_data_2_in1[11]), .B(exu_n16305), .Y(exu_n24963));
INVX1 exu_U13411(.A(exu_n24963), .Y(exu_n2112));
AND2X1 exu_U13412(.A(lsu_exu_dfill_data_g[10]), .B(exu_n16304), .Y(exu_n24967));
INVX1 exu_U13413(.A(exu_n24967), .Y(exu_n2113));
AND2X1 exu_U13414(.A(bypass_mux_rcc_data_2_in1[10]), .B(exu_n16305), .Y(exu_n24969));
INVX1 exu_U13415(.A(exu_n24969), .Y(exu_n2114));
AND2X1 exu_U13416(.A(lsu_exu_dfill_data_g[0]), .B(exu_n16304), .Y(exu_n24973));
INVX1 exu_U13417(.A(exu_n24973), .Y(exu_n2115));
AND2X1 exu_U13418(.A(bypass_mux_rcc_data_2_in1[0]), .B(exu_n16305), .Y(exu_n24975));
INVX1 exu_U13419(.A(exu_n24975), .Y(exu_n2116));
AND2X1 exu_U13420(.A(ecl_byplog_rs2_n14), .B(ifu_exu_imm_data_d[9]), .Y(exu_n24979));
INVX1 exu_U13421(.A(exu_n24979), .Y(exu_n2117));
AND2X1 exu_U13422(.A(exu_n16293), .B(byp_irf_rd_data_w[9]), .Y(exu_n24981));
INVX1 exu_U13423(.A(exu_n24981), .Y(exu_n2118));
AND2X1 exu_U13424(.A(ifu_exu_imm_data_d[8]), .B(ecl_byplog_rs2_n14), .Y(exu_n24985));
INVX1 exu_U13425(.A(exu_n24985), .Y(exu_n2119));
AND2X1 exu_U13426(.A(byp_irf_rd_data_w[8]), .B(exu_n16293), .Y(exu_n24987));
INVX1 exu_U13427(.A(exu_n24987), .Y(exu_n2120));
AND2X1 exu_U13428(.A(ifu_exu_imm_data_d[7]), .B(ecl_byplog_rs2_n14), .Y(exu_n24991));
INVX1 exu_U13429(.A(exu_n24991), .Y(exu_n2121));
AND2X1 exu_U13430(.A(byp_irf_rd_data_w[7]), .B(exu_n16293), .Y(exu_n24993));
INVX1 exu_U13431(.A(exu_n24993), .Y(exu_n2122));
AND2X1 exu_U13432(.A(ifu_exu_imm_data_d[6]), .B(ecl_byplog_rs2_n14), .Y(exu_n24997));
INVX1 exu_U13433(.A(exu_n24997), .Y(exu_n2123));
AND2X1 exu_U13434(.A(byp_irf_rd_data_w[6]), .B(exu_n16293), .Y(exu_n24999));
INVX1 exu_U13435(.A(exu_n24999), .Y(exu_n2124));
AND2X1 exu_U13436(.A(byp_irf_rd_data_w[63]), .B(exu_n16293), .Y(exu_n25004));
INVX1 exu_U13437(.A(exu_n25004), .Y(exu_n2125));
INVX1 exu_U13438(.A(exu_n2130), .Y(exu_n2126));
INVX1 exu_U13439(.A(exu_n2126), .Y(exu_n2127));
AND2X1 exu_U13440(.A(byp_irf_rd_data_w[62]), .B(exu_n16293), .Y(exu_n25009));
INVX1 exu_U13441(.A(exu_n25009), .Y(exu_n2128));
INVX1 exu_U13442(.A(exu_n2133), .Y(exu_n2129));
INVX1 exu_U13443(.A(exu_n2129), .Y(exu_n2130));
AND2X1 exu_U13444(.A(byp_irf_rd_data_w[61]), .B(exu_n16293), .Y(exu_n25014));
INVX1 exu_U13445(.A(exu_n25014), .Y(exu_n2131));
INVX1 exu_U13446(.A(exu_n2138), .Y(exu_n2132));
INVX1 exu_U13447(.A(exu_n2132), .Y(exu_n2133));
AND2X1 exu_U13448(.A(byp_irf_rd_data_w[60]), .B(exu_n16293), .Y(exu_n25019));
INVX1 exu_U13449(.A(exu_n25019), .Y(exu_n2134));
AND2X1 exu_U13450(.A(ifu_exu_imm_data_d[5]), .B(ecl_byplog_rs2_n14), .Y(exu_n25023));
INVX1 exu_U13451(.A(exu_n25023), .Y(exu_n2135));
AND2X1 exu_U13452(.A(byp_irf_rd_data_w[5]), .B(exu_n16293), .Y(exu_n25025));
INVX1 exu_U13453(.A(exu_n25025), .Y(exu_n2136));
INVX1 exu_U13454(.A(exu_n2141), .Y(exu_n2137));
INVX1 exu_U13455(.A(exu_n2137), .Y(exu_n2138));
AND2X1 exu_U13456(.A(byp_irf_rd_data_w[59]), .B(exu_n16293), .Y(exu_n25030));
INVX1 exu_U13457(.A(exu_n25030), .Y(exu_n2139));
INVX1 exu_U13458(.A(exu_n2144), .Y(exu_n2140));
INVX1 exu_U13459(.A(exu_n2140), .Y(exu_n2141));
AND2X1 exu_U13460(.A(byp_irf_rd_data_w[58]), .B(exu_n16293), .Y(exu_n25035));
INVX1 exu_U13461(.A(exu_n25035), .Y(exu_n2142));
INVX1 exu_U13462(.A(exu_n2147), .Y(exu_n2143));
INVX1 exu_U13463(.A(exu_n2143), .Y(exu_n2144));
AND2X1 exu_U13464(.A(byp_irf_rd_data_w[57]), .B(exu_n16293), .Y(exu_n25040));
INVX1 exu_U13465(.A(exu_n25040), .Y(exu_n2145));
INVX1 exu_U13466(.A(exu_n2150), .Y(exu_n2146));
INVX1 exu_U13467(.A(exu_n2146), .Y(exu_n2147));
AND2X1 exu_U13468(.A(byp_irf_rd_data_w[56]), .B(exu_n16293), .Y(exu_n25045));
INVX1 exu_U13469(.A(exu_n25045), .Y(exu_n2148));
INVX1 exu_U13470(.A(exu_n2153), .Y(exu_n2149));
INVX1 exu_U13471(.A(exu_n2149), .Y(exu_n2150));
AND2X1 exu_U13472(.A(byp_irf_rd_data_w[55]), .B(exu_n16293), .Y(exu_n25050));
INVX1 exu_U13473(.A(exu_n25050), .Y(exu_n2151));
INVX1 exu_U13474(.A(exu_n2156), .Y(exu_n2152));
INVX1 exu_U13475(.A(exu_n2152), .Y(exu_n2153));
AND2X1 exu_U13476(.A(byp_irf_rd_data_w[54]), .B(exu_n16293), .Y(exu_n25055));
INVX1 exu_U13477(.A(exu_n25055), .Y(exu_n2154));
INVX1 exu_U13478(.A(exu_n2159), .Y(exu_n2155));
INVX1 exu_U13479(.A(exu_n2155), .Y(exu_n2156));
AND2X1 exu_U13480(.A(byp_irf_rd_data_w[53]), .B(exu_n16293), .Y(exu_n25060));
INVX1 exu_U13481(.A(exu_n25060), .Y(exu_n2157));
INVX1 exu_U13482(.A(exu_n2162), .Y(exu_n2158));
INVX1 exu_U13483(.A(exu_n2158), .Y(exu_n2159));
AND2X1 exu_U13484(.A(byp_irf_rd_data_w[52]), .B(exu_n16293), .Y(exu_n25065));
INVX1 exu_U13485(.A(exu_n25065), .Y(exu_n2160));
INVX1 exu_U13486(.A(exu_n2165), .Y(exu_n2161));
INVX1 exu_U13487(.A(exu_n2161), .Y(exu_n2162));
AND2X1 exu_U13488(.A(byp_irf_rd_data_w[51]), .B(exu_n16293), .Y(exu_n25070));
INVX1 exu_U13489(.A(exu_n25070), .Y(exu_n2163));
INVX1 exu_U13490(.A(exu_n2170), .Y(exu_n2164));
INVX1 exu_U13491(.A(exu_n2164), .Y(exu_n2165));
AND2X1 exu_U13492(.A(byp_irf_rd_data_w[50]), .B(exu_n16293), .Y(exu_n25075));
INVX1 exu_U13493(.A(exu_n25075), .Y(exu_n2166));
AND2X1 exu_U13494(.A(ifu_exu_imm_data_d[4]), .B(ecl_byplog_rs2_n14), .Y(exu_n25079));
INVX1 exu_U13495(.A(exu_n25079), .Y(exu_n2167));
AND2X1 exu_U13496(.A(byp_irf_rd_data_w[4]), .B(exu_n16293), .Y(exu_n25081));
INVX1 exu_U13497(.A(exu_n25081), .Y(exu_n2168));
INVX1 exu_U13498(.A(exu_n2173), .Y(exu_n2169));
INVX1 exu_U13499(.A(exu_n2169), .Y(exu_n2170));
AND2X1 exu_U13500(.A(byp_irf_rd_data_w[49]), .B(exu_n16293), .Y(exu_n25086));
INVX1 exu_U13501(.A(exu_n25086), .Y(exu_n2171));
INVX1 exu_U13502(.A(exu_n2176), .Y(exu_n2172));
INVX1 exu_U13503(.A(exu_n2172), .Y(exu_n2173));
AND2X1 exu_U13504(.A(byp_irf_rd_data_w[48]), .B(exu_n16293), .Y(exu_n25091));
INVX1 exu_U13505(.A(exu_n25091), .Y(exu_n2174));
INVX1 exu_U13506(.A(exu_n2179), .Y(exu_n2175));
INVX1 exu_U13507(.A(exu_n2175), .Y(exu_n2176));
AND2X1 exu_U13508(.A(byp_irf_rd_data_w[47]), .B(exu_n16293), .Y(exu_n25096));
INVX1 exu_U13509(.A(exu_n25096), .Y(exu_n2177));
INVX1 exu_U13510(.A(exu_n2197), .Y(exu_n2178));
INVX1 exu_U13511(.A(exu_n2178), .Y(exu_n2179));
AND2X1 exu_U13512(.A(byp_irf_rd_data_w[46]), .B(exu_n16293), .Y(exu_n25101));
INVX1 exu_U13513(.A(exu_n25101), .Y(exu_n2180));
AND2X1 exu_U13514(.A(byp_irf_rd_data_w[45]), .B(exu_n16293), .Y(exu_n25106));
INVX1 exu_U13515(.A(exu_n25106), .Y(exu_n2181));
AND2X1 exu_U13516(.A(byp_irf_rd_data_w[44]), .B(exu_n16293), .Y(exu_n25111));
INVX1 exu_U13517(.A(exu_n25111), .Y(exu_n2182));
AND2X1 exu_U13518(.A(byp_irf_rd_data_w[43]), .B(exu_n16293), .Y(exu_n25116));
INVX1 exu_U13519(.A(exu_n25116), .Y(exu_n2183));
AND2X1 exu_U13520(.A(byp_irf_rd_data_w[42]), .B(exu_n16293), .Y(exu_n25121));
INVX1 exu_U13521(.A(exu_n25121), .Y(exu_n2184));
AND2X1 exu_U13522(.A(byp_irf_rd_data_w[41]), .B(exu_n16293), .Y(exu_n25126));
INVX1 exu_U13523(.A(exu_n25126), .Y(exu_n2185));
AND2X1 exu_U13524(.A(byp_irf_rd_data_w[40]), .B(exu_n16293), .Y(exu_n25131));
INVX1 exu_U13525(.A(exu_n25131), .Y(exu_n2186));
AND2X1 exu_U13526(.A(ifu_exu_imm_data_d[3]), .B(ecl_byplog_rs2_n14), .Y(exu_n25135));
INVX1 exu_U13527(.A(exu_n25135), .Y(exu_n2187));
AND2X1 exu_U13528(.A(byp_irf_rd_data_w[3]), .B(exu_n16293), .Y(exu_n25137));
INVX1 exu_U13529(.A(exu_n25137), .Y(exu_n2188));
AND2X1 exu_U13530(.A(byp_irf_rd_data_w[39]), .B(exu_n16293), .Y(exu_n25142));
INVX1 exu_U13531(.A(exu_n25142), .Y(exu_n2189));
AND2X1 exu_U13532(.A(byp_irf_rd_data_w[38]), .B(exu_n16293), .Y(exu_n25147));
INVX1 exu_U13533(.A(exu_n25147), .Y(exu_n2190));
AND2X1 exu_U13534(.A(byp_irf_rd_data_w[37]), .B(exu_n16293), .Y(exu_n25152));
INVX1 exu_U13535(.A(exu_n25152), .Y(exu_n2191));
AND2X1 exu_U13536(.A(byp_irf_rd_data_w[36]), .B(exu_n16293), .Y(exu_n25157));
INVX1 exu_U13537(.A(exu_n25157), .Y(exu_n2192));
AND2X1 exu_U13538(.A(byp_irf_rd_data_w[35]), .B(exu_n16293), .Y(exu_n25162));
INVX1 exu_U13539(.A(exu_n25162), .Y(exu_n2193));
AND2X1 exu_U13540(.A(byp_irf_rd_data_w[34]), .B(exu_n16293), .Y(exu_n25167));
INVX1 exu_U13541(.A(exu_n25167), .Y(exu_n2194));
AND2X1 exu_U13542(.A(byp_irf_rd_data_w[33]), .B(exu_n16293), .Y(exu_n25172));
INVX1 exu_U13543(.A(exu_n25172), .Y(exu_n2195));
AND2X1 exu_U13544(.A(byp_irf_rd_data_w[32]), .B(exu_n16293), .Y(exu_n25177));
INVX1 exu_U13545(.A(exu_n25177), .Y(exu_n2196));
AND2X1 exu_U13546(.A(ifu_exu_imm_data_d[31]), .B(exu_n15964), .Y(exu_n25181));
INVX1 exu_U13547(.A(exu_n25181), .Y(exu_n2197));
AND2X1 exu_U13548(.A(byp_irf_rd_data_w[31]), .B(exu_n16293), .Y(exu_n25183));
INVX1 exu_U13549(.A(exu_n25183), .Y(exu_n2198));
AND2X1 exu_U13550(.A(ifu_exu_imm_data_d[30]), .B(exu_n15964), .Y(exu_n25187));
INVX1 exu_U13551(.A(exu_n25187), .Y(exu_n2199));
AND2X1 exu_U13552(.A(byp_irf_rd_data_w[30]), .B(exu_n16293), .Y(exu_n25189));
INVX1 exu_U13553(.A(exu_n25189), .Y(exu_n2200));
AND2X1 exu_U13554(.A(ifu_exu_imm_data_d[2]), .B(exu_n15964), .Y(exu_n25193));
INVX1 exu_U13555(.A(exu_n25193), .Y(exu_n2201));
AND2X1 exu_U13556(.A(byp_irf_rd_data_w[2]), .B(exu_n16293), .Y(exu_n25195));
INVX1 exu_U13557(.A(exu_n25195), .Y(exu_n2202));
AND2X1 exu_U13558(.A(ifu_exu_imm_data_d[29]), .B(exu_n15964), .Y(exu_n25199));
INVX1 exu_U13559(.A(exu_n25199), .Y(exu_n2203));
AND2X1 exu_U13560(.A(byp_irf_rd_data_w[29]), .B(exu_n16293), .Y(exu_n25201));
INVX1 exu_U13561(.A(exu_n25201), .Y(exu_n2204));
AND2X1 exu_U13562(.A(ifu_exu_imm_data_d[28]), .B(exu_n15964), .Y(exu_n25205));
INVX1 exu_U13563(.A(exu_n25205), .Y(exu_n2205));
AND2X1 exu_U13564(.A(byp_irf_rd_data_w[28]), .B(exu_n16293), .Y(exu_n25207));
INVX1 exu_U13565(.A(exu_n25207), .Y(exu_n2206));
AND2X1 exu_U13566(.A(ifu_exu_imm_data_d[27]), .B(exu_n15964), .Y(exu_n25211));
INVX1 exu_U13567(.A(exu_n25211), .Y(exu_n2207));
AND2X1 exu_U13568(.A(byp_irf_rd_data_w[27]), .B(exu_n16293), .Y(exu_n25213));
INVX1 exu_U13569(.A(exu_n25213), .Y(exu_n2208));
AND2X1 exu_U13570(.A(ifu_exu_imm_data_d[26]), .B(exu_n15964), .Y(exu_n25217));
INVX1 exu_U13571(.A(exu_n25217), .Y(exu_n2209));
AND2X1 exu_U13572(.A(byp_irf_rd_data_w[26]), .B(exu_n16293), .Y(exu_n25219));
INVX1 exu_U13573(.A(exu_n25219), .Y(exu_n2210));
AND2X1 exu_U13574(.A(ifu_exu_imm_data_d[25]), .B(exu_n15964), .Y(exu_n25223));
INVX1 exu_U13575(.A(exu_n25223), .Y(exu_n2211));
AND2X1 exu_U13576(.A(byp_irf_rd_data_w[25]), .B(exu_n16293), .Y(exu_n25225));
INVX1 exu_U13577(.A(exu_n25225), .Y(exu_n2212));
AND2X1 exu_U13578(.A(ifu_exu_imm_data_d[24]), .B(exu_n15964), .Y(exu_n25229));
INVX1 exu_U13579(.A(exu_n25229), .Y(exu_n2213));
AND2X1 exu_U13580(.A(byp_irf_rd_data_w[24]), .B(exu_n16293), .Y(exu_n25231));
INVX1 exu_U13581(.A(exu_n25231), .Y(exu_n2214));
AND2X1 exu_U13582(.A(ifu_exu_imm_data_d[23]), .B(exu_n15964), .Y(exu_n25235));
INVX1 exu_U13583(.A(exu_n25235), .Y(exu_n2215));
AND2X1 exu_U13584(.A(byp_irf_rd_data_w[23]), .B(exu_n16293), .Y(exu_n25237));
INVX1 exu_U13585(.A(exu_n25237), .Y(exu_n2216));
AND2X1 exu_U13586(.A(ifu_exu_imm_data_d[22]), .B(exu_n15964), .Y(exu_n25241));
INVX1 exu_U13587(.A(exu_n25241), .Y(exu_n2217));
AND2X1 exu_U13588(.A(byp_irf_rd_data_w[22]), .B(exu_n16293), .Y(exu_n25243));
INVX1 exu_U13589(.A(exu_n25243), .Y(exu_n2218));
AND2X1 exu_U13590(.A(ifu_exu_imm_data_d[21]), .B(exu_n15964), .Y(exu_n25247));
INVX1 exu_U13591(.A(exu_n25247), .Y(exu_n2219));
AND2X1 exu_U13592(.A(byp_irf_rd_data_w[21]), .B(exu_n16293), .Y(exu_n25249));
INVX1 exu_U13593(.A(exu_n25249), .Y(exu_n2220));
AND2X1 exu_U13594(.A(ifu_exu_imm_data_d[20]), .B(exu_n15964), .Y(exu_n25253));
INVX1 exu_U13595(.A(exu_n25253), .Y(exu_n2221));
AND2X1 exu_U13596(.A(byp_irf_rd_data_w[20]), .B(exu_n16293), .Y(exu_n25255));
INVX1 exu_U13597(.A(exu_n25255), .Y(exu_n2222));
AND2X1 exu_U13598(.A(ifu_exu_imm_data_d[1]), .B(ecl_byplog_rs2_n14), .Y(exu_n25259));
INVX1 exu_U13599(.A(exu_n25259), .Y(exu_n2223));
AND2X1 exu_U13600(.A(byp_irf_rd_data_w[1]), .B(exu_n16293), .Y(exu_n25261));
INVX1 exu_U13601(.A(exu_n25261), .Y(exu_n2224));
AND2X1 exu_U13602(.A(ifu_exu_imm_data_d[19]), .B(ecl_byplog_rs2_n14), .Y(exu_n25265));
INVX1 exu_U13603(.A(exu_n25265), .Y(exu_n2225));
AND2X1 exu_U13604(.A(byp_irf_rd_data_w[19]), .B(exu_n16293), .Y(exu_n25267));
INVX1 exu_U13605(.A(exu_n25267), .Y(exu_n2226));
AND2X1 exu_U13606(.A(ifu_exu_imm_data_d[18]), .B(ecl_byplog_rs2_n14), .Y(exu_n25271));
INVX1 exu_U13607(.A(exu_n25271), .Y(exu_n2227));
AND2X1 exu_U13608(.A(byp_irf_rd_data_w[18]), .B(exu_n16293), .Y(exu_n25273));
INVX1 exu_U13609(.A(exu_n25273), .Y(exu_n2228));
AND2X1 exu_U13610(.A(ifu_exu_imm_data_d[17]), .B(ecl_byplog_rs2_n14), .Y(exu_n25277));
INVX1 exu_U13611(.A(exu_n25277), .Y(exu_n2229));
AND2X1 exu_U13612(.A(byp_irf_rd_data_w[17]), .B(exu_n16293), .Y(exu_n25279));
INVX1 exu_U13613(.A(exu_n25279), .Y(exu_n2230));
AND2X1 exu_U13614(.A(ifu_exu_imm_data_d[16]), .B(ecl_byplog_rs2_n14), .Y(exu_n25283));
INVX1 exu_U13615(.A(exu_n25283), .Y(exu_n2231));
AND2X1 exu_U13616(.A(byp_irf_rd_data_w[16]), .B(exu_n16293), .Y(exu_n25285));
INVX1 exu_U13617(.A(exu_n25285), .Y(exu_n2232));
AND2X1 exu_U13618(.A(ifu_exu_imm_data_d[15]), .B(exu_n15964), .Y(exu_n25289));
INVX1 exu_U13619(.A(exu_n25289), .Y(exu_n2233));
AND2X1 exu_U13620(.A(byp_irf_rd_data_w[15]), .B(exu_n16293), .Y(exu_n25291));
INVX1 exu_U13621(.A(exu_n25291), .Y(exu_n2234));
AND2X1 exu_U13622(.A(ifu_exu_imm_data_d[14]), .B(ecl_byplog_rs2_n14), .Y(exu_n25295));
INVX1 exu_U13623(.A(exu_n25295), .Y(exu_n2235));
AND2X1 exu_U13624(.A(byp_irf_rd_data_w[14]), .B(exu_n16293), .Y(exu_n25297));
INVX1 exu_U13625(.A(exu_n25297), .Y(exu_n2236));
AND2X1 exu_U13626(.A(ifu_exu_imm_data_d[13]), .B(exu_n15964), .Y(exu_n25301));
INVX1 exu_U13627(.A(exu_n25301), .Y(exu_n2237));
AND2X1 exu_U13628(.A(byp_irf_rd_data_w[13]), .B(exu_n16293), .Y(exu_n25303));
INVX1 exu_U13629(.A(exu_n25303), .Y(exu_n2238));
AND2X1 exu_U13630(.A(ifu_exu_imm_data_d[12]), .B(ecl_byplog_rs2_n14), .Y(exu_n25307));
INVX1 exu_U13631(.A(exu_n25307), .Y(exu_n2239));
AND2X1 exu_U13632(.A(byp_irf_rd_data_w[12]), .B(exu_n16293), .Y(exu_n25309));
INVX1 exu_U13633(.A(exu_n25309), .Y(exu_n2240));
AND2X1 exu_U13634(.A(ifu_exu_imm_data_d[11]), .B(exu_n15964), .Y(exu_n25313));
INVX1 exu_U13635(.A(exu_n25313), .Y(exu_n2241));
AND2X1 exu_U13636(.A(byp_irf_rd_data_w[11]), .B(exu_n16293), .Y(exu_n25315));
INVX1 exu_U13637(.A(exu_n25315), .Y(exu_n2242));
AND2X1 exu_U13638(.A(ifu_exu_imm_data_d[10]), .B(ecl_byplog_rs2_n14), .Y(exu_n25319));
INVX1 exu_U13639(.A(exu_n25319), .Y(exu_n2243));
AND2X1 exu_U13640(.A(byp_irf_rd_data_w[10]), .B(exu_n16293), .Y(exu_n25321));
INVX1 exu_U13641(.A(exu_n25321), .Y(exu_n2244));
AND2X1 exu_U13642(.A(ifu_exu_imm_data_d[0]), .B(exu_n15964), .Y(exu_n25325));
INVX1 exu_U13643(.A(exu_n25325), .Y(exu_n2245));
AND2X1 exu_U13644(.A(byp_irf_rd_data_w[0]), .B(exu_n16293), .Y(exu_n25327));
INVX1 exu_U13645(.A(exu_n25327), .Y(exu_n2246));
AND2X1 exu_U13646(.A(exu_n16296), .B(lsu_exu_dfill_data_g[9]), .Y(exu_n25331));
INVX1 exu_U13647(.A(exu_n25331), .Y(exu_n2247));
AND2X1 exu_U13648(.A(exu_n16297), .B(bypass_mux_rs2_data_2_in1[9]), .Y(exu_n25333));
INVX1 exu_U13649(.A(exu_n25333), .Y(exu_n2248));
AND2X1 exu_U13650(.A(lsu_exu_dfill_data_g[8]), .B(exu_n16296), .Y(exu_n25337));
INVX1 exu_U13651(.A(exu_n25337), .Y(exu_n2249));
AND2X1 exu_U13652(.A(bypass_mux_rs2_data_2_in1[8]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25339));
INVX1 exu_U13653(.A(exu_n25339), .Y(exu_n2250));
AND2X1 exu_U13654(.A(lsu_exu_dfill_data_g[7]), .B(exu_n16296), .Y(exu_n25343));
INVX1 exu_U13655(.A(exu_n25343), .Y(exu_n2251));
AND2X1 exu_U13656(.A(bypass_mux_rs2_data_2_in1[7]), .B(exu_n16297), .Y(exu_n25345));
INVX1 exu_U13657(.A(exu_n25345), .Y(exu_n2252));
AND2X1 exu_U13658(.A(lsu_exu_dfill_data_g[6]), .B(exu_n16296), .Y(exu_n25349));
INVX1 exu_U13659(.A(exu_n25349), .Y(exu_n2253));
AND2X1 exu_U13660(.A(bypass_mux_rs2_data_2_in1[6]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25351));
INVX1 exu_U13661(.A(exu_n25351), .Y(exu_n2254));
AND2X1 exu_U13662(.A(lsu_exu_dfill_data_g[63]), .B(exu_n16296), .Y(exu_n25355));
INVX1 exu_U13663(.A(exu_n25355), .Y(exu_n2255));
AND2X1 exu_U13664(.A(bypass_mux_rs2_data_2_in1[63]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25357));
INVX1 exu_U13665(.A(exu_n25357), .Y(exu_n2256));
AND2X1 exu_U13666(.A(lsu_exu_dfill_data_g[62]), .B(exu_n16296), .Y(exu_n25361));
INVX1 exu_U13667(.A(exu_n25361), .Y(exu_n2257));
AND2X1 exu_U13668(.A(bypass_mux_rs2_data_2_in1[62]), .B(exu_n16297), .Y(exu_n25363));
INVX1 exu_U13669(.A(exu_n25363), .Y(exu_n2258));
AND2X1 exu_U13670(.A(lsu_exu_dfill_data_g[61]), .B(exu_n16296), .Y(exu_n25367));
INVX1 exu_U13671(.A(exu_n25367), .Y(exu_n2259));
AND2X1 exu_U13672(.A(bypass_mux_rs2_data_2_in1[61]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25369));
INVX1 exu_U13673(.A(exu_n25369), .Y(exu_n2260));
AND2X1 exu_U13674(.A(lsu_exu_dfill_data_g[60]), .B(exu_n16296), .Y(exu_n25373));
INVX1 exu_U13675(.A(exu_n25373), .Y(exu_n2261));
AND2X1 exu_U13676(.A(bypass_mux_rs2_data_2_in1[60]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25375));
INVX1 exu_U13677(.A(exu_n25375), .Y(exu_n2262));
AND2X1 exu_U13678(.A(lsu_exu_dfill_data_g[5]), .B(exu_n16296), .Y(exu_n25379));
INVX1 exu_U13679(.A(exu_n25379), .Y(exu_n2263));
AND2X1 exu_U13680(.A(bypass_mux_rs2_data_2_in1[5]), .B(exu_n16297), .Y(exu_n25381));
INVX1 exu_U13681(.A(exu_n25381), .Y(exu_n2264));
AND2X1 exu_U13682(.A(lsu_exu_dfill_data_g[59]), .B(exu_n16296), .Y(exu_n25385));
INVX1 exu_U13683(.A(exu_n25385), .Y(exu_n2265));
AND2X1 exu_U13684(.A(bypass_mux_rs2_data_2_in1[59]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25387));
INVX1 exu_U13685(.A(exu_n25387), .Y(exu_n2266));
AND2X1 exu_U13686(.A(lsu_exu_dfill_data_g[58]), .B(exu_n16296), .Y(exu_n25391));
INVX1 exu_U13687(.A(exu_n25391), .Y(exu_n2267));
AND2X1 exu_U13688(.A(bypass_mux_rs2_data_2_in1[58]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25393));
INVX1 exu_U13689(.A(exu_n25393), .Y(exu_n2268));
AND2X1 exu_U13690(.A(lsu_exu_dfill_data_g[57]), .B(exu_n16296), .Y(exu_n25397));
INVX1 exu_U13691(.A(exu_n25397), .Y(exu_n2269));
AND2X1 exu_U13692(.A(bypass_mux_rs2_data_2_in1[57]), .B(exu_n16297), .Y(exu_n25399));
INVX1 exu_U13693(.A(exu_n25399), .Y(exu_n2270));
AND2X1 exu_U13694(.A(lsu_exu_dfill_data_g[56]), .B(exu_n16296), .Y(exu_n25403));
INVX1 exu_U13695(.A(exu_n25403), .Y(exu_n2271));
AND2X1 exu_U13696(.A(bypass_mux_rs2_data_2_in1[56]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25405));
INVX1 exu_U13697(.A(exu_n25405), .Y(exu_n2272));
AND2X1 exu_U13698(.A(lsu_exu_dfill_data_g[55]), .B(exu_n16296), .Y(exu_n25409));
INVX1 exu_U13699(.A(exu_n25409), .Y(exu_n2273));
AND2X1 exu_U13700(.A(bypass_mux_rs2_data_2_in1[55]), .B(exu_n16297), .Y(exu_n25411));
INVX1 exu_U13701(.A(exu_n25411), .Y(exu_n2274));
AND2X1 exu_U13702(.A(lsu_exu_dfill_data_g[54]), .B(exu_n16296), .Y(exu_n25415));
INVX1 exu_U13703(.A(exu_n25415), .Y(exu_n2275));
AND2X1 exu_U13704(.A(bypass_mux_rs2_data_2_in1[54]), .B(exu_n16297), .Y(exu_n25417));
INVX1 exu_U13705(.A(exu_n25417), .Y(exu_n2276));
AND2X1 exu_U13706(.A(lsu_exu_dfill_data_g[53]), .B(exu_n16296), .Y(exu_n25421));
INVX1 exu_U13707(.A(exu_n25421), .Y(exu_n2277));
AND2X1 exu_U13708(.A(bypass_mux_rs2_data_2_in1[53]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25423));
INVX1 exu_U13709(.A(exu_n25423), .Y(exu_n2278));
AND2X1 exu_U13710(.A(lsu_exu_dfill_data_g[52]), .B(exu_n16296), .Y(exu_n25427));
INVX1 exu_U13711(.A(exu_n25427), .Y(exu_n2279));
AND2X1 exu_U13712(.A(bypass_mux_rs2_data_2_in1[52]), .B(exu_n16297), .Y(exu_n25429));
INVX1 exu_U13713(.A(exu_n25429), .Y(exu_n2280));
AND2X1 exu_U13714(.A(lsu_exu_dfill_data_g[51]), .B(exu_n16296), .Y(exu_n25433));
INVX1 exu_U13715(.A(exu_n25433), .Y(exu_n2281));
AND2X1 exu_U13716(.A(bypass_mux_rs2_data_2_in1[51]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25435));
INVX1 exu_U13717(.A(exu_n25435), .Y(exu_n2282));
AND2X1 exu_U13718(.A(lsu_exu_dfill_data_g[50]), .B(exu_n16296), .Y(exu_n25439));
INVX1 exu_U13719(.A(exu_n25439), .Y(exu_n2283));
AND2X1 exu_U13720(.A(bypass_mux_rs2_data_2_in1[50]), .B(exu_n16297), .Y(exu_n25441));
INVX1 exu_U13721(.A(exu_n25441), .Y(exu_n2284));
AND2X1 exu_U13722(.A(lsu_exu_dfill_data_g[4]), .B(exu_n16296), .Y(exu_n25445));
INVX1 exu_U13723(.A(exu_n25445), .Y(exu_n2285));
AND2X1 exu_U13724(.A(bypass_mux_rs2_data_2_in1[4]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25447));
INVX1 exu_U13725(.A(exu_n25447), .Y(exu_n2286));
AND2X1 exu_U13726(.A(lsu_exu_dfill_data_g[49]), .B(exu_n16296), .Y(exu_n25451));
INVX1 exu_U13727(.A(exu_n25451), .Y(exu_n2287));
AND2X1 exu_U13728(.A(bypass_mux_rs2_data_2_in1[49]), .B(exu_n16297), .Y(exu_n25453));
INVX1 exu_U13729(.A(exu_n25453), .Y(exu_n2288));
AND2X1 exu_U13730(.A(lsu_exu_dfill_data_g[48]), .B(exu_n16296), .Y(exu_n25457));
INVX1 exu_U13731(.A(exu_n25457), .Y(exu_n2289));
AND2X1 exu_U13732(.A(bypass_mux_rs2_data_2_in1[48]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25459));
INVX1 exu_U13733(.A(exu_n25459), .Y(exu_n2290));
AND2X1 exu_U13734(.A(lsu_exu_dfill_data_g[47]), .B(exu_n16296), .Y(exu_n25463));
INVX1 exu_U13735(.A(exu_n25463), .Y(exu_n2291));
AND2X1 exu_U13736(.A(bypass_mux_rs2_data_2_in1[47]), .B(exu_n16297), .Y(exu_n25465));
INVX1 exu_U13737(.A(exu_n25465), .Y(exu_n2292));
AND2X1 exu_U13738(.A(lsu_exu_dfill_data_g[46]), .B(exu_n16296), .Y(exu_n25469));
INVX1 exu_U13739(.A(exu_n25469), .Y(exu_n2293));
AND2X1 exu_U13740(.A(bypass_mux_rs2_data_2_in1[46]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25471));
INVX1 exu_U13741(.A(exu_n25471), .Y(exu_n2294));
AND2X1 exu_U13742(.A(lsu_exu_dfill_data_g[45]), .B(exu_n16296), .Y(exu_n25475));
INVX1 exu_U13743(.A(exu_n25475), .Y(exu_n2295));
AND2X1 exu_U13744(.A(bypass_mux_rs2_data_2_in1[45]), .B(exu_n16297), .Y(exu_n25477));
INVX1 exu_U13745(.A(exu_n25477), .Y(exu_n2296));
AND2X1 exu_U13746(.A(lsu_exu_dfill_data_g[44]), .B(exu_n16296), .Y(exu_n25481));
INVX1 exu_U13747(.A(exu_n25481), .Y(exu_n2297));
AND2X1 exu_U13748(.A(bypass_mux_rs2_data_2_in1[44]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25483));
INVX1 exu_U13749(.A(exu_n25483), .Y(exu_n2298));
AND2X1 exu_U13750(.A(lsu_exu_dfill_data_g[43]), .B(exu_n16296), .Y(exu_n25487));
INVX1 exu_U13751(.A(exu_n25487), .Y(exu_n2299));
AND2X1 exu_U13752(.A(bypass_mux_rs2_data_2_in1[43]), .B(exu_n16297), .Y(exu_n25489));
INVX1 exu_U13753(.A(exu_n25489), .Y(exu_n2300));
AND2X1 exu_U13754(.A(lsu_exu_dfill_data_g[42]), .B(exu_n16296), .Y(exu_n25493));
INVX1 exu_U13755(.A(exu_n25493), .Y(exu_n2301));
AND2X1 exu_U13756(.A(bypass_mux_rs2_data_2_in1[42]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25495));
INVX1 exu_U13757(.A(exu_n25495), .Y(exu_n2302));
AND2X1 exu_U13758(.A(lsu_exu_dfill_data_g[41]), .B(exu_n16296), .Y(exu_n25499));
INVX1 exu_U13759(.A(exu_n25499), .Y(exu_n2303));
AND2X1 exu_U13760(.A(bypass_mux_rs2_data_2_in1[41]), .B(exu_n16297), .Y(exu_n25501));
INVX1 exu_U13761(.A(exu_n25501), .Y(exu_n2304));
AND2X1 exu_U13762(.A(lsu_exu_dfill_data_g[40]), .B(exu_n16296), .Y(exu_n25505));
INVX1 exu_U13763(.A(exu_n25505), .Y(exu_n2305));
AND2X1 exu_U13764(.A(bypass_mux_rs2_data_2_in1[40]), .B(exu_n16297), .Y(exu_n25507));
INVX1 exu_U13765(.A(exu_n25507), .Y(exu_n2306));
AND2X1 exu_U13766(.A(lsu_exu_dfill_data_g[3]), .B(exu_n16296), .Y(exu_n25511));
INVX1 exu_U13767(.A(exu_n25511), .Y(exu_n2307));
AND2X1 exu_U13768(.A(bypass_mux_rs2_data_2_in1[3]), .B(exu_n16297), .Y(exu_n25513));
INVX1 exu_U13769(.A(exu_n25513), .Y(exu_n2308));
AND2X1 exu_U13770(.A(lsu_exu_dfill_data_g[39]), .B(exu_n16296), .Y(exu_n25517));
INVX1 exu_U13771(.A(exu_n25517), .Y(exu_n2309));
AND2X1 exu_U13772(.A(bypass_mux_rs2_data_2_in1[39]), .B(exu_n16297), .Y(exu_n25519));
INVX1 exu_U13773(.A(exu_n25519), .Y(exu_n2310));
AND2X1 exu_U13774(.A(lsu_exu_dfill_data_g[38]), .B(exu_n16296), .Y(exu_n25523));
INVX1 exu_U13775(.A(exu_n25523), .Y(exu_n2311));
AND2X1 exu_U13776(.A(bypass_mux_rs2_data_2_in1[38]), .B(exu_n16297), .Y(exu_n25525));
INVX1 exu_U13777(.A(exu_n25525), .Y(exu_n2312));
AND2X1 exu_U13778(.A(lsu_exu_dfill_data_g[37]), .B(exu_n16296), .Y(exu_n25529));
INVX1 exu_U13779(.A(exu_n25529), .Y(exu_n2313));
AND2X1 exu_U13780(.A(bypass_mux_rs2_data_2_in1[37]), .B(exu_n16297), .Y(exu_n25531));
INVX1 exu_U13781(.A(exu_n25531), .Y(exu_n2314));
AND2X1 exu_U13782(.A(lsu_exu_dfill_data_g[36]), .B(exu_n16296), .Y(exu_n25535));
INVX1 exu_U13783(.A(exu_n25535), .Y(exu_n2315));
AND2X1 exu_U13784(.A(bypass_mux_rs2_data_2_in1[36]), .B(exu_n16297), .Y(exu_n25537));
INVX1 exu_U13785(.A(exu_n25537), .Y(exu_n2316));
AND2X1 exu_U13786(.A(lsu_exu_dfill_data_g[35]), .B(exu_n16296), .Y(exu_n25541));
INVX1 exu_U13787(.A(exu_n25541), .Y(exu_n2317));
AND2X1 exu_U13788(.A(bypass_mux_rs2_data_2_in1[35]), .B(exu_n16297), .Y(exu_n25543));
INVX1 exu_U13789(.A(exu_n25543), .Y(exu_n2318));
AND2X1 exu_U13790(.A(lsu_exu_dfill_data_g[34]), .B(exu_n16296), .Y(exu_n25547));
INVX1 exu_U13791(.A(exu_n25547), .Y(exu_n2319));
AND2X1 exu_U13792(.A(bypass_mux_rs2_data_2_in1[34]), .B(exu_n16297), .Y(exu_n25549));
INVX1 exu_U13793(.A(exu_n25549), .Y(exu_n2320));
AND2X1 exu_U13794(.A(lsu_exu_dfill_data_g[33]), .B(exu_n16296), .Y(exu_n25553));
INVX1 exu_U13795(.A(exu_n25553), .Y(exu_n2321));
AND2X1 exu_U13796(.A(bypass_mux_rs2_data_2_in1[33]), .B(exu_n16297), .Y(exu_n25555));
INVX1 exu_U13797(.A(exu_n25555), .Y(exu_n2322));
AND2X1 exu_U13798(.A(lsu_exu_dfill_data_g[32]), .B(exu_n16296), .Y(exu_n25559));
INVX1 exu_U13799(.A(exu_n25559), .Y(exu_n2323));
AND2X1 exu_U13800(.A(bypass_mux_rs2_data_2_in1[32]), .B(exu_n16297), .Y(exu_n25561));
INVX1 exu_U13801(.A(exu_n25561), .Y(exu_n2324));
AND2X1 exu_U13802(.A(lsu_exu_dfill_data_g[31]), .B(exu_n16296), .Y(exu_n25565));
INVX1 exu_U13803(.A(exu_n25565), .Y(exu_n2325));
AND2X1 exu_U13804(.A(bypass_mux_rs2_data_2_in1[31]), .B(exu_n16297), .Y(exu_n25567));
INVX1 exu_U13805(.A(exu_n25567), .Y(exu_n2326));
AND2X1 exu_U13806(.A(lsu_exu_dfill_data_g[30]), .B(exu_n16296), .Y(exu_n25571));
INVX1 exu_U13807(.A(exu_n25571), .Y(exu_n2327));
AND2X1 exu_U13808(.A(bypass_mux_rs2_data_2_in1[30]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25573));
INVX1 exu_U13809(.A(exu_n25573), .Y(exu_n2328));
AND2X1 exu_U13810(.A(lsu_exu_dfill_data_g[2]), .B(exu_n16296), .Y(exu_n25577));
INVX1 exu_U13811(.A(exu_n25577), .Y(exu_n2329));
AND2X1 exu_U13812(.A(bypass_mux_rs2_data_2_in1[2]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25579));
INVX1 exu_U13813(.A(exu_n25579), .Y(exu_n2330));
AND2X1 exu_U13814(.A(lsu_exu_dfill_data_g[29]), .B(exu_n16296), .Y(exu_n25583));
INVX1 exu_U13815(.A(exu_n25583), .Y(exu_n2331));
AND2X1 exu_U13816(.A(bypass_mux_rs2_data_2_in1[29]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25585));
INVX1 exu_U13817(.A(exu_n25585), .Y(exu_n2332));
AND2X1 exu_U13818(.A(lsu_exu_dfill_data_g[28]), .B(exu_n16296), .Y(exu_n25589));
INVX1 exu_U13819(.A(exu_n25589), .Y(exu_n2333));
AND2X1 exu_U13820(.A(bypass_mux_rs2_data_2_in1[28]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25591));
INVX1 exu_U13821(.A(exu_n25591), .Y(exu_n2334));
AND2X1 exu_U13822(.A(lsu_exu_dfill_data_g[27]), .B(exu_n16296), .Y(exu_n25595));
INVX1 exu_U13823(.A(exu_n25595), .Y(exu_n2335));
AND2X1 exu_U13824(.A(bypass_mux_rs2_data_2_in1[27]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25597));
INVX1 exu_U13825(.A(exu_n25597), .Y(exu_n2336));
AND2X1 exu_U13826(.A(lsu_exu_dfill_data_g[26]), .B(exu_n16296), .Y(exu_n25601));
INVX1 exu_U13827(.A(exu_n25601), .Y(exu_n2337));
AND2X1 exu_U13828(.A(bypass_mux_rs2_data_2_in1[26]), .B(exu_n16297), .Y(exu_n25603));
INVX1 exu_U13829(.A(exu_n25603), .Y(exu_n2338));
AND2X1 exu_U13830(.A(lsu_exu_dfill_data_g[25]), .B(exu_n16296), .Y(exu_n25607));
INVX1 exu_U13831(.A(exu_n25607), .Y(exu_n2339));
AND2X1 exu_U13832(.A(bypass_mux_rs2_data_2_in1[25]), .B(exu_n16297), .Y(exu_n25609));
INVX1 exu_U13833(.A(exu_n25609), .Y(exu_n2340));
AND2X1 exu_U13834(.A(lsu_exu_dfill_data_g[24]), .B(exu_n16296), .Y(exu_n25613));
INVX1 exu_U13835(.A(exu_n25613), .Y(exu_n2341));
AND2X1 exu_U13836(.A(bypass_mux_rs2_data_2_in1[24]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25615));
INVX1 exu_U13837(.A(exu_n25615), .Y(exu_n2342));
AND2X1 exu_U13838(.A(lsu_exu_dfill_data_g[23]), .B(exu_n16296), .Y(exu_n25619));
INVX1 exu_U13839(.A(exu_n25619), .Y(exu_n2343));
AND2X1 exu_U13840(.A(bypass_mux_rs2_data_2_in1[23]), .B(exu_n16297), .Y(exu_n25621));
INVX1 exu_U13841(.A(exu_n25621), .Y(exu_n2344));
AND2X1 exu_U13842(.A(lsu_exu_dfill_data_g[22]), .B(exu_n16296), .Y(exu_n25625));
INVX1 exu_U13843(.A(exu_n25625), .Y(exu_n2345));
AND2X1 exu_U13844(.A(bypass_mux_rs2_data_2_in1[22]), .B(exu_n16297), .Y(exu_n25627));
INVX1 exu_U13845(.A(exu_n25627), .Y(exu_n2346));
AND2X1 exu_U13846(.A(lsu_exu_dfill_data_g[21]), .B(exu_n16296), .Y(exu_n25631));
INVX1 exu_U13847(.A(exu_n25631), .Y(exu_n2347));
AND2X1 exu_U13848(.A(bypass_mux_rs2_data_2_in1[21]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25633));
INVX1 exu_U13849(.A(exu_n25633), .Y(exu_n2348));
AND2X1 exu_U13850(.A(lsu_exu_dfill_data_g[20]), .B(exu_n16296), .Y(exu_n25637));
INVX1 exu_U13851(.A(exu_n25637), .Y(exu_n2349));
AND2X1 exu_U13852(.A(bypass_mux_rs2_data_2_in1[20]), .B(exu_n16297), .Y(exu_n25639));
INVX1 exu_U13853(.A(exu_n25639), .Y(exu_n2350));
AND2X1 exu_U13854(.A(lsu_exu_dfill_data_g[1]), .B(exu_n16296), .Y(exu_n25643));
INVX1 exu_U13855(.A(exu_n25643), .Y(exu_n2351));
AND2X1 exu_U13856(.A(bypass_mux_rs2_data_2_in1[1]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25645));
INVX1 exu_U13857(.A(exu_n25645), .Y(exu_n2352));
AND2X1 exu_U13858(.A(lsu_exu_dfill_data_g[19]), .B(exu_n16296), .Y(exu_n25649));
INVX1 exu_U13859(.A(exu_n25649), .Y(exu_n2353));
AND2X1 exu_U13860(.A(bypass_mux_rs2_data_2_in1[19]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25651));
INVX1 exu_U13861(.A(exu_n25651), .Y(exu_n2354));
AND2X1 exu_U13862(.A(lsu_exu_dfill_data_g[18]), .B(exu_n16296), .Y(exu_n25655));
INVX1 exu_U13863(.A(exu_n25655), .Y(exu_n2355));
AND2X1 exu_U13864(.A(bypass_mux_rs2_data_2_in1[18]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25657));
INVX1 exu_U13865(.A(exu_n25657), .Y(exu_n2356));
AND2X1 exu_U13866(.A(lsu_exu_dfill_data_g[17]), .B(exu_n16296), .Y(exu_n25661));
INVX1 exu_U13867(.A(exu_n25661), .Y(exu_n2357));
AND2X1 exu_U13868(.A(bypass_mux_rs2_data_2_in1[17]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25663));
INVX1 exu_U13869(.A(exu_n25663), .Y(exu_n2358));
AND2X1 exu_U13870(.A(lsu_exu_dfill_data_g[16]), .B(exu_n16296), .Y(exu_n25667));
INVX1 exu_U13871(.A(exu_n25667), .Y(exu_n2359));
AND2X1 exu_U13872(.A(bypass_mux_rs2_data_2_in1[16]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25669));
INVX1 exu_U13873(.A(exu_n25669), .Y(exu_n2360));
AND2X1 exu_U13874(.A(lsu_exu_dfill_data_g[15]), .B(exu_n16296), .Y(exu_n25673));
INVX1 exu_U13875(.A(exu_n25673), .Y(exu_n2361));
AND2X1 exu_U13876(.A(bypass_mux_rs2_data_2_in1[15]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25675));
INVX1 exu_U13877(.A(exu_n25675), .Y(exu_n2362));
AND2X1 exu_U13878(.A(lsu_exu_dfill_data_g[14]), .B(exu_n16296), .Y(exu_n25679));
INVX1 exu_U13879(.A(exu_n25679), .Y(exu_n2363));
AND2X1 exu_U13880(.A(bypass_mux_rs2_data_2_in1[14]), .B(exu_n16297), .Y(exu_n25681));
INVX1 exu_U13881(.A(exu_n25681), .Y(exu_n2364));
AND2X1 exu_U13882(.A(lsu_exu_dfill_data_g[13]), .B(exu_n16296), .Y(exu_n25685));
INVX1 exu_U13883(.A(exu_n25685), .Y(exu_n2365));
AND2X1 exu_U13884(.A(bypass_mux_rs2_data_2_in1[13]), .B(exu_n16297), .Y(exu_n25687));
INVX1 exu_U13885(.A(exu_n25687), .Y(exu_n2366));
AND2X1 exu_U13886(.A(lsu_exu_dfill_data_g[12]), .B(exu_n16296), .Y(exu_n25691));
INVX1 exu_U13887(.A(exu_n25691), .Y(exu_n2367));
AND2X1 exu_U13888(.A(bypass_mux_rs2_data_2_in1[12]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25693));
INVX1 exu_U13889(.A(exu_n25693), .Y(exu_n2368));
AND2X1 exu_U13890(.A(lsu_exu_dfill_data_g[11]), .B(exu_n16296), .Y(exu_n25697));
INVX1 exu_U13891(.A(exu_n25697), .Y(exu_n2369));
AND2X1 exu_U13892(.A(bypass_mux_rs2_data_2_in1[11]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25699));
INVX1 exu_U13893(.A(exu_n25699), .Y(exu_n2370));
AND2X1 exu_U13894(.A(lsu_exu_dfill_data_g[10]), .B(exu_n16296), .Y(exu_n25703));
INVX1 exu_U13895(.A(exu_n25703), .Y(exu_n2371));
AND2X1 exu_U13896(.A(bypass_mux_rs2_data_2_in1[10]), .B(ecl_byp_rs2_mux2_sel_rf), .Y(exu_n25705));
INVX1 exu_U13897(.A(exu_n25705), .Y(exu_n2372));
AND2X1 exu_U13898(.A(lsu_exu_dfill_data_g[0]), .B(exu_n16296), .Y(exu_n25709));
INVX1 exu_U13899(.A(exu_n25709), .Y(exu_n2373));
AND2X1 exu_U13900(.A(bypass_mux_rs2_data_2_in1[0]), .B(exu_n16297), .Y(exu_n25711));
INVX1 exu_U13901(.A(exu_n25711), .Y(exu_n2374));
AND2X1 exu_U13902(.A(exu_n16289), .B(byp_irf_rd_data_w[9]), .Y(exu_n25715));
INVX1 exu_U13903(.A(exu_n25715), .Y(exu_n2375));
AND2X1 exu_U13904(.A(byp_irf_rd_data_w[8]), .B(exu_n16289), .Y(exu_n25719));
INVX1 exu_U13905(.A(exu_n25719), .Y(exu_n2376));
AND2X1 exu_U13906(.A(byp_irf_rd_data_w[7]), .B(exu_n16289), .Y(exu_n25723));
INVX1 exu_U13907(.A(exu_n25723), .Y(exu_n2377));
AND2X1 exu_U13908(.A(byp_irf_rd_data_w[6]), .B(exu_n16289), .Y(exu_n25727));
INVX1 exu_U13909(.A(exu_n25727), .Y(exu_n2378));
AND2X1 exu_U13910(.A(byp_irf_rd_data_w[63]), .B(exu_n16289), .Y(exu_n25731));
INVX1 exu_U13911(.A(exu_n25731), .Y(exu_n2379));
AND2X1 exu_U13912(.A(byp_irf_rd_data_w[62]), .B(exu_n16289), .Y(exu_n25735));
INVX1 exu_U13913(.A(exu_n25735), .Y(exu_n2380));
AND2X1 exu_U13914(.A(byp_irf_rd_data_w[61]), .B(exu_n16289), .Y(exu_n25739));
INVX1 exu_U13915(.A(exu_n25739), .Y(exu_n2381));
AND2X1 exu_U13916(.A(byp_irf_rd_data_w[60]), .B(exu_n16289), .Y(exu_n25743));
INVX1 exu_U13917(.A(exu_n25743), .Y(exu_n2382));
AND2X1 exu_U13918(.A(byp_irf_rd_data_w[5]), .B(exu_n16289), .Y(exu_n25747));
INVX1 exu_U13919(.A(exu_n25747), .Y(exu_n2383));
AND2X1 exu_U13920(.A(byp_irf_rd_data_w[59]), .B(exu_n16289), .Y(exu_n25751));
INVX1 exu_U13921(.A(exu_n25751), .Y(exu_n2384));
AND2X1 exu_U13922(.A(byp_irf_rd_data_w[58]), .B(exu_n16289), .Y(exu_n25755));
INVX1 exu_U13923(.A(exu_n25755), .Y(exu_n2385));
AND2X1 exu_U13924(.A(byp_irf_rd_data_w[57]), .B(exu_n16289), .Y(exu_n25759));
INVX1 exu_U13925(.A(exu_n25759), .Y(exu_n2386));
AND2X1 exu_U13926(.A(byp_irf_rd_data_w[56]), .B(exu_n16289), .Y(exu_n25763));
INVX1 exu_U13927(.A(exu_n25763), .Y(exu_n2387));
AND2X1 exu_U13928(.A(byp_irf_rd_data_w[55]), .B(exu_n16289), .Y(exu_n25767));
INVX1 exu_U13929(.A(exu_n25767), .Y(exu_n2388));
AND2X1 exu_U13930(.A(byp_irf_rd_data_w[54]), .B(exu_n16289), .Y(exu_n25771));
INVX1 exu_U13931(.A(exu_n25771), .Y(exu_n2389));
AND2X1 exu_U13932(.A(byp_irf_rd_data_w[53]), .B(exu_n16289), .Y(exu_n25775));
INVX1 exu_U13933(.A(exu_n25775), .Y(exu_n2390));
AND2X1 exu_U13934(.A(byp_irf_rd_data_w[52]), .B(exu_n16289), .Y(exu_n25779));
INVX1 exu_U13935(.A(exu_n25779), .Y(exu_n2391));
AND2X1 exu_U13936(.A(byp_irf_rd_data_w[51]), .B(exu_n16289), .Y(exu_n25783));
INVX1 exu_U13937(.A(exu_n25783), .Y(exu_n2392));
AND2X1 exu_U13938(.A(byp_irf_rd_data_w[50]), .B(exu_n16289), .Y(exu_n25787));
INVX1 exu_U13939(.A(exu_n25787), .Y(exu_n2393));
AND2X1 exu_U13940(.A(byp_irf_rd_data_w[4]), .B(exu_n16289), .Y(exu_n25791));
INVX1 exu_U13941(.A(exu_n25791), .Y(exu_n2394));
AND2X1 exu_U13942(.A(byp_irf_rd_data_w[49]), .B(exu_n16289), .Y(exu_n25795));
INVX1 exu_U13943(.A(exu_n25795), .Y(exu_n2395));
AND2X1 exu_U13944(.A(byp_irf_rd_data_w[48]), .B(exu_n16289), .Y(exu_n25799));
INVX1 exu_U13945(.A(exu_n25799), .Y(exu_n2396));
AND2X1 exu_U13946(.A(byp_irf_rd_data_w[47]), .B(exu_n16289), .Y(exu_n25803));
INVX1 exu_U13947(.A(exu_n25803), .Y(exu_n2397));
AND2X1 exu_U13948(.A(byp_irf_rd_data_w[46]), .B(exu_n16289), .Y(exu_n25807));
INVX1 exu_U13949(.A(exu_n25807), .Y(exu_n2398));
AND2X1 exu_U13950(.A(byp_irf_rd_data_w[45]), .B(exu_n16289), .Y(exu_n25811));
INVX1 exu_U13951(.A(exu_n25811), .Y(exu_n2399));
AND2X1 exu_U13952(.A(byp_irf_rd_data_w[44]), .B(exu_n16289), .Y(exu_n25815));
INVX1 exu_U13953(.A(exu_n25815), .Y(exu_n2400));
AND2X1 exu_U13954(.A(byp_irf_rd_data_w[43]), .B(exu_n16289), .Y(exu_n25819));
INVX1 exu_U13955(.A(exu_n25819), .Y(exu_n2401));
AND2X1 exu_U13956(.A(byp_irf_rd_data_w[42]), .B(exu_n16289), .Y(exu_n25823));
INVX1 exu_U13957(.A(exu_n25823), .Y(exu_n2402));
AND2X1 exu_U13958(.A(byp_irf_rd_data_w[41]), .B(exu_n16289), .Y(exu_n25827));
INVX1 exu_U13959(.A(exu_n25827), .Y(exu_n2403));
AND2X1 exu_U13960(.A(byp_irf_rd_data_w[40]), .B(exu_n16289), .Y(exu_n25831));
INVX1 exu_U13961(.A(exu_n25831), .Y(exu_n2404));
AND2X1 exu_U13962(.A(byp_irf_rd_data_w[3]), .B(exu_n16289), .Y(exu_n25835));
INVX1 exu_U13963(.A(exu_n25835), .Y(exu_n2405));
AND2X1 exu_U13964(.A(byp_irf_rd_data_w[39]), .B(exu_n16289), .Y(exu_n25839));
INVX1 exu_U13965(.A(exu_n25839), .Y(exu_n2406));
AND2X1 exu_U13966(.A(byp_irf_rd_data_w[38]), .B(exu_n16289), .Y(exu_n25843));
INVX1 exu_U13967(.A(exu_n25843), .Y(exu_n2407));
AND2X1 exu_U13968(.A(byp_irf_rd_data_w[37]), .B(exu_n16289), .Y(exu_n25847));
INVX1 exu_U13969(.A(exu_n25847), .Y(exu_n2408));
AND2X1 exu_U13970(.A(byp_irf_rd_data_w[36]), .B(exu_n16289), .Y(exu_n25851));
INVX1 exu_U13971(.A(exu_n25851), .Y(exu_n2409));
AND2X1 exu_U13972(.A(byp_irf_rd_data_w[35]), .B(exu_n16289), .Y(exu_n25855));
INVX1 exu_U13973(.A(exu_n25855), .Y(exu_n2410));
AND2X1 exu_U13974(.A(byp_irf_rd_data_w[34]), .B(exu_n16289), .Y(exu_n25859));
INVX1 exu_U13975(.A(exu_n25859), .Y(exu_n2411));
AND2X1 exu_U13976(.A(byp_irf_rd_data_w[33]), .B(exu_n16289), .Y(exu_n25863));
INVX1 exu_U13977(.A(exu_n25863), .Y(exu_n2412));
AND2X1 exu_U13978(.A(byp_irf_rd_data_w[32]), .B(exu_n16289), .Y(exu_n25867));
INVX1 exu_U13979(.A(exu_n25867), .Y(exu_n2413));
AND2X1 exu_U13980(.A(byp_irf_rd_data_w[31]), .B(exu_n16289), .Y(exu_n25871));
INVX1 exu_U13981(.A(exu_n25871), .Y(exu_n2414));
AND2X1 exu_U13982(.A(byp_irf_rd_data_w[30]), .B(exu_n16289), .Y(exu_n25875));
INVX1 exu_U13983(.A(exu_n25875), .Y(exu_n2415));
AND2X1 exu_U13984(.A(byp_irf_rd_data_w[2]), .B(exu_n16289), .Y(exu_n25879));
INVX1 exu_U13985(.A(exu_n25879), .Y(exu_n2416));
AND2X1 exu_U13986(.A(byp_irf_rd_data_w[29]), .B(exu_n16289), .Y(exu_n25883));
INVX1 exu_U13987(.A(exu_n25883), .Y(exu_n2417));
AND2X1 exu_U13988(.A(byp_irf_rd_data_w[28]), .B(exu_n16289), .Y(exu_n25887));
INVX1 exu_U13989(.A(exu_n25887), .Y(exu_n2418));
AND2X1 exu_U13990(.A(byp_irf_rd_data_w[27]), .B(exu_n16289), .Y(exu_n25891));
INVX1 exu_U13991(.A(exu_n25891), .Y(exu_n2419));
AND2X1 exu_U13992(.A(byp_irf_rd_data_w[26]), .B(exu_n16289), .Y(exu_n25895));
INVX1 exu_U13993(.A(exu_n25895), .Y(exu_n2420));
AND2X1 exu_U13994(.A(byp_irf_rd_data_w[25]), .B(exu_n16289), .Y(exu_n25899));
INVX1 exu_U13995(.A(exu_n25899), .Y(exu_n2421));
AND2X1 exu_U13996(.A(byp_irf_rd_data_w[24]), .B(exu_n16289), .Y(exu_n25903));
INVX1 exu_U13997(.A(exu_n25903), .Y(exu_n2422));
AND2X1 exu_U13998(.A(byp_irf_rd_data_w[23]), .B(exu_n16289), .Y(exu_n25907));
INVX1 exu_U13999(.A(exu_n25907), .Y(exu_n2423));
AND2X1 exu_U14000(.A(byp_irf_rd_data_w[22]), .B(exu_n16289), .Y(exu_n25911));
INVX1 exu_U14001(.A(exu_n25911), .Y(exu_n2424));
AND2X1 exu_U14002(.A(byp_irf_rd_data_w[21]), .B(exu_n16289), .Y(exu_n25915));
INVX1 exu_U14003(.A(exu_n25915), .Y(exu_n2425));
AND2X1 exu_U14004(.A(byp_irf_rd_data_w[20]), .B(exu_n16289), .Y(exu_n25919));
INVX1 exu_U14005(.A(exu_n25919), .Y(exu_n2426));
AND2X1 exu_U14006(.A(byp_irf_rd_data_w[1]), .B(exu_n16289), .Y(exu_n25923));
INVX1 exu_U14007(.A(exu_n25923), .Y(exu_n2427));
AND2X1 exu_U14008(.A(byp_irf_rd_data_w[19]), .B(exu_n16289), .Y(exu_n25927));
INVX1 exu_U14009(.A(exu_n25927), .Y(exu_n2428));
AND2X1 exu_U14010(.A(byp_irf_rd_data_w[18]), .B(exu_n16289), .Y(exu_n25931));
INVX1 exu_U14011(.A(exu_n25931), .Y(exu_n2429));
AND2X1 exu_U14012(.A(byp_irf_rd_data_w[17]), .B(exu_n16289), .Y(exu_n25935));
INVX1 exu_U14013(.A(exu_n25935), .Y(exu_n2430));
AND2X1 exu_U14014(.A(byp_irf_rd_data_w[16]), .B(exu_n16289), .Y(exu_n25939));
INVX1 exu_U14015(.A(exu_n25939), .Y(exu_n2431));
AND2X1 exu_U14016(.A(byp_irf_rd_data_w[15]), .B(exu_n16289), .Y(exu_n25943));
INVX1 exu_U14017(.A(exu_n25943), .Y(exu_n2432));
AND2X1 exu_U14018(.A(byp_irf_rd_data_w[14]), .B(exu_n16289), .Y(exu_n25947));
INVX1 exu_U14019(.A(exu_n25947), .Y(exu_n2433));
AND2X1 exu_U14020(.A(byp_irf_rd_data_w[13]), .B(exu_n16289), .Y(exu_n25951));
INVX1 exu_U14021(.A(exu_n25951), .Y(exu_n2434));
AND2X1 exu_U14022(.A(byp_irf_rd_data_w[12]), .B(exu_n16289), .Y(exu_n25955));
INVX1 exu_U14023(.A(exu_n25955), .Y(exu_n2435));
AND2X1 exu_U14024(.A(byp_irf_rd_data_w[11]), .B(exu_n16289), .Y(exu_n25959));
INVX1 exu_U14025(.A(exu_n25959), .Y(exu_n2436));
AND2X1 exu_U14026(.A(byp_irf_rd_data_w[10]), .B(exu_n16289), .Y(exu_n25963));
INVX1 exu_U14027(.A(exu_n25963), .Y(exu_n2437));
AND2X1 exu_U14028(.A(byp_irf_rd_data_w[0]), .B(exu_n16289), .Y(exu_n25967));
INVX1 exu_U14029(.A(exu_n25967), .Y(exu_n2438));
AND2X1 exu_U14030(.A(exu_n16291), .B(lsu_exu_dfill_data_g[9]), .Y(exu_n25971));
INVX1 exu_U14031(.A(exu_n25971), .Y(exu_n2439));
AND2X1 exu_U14032(.A(exu_n16004), .B(bypass_mux_rs3_data_2_in1[9]), .Y(exu_n25973));
INVX1 exu_U14033(.A(exu_n25973), .Y(exu_n2440));
AND2X1 exu_U14034(.A(lsu_exu_dfill_data_g[8]), .B(exu_n16291), .Y(exu_n25977));
INVX1 exu_U14035(.A(exu_n25977), .Y(exu_n2441));
AND2X1 exu_U14036(.A(bypass_mux_rs3_data_2_in1[8]), .B(exu_n16004), .Y(exu_n25979));
INVX1 exu_U14037(.A(exu_n25979), .Y(exu_n2442));
AND2X1 exu_U14038(.A(lsu_exu_dfill_data_g[7]), .B(exu_n16291), .Y(exu_n25983));
INVX1 exu_U14039(.A(exu_n25983), .Y(exu_n2443));
AND2X1 exu_U14040(.A(bypass_mux_rs3_data_2_in1[7]), .B(exu_n16004), .Y(exu_n25985));
INVX1 exu_U14041(.A(exu_n25985), .Y(exu_n2444));
AND2X1 exu_U14042(.A(lsu_exu_dfill_data_g[6]), .B(exu_n16291), .Y(exu_n25989));
INVX1 exu_U14043(.A(exu_n25989), .Y(exu_n2445));
AND2X1 exu_U14044(.A(bypass_mux_rs3_data_2_in1[6]), .B(exu_n16004), .Y(exu_n25991));
INVX1 exu_U14045(.A(exu_n25991), .Y(exu_n2446));
AND2X1 exu_U14046(.A(lsu_exu_dfill_data_g[63]), .B(exu_n16291), .Y(exu_n25995));
INVX1 exu_U14047(.A(exu_n25995), .Y(exu_n2447));
AND2X1 exu_U14048(.A(bypass_mux_rs3_data_2_in1[63]), .B(exu_n16004), .Y(exu_n25997));
INVX1 exu_U14049(.A(exu_n25997), .Y(exu_n2448));
AND2X1 exu_U14050(.A(lsu_exu_dfill_data_g[62]), .B(exu_n16291), .Y(exu_n26001));
INVX1 exu_U14051(.A(exu_n26001), .Y(exu_n2449));
AND2X1 exu_U14052(.A(bypass_mux_rs3_data_2_in1[62]), .B(exu_n16004), .Y(exu_n26003));
INVX1 exu_U14053(.A(exu_n26003), .Y(exu_n2450));
AND2X1 exu_U14054(.A(lsu_exu_dfill_data_g[61]), .B(exu_n16291), .Y(exu_n26007));
INVX1 exu_U14055(.A(exu_n26007), .Y(exu_n2451));
AND2X1 exu_U14056(.A(bypass_mux_rs3_data_2_in1[61]), .B(exu_n16004), .Y(exu_n26009));
INVX1 exu_U14057(.A(exu_n26009), .Y(exu_n2452));
AND2X1 exu_U14058(.A(lsu_exu_dfill_data_g[60]), .B(exu_n16291), .Y(exu_n26013));
INVX1 exu_U14059(.A(exu_n26013), .Y(exu_n2453));
AND2X1 exu_U14060(.A(bypass_mux_rs3_data_2_in1[60]), .B(exu_n16004), .Y(exu_n26015));
INVX1 exu_U14061(.A(exu_n26015), .Y(exu_n2454));
AND2X1 exu_U14062(.A(lsu_exu_dfill_data_g[5]), .B(exu_n16291), .Y(exu_n26019));
INVX1 exu_U14063(.A(exu_n26019), .Y(exu_n2455));
AND2X1 exu_U14064(.A(bypass_mux_rs3_data_2_in1[5]), .B(exu_n16004), .Y(exu_n26021));
INVX1 exu_U14065(.A(exu_n26021), .Y(exu_n2456));
AND2X1 exu_U14066(.A(lsu_exu_dfill_data_g[59]), .B(exu_n16291), .Y(exu_n26025));
INVX1 exu_U14067(.A(exu_n26025), .Y(exu_n2457));
AND2X1 exu_U14068(.A(bypass_mux_rs3_data_2_in1[59]), .B(exu_n16004), .Y(exu_n26027));
INVX1 exu_U14069(.A(exu_n26027), .Y(exu_n2458));
AND2X1 exu_U14070(.A(lsu_exu_dfill_data_g[58]), .B(exu_n16291), .Y(exu_n26031));
INVX1 exu_U14071(.A(exu_n26031), .Y(exu_n2459));
AND2X1 exu_U14072(.A(bypass_mux_rs3_data_2_in1[58]), .B(exu_n16004), .Y(exu_n26033));
INVX1 exu_U14073(.A(exu_n26033), .Y(exu_n2460));
AND2X1 exu_U14074(.A(lsu_exu_dfill_data_g[57]), .B(exu_n16291), .Y(exu_n26037));
INVX1 exu_U14075(.A(exu_n26037), .Y(exu_n2461));
AND2X1 exu_U14076(.A(bypass_mux_rs3_data_2_in1[57]), .B(exu_n16004), .Y(exu_n26039));
INVX1 exu_U14077(.A(exu_n26039), .Y(exu_n2462));
AND2X1 exu_U14078(.A(lsu_exu_dfill_data_g[56]), .B(exu_n16291), .Y(exu_n26043));
INVX1 exu_U14079(.A(exu_n26043), .Y(exu_n2463));
AND2X1 exu_U14080(.A(bypass_mux_rs3_data_2_in1[56]), .B(exu_n16004), .Y(exu_n26045));
INVX1 exu_U14081(.A(exu_n26045), .Y(exu_n2464));
AND2X1 exu_U14082(.A(lsu_exu_dfill_data_g[55]), .B(exu_n16291), .Y(exu_n26049));
INVX1 exu_U14083(.A(exu_n26049), .Y(exu_n2465));
AND2X1 exu_U14084(.A(bypass_mux_rs3_data_2_in1[55]), .B(exu_n16004), .Y(exu_n26051));
INVX1 exu_U14085(.A(exu_n26051), .Y(exu_n2466));
AND2X1 exu_U14086(.A(lsu_exu_dfill_data_g[54]), .B(exu_n16291), .Y(exu_n26055));
INVX1 exu_U14087(.A(exu_n26055), .Y(exu_n2467));
AND2X1 exu_U14088(.A(bypass_mux_rs3_data_2_in1[54]), .B(exu_n16004), .Y(exu_n26057));
INVX1 exu_U14089(.A(exu_n26057), .Y(exu_n2468));
AND2X1 exu_U14090(.A(lsu_exu_dfill_data_g[53]), .B(exu_n16291), .Y(exu_n26061));
INVX1 exu_U14091(.A(exu_n26061), .Y(exu_n2469));
AND2X1 exu_U14092(.A(bypass_mux_rs3_data_2_in1[53]), .B(exu_n16004), .Y(exu_n26063));
INVX1 exu_U14093(.A(exu_n26063), .Y(exu_n2470));
AND2X1 exu_U14094(.A(lsu_exu_dfill_data_g[52]), .B(exu_n16291), .Y(exu_n26067));
INVX1 exu_U14095(.A(exu_n26067), .Y(exu_n2471));
AND2X1 exu_U14096(.A(bypass_mux_rs3_data_2_in1[52]), .B(exu_n16004), .Y(exu_n26069));
INVX1 exu_U14097(.A(exu_n26069), .Y(exu_n2472));
AND2X1 exu_U14098(.A(lsu_exu_dfill_data_g[51]), .B(exu_n16291), .Y(exu_n26073));
INVX1 exu_U14099(.A(exu_n26073), .Y(exu_n2473));
AND2X1 exu_U14100(.A(bypass_mux_rs3_data_2_in1[51]), .B(exu_n16004), .Y(exu_n26075));
INVX1 exu_U14101(.A(exu_n26075), .Y(exu_n2474));
AND2X1 exu_U14102(.A(lsu_exu_dfill_data_g[50]), .B(exu_n16291), .Y(exu_n26079));
INVX1 exu_U14103(.A(exu_n26079), .Y(exu_n2475));
AND2X1 exu_U14104(.A(bypass_mux_rs3_data_2_in1[50]), .B(exu_n16004), .Y(exu_n26081));
INVX1 exu_U14105(.A(exu_n26081), .Y(exu_n2476));
AND2X1 exu_U14106(.A(lsu_exu_dfill_data_g[4]), .B(exu_n16291), .Y(exu_n26085));
INVX1 exu_U14107(.A(exu_n26085), .Y(exu_n2477));
AND2X1 exu_U14108(.A(bypass_mux_rs3_data_2_in1[4]), .B(exu_n16004), .Y(exu_n26087));
INVX1 exu_U14109(.A(exu_n26087), .Y(exu_n2478));
AND2X1 exu_U14110(.A(lsu_exu_dfill_data_g[49]), .B(exu_n16291), .Y(exu_n26091));
INVX1 exu_U14111(.A(exu_n26091), .Y(exu_n2479));
AND2X1 exu_U14112(.A(bypass_mux_rs3_data_2_in1[49]), .B(exu_n16004), .Y(exu_n26093));
INVX1 exu_U14113(.A(exu_n26093), .Y(exu_n2480));
AND2X1 exu_U14114(.A(lsu_exu_dfill_data_g[48]), .B(exu_n16291), .Y(exu_n26097));
INVX1 exu_U14115(.A(exu_n26097), .Y(exu_n2481));
AND2X1 exu_U14116(.A(bypass_mux_rs3_data_2_in1[48]), .B(exu_n16004), .Y(exu_n26099));
INVX1 exu_U14117(.A(exu_n26099), .Y(exu_n2482));
AND2X1 exu_U14118(.A(lsu_exu_dfill_data_g[47]), .B(exu_n16291), .Y(exu_n26103));
INVX1 exu_U14119(.A(exu_n26103), .Y(exu_n2483));
AND2X1 exu_U14120(.A(bypass_mux_rs3_data_2_in1[47]), .B(exu_n16004), .Y(exu_n26105));
INVX1 exu_U14121(.A(exu_n26105), .Y(exu_n2484));
AND2X1 exu_U14122(.A(lsu_exu_dfill_data_g[46]), .B(exu_n16291), .Y(exu_n26109));
INVX1 exu_U14123(.A(exu_n26109), .Y(exu_n2485));
AND2X1 exu_U14124(.A(bypass_mux_rs3_data_2_in1[46]), .B(exu_n16004), .Y(exu_n26111));
INVX1 exu_U14125(.A(exu_n26111), .Y(exu_n2486));
AND2X1 exu_U14126(.A(lsu_exu_dfill_data_g[45]), .B(exu_n16291), .Y(exu_n26115));
INVX1 exu_U14127(.A(exu_n26115), .Y(exu_n2487));
AND2X1 exu_U14128(.A(bypass_mux_rs3_data_2_in1[45]), .B(exu_n16004), .Y(exu_n26117));
INVX1 exu_U14129(.A(exu_n26117), .Y(exu_n2488));
AND2X1 exu_U14130(.A(lsu_exu_dfill_data_g[44]), .B(exu_n16291), .Y(exu_n26121));
INVX1 exu_U14131(.A(exu_n26121), .Y(exu_n2489));
AND2X1 exu_U14132(.A(bypass_mux_rs3_data_2_in1[44]), .B(exu_n16004), .Y(exu_n26123));
INVX1 exu_U14133(.A(exu_n26123), .Y(exu_n2490));
AND2X1 exu_U14134(.A(lsu_exu_dfill_data_g[43]), .B(exu_n16291), .Y(exu_n26127));
INVX1 exu_U14135(.A(exu_n26127), .Y(exu_n2491));
AND2X1 exu_U14136(.A(bypass_mux_rs3_data_2_in1[43]), .B(exu_n16004), .Y(exu_n26129));
INVX1 exu_U14137(.A(exu_n26129), .Y(exu_n2492));
AND2X1 exu_U14138(.A(lsu_exu_dfill_data_g[42]), .B(exu_n16291), .Y(exu_n26133));
INVX1 exu_U14139(.A(exu_n26133), .Y(exu_n2493));
AND2X1 exu_U14140(.A(bypass_mux_rs3_data_2_in1[42]), .B(exu_n16004), .Y(exu_n26135));
INVX1 exu_U14141(.A(exu_n26135), .Y(exu_n2494));
AND2X1 exu_U14142(.A(lsu_exu_dfill_data_g[41]), .B(exu_n16291), .Y(exu_n26139));
INVX1 exu_U14143(.A(exu_n26139), .Y(exu_n2495));
AND2X1 exu_U14144(.A(bypass_mux_rs3_data_2_in1[41]), .B(exu_n16004), .Y(exu_n26141));
INVX1 exu_U14145(.A(exu_n26141), .Y(exu_n2496));
AND2X1 exu_U14146(.A(lsu_exu_dfill_data_g[40]), .B(exu_n16291), .Y(exu_n26145));
INVX1 exu_U14147(.A(exu_n26145), .Y(exu_n2497));
AND2X1 exu_U14148(.A(bypass_mux_rs3_data_2_in1[40]), .B(exu_n16004), .Y(exu_n26147));
INVX1 exu_U14149(.A(exu_n26147), .Y(exu_n2498));
AND2X1 exu_U14150(.A(lsu_exu_dfill_data_g[3]), .B(exu_n16291), .Y(exu_n26151));
INVX1 exu_U14151(.A(exu_n26151), .Y(exu_n2499));
AND2X1 exu_U14152(.A(bypass_mux_rs3_data_2_in1[3]), .B(exu_n16004), .Y(exu_n26153));
INVX1 exu_U14153(.A(exu_n26153), .Y(exu_n2500));
AND2X1 exu_U14154(.A(lsu_exu_dfill_data_g[39]), .B(exu_n16291), .Y(exu_n26157));
INVX1 exu_U14155(.A(exu_n26157), .Y(exu_n2501));
AND2X1 exu_U14156(.A(bypass_mux_rs3_data_2_in1[39]), .B(exu_n16004), .Y(exu_n26159));
INVX1 exu_U14157(.A(exu_n26159), .Y(exu_n2502));
AND2X1 exu_U14158(.A(lsu_exu_dfill_data_g[38]), .B(exu_n16291), .Y(exu_n26163));
INVX1 exu_U14159(.A(exu_n26163), .Y(exu_n2503));
AND2X1 exu_U14160(.A(bypass_mux_rs3_data_2_in1[38]), .B(exu_n16004), .Y(exu_n26165));
INVX1 exu_U14161(.A(exu_n26165), .Y(exu_n2504));
AND2X1 exu_U14162(.A(lsu_exu_dfill_data_g[37]), .B(exu_n16291), .Y(exu_n26169));
INVX1 exu_U14163(.A(exu_n26169), .Y(exu_n2505));
AND2X1 exu_U14164(.A(bypass_mux_rs3_data_2_in1[37]), .B(exu_n16004), .Y(exu_n26171));
INVX1 exu_U14165(.A(exu_n26171), .Y(exu_n2506));
AND2X1 exu_U14166(.A(lsu_exu_dfill_data_g[36]), .B(exu_n16291), .Y(exu_n26175));
INVX1 exu_U14167(.A(exu_n26175), .Y(exu_n2507));
AND2X1 exu_U14168(.A(bypass_mux_rs3_data_2_in1[36]), .B(exu_n16004), .Y(exu_n26177));
INVX1 exu_U14169(.A(exu_n26177), .Y(exu_n2508));
AND2X1 exu_U14170(.A(lsu_exu_dfill_data_g[35]), .B(exu_n16291), .Y(exu_n26181));
INVX1 exu_U14171(.A(exu_n26181), .Y(exu_n2509));
AND2X1 exu_U14172(.A(bypass_mux_rs3_data_2_in1[35]), .B(exu_n16004), .Y(exu_n26183));
INVX1 exu_U14173(.A(exu_n26183), .Y(exu_n2510));
AND2X1 exu_U14174(.A(lsu_exu_dfill_data_g[34]), .B(exu_n16291), .Y(exu_n26187));
INVX1 exu_U14175(.A(exu_n26187), .Y(exu_n2511));
AND2X1 exu_U14176(.A(bypass_mux_rs3_data_2_in1[34]), .B(exu_n16004), .Y(exu_n26189));
INVX1 exu_U14177(.A(exu_n26189), .Y(exu_n2512));
AND2X1 exu_U14178(.A(lsu_exu_dfill_data_g[33]), .B(exu_n16291), .Y(exu_n26193));
INVX1 exu_U14179(.A(exu_n26193), .Y(exu_n2513));
AND2X1 exu_U14180(.A(bypass_mux_rs3_data_2_in1[33]), .B(exu_n16004), .Y(exu_n26195));
INVX1 exu_U14181(.A(exu_n26195), .Y(exu_n2514));
AND2X1 exu_U14182(.A(lsu_exu_dfill_data_g[32]), .B(exu_n16291), .Y(exu_n26199));
INVX1 exu_U14183(.A(exu_n26199), .Y(exu_n2515));
AND2X1 exu_U14184(.A(bypass_mux_rs3_data_2_in1[32]), .B(exu_n16004), .Y(exu_n26201));
INVX1 exu_U14185(.A(exu_n26201), .Y(exu_n2516));
AND2X1 exu_U14186(.A(lsu_exu_dfill_data_g[31]), .B(exu_n16291), .Y(exu_n26205));
INVX1 exu_U14187(.A(exu_n26205), .Y(exu_n2517));
AND2X1 exu_U14188(.A(bypass_mux_rs3_data_2_in1[31]), .B(exu_n16004), .Y(exu_n26207));
INVX1 exu_U14189(.A(exu_n26207), .Y(exu_n2518));
AND2X1 exu_U14190(.A(lsu_exu_dfill_data_g[30]), .B(exu_n16291), .Y(exu_n26211));
INVX1 exu_U14191(.A(exu_n26211), .Y(exu_n2519));
AND2X1 exu_U14192(.A(bypass_mux_rs3_data_2_in1[30]), .B(exu_n16004), .Y(exu_n26213));
INVX1 exu_U14193(.A(exu_n26213), .Y(exu_n2520));
AND2X1 exu_U14194(.A(lsu_exu_dfill_data_g[2]), .B(exu_n16291), .Y(exu_n26217));
INVX1 exu_U14195(.A(exu_n26217), .Y(exu_n2521));
AND2X1 exu_U14196(.A(bypass_mux_rs3_data_2_in1[2]), .B(exu_n16004), .Y(exu_n26219));
INVX1 exu_U14197(.A(exu_n26219), .Y(exu_n2522));
AND2X1 exu_U14198(.A(lsu_exu_dfill_data_g[29]), .B(exu_n16291), .Y(exu_n26223));
INVX1 exu_U14199(.A(exu_n26223), .Y(exu_n2523));
AND2X1 exu_U14200(.A(bypass_mux_rs3_data_2_in1[29]), .B(exu_n16004), .Y(exu_n26225));
INVX1 exu_U14201(.A(exu_n26225), .Y(exu_n2524));
AND2X1 exu_U14202(.A(lsu_exu_dfill_data_g[28]), .B(exu_n16291), .Y(exu_n26229));
INVX1 exu_U14203(.A(exu_n26229), .Y(exu_n2525));
AND2X1 exu_U14204(.A(bypass_mux_rs3_data_2_in1[28]), .B(exu_n16004), .Y(exu_n26231));
INVX1 exu_U14205(.A(exu_n26231), .Y(exu_n2526));
AND2X1 exu_U14206(.A(lsu_exu_dfill_data_g[27]), .B(exu_n16291), .Y(exu_n26235));
INVX1 exu_U14207(.A(exu_n26235), .Y(exu_n2527));
AND2X1 exu_U14208(.A(bypass_mux_rs3_data_2_in1[27]), .B(exu_n16004), .Y(exu_n26237));
INVX1 exu_U14209(.A(exu_n26237), .Y(exu_n2528));
AND2X1 exu_U14210(.A(lsu_exu_dfill_data_g[26]), .B(exu_n16291), .Y(exu_n26241));
INVX1 exu_U14211(.A(exu_n26241), .Y(exu_n2529));
AND2X1 exu_U14212(.A(bypass_mux_rs3_data_2_in1[26]), .B(exu_n16004), .Y(exu_n26243));
INVX1 exu_U14213(.A(exu_n26243), .Y(exu_n2530));
AND2X1 exu_U14214(.A(lsu_exu_dfill_data_g[25]), .B(exu_n16291), .Y(exu_n26247));
INVX1 exu_U14215(.A(exu_n26247), .Y(exu_n2531));
AND2X1 exu_U14216(.A(bypass_mux_rs3_data_2_in1[25]), .B(exu_n16004), .Y(exu_n26249));
INVX1 exu_U14217(.A(exu_n26249), .Y(exu_n2532));
AND2X1 exu_U14218(.A(lsu_exu_dfill_data_g[24]), .B(exu_n16291), .Y(exu_n26253));
INVX1 exu_U14219(.A(exu_n26253), .Y(exu_n2533));
AND2X1 exu_U14220(.A(bypass_mux_rs3_data_2_in1[24]), .B(exu_n16004), .Y(exu_n26255));
INVX1 exu_U14221(.A(exu_n26255), .Y(exu_n2534));
AND2X1 exu_U14222(.A(lsu_exu_dfill_data_g[23]), .B(exu_n16291), .Y(exu_n26259));
INVX1 exu_U14223(.A(exu_n26259), .Y(exu_n2535));
AND2X1 exu_U14224(.A(bypass_mux_rs3_data_2_in1[23]), .B(exu_n16004), .Y(exu_n26261));
INVX1 exu_U14225(.A(exu_n26261), .Y(exu_n2536));
AND2X1 exu_U14226(.A(lsu_exu_dfill_data_g[22]), .B(exu_n16291), .Y(exu_n26265));
INVX1 exu_U14227(.A(exu_n26265), .Y(exu_n2537));
AND2X1 exu_U14228(.A(bypass_mux_rs3_data_2_in1[22]), .B(exu_n16004), .Y(exu_n26267));
INVX1 exu_U14229(.A(exu_n26267), .Y(exu_n2538));
AND2X1 exu_U14230(.A(lsu_exu_dfill_data_g[21]), .B(exu_n16291), .Y(exu_n26271));
INVX1 exu_U14231(.A(exu_n26271), .Y(exu_n2539));
AND2X1 exu_U14232(.A(bypass_mux_rs3_data_2_in1[21]), .B(exu_n16004), .Y(exu_n26273));
INVX1 exu_U14233(.A(exu_n26273), .Y(exu_n2540));
AND2X1 exu_U14234(.A(lsu_exu_dfill_data_g[20]), .B(exu_n16291), .Y(exu_n26277));
INVX1 exu_U14235(.A(exu_n26277), .Y(exu_n2541));
AND2X1 exu_U14236(.A(bypass_mux_rs3_data_2_in1[20]), .B(exu_n16004), .Y(exu_n26279));
INVX1 exu_U14237(.A(exu_n26279), .Y(exu_n2542));
AND2X1 exu_U14238(.A(lsu_exu_dfill_data_g[1]), .B(exu_n16291), .Y(exu_n26283));
INVX1 exu_U14239(.A(exu_n26283), .Y(exu_n2543));
AND2X1 exu_U14240(.A(bypass_mux_rs3_data_2_in1[1]), .B(exu_n16004), .Y(exu_n26285));
INVX1 exu_U14241(.A(exu_n26285), .Y(exu_n2544));
AND2X1 exu_U14242(.A(lsu_exu_dfill_data_g[19]), .B(exu_n16291), .Y(exu_n26289));
INVX1 exu_U14243(.A(exu_n26289), .Y(exu_n2545));
AND2X1 exu_U14244(.A(bypass_mux_rs3_data_2_in1[19]), .B(exu_n16004), .Y(exu_n26291));
INVX1 exu_U14245(.A(exu_n26291), .Y(exu_n2546));
AND2X1 exu_U14246(.A(lsu_exu_dfill_data_g[18]), .B(exu_n16291), .Y(exu_n26295));
INVX1 exu_U14247(.A(exu_n26295), .Y(exu_n2547));
AND2X1 exu_U14248(.A(bypass_mux_rs3_data_2_in1[18]), .B(exu_n16004), .Y(exu_n26297));
INVX1 exu_U14249(.A(exu_n26297), .Y(exu_n2548));
AND2X1 exu_U14250(.A(lsu_exu_dfill_data_g[17]), .B(exu_n16291), .Y(exu_n26301));
INVX1 exu_U14251(.A(exu_n26301), .Y(exu_n2549));
AND2X1 exu_U14252(.A(bypass_mux_rs3_data_2_in1[17]), .B(exu_n16004), .Y(exu_n26303));
INVX1 exu_U14253(.A(exu_n26303), .Y(exu_n2550));
AND2X1 exu_U14254(.A(lsu_exu_dfill_data_g[16]), .B(exu_n16291), .Y(exu_n26307));
INVX1 exu_U14255(.A(exu_n26307), .Y(exu_n2551));
AND2X1 exu_U14256(.A(bypass_mux_rs3_data_2_in1[16]), .B(exu_n16004), .Y(exu_n26309));
INVX1 exu_U14257(.A(exu_n26309), .Y(exu_n2552));
AND2X1 exu_U14258(.A(lsu_exu_dfill_data_g[15]), .B(exu_n16291), .Y(exu_n26313));
INVX1 exu_U14259(.A(exu_n26313), .Y(exu_n2553));
AND2X1 exu_U14260(.A(bypass_mux_rs3_data_2_in1[15]), .B(exu_n16004), .Y(exu_n26315));
INVX1 exu_U14261(.A(exu_n26315), .Y(exu_n2554));
AND2X1 exu_U14262(.A(lsu_exu_dfill_data_g[14]), .B(exu_n16291), .Y(exu_n26319));
INVX1 exu_U14263(.A(exu_n26319), .Y(exu_n2555));
AND2X1 exu_U14264(.A(bypass_mux_rs3_data_2_in1[14]), .B(exu_n16004), .Y(exu_n26321));
INVX1 exu_U14265(.A(exu_n26321), .Y(exu_n2556));
AND2X1 exu_U14266(.A(lsu_exu_dfill_data_g[13]), .B(exu_n16291), .Y(exu_n26325));
INVX1 exu_U14267(.A(exu_n26325), .Y(exu_n2557));
AND2X1 exu_U14268(.A(bypass_mux_rs3_data_2_in1[13]), .B(exu_n16004), .Y(exu_n26327));
INVX1 exu_U14269(.A(exu_n26327), .Y(exu_n2558));
AND2X1 exu_U14270(.A(lsu_exu_dfill_data_g[12]), .B(exu_n16291), .Y(exu_n26331));
INVX1 exu_U14271(.A(exu_n26331), .Y(exu_n2559));
AND2X1 exu_U14272(.A(bypass_mux_rs3_data_2_in1[12]), .B(exu_n16004), .Y(exu_n26333));
INVX1 exu_U14273(.A(exu_n26333), .Y(exu_n2560));
AND2X1 exu_U14274(.A(lsu_exu_dfill_data_g[11]), .B(exu_n16291), .Y(exu_n26337));
INVX1 exu_U14275(.A(exu_n26337), .Y(exu_n2561));
AND2X1 exu_U14276(.A(bypass_mux_rs3_data_2_in1[11]), .B(exu_n16004), .Y(exu_n26339));
INVX1 exu_U14277(.A(exu_n26339), .Y(exu_n2562));
AND2X1 exu_U14278(.A(lsu_exu_dfill_data_g[10]), .B(exu_n16291), .Y(exu_n26343));
INVX1 exu_U14279(.A(exu_n26343), .Y(exu_n2563));
AND2X1 exu_U14280(.A(bypass_mux_rs3_data_2_in1[10]), .B(exu_n16004), .Y(exu_n26345));
INVX1 exu_U14281(.A(exu_n26345), .Y(exu_n2564));
AND2X1 exu_U14282(.A(lsu_exu_dfill_data_g[0]), .B(exu_n16291), .Y(exu_n26349));
INVX1 exu_U14283(.A(exu_n26349), .Y(exu_n2565));
AND2X1 exu_U14284(.A(bypass_mux_rs3_data_2_in1[0]), .B(exu_n16004), .Y(exu_n26351));
INVX1 exu_U14285(.A(exu_n26351), .Y(exu_n2566));
AND2X1 exu_U14286(.A(exu_n15969), .B(alu_logic_out_9), .Y(exu_n26355));
INVX1 exu_U14287(.A(exu_n26355), .Y(exu_n2567));
AND2X1 exu_U14288(.A(exu_n15971), .B(exu_lsu_rs3_data_e[9]), .Y(exu_n26357));
INVX1 exu_U14289(.A(exu_n26357), .Y(exu_n2568));
AND2X1 exu_U14290(.A(alu_logic_out_8), .B(exu_n15969), .Y(exu_n26361));
INVX1 exu_U14291(.A(exu_n26361), .Y(exu_n2569));
AND2X1 exu_U14292(.A(exu_lsu_rs3_data_e[8]), .B(exu_n15971), .Y(exu_n26363));
INVX1 exu_U14293(.A(exu_n26363), .Y(exu_n2570));
AND2X1 exu_U14294(.A(alu_logic_out_7), .B(exu_n15969), .Y(exu_n26367));
INVX1 exu_U14295(.A(exu_n26367), .Y(exu_n2571));
AND2X1 exu_U14296(.A(exu_lsu_rs3_data_e[7]), .B(exu_n15971), .Y(exu_n26369));
INVX1 exu_U14297(.A(exu_n26369), .Y(exu_n2572));
AND2X1 exu_U14298(.A(alu_logic_out_6), .B(exu_n15969), .Y(exu_n26373));
INVX1 exu_U14299(.A(exu_n26373), .Y(exu_n2573));
AND2X1 exu_U14300(.A(exu_lsu_rs3_data_e[6]), .B(exu_n15971), .Y(exu_n26375));
INVX1 exu_U14301(.A(exu_n26375), .Y(exu_n2574));
AND2X1 exu_U14302(.A(alu_ecl_log_n64_e), .B(exu_n15969), .Y(exu_n26379));
INVX1 exu_U14303(.A(exu_n26379), .Y(exu_n2575));
AND2X1 exu_U14304(.A(exu_lsu_rs3_data_e[63]), .B(exu_n15971), .Y(exu_n26381));
INVX1 exu_U14305(.A(exu_n26381), .Y(exu_n2576));
AND2X1 exu_U14306(.A(alu_logic_out[62]), .B(exu_n15969), .Y(exu_n26384));
INVX1 exu_U14307(.A(exu_n26384), .Y(exu_n2577));
AND2X1 exu_U14308(.A(exu_lsu_rs3_data_e[62]), .B(exu_n15971), .Y(exu_n26386));
INVX1 exu_U14309(.A(exu_n26386), .Y(exu_n2578));
AND2X1 exu_U14310(.A(alu_logic_out[61]), .B(exu_n15969), .Y(exu_n26390));
INVX1 exu_U14311(.A(exu_n26390), .Y(exu_n2579));
AND2X1 exu_U14312(.A(exu_lsu_rs3_data_e[61]), .B(exu_n15971), .Y(exu_n26392));
INVX1 exu_U14313(.A(exu_n26392), .Y(exu_n2580));
AND2X1 exu_U14314(.A(alu_logic_out[60]), .B(exu_n15969), .Y(exu_n26396));
INVX1 exu_U14315(.A(exu_n26396), .Y(exu_n2581));
AND2X1 exu_U14316(.A(exu_lsu_rs3_data_e[60]), .B(exu_n15971), .Y(exu_n26398));
INVX1 exu_U14317(.A(exu_n26398), .Y(exu_n2582));
AND2X1 exu_U14318(.A(alu_logic_out_5), .B(exu_n15969), .Y(exu_n26402));
INVX1 exu_U14319(.A(exu_n26402), .Y(exu_n2583));
AND2X1 exu_U14320(.A(exu_lsu_rs3_data_e[5]), .B(exu_n15971), .Y(exu_n26404));
INVX1 exu_U14321(.A(exu_n26404), .Y(exu_n2584));
AND2X1 exu_U14322(.A(alu_logic_out[59]), .B(exu_n15969), .Y(exu_n26408));
INVX1 exu_U14323(.A(exu_n26408), .Y(exu_n2585));
AND2X1 exu_U14324(.A(exu_lsu_rs3_data_e[59]), .B(exu_n15971), .Y(exu_n26410));
INVX1 exu_U14325(.A(exu_n26410), .Y(exu_n2586));
AND2X1 exu_U14326(.A(alu_logic_out[58]), .B(exu_n15969), .Y(exu_n26414));
INVX1 exu_U14327(.A(exu_n26414), .Y(exu_n2587));
AND2X1 exu_U14328(.A(exu_lsu_rs3_data_e[58]), .B(exu_n15971), .Y(exu_n26416));
INVX1 exu_U14329(.A(exu_n26416), .Y(exu_n2588));
AND2X1 exu_U14330(.A(alu_logic_out[57]), .B(exu_n15969), .Y(exu_n26420));
INVX1 exu_U14331(.A(exu_n26420), .Y(exu_n2589));
AND2X1 exu_U14332(.A(exu_lsu_rs3_data_e[57]), .B(exu_n15971), .Y(exu_n26422));
INVX1 exu_U14333(.A(exu_n26422), .Y(exu_n2590));
AND2X1 exu_U14334(.A(alu_logic_out[56]), .B(exu_n15969), .Y(exu_n26426));
INVX1 exu_U14335(.A(exu_n26426), .Y(exu_n2591));
AND2X1 exu_U14336(.A(exu_lsu_rs3_data_e[56]), .B(exu_n15971), .Y(exu_n26428));
INVX1 exu_U14337(.A(exu_n26428), .Y(exu_n2592));
AND2X1 exu_U14338(.A(alu_logic_out[55]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26432));
INVX1 exu_U14339(.A(exu_n26432), .Y(exu_n2593));
AND2X1 exu_U14340(.A(exu_lsu_rs3_data_e[55]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26434));
INVX1 exu_U14341(.A(exu_n26434), .Y(exu_n2594));
AND2X1 exu_U14342(.A(alu_logic_out[54]), .B(exu_n15969), .Y(exu_n26438));
INVX1 exu_U14343(.A(exu_n26438), .Y(exu_n2595));
AND2X1 exu_U14344(.A(exu_lsu_rs3_data_e[54]), .B(exu_n15971), .Y(exu_n26440));
INVX1 exu_U14345(.A(exu_n26440), .Y(exu_n2596));
AND2X1 exu_U14346(.A(alu_logic_out[53]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26444));
INVX1 exu_U14347(.A(exu_n26444), .Y(exu_n2597));
AND2X1 exu_U14348(.A(exu_lsu_rs3_data_e[53]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26446));
INVX1 exu_U14349(.A(exu_n26446), .Y(exu_n2598));
AND2X1 exu_U14350(.A(alu_logic_out[52]), .B(exu_n15969), .Y(exu_n26450));
INVX1 exu_U14351(.A(exu_n26450), .Y(exu_n2599));
AND2X1 exu_U14352(.A(exu_lsu_rs3_data_e[52]), .B(exu_n15971), .Y(exu_n26452));
INVX1 exu_U14353(.A(exu_n26452), .Y(exu_n2600));
AND2X1 exu_U14354(.A(alu_logic_out[51]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26456));
INVX1 exu_U14355(.A(exu_n26456), .Y(exu_n2601));
AND2X1 exu_U14356(.A(exu_lsu_rs3_data_e[51]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26458));
INVX1 exu_U14357(.A(exu_n26458), .Y(exu_n2602));
AND2X1 exu_U14358(.A(alu_logic_out[50]), .B(exu_n15969), .Y(exu_n26462));
INVX1 exu_U14359(.A(exu_n26462), .Y(exu_n2603));
AND2X1 exu_U14360(.A(exu_lsu_rs3_data_e[50]), .B(exu_n15971), .Y(exu_n26464));
INVX1 exu_U14361(.A(exu_n26464), .Y(exu_n2604));
AND2X1 exu_U14362(.A(alu_logic_out_4), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26468));
INVX1 exu_U14363(.A(exu_n26468), .Y(exu_n2605));
AND2X1 exu_U14364(.A(exu_lsu_rs3_data_e[4]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26470));
INVX1 exu_U14365(.A(exu_n26470), .Y(exu_n2606));
AND2X1 exu_U14366(.A(alu_logic_out[49]), .B(exu_n15969), .Y(exu_n26474));
INVX1 exu_U14367(.A(exu_n26474), .Y(exu_n2607));
AND2X1 exu_U14368(.A(exu_lsu_rs3_data_e[49]), .B(exu_n15971), .Y(exu_n26476));
INVX1 exu_U14369(.A(exu_n26476), .Y(exu_n2608));
AND2X1 exu_U14370(.A(alu_logic_out[48]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26480));
INVX1 exu_U14371(.A(exu_n26480), .Y(exu_n2609));
AND2X1 exu_U14372(.A(exu_lsu_rs3_data_e[48]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26482));
INVX1 exu_U14373(.A(exu_n26482), .Y(exu_n2610));
AND2X1 exu_U14374(.A(alu_logic_out[47]), .B(exu_n15969), .Y(exu_n26486));
INVX1 exu_U14375(.A(exu_n26486), .Y(exu_n2611));
AND2X1 exu_U14376(.A(exu_lsu_rs3_data_e[47]), .B(exu_n15971), .Y(exu_n26488));
INVX1 exu_U14377(.A(exu_n26488), .Y(exu_n2612));
AND2X1 exu_U14378(.A(alu_logic_out[46]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26492));
INVX1 exu_U14379(.A(exu_n26492), .Y(exu_n2613));
AND2X1 exu_U14380(.A(exu_lsu_rs3_data_e[46]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26494));
INVX1 exu_U14381(.A(exu_n26494), .Y(exu_n2614));
AND2X1 exu_U14382(.A(alu_logic_out[45]), .B(exu_n15969), .Y(exu_n26498));
INVX1 exu_U14383(.A(exu_n26498), .Y(exu_n2615));
AND2X1 exu_U14384(.A(exu_lsu_rs3_data_e[45]), .B(exu_n15971), .Y(exu_n26500));
INVX1 exu_U14385(.A(exu_n26500), .Y(exu_n2616));
AND2X1 exu_U14386(.A(alu_logic_out[44]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26504));
INVX1 exu_U14387(.A(exu_n26504), .Y(exu_n2617));
AND2X1 exu_U14388(.A(exu_lsu_rs3_data_e[44]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26506));
INVX1 exu_U14389(.A(exu_n26506), .Y(exu_n2618));
AND2X1 exu_U14390(.A(alu_logic_out[43]), .B(exu_n15969), .Y(exu_n26510));
INVX1 exu_U14391(.A(exu_n26510), .Y(exu_n2619));
AND2X1 exu_U14392(.A(exu_lsu_rs3_data_e[43]), .B(exu_n15971), .Y(exu_n26512));
INVX1 exu_U14393(.A(exu_n26512), .Y(exu_n2620));
AND2X1 exu_U14394(.A(alu_logic_out[42]), .B(exu_n15969), .Y(exu_n26516));
INVX1 exu_U14395(.A(exu_n26516), .Y(exu_n2621));
AND2X1 exu_U14396(.A(exu_lsu_rs3_data_e[42]), .B(exu_n15971), .Y(exu_n26518));
INVX1 exu_U14397(.A(exu_n26518), .Y(exu_n2622));
AND2X1 exu_U14398(.A(alu_logic_out[41]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26522));
INVX1 exu_U14399(.A(exu_n26522), .Y(exu_n2623));
AND2X1 exu_U14400(.A(exu_lsu_rs3_data_e[41]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26524));
INVX1 exu_U14401(.A(exu_n26524), .Y(exu_n2624));
AND2X1 exu_U14402(.A(alu_logic_out[40]), .B(exu_n15969), .Y(exu_n26528));
INVX1 exu_U14403(.A(exu_n26528), .Y(exu_n2625));
AND2X1 exu_U14404(.A(exu_lsu_rs3_data_e[40]), .B(exu_n15971), .Y(exu_n26530));
INVX1 exu_U14405(.A(exu_n26530), .Y(exu_n2626));
AND2X1 exu_U14406(.A(alu_logic_out_3), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26534));
INVX1 exu_U14407(.A(exu_n26534), .Y(exu_n2627));
AND2X1 exu_U14408(.A(exu_lsu_rs3_data_e[3]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26536));
INVX1 exu_U14409(.A(exu_n26536), .Y(exu_n2628));
AND2X1 exu_U14410(.A(alu_logic_out[39]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26540));
INVX1 exu_U14411(.A(exu_n26540), .Y(exu_n2629));
AND2X1 exu_U14412(.A(exu_lsu_rs3_data_e[39]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26542));
INVX1 exu_U14413(.A(exu_n26542), .Y(exu_n2630));
AND2X1 exu_U14414(.A(alu_logic_out[38]), .B(exu_n15969), .Y(exu_n26546));
INVX1 exu_U14415(.A(exu_n26546), .Y(exu_n2631));
AND2X1 exu_U14416(.A(exu_lsu_rs3_data_e[38]), .B(exu_n15971), .Y(exu_n26548));
INVX1 exu_U14417(.A(exu_n26548), .Y(exu_n2632));
AND2X1 exu_U14418(.A(alu_logic_out[37]), .B(exu_n15969), .Y(exu_n26552));
INVX1 exu_U14419(.A(exu_n26552), .Y(exu_n2633));
AND2X1 exu_U14420(.A(exu_lsu_rs3_data_e[37]), .B(exu_n15971), .Y(exu_n26554));
INVX1 exu_U14421(.A(exu_n26554), .Y(exu_n2634));
AND2X1 exu_U14422(.A(alu_logic_out[36]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26558));
INVX1 exu_U14423(.A(exu_n26558), .Y(exu_n2635));
AND2X1 exu_U14424(.A(exu_lsu_rs3_data_e[36]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26560));
INVX1 exu_U14425(.A(exu_n26560), .Y(exu_n2636));
AND2X1 exu_U14426(.A(alu_logic_out[35]), .B(exu_n15969), .Y(exu_n26564));
INVX1 exu_U14427(.A(exu_n26564), .Y(exu_n2637));
AND2X1 exu_U14428(.A(exu_lsu_rs3_data_e[35]), .B(exu_n15971), .Y(exu_n26566));
INVX1 exu_U14429(.A(exu_n26566), .Y(exu_n2638));
AND2X1 exu_U14430(.A(alu_logic_out[34]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26570));
INVX1 exu_U14431(.A(exu_n26570), .Y(exu_n2639));
AND2X1 exu_U14432(.A(exu_lsu_rs3_data_e[34]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26572));
INVX1 exu_U14433(.A(exu_n26572), .Y(exu_n2640));
AND2X1 exu_U14434(.A(alu_logic_out[33]), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26576));
INVX1 exu_U14435(.A(exu_n26576), .Y(exu_n2641));
AND2X1 exu_U14436(.A(exu_lsu_rs3_data_e[33]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26578));
INVX1 exu_U14437(.A(exu_n26578), .Y(exu_n2642));
AND2X1 exu_U14438(.A(alu_logic_out[32]), .B(exu_n15969), .Y(exu_n26582));
INVX1 exu_U14439(.A(exu_n26582), .Y(exu_n2643));
AND2X1 exu_U14440(.A(exu_lsu_rs3_data_e[32]), .B(exu_n15971), .Y(exu_n26584));
INVX1 exu_U14441(.A(exu_n26584), .Y(exu_n2644));
AND2X1 exu_U14442(.A(alu_ecl_log_n32_e), .B(exu_n15969), .Y(exu_n26588));
INVX1 exu_U14443(.A(exu_n26588), .Y(exu_n2645));
AND2X1 exu_U14444(.A(exu_lsu_rs3_data_e[31]), .B(exu_n15971), .Y(exu_n26590));
INVX1 exu_U14445(.A(exu_n26590), .Y(exu_n2646));
AND2X1 exu_U14446(.A(alu_logic_out_30), .B(exu_n15969), .Y(exu_n26593));
INVX1 exu_U14447(.A(exu_n26593), .Y(exu_n2647));
AND2X1 exu_U14448(.A(exu_lsu_rs3_data_e[30]), .B(exu_n15971), .Y(exu_n26595));
INVX1 exu_U14449(.A(exu_n26595), .Y(exu_n2648));
AND2X1 exu_U14450(.A(alu_logic_out_2), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26599));
INVX1 exu_U14451(.A(exu_n26599), .Y(exu_n2649));
AND2X1 exu_U14452(.A(exu_lsu_rs3_data_e[2]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26601));
INVX1 exu_U14453(.A(exu_n26601), .Y(exu_n2650));
AND2X1 exu_U14454(.A(alu_logic_out_29), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26605));
INVX1 exu_U14455(.A(exu_n26605), .Y(exu_n2651));
AND2X1 exu_U14456(.A(exu_lsu_rs3_data_e[29]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26607));
INVX1 exu_U14457(.A(exu_n26607), .Y(exu_n2652));
AND2X1 exu_U14458(.A(alu_logic_out_28), .B(exu_n15969), .Y(exu_n26611));
INVX1 exu_U14459(.A(exu_n26611), .Y(exu_n2653));
AND2X1 exu_U14460(.A(exu_lsu_rs3_data_e[28]), .B(exu_n15971), .Y(exu_n26613));
INVX1 exu_U14461(.A(exu_n26613), .Y(exu_n2654));
AND2X1 exu_U14462(.A(alu_logic_out_27), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26617));
INVX1 exu_U14463(.A(exu_n26617), .Y(exu_n2655));
AND2X1 exu_U14464(.A(exu_lsu_rs3_data_e[27]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26619));
INVX1 exu_U14465(.A(exu_n26619), .Y(exu_n2656));
AND2X1 exu_U14466(.A(alu_logic_out_26), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26623));
INVX1 exu_U14467(.A(exu_n26623), .Y(exu_n2657));
AND2X1 exu_U14468(.A(exu_lsu_rs3_data_e[26]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26625));
INVX1 exu_U14469(.A(exu_n26625), .Y(exu_n2658));
AND2X1 exu_U14470(.A(alu_logic_out_25), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26629));
INVX1 exu_U14471(.A(exu_n26629), .Y(exu_n2659));
AND2X1 exu_U14472(.A(exu_lsu_rs3_data_e[25]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26631));
INVX1 exu_U14473(.A(exu_n26631), .Y(exu_n2660));
AND2X1 exu_U14474(.A(alu_logic_out_24), .B(exu_n15969), .Y(exu_n26635));
INVX1 exu_U14475(.A(exu_n26635), .Y(exu_n2661));
AND2X1 exu_U14476(.A(exu_lsu_rs3_data_e[24]), .B(exu_n15971), .Y(exu_n26637));
INVX1 exu_U14477(.A(exu_n26637), .Y(exu_n2662));
AND2X1 exu_U14478(.A(alu_logic_out_23), .B(exu_n15969), .Y(exu_n26641));
INVX1 exu_U14479(.A(exu_n26641), .Y(exu_n2663));
AND2X1 exu_U14480(.A(exu_lsu_rs3_data_e[23]), .B(exu_n15971), .Y(exu_n26643));
INVX1 exu_U14481(.A(exu_n26643), .Y(exu_n2664));
AND2X1 exu_U14482(.A(alu_logic_out_22), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26647));
INVX1 exu_U14483(.A(exu_n26647), .Y(exu_n2665));
AND2X1 exu_U14484(.A(exu_lsu_rs3_data_e[22]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26649));
INVX1 exu_U14485(.A(exu_n26649), .Y(exu_n2666));
AND2X1 exu_U14486(.A(alu_logic_out_21), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26653));
INVX1 exu_U14487(.A(exu_n26653), .Y(exu_n2667));
AND2X1 exu_U14488(.A(exu_lsu_rs3_data_e[21]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26655));
INVX1 exu_U14489(.A(exu_n26655), .Y(exu_n2668));
AND2X1 exu_U14490(.A(alu_logic_out_20), .B(exu_n15969), .Y(exu_n26659));
INVX1 exu_U14491(.A(exu_n26659), .Y(exu_n2669));
AND2X1 exu_U14492(.A(exu_lsu_rs3_data_e[20]), .B(exu_n15971), .Y(exu_n26661));
INVX1 exu_U14493(.A(exu_n26661), .Y(exu_n2670));
AND2X1 exu_U14494(.A(alu_logic_out_1), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26665));
INVX1 exu_U14495(.A(exu_n26665), .Y(exu_n2671));
AND2X1 exu_U14496(.A(exu_lsu_rs3_data_e[1]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26667));
INVX1 exu_U14497(.A(exu_n26667), .Y(exu_n2672));
AND2X1 exu_U14498(.A(alu_logic_out_19), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26671));
INVX1 exu_U14499(.A(exu_n26671), .Y(exu_n2673));
AND2X1 exu_U14500(.A(exu_lsu_rs3_data_e[19]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26673));
INVX1 exu_U14501(.A(exu_n26673), .Y(exu_n2674));
AND2X1 exu_U14502(.A(alu_logic_out_18), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26677));
INVX1 exu_U14503(.A(exu_n26677), .Y(exu_n2675));
AND2X1 exu_U14504(.A(exu_lsu_rs3_data_e[18]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26679));
INVX1 exu_U14505(.A(exu_n26679), .Y(exu_n2676));
AND2X1 exu_U14506(.A(alu_logic_out_17), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26683));
INVX1 exu_U14507(.A(exu_n26683), .Y(exu_n2677));
AND2X1 exu_U14508(.A(exu_lsu_rs3_data_e[17]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26685));
INVX1 exu_U14509(.A(exu_n26685), .Y(exu_n2678));
AND2X1 exu_U14510(.A(alu_logic_out_16), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26689));
INVX1 exu_U14511(.A(exu_n26689), .Y(exu_n2679));
AND2X1 exu_U14512(.A(exu_lsu_rs3_data_e[16]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26691));
INVX1 exu_U14513(.A(exu_n26691), .Y(exu_n2680));
AND2X1 exu_U14514(.A(alu_logic_out_15), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26695));
INVX1 exu_U14515(.A(exu_n26695), .Y(exu_n2681));
AND2X1 exu_U14516(.A(exu_lsu_rs3_data_e[15]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26697));
INVX1 exu_U14517(.A(exu_n26697), .Y(exu_n2682));
AND2X1 exu_U14518(.A(alu_logic_out_14), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26701));
INVX1 exu_U14519(.A(exu_n26701), .Y(exu_n2683));
AND2X1 exu_U14520(.A(exu_lsu_rs3_data_e[14]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26703));
INVX1 exu_U14521(.A(exu_n26703), .Y(exu_n2684));
AND2X1 exu_U14522(.A(alu_logic_out_13), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26707));
INVX1 exu_U14523(.A(exu_n26707), .Y(exu_n2685));
AND2X1 exu_U14524(.A(exu_lsu_rs3_data_e[13]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26709));
INVX1 exu_U14525(.A(exu_n26709), .Y(exu_n2686));
AND2X1 exu_U14526(.A(alu_logic_out_12), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26713));
INVX1 exu_U14527(.A(exu_n26713), .Y(exu_n2687));
AND2X1 exu_U14528(.A(exu_lsu_rs3_data_e[12]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26715));
INVX1 exu_U14529(.A(exu_n26715), .Y(exu_n2688));
AND2X1 exu_U14530(.A(alu_logic_out_11), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26719));
INVX1 exu_U14531(.A(exu_n26719), .Y(exu_n2689));
AND2X1 exu_U14532(.A(exu_lsu_rs3_data_e[11]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26721));
INVX1 exu_U14533(.A(exu_n26721), .Y(exu_n2690));
AND2X1 exu_U14534(.A(alu_logic_out_10), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26725));
INVX1 exu_U14535(.A(exu_n26725), .Y(exu_n2691));
AND2X1 exu_U14536(.A(exu_lsu_rs3_data_e[10]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26727));
INVX1 exu_U14537(.A(exu_n26727), .Y(exu_n2692));
AND2X1 exu_U14538(.A(alu_logic_out_0), .B(ecl_alu_out_sel_logic_e_l), .Y(exu_n26731));
INVX1 exu_U14539(.A(exu_n26731), .Y(exu_n2693));
AND2X1 exu_U14540(.A(exu_lsu_rs3_data_e[0]), .B(ecl_alu_out_sel_rs3_e_l), .Y(exu_n26733));
INVX1 exu_U14541(.A(exu_n26733), .Y(exu_n2694));
AND2X1 exu_U14542(.A(exu_n16145), .B(exu_n15438), .Y(exu_n26738));
INVX1 exu_U14543(.A(exu_n26738), .Y(exu_n2695));
AND2X1 exu_U14544(.A(exu_n15442), .B(exu_n16145), .Y(exu_n26742));
INVX1 exu_U14545(.A(exu_n26742), .Y(exu_n2696));
AND2X1 exu_U14546(.A(exu_n15443), .B(exu_n16145), .Y(exu_n26746));
INVX1 exu_U14547(.A(exu_n26746), .Y(exu_n2697));
AND2X1 exu_U14548(.A(exu_n15444), .B(exu_n16145), .Y(exu_n26750));
INVX1 exu_U14549(.A(exu_n26750), .Y(exu_n2698));
AND2X1 exu_U14550(.A(exu_n15721), .B(shft_shift16_e[0]), .Y(exu_n26754));
INVX1 exu_U14551(.A(exu_n26754), .Y(exu_n2699));
AND2X1 exu_U14552(.A(exu_n15722), .B(shft_shift16_e[0]), .Y(exu_n26758));
INVX1 exu_U14553(.A(exu_n26758), .Y(exu_n2700));
INVX1 exu_U14554(.A(exu_n2705), .Y(exu_n2701));
INVX1 exu_U14555(.A(exu_n2701), .Y(exu_n2702));
AND2X1 exu_U14556(.A(exu_n15723), .B(exu_n16148), .Y(exu_n26762));
INVX1 exu_U14557(.A(exu_n26762), .Y(exu_n2703));
INVX1 exu_U14558(.A(exu_n2708), .Y(exu_n2704));
INVX1 exu_U14559(.A(exu_n2704), .Y(exu_n2705));
AND2X1 exu_U14560(.A(exu_n15724), .B(shft_shift16_e[0]), .Y(exu_n26766));
INVX1 exu_U14561(.A(exu_n26766), .Y(exu_n2706));
INVX1 exu_U14562(.A(exu_n2712), .Y(exu_n2707));
INVX1 exu_U14563(.A(exu_n2707), .Y(exu_n2708));
AND2X1 exu_U14564(.A(exu_n15445), .B(exu_n16145), .Y(exu_n26770));
INVX1 exu_U14565(.A(exu_n26770), .Y(exu_n2709));
AND2X1 exu_U14566(.A(exu_n15725), .B(exu_n16148), .Y(exu_n26774));
INVX1 exu_U14567(.A(exu_n26774), .Y(exu_n2710));
INVX1 exu_U14568(.A(exu_n2715), .Y(exu_n2711));
INVX1 exu_U14569(.A(exu_n2711), .Y(exu_n2712));
AND2X1 exu_U14570(.A(exu_n15726), .B(exu_n16148), .Y(exu_n26778));
INVX1 exu_U14571(.A(exu_n26778), .Y(exu_n2713));
INVX1 exu_U14572(.A(exu_n2718), .Y(exu_n2714));
INVX1 exu_U14573(.A(exu_n2714), .Y(exu_n2715));
AND2X1 exu_U14574(.A(exu_n15694), .B(shft_shift16_e[0]), .Y(exu_n26782));
INVX1 exu_U14575(.A(exu_n26782), .Y(exu_n2716));
INVX1 exu_U14576(.A(exu_n2721), .Y(exu_n2717));
INVX1 exu_U14577(.A(exu_n2717), .Y(exu_n2718));
AND2X1 exu_U14578(.A(exu_n15727), .B(shft_shift16_e[0]), .Y(exu_n26786));
INVX1 exu_U14579(.A(exu_n26786), .Y(exu_n2719));
INVX1 exu_U14580(.A(exu_n2724), .Y(exu_n2720));
INVX1 exu_U14581(.A(exu_n2720), .Y(exu_n2721));
AND2X1 exu_U14582(.A(exu_n15728), .B(shft_shift16_e[0]), .Y(exu_n26790));
INVX1 exu_U14583(.A(exu_n26790), .Y(exu_n2722));
INVX1 exu_U14584(.A(exu_n2727), .Y(exu_n2723));
INVX1 exu_U14585(.A(exu_n2723), .Y(exu_n2724));
AND2X1 exu_U14586(.A(exu_n15729), .B(shft_shift16_e[0]), .Y(exu_n26794));
INVX1 exu_U14587(.A(exu_n26794), .Y(exu_n2725));
INVX1 exu_U14588(.A(exu_n2730), .Y(exu_n2726));
INVX1 exu_U14589(.A(exu_n2726), .Y(exu_n2727));
AND2X1 exu_U14590(.A(exu_n15730), .B(shft_shift16_e[0]), .Y(exu_n26798));
INVX1 exu_U14591(.A(exu_n26798), .Y(exu_n2728));
INVX1 exu_U14592(.A(exu_n2733), .Y(exu_n2729));
INVX1 exu_U14593(.A(exu_n2729), .Y(exu_n2730));
AND2X1 exu_U14594(.A(exu_n15731), .B(shft_shift16_e[0]), .Y(exu_n26802));
INVX1 exu_U14595(.A(exu_n26802), .Y(exu_n2731));
INVX1 exu_U14596(.A(exu_n2736), .Y(exu_n2732));
INVX1 exu_U14597(.A(exu_n2732), .Y(exu_n2733));
AND2X1 exu_U14598(.A(exu_n15732), .B(shft_shift16_e[0]), .Y(exu_n26806));
INVX1 exu_U14599(.A(exu_n26806), .Y(exu_n2734));
INVX1 exu_U14600(.A(exu_n2739), .Y(exu_n2735));
INVX1 exu_U14601(.A(exu_n2735), .Y(exu_n2736));
AND2X1 exu_U14602(.A(exu_n15733), .B(shft_shift16_e[0]), .Y(exu_n26810));
INVX1 exu_U14603(.A(exu_n26810), .Y(exu_n2737));
INVX1 exu_U14604(.A(exu_n2743), .Y(exu_n2738));
INVX1 exu_U14605(.A(exu_n2738), .Y(exu_n2739));
AND2X1 exu_U14606(.A(exu_n15446), .B(exu_n16145), .Y(exu_n26814));
INVX1 exu_U14607(.A(exu_n26814), .Y(exu_n2740));
AND2X1 exu_U14608(.A(exu_n15734), .B(shft_shift16_e[0]), .Y(exu_n26818));
INVX1 exu_U14609(.A(exu_n26818), .Y(exu_n2741));
INVX1 exu_U14610(.A(exu_n2746), .Y(exu_n2742));
INVX1 exu_U14611(.A(exu_n2742), .Y(exu_n2743));
AND2X1 exu_U14612(.A(exu_n15735), .B(shft_shift16_e[0]), .Y(exu_n26822));
INVX1 exu_U14613(.A(exu_n26822), .Y(exu_n2744));
INVX1 exu_U14614(.A(exu_n2749), .Y(exu_n2745));
INVX1 exu_U14615(.A(exu_n2745), .Y(exu_n2746));
AND2X1 exu_U14616(.A(exu_n15450), .B(shft_shift16_e[0]), .Y(exu_n26827));
INVX1 exu_U14617(.A(exu_n26827), .Y(exu_n2747));
INVX1 exu_U14618(.A(exu_n2766), .Y(exu_n2748));
INVX1 exu_U14619(.A(exu_n2748), .Y(exu_n2749));
AND2X1 exu_U14620(.A(exu_n15451), .B(exu_n16148), .Y(exu_n26832));
INVX1 exu_U14621(.A(exu_n26832), .Y(exu_n2750));
AND2X1 exu_U14622(.A(exu_n15452), .B(shft_shift16_e[0]), .Y(exu_n26837));
INVX1 exu_U14623(.A(exu_n26837), .Y(exu_n2751));
AND2X1 exu_U14624(.A(exu_n15453), .B(exu_n16148), .Y(exu_n26842));
INVX1 exu_U14625(.A(exu_n26842), .Y(exu_n2752));
AND2X1 exu_U14626(.A(exu_n15454), .B(exu_n16148), .Y(exu_n26847));
INVX1 exu_U14627(.A(exu_n26847), .Y(exu_n2753));
AND2X1 exu_U14628(.A(exu_n15455), .B(exu_n16148), .Y(exu_n26852));
INVX1 exu_U14629(.A(exu_n26852), .Y(exu_n2754));
AND2X1 exu_U14630(.A(exu_n15438), .B(shft_shift16_e[0]), .Y(exu_n26857));
INVX1 exu_U14631(.A(exu_n26857), .Y(exu_n2755));
AND2X1 exu_U14632(.A(exu_n15442), .B(exu_n16148), .Y(exu_n26862));
INVX1 exu_U14633(.A(exu_n26862), .Y(exu_n2756));
AND2X1 exu_U14634(.A(exu_n15447), .B(exu_n16145), .Y(exu_n26867));
INVX1 exu_U14635(.A(exu_n26867), .Y(exu_n2757));
AND2X1 exu_U14636(.A(exu_n15443), .B(exu_n16148), .Y(exu_n26871));
INVX1 exu_U14637(.A(exu_n26871), .Y(exu_n2758));
AND2X1 exu_U14638(.A(exu_n15444), .B(shft_shift16_e[0]), .Y(exu_n26876));
INVX1 exu_U14639(.A(exu_n26876), .Y(exu_n2759));
AND2X1 exu_U14640(.A(exu_n15445), .B(shft_shift16_e[0]), .Y(exu_n26881));
INVX1 exu_U14641(.A(exu_n26881), .Y(exu_n2760));
AND2X1 exu_U14642(.A(exu_n15446), .B(shft_shift16_e[0]), .Y(exu_n26886));
INVX1 exu_U14643(.A(exu_n26886), .Y(exu_n2761));
AND2X1 exu_U14644(.A(exu_n15447), .B(exu_n16148), .Y(exu_n26891));
INVX1 exu_U14645(.A(exu_n26891), .Y(exu_n2762));
AND2X1 exu_U14646(.A(exu_n15448), .B(exu_n16148), .Y(exu_n26896));
INVX1 exu_U14647(.A(exu_n26896), .Y(exu_n2763));
AND2X1 exu_U14648(.A(exu_n15449), .B(shft_shift16_e[0]), .Y(exu_n26901));
INVX1 exu_U14649(.A(exu_n26901), .Y(exu_n2764));
AND2X1 exu_U14650(.A(exu_n15456), .B(exu_n16148), .Y(exu_n26906));
INVX1 exu_U14651(.A(exu_n26906), .Y(exu_n2765));
AND2X1 exu_U14652(.A(exu_n16189), .B(exu_n16145), .Y(exu_n26908));
INVX1 exu_U14653(.A(exu_n26908), .Y(exu_n2766));
AND2X1 exu_U14654(.A(exu_n15721), .B(exu_n16145), .Y(exu_n26913));
INVX1 exu_U14655(.A(exu_n26913), .Y(exu_n2767));
AND2X1 exu_U14656(.A(exu_n15722), .B(exu_n16145), .Y(exu_n26917));
INVX1 exu_U14657(.A(exu_n26917), .Y(exu_n2768));
AND2X1 exu_U14658(.A(exu_n15448), .B(exu_n16145), .Y(exu_n26920));
INVX1 exu_U14659(.A(exu_n26920), .Y(exu_n2769));
AND2X1 exu_U14660(.A(exu_n15723), .B(exu_n16145), .Y(exu_n26925));
INVX1 exu_U14661(.A(exu_n26925), .Y(exu_n2770));
AND2X1 exu_U14662(.A(exu_n15724), .B(exu_n16145), .Y(exu_n26929));
INVX1 exu_U14663(.A(exu_n26929), .Y(exu_n2771));
AND2X1 exu_U14664(.A(exu_n15725), .B(exu_n16145), .Y(exu_n26933));
INVX1 exu_U14665(.A(exu_n26933), .Y(exu_n2772));
AND2X1 exu_U14666(.A(exu_n15726), .B(exu_n16145), .Y(exu_n26937));
INVX1 exu_U14667(.A(exu_n26937), .Y(exu_n2773));
AND2X1 exu_U14668(.A(exu_n15694), .B(exu_n16145), .Y(exu_n26941));
INVX1 exu_U14669(.A(exu_n26941), .Y(exu_n2774));
AND2X1 exu_U14670(.A(exu_n15727), .B(exu_n16145), .Y(exu_n26945));
INVX1 exu_U14671(.A(exu_n26945), .Y(exu_n2775));
AND2X1 exu_U14672(.A(exu_n15728), .B(exu_n16145), .Y(exu_n26949));
INVX1 exu_U14673(.A(exu_n26949), .Y(exu_n2776));
AND2X1 exu_U14674(.A(exu_n15729), .B(exu_n16145), .Y(exu_n26953));
INVX1 exu_U14675(.A(exu_n26953), .Y(exu_n2777));
AND2X1 exu_U14676(.A(exu_n15730), .B(exu_n16145), .Y(exu_n26957));
INVX1 exu_U14677(.A(exu_n26957), .Y(exu_n2778));
AND2X1 exu_U14678(.A(exu_n15731), .B(exu_n16145), .Y(exu_n26961));
INVX1 exu_U14679(.A(exu_n26961), .Y(exu_n2779));
AND2X1 exu_U14680(.A(exu_n15449), .B(exu_n16145), .Y(exu_n26964));
INVX1 exu_U14681(.A(exu_n26964), .Y(exu_n2780));
AND2X1 exu_U14682(.A(exu_n15732), .B(exu_n16145), .Y(exu_n26969));
INVX1 exu_U14683(.A(exu_n26969), .Y(exu_n2781));
AND2X1 exu_U14684(.A(exu_n15733), .B(exu_n16145), .Y(exu_n26973));
INVX1 exu_U14685(.A(exu_n26973), .Y(exu_n2782));
AND2X1 exu_U14686(.A(exu_n15734), .B(exu_n16145), .Y(exu_n26977));
INVX1 exu_U14687(.A(exu_n26977), .Y(exu_n2783));
AND2X1 exu_U14688(.A(exu_n15735), .B(exu_n16145), .Y(exu_n26981));
INVX1 exu_U14689(.A(exu_n26981), .Y(exu_n2784));
AND2X1 exu_U14690(.A(exu_n15450), .B(exu_n16145), .Y(exu_n26985));
INVX1 exu_U14691(.A(exu_n26985), .Y(exu_n2785));
AND2X1 exu_U14692(.A(exu_n15451), .B(exu_n16145), .Y(exu_n26989));
INVX1 exu_U14693(.A(exu_n26989), .Y(exu_n2786));
AND2X1 exu_U14694(.A(exu_n15452), .B(exu_n16145), .Y(exu_n26993));
INVX1 exu_U14695(.A(exu_n26993), .Y(exu_n2787));
AND2X1 exu_U14696(.A(exu_n15453), .B(exu_n16145), .Y(exu_n26997));
INVX1 exu_U14697(.A(exu_n26997), .Y(exu_n2788));
AND2X1 exu_U14698(.A(exu_n15454), .B(exu_n16145), .Y(exu_n27001));
INVX1 exu_U14699(.A(exu_n27001), .Y(exu_n2789));
AND2X1 exu_U14700(.A(exu_n15455), .B(exu_n16145), .Y(exu_n27005));
INVX1 exu_U14701(.A(exu_n27005), .Y(exu_n2790));
AND2X1 exu_U14702(.A(exu_n15456), .B(exu_n16145), .Y(exu_n27009));
INVX1 exu_U14703(.A(exu_n27009), .Y(exu_n2791));
AND2X1 exu_U14704(.A(exu_n16230), .B(shft_rshift16_b1[9]), .Y(exu_n27013));
INVX1 exu_U14705(.A(exu_n27013), .Y(exu_n2792));
AND2X1 exu_U14706(.A(exu_n16232), .B(shft_rshift16_b1[17]), .Y(exu_n27015));
INVX1 exu_U14707(.A(exu_n27015), .Y(exu_n2793));
AND2X1 exu_U14708(.A(shft_rshift16_b1[8]), .B(exu_n16230), .Y(exu_n27019));
INVX1 exu_U14709(.A(exu_n27019), .Y(exu_n2794));
AND2X1 exu_U14710(.A(shft_rshift16_b1[16]), .B(exu_n16233), .Y(exu_n27021));
INVX1 exu_U14711(.A(exu_n27021), .Y(exu_n2795));
AND2X1 exu_U14712(.A(shft_rshift16_b1[7]), .B(exu_n16230), .Y(exu_n27025));
INVX1 exu_U14713(.A(exu_n27025), .Y(exu_n2796));
AND2X1 exu_U14714(.A(shft_rshift16_b1[15]), .B(exu_n16233), .Y(exu_n27027));
INVX1 exu_U14715(.A(exu_n27027), .Y(exu_n2797));
AND2X1 exu_U14716(.A(shft_rshift16_b1[6]), .B(exu_n16230), .Y(exu_n27031));
INVX1 exu_U14717(.A(exu_n27031), .Y(exu_n2798));
AND2X1 exu_U14718(.A(shft_rshift16_b1[14]), .B(exu_n16233), .Y(exu_n27033));
INVX1 exu_U14719(.A(exu_n27033), .Y(exu_n2799));
AND2X1 exu_U14720(.A(shft_rshift16_b1[63]), .B(exu_n16230), .Y(exu_n27036));
INVX1 exu_U14721(.A(exu_n27036), .Y(exu_n2800));
AND2X1 exu_U14722(.A(shft_rshift16_b1[62]), .B(exu_n16230), .Y(exu_n27039));
INVX1 exu_U14723(.A(exu_n27039), .Y(exu_n2801));
AND2X1 exu_U14724(.A(shft_rshift16_b1[61]), .B(exu_n16230), .Y(exu_n27042));
INVX1 exu_U14725(.A(exu_n27042), .Y(exu_n2802));
AND2X1 exu_U14726(.A(shft_rshift16_b1[60]), .B(exu_n16230), .Y(exu_n27045));
INVX1 exu_U14727(.A(exu_n27045), .Y(exu_n2803));
AND2X1 exu_U14728(.A(shft_rshift16_b1[5]), .B(exu_n16230), .Y(exu_n27050));
INVX1 exu_U14729(.A(exu_n27050), .Y(exu_n2804));
AND2X1 exu_U14730(.A(shft_rshift16_b1[13]), .B(exu_n16233), .Y(exu_n27052));
INVX1 exu_U14731(.A(exu_n27052), .Y(exu_n2805));
AND2X1 exu_U14732(.A(shft_rshift16_b1[59]), .B(exu_n16230), .Y(exu_n27056));
INVX1 exu_U14733(.A(exu_n27056), .Y(exu_n2806));
AND2X1 exu_U14734(.A(shft_rshift16_b1[58]), .B(exu_n16230), .Y(exu_n27061));
INVX1 exu_U14735(.A(exu_n27061), .Y(exu_n2807));
AND2X1 exu_U14736(.A(shft_rshift16_b1[57]), .B(exu_n16230), .Y(exu_n27065));
INVX1 exu_U14737(.A(exu_n27065), .Y(exu_n2808));
AND2X1 exu_U14738(.A(shft_rshift16_b1[56]), .B(exu_n16230), .Y(exu_n27069));
INVX1 exu_U14739(.A(exu_n27069), .Y(exu_n2809));
AND2X1 exu_U14740(.A(exu_n15403), .B(exu_n16232), .Y(exu_n27071));
INVX1 exu_U14741(.A(exu_n27071), .Y(exu_n2810));
AND2X1 exu_U14742(.A(shft_rshift16_b1[55]), .B(exu_n15401), .Y(exu_n27074));
INVX1 exu_U14743(.A(exu_n27074), .Y(exu_n2811));
AND2X1 exu_U14744(.A(shft_rshift16_b1[63]), .B(exu_n16233), .Y(exu_n27076));
INVX1 exu_U14745(.A(exu_n27076), .Y(exu_n2812));
AND2X1 exu_U14746(.A(shft_rshift16_b1[54]), .B(exu_n15401), .Y(exu_n27079));
INVX1 exu_U14747(.A(exu_n27079), .Y(exu_n2813));
AND2X1 exu_U14748(.A(shft_rshift16_b1[62]), .B(exu_n16233), .Y(exu_n27081));
INVX1 exu_U14749(.A(exu_n27081), .Y(exu_n2814));
AND2X1 exu_U14750(.A(shft_rshift16_b1[53]), .B(exu_n15401), .Y(exu_n27084));
INVX1 exu_U14751(.A(exu_n27084), .Y(exu_n2815));
AND2X1 exu_U14752(.A(shft_rshift16_b1[61]), .B(exu_n16232), .Y(exu_n27086));
INVX1 exu_U14753(.A(exu_n27086), .Y(exu_n2816));
AND2X1 exu_U14754(.A(shft_rshift16_b1[52]), .B(exu_n16230), .Y(exu_n27089));
INVX1 exu_U14755(.A(exu_n27089), .Y(exu_n2817));
AND2X1 exu_U14756(.A(shft_rshift16_b1[60]), .B(exu_n16232), .Y(exu_n27091));
INVX1 exu_U14757(.A(exu_n27091), .Y(exu_n2818));
AND2X1 exu_U14758(.A(shft_rshift16_b1[51]), .B(exu_n16230), .Y(exu_n27094));
INVX1 exu_U14759(.A(exu_n27094), .Y(exu_n2819));
AND2X1 exu_U14760(.A(shft_rshift16_b1[59]), .B(exu_n16233), .Y(exu_n27096));
INVX1 exu_U14761(.A(exu_n27096), .Y(exu_n2820));
AND2X1 exu_U14762(.A(shft_rshift16_b1[50]), .B(exu_n15401), .Y(exu_n27100));
INVX1 exu_U14763(.A(exu_n27100), .Y(exu_n2821));
AND2X1 exu_U14764(.A(shft_rshift16_b1[58]), .B(exu_n16233), .Y(exu_n27102));
INVX1 exu_U14765(.A(exu_n27102), .Y(exu_n2822));
AND2X1 exu_U14766(.A(shft_rshift16_b1[4]), .B(exu_n16230), .Y(exu_n27106));
INVX1 exu_U14767(.A(exu_n27106), .Y(exu_n2823));
AND2X1 exu_U14768(.A(shft_rshift16_b1[12]), .B(exu_n16233), .Y(exu_n27108));
INVX1 exu_U14769(.A(exu_n27108), .Y(exu_n2824));
AND2X1 exu_U14770(.A(shft_rshift16_b1[49]), .B(exu_n16230), .Y(exu_n27112));
INVX1 exu_U14771(.A(exu_n27112), .Y(exu_n2825));
AND2X1 exu_U14772(.A(shft_rshift16_b1[57]), .B(exu_n16232), .Y(exu_n27114));
INVX1 exu_U14773(.A(exu_n27114), .Y(exu_n2826));
AND2X1 exu_U14774(.A(shft_rshift16_b1[48]), .B(exu_n15401), .Y(exu_n27118));
INVX1 exu_U14775(.A(exu_n27118), .Y(exu_n2827));
AND2X1 exu_U14776(.A(shft_rshift16_b1[56]), .B(exu_n16232), .Y(exu_n27120));
INVX1 exu_U14777(.A(exu_n27120), .Y(exu_n2828));
AND2X1 exu_U14778(.A(shft_rshift16_b1[47]), .B(exu_n15401), .Y(exu_n27124));
INVX1 exu_U14779(.A(exu_n27124), .Y(exu_n2829));
AND2X1 exu_U14780(.A(shft_rshift16_b1[55]), .B(exu_n16232), .Y(exu_n27126));
INVX1 exu_U14781(.A(exu_n27126), .Y(exu_n2830));
AND2X1 exu_U14782(.A(shft_rshift16_b1[46]), .B(exu_n15401), .Y(exu_n27130));
INVX1 exu_U14783(.A(exu_n27130), .Y(exu_n2831));
AND2X1 exu_U14784(.A(shft_rshift16_b1[54]), .B(exu_n16233), .Y(exu_n27132));
INVX1 exu_U14785(.A(exu_n27132), .Y(exu_n2832));
AND2X1 exu_U14786(.A(shft_rshift16_b1[45]), .B(exu_n15401), .Y(exu_n27136));
INVX1 exu_U14787(.A(exu_n27136), .Y(exu_n2833));
AND2X1 exu_U14788(.A(shft_rshift16_b1[53]), .B(exu_n16232), .Y(exu_n27138));
INVX1 exu_U14789(.A(exu_n27138), .Y(exu_n2834));
AND2X1 exu_U14790(.A(shft_rshift16_b1[44]), .B(exu_n16230), .Y(exu_n27142));
INVX1 exu_U14791(.A(exu_n27142), .Y(exu_n2835));
AND2X1 exu_U14792(.A(shft_rshift16_b1[52]), .B(exu_n16232), .Y(exu_n27144));
INVX1 exu_U14793(.A(exu_n27144), .Y(exu_n2836));
AND2X1 exu_U14794(.A(shft_rshift16_b1[43]), .B(exu_n16230), .Y(exu_n27148));
INVX1 exu_U14795(.A(exu_n27148), .Y(exu_n2837));
AND2X1 exu_U14796(.A(shft_rshift16_b1[51]), .B(exu_n16233), .Y(exu_n27150));
INVX1 exu_U14797(.A(exu_n27150), .Y(exu_n2838));
AND2X1 exu_U14798(.A(shft_rshift16_b1[42]), .B(exu_n15401), .Y(exu_n27154));
INVX1 exu_U14799(.A(exu_n27154), .Y(exu_n2839));
AND2X1 exu_U14800(.A(shft_rshift16_b1[50]), .B(exu_n16233), .Y(exu_n27156));
INVX1 exu_U14801(.A(exu_n27156), .Y(exu_n2840));
AND2X1 exu_U14802(.A(shft_rshift16_b1[41]), .B(exu_n15401), .Y(exu_n27160));
INVX1 exu_U14803(.A(exu_n27160), .Y(exu_n2841));
AND2X1 exu_U14804(.A(shft_rshift16_b1[49]), .B(exu_n16233), .Y(exu_n27162));
INVX1 exu_U14805(.A(exu_n27162), .Y(exu_n2842));
AND2X1 exu_U14806(.A(shft_rshift16_b1[40]), .B(exu_n16230), .Y(exu_n27166));
INVX1 exu_U14807(.A(exu_n27166), .Y(exu_n2843));
AND2X1 exu_U14808(.A(shft_rshift16_b1[48]), .B(exu_n16233), .Y(exu_n27168));
INVX1 exu_U14809(.A(exu_n27168), .Y(exu_n2844));
AND2X1 exu_U14810(.A(shft_rshift16_b1[3]), .B(exu_n15401), .Y(exu_n27172));
INVX1 exu_U14811(.A(exu_n27172), .Y(exu_n2845));
AND2X1 exu_U14812(.A(shft_rshift16_b1[11]), .B(exu_n16232), .Y(exu_n27174));
INVX1 exu_U14813(.A(exu_n27174), .Y(exu_n2846));
AND2X1 exu_U14814(.A(shft_rshift16_b1[39]), .B(exu_n15401), .Y(exu_n27178));
INVX1 exu_U14815(.A(exu_n27178), .Y(exu_n2847));
AND2X1 exu_U14816(.A(shft_rshift16_b1[47]), .B(exu_n16232), .Y(exu_n27180));
INVX1 exu_U14817(.A(exu_n27180), .Y(exu_n2848));
AND2X1 exu_U14818(.A(shft_rshift16_b1[38]), .B(exu_n16230), .Y(exu_n27184));
INVX1 exu_U14819(.A(exu_n27184), .Y(exu_n2849));
AND2X1 exu_U14820(.A(shft_rshift16_b1[46]), .B(exu_n16233), .Y(exu_n27186));
INVX1 exu_U14821(.A(exu_n27186), .Y(exu_n2850));
AND2X1 exu_U14822(.A(shft_rshift16_b1[37]), .B(exu_n16230), .Y(exu_n27190));
INVX1 exu_U14823(.A(exu_n27190), .Y(exu_n2851));
AND2X1 exu_U14824(.A(shft_rshift16_b1[45]), .B(exu_n16233), .Y(exu_n27192));
INVX1 exu_U14825(.A(exu_n27192), .Y(exu_n2852));
AND2X1 exu_U14826(.A(shft_rshift16_b1[36]), .B(exu_n16230), .Y(exu_n27196));
INVX1 exu_U14827(.A(exu_n27196), .Y(exu_n2853));
AND2X1 exu_U14828(.A(shft_rshift16_b1[44]), .B(exu_n16233), .Y(exu_n27198));
INVX1 exu_U14829(.A(exu_n27198), .Y(exu_n2854));
AND2X1 exu_U14830(.A(shft_rshift16_b1[35]), .B(exu_n15401), .Y(exu_n27202));
INVX1 exu_U14831(.A(exu_n27202), .Y(exu_n2855));
AND2X1 exu_U14832(.A(shft_rshift16_b1[43]), .B(exu_n16233), .Y(exu_n27204));
INVX1 exu_U14833(.A(exu_n27204), .Y(exu_n2856));
AND2X1 exu_U14834(.A(shft_rshift16_b1[34]), .B(exu_n16230), .Y(exu_n27208));
INVX1 exu_U14835(.A(exu_n27208), .Y(exu_n2857));
AND2X1 exu_U14836(.A(shft_rshift16_b1[42]), .B(exu_n16232), .Y(exu_n27210));
INVX1 exu_U14837(.A(exu_n27210), .Y(exu_n2858));
AND2X1 exu_U14838(.A(shft_rshift16_b1[33]), .B(exu_n16230), .Y(exu_n27214));
INVX1 exu_U14839(.A(exu_n27214), .Y(exu_n2859));
AND2X1 exu_U14840(.A(shft_rshift16_b1[41]), .B(exu_n16233), .Y(exu_n27216));
INVX1 exu_U14841(.A(exu_n27216), .Y(exu_n2860));
AND2X1 exu_U14842(.A(shft_rshift16_b1[32]), .B(exu_n15401), .Y(exu_n27220));
INVX1 exu_U14843(.A(exu_n27220), .Y(exu_n2861));
AND2X1 exu_U14844(.A(shft_rshift16_b1[40]), .B(exu_n16233), .Y(exu_n27222));
INVX1 exu_U14845(.A(exu_n27222), .Y(exu_n2862));
AND2X1 exu_U14846(.A(shft_rshift16_b1[31]), .B(exu_n16230), .Y(exu_n27226));
INVX1 exu_U14847(.A(exu_n27226), .Y(exu_n2863));
AND2X1 exu_U14848(.A(shft_rshift16_b1[39]), .B(exu_n16232), .Y(exu_n27228));
INVX1 exu_U14849(.A(exu_n27228), .Y(exu_n2864));
AND2X1 exu_U14850(.A(shft_rshift16_b1[30]), .B(exu_n15401), .Y(exu_n27232));
INVX1 exu_U14851(.A(exu_n27232), .Y(exu_n2865));
AND2X1 exu_U14852(.A(shft_rshift16_b1[38]), .B(exu_n16232), .Y(exu_n27234));
INVX1 exu_U14853(.A(exu_n27234), .Y(exu_n2866));
AND2X1 exu_U14854(.A(shft_rshift16_b1[2]), .B(exu_n16230), .Y(exu_n27238));
INVX1 exu_U14855(.A(exu_n27238), .Y(exu_n2867));
AND2X1 exu_U14856(.A(shft_rshift16_b1[10]), .B(exu_n16232), .Y(exu_n27240));
INVX1 exu_U14857(.A(exu_n27240), .Y(exu_n2868));
AND2X1 exu_U14858(.A(shft_rshift16_b1[29]), .B(exu_n16230), .Y(exu_n27244));
INVX1 exu_U14859(.A(exu_n27244), .Y(exu_n2869));
AND2X1 exu_U14860(.A(shft_rshift16_b1[37]), .B(exu_n16233), .Y(exu_n27246));
INVX1 exu_U14861(.A(exu_n27246), .Y(exu_n2870));
AND2X1 exu_U14862(.A(shft_rshift16_b1[28]), .B(exu_n15401), .Y(exu_n27250));
INVX1 exu_U14863(.A(exu_n27250), .Y(exu_n2871));
AND2X1 exu_U14864(.A(shft_rshift16_b1[36]), .B(exu_n16232), .Y(exu_n27252));
INVX1 exu_U14865(.A(exu_n27252), .Y(exu_n2872));
AND2X1 exu_U14866(.A(shft_rshift16_b1[27]), .B(exu_n16230), .Y(exu_n27256));
INVX1 exu_U14867(.A(exu_n27256), .Y(exu_n2873));
AND2X1 exu_U14868(.A(shft_rshift16_b1[35]), .B(exu_n16232), .Y(exu_n27258));
INVX1 exu_U14869(.A(exu_n27258), .Y(exu_n2874));
AND2X1 exu_U14870(.A(shft_rshift16_b1[26]), .B(exu_n15401), .Y(exu_n27262));
INVX1 exu_U14871(.A(exu_n27262), .Y(exu_n2875));
AND2X1 exu_U14872(.A(shft_rshift16_b1[34]), .B(exu_n16233), .Y(exu_n27264));
INVX1 exu_U14873(.A(exu_n27264), .Y(exu_n2876));
AND2X1 exu_U14874(.A(shft_rshift16_b1[25]), .B(exu_n15401), .Y(exu_n27268));
INVX1 exu_U14875(.A(exu_n27268), .Y(exu_n2877));
AND2X1 exu_U14876(.A(shft_rshift16_b1[33]), .B(exu_n16233), .Y(exu_n27270));
INVX1 exu_U14877(.A(exu_n27270), .Y(exu_n2878));
AND2X1 exu_U14878(.A(shft_rshift16_b1[24]), .B(exu_n16230), .Y(exu_n27274));
INVX1 exu_U14879(.A(exu_n27274), .Y(exu_n2879));
AND2X1 exu_U14880(.A(shft_rshift16_b1[32]), .B(exu_n16232), .Y(exu_n27276));
INVX1 exu_U14881(.A(exu_n27276), .Y(exu_n2880));
AND2X1 exu_U14882(.A(shft_rshift16_b1[23]), .B(exu_n15401), .Y(exu_n27280));
INVX1 exu_U14883(.A(exu_n27280), .Y(exu_n2881));
AND2X1 exu_U14884(.A(shft_rshift16_b1[31]), .B(exu_n16232), .Y(exu_n27282));
INVX1 exu_U14885(.A(exu_n27282), .Y(exu_n2882));
AND2X1 exu_U14886(.A(shft_rshift16_b1[22]), .B(exu_n15401), .Y(exu_n27286));
INVX1 exu_U14887(.A(exu_n27286), .Y(exu_n2883));
AND2X1 exu_U14888(.A(shft_rshift16_b1[30]), .B(exu_n16232), .Y(exu_n27288));
INVX1 exu_U14889(.A(exu_n27288), .Y(exu_n2884));
AND2X1 exu_U14890(.A(shft_rshift16_b1[21]), .B(exu_n15401), .Y(exu_n27292));
INVX1 exu_U14891(.A(exu_n27292), .Y(exu_n2885));
AND2X1 exu_U14892(.A(shft_rshift16_b1[29]), .B(exu_n16232), .Y(exu_n27294));
INVX1 exu_U14893(.A(exu_n27294), .Y(exu_n2886));
AND2X1 exu_U14894(.A(shft_rshift16_b1[20]), .B(exu_n16230), .Y(exu_n27298));
INVX1 exu_U14895(.A(exu_n27298), .Y(exu_n2887));
AND2X1 exu_U14896(.A(shft_rshift16_b1[28]), .B(exu_n16232), .Y(exu_n27300));
INVX1 exu_U14897(.A(exu_n27300), .Y(exu_n2888));
AND2X1 exu_U14898(.A(shft_rshift16_b1[1]), .B(exu_n15401), .Y(exu_n27304));
INVX1 exu_U14899(.A(exu_n27304), .Y(exu_n2889));
AND2X1 exu_U14900(.A(shft_rshift16_b1[9]), .B(exu_n16232), .Y(exu_n27306));
INVX1 exu_U14901(.A(exu_n27306), .Y(exu_n2890));
AND2X1 exu_U14902(.A(shft_rshift16_b1[19]), .B(exu_n15401), .Y(exu_n27310));
INVX1 exu_U14903(.A(exu_n27310), .Y(exu_n2891));
AND2X1 exu_U14904(.A(shft_rshift16_b1[27]), .B(exu_n16232), .Y(exu_n27312));
INVX1 exu_U14905(.A(exu_n27312), .Y(exu_n2892));
AND2X1 exu_U14906(.A(shft_rshift16_b1[18]), .B(exu_n15401), .Y(exu_n27316));
INVX1 exu_U14907(.A(exu_n27316), .Y(exu_n2893));
AND2X1 exu_U14908(.A(shft_rshift16_b1[26]), .B(exu_n16232), .Y(exu_n27318));
INVX1 exu_U14909(.A(exu_n27318), .Y(exu_n2894));
AND2X1 exu_U14910(.A(shft_rshift16_b1[17]), .B(exu_n15401), .Y(exu_n27322));
INVX1 exu_U14911(.A(exu_n27322), .Y(exu_n2895));
AND2X1 exu_U14912(.A(shft_rshift16_b1[25]), .B(exu_n16232), .Y(exu_n27324));
INVX1 exu_U14913(.A(exu_n27324), .Y(exu_n2896));
AND2X1 exu_U14914(.A(shft_rshift16_b1[16]), .B(exu_n16230), .Y(exu_n27328));
INVX1 exu_U14915(.A(exu_n27328), .Y(exu_n2897));
AND2X1 exu_U14916(.A(shft_rshift16_b1[24]), .B(exu_n16232), .Y(exu_n27330));
INVX1 exu_U14917(.A(exu_n27330), .Y(exu_n2898));
AND2X1 exu_U14918(.A(shft_rshift16_b1[15]), .B(exu_n15401), .Y(exu_n27334));
INVX1 exu_U14919(.A(exu_n27334), .Y(exu_n2899));
AND2X1 exu_U14920(.A(shft_rshift16_b1[23]), .B(exu_n16232), .Y(exu_n27336));
INVX1 exu_U14921(.A(exu_n27336), .Y(exu_n2900));
AND2X1 exu_U14922(.A(shft_rshift16_b1[14]), .B(exu_n15401), .Y(exu_n27340));
INVX1 exu_U14923(.A(exu_n27340), .Y(exu_n2901));
AND2X1 exu_U14924(.A(shft_rshift16_b1[22]), .B(exu_n16232), .Y(exu_n27342));
INVX1 exu_U14925(.A(exu_n27342), .Y(exu_n2902));
AND2X1 exu_U14926(.A(shft_rshift16_b1[13]), .B(exu_n15401), .Y(exu_n27346));
INVX1 exu_U14927(.A(exu_n27346), .Y(exu_n2903));
AND2X1 exu_U14928(.A(shft_rshift16_b1[21]), .B(exu_n16232), .Y(exu_n27348));
INVX1 exu_U14929(.A(exu_n27348), .Y(exu_n2904));
AND2X1 exu_U14930(.A(shft_rshift16_b1[12]), .B(exu_n16230), .Y(exu_n27352));
INVX1 exu_U14931(.A(exu_n27352), .Y(exu_n2905));
AND2X1 exu_U14932(.A(shft_rshift16_b1[20]), .B(exu_n16232), .Y(exu_n27354));
INVX1 exu_U14933(.A(exu_n27354), .Y(exu_n2906));
AND2X1 exu_U14934(.A(shft_rshift16_b1[11]), .B(exu_n15401), .Y(exu_n27358));
INVX1 exu_U14935(.A(exu_n27358), .Y(exu_n2907));
AND2X1 exu_U14936(.A(shft_rshift16_b1[19]), .B(exu_n16233), .Y(exu_n27360));
INVX1 exu_U14937(.A(exu_n27360), .Y(exu_n2908));
AND2X1 exu_U14938(.A(shft_rshift16_b1[10]), .B(exu_n15401), .Y(exu_n27364));
INVX1 exu_U14939(.A(exu_n27364), .Y(exu_n2909));
AND2X1 exu_U14940(.A(shft_rshift16_b1[18]), .B(exu_n16233), .Y(exu_n27366));
INVX1 exu_U14941(.A(exu_n27366), .Y(exu_n2910));
AND2X1 exu_U14942(.A(shft_rshift16_b1[0]), .B(exu_n16230), .Y(exu_n27370));
INVX1 exu_U14943(.A(exu_n27370), .Y(exu_n2911));
AND2X1 exu_U14944(.A(shft_rshift16_b1[8]), .B(exu_n16232), .Y(exu_n27372));
INVX1 exu_U14945(.A(exu_n27372), .Y(exu_n2912));
AND2X1 exu_U14946(.A(exu_n16224), .B(shft_rshift4_b1[9]), .Y(exu_n27376));
INVX1 exu_U14947(.A(exu_n27376), .Y(exu_n2913));
AND2X1 exu_U14948(.A(exu_n15402), .B(shft_rshift4_b1[11]), .Y(exu_n27378));
INVX1 exu_U14949(.A(exu_n27378), .Y(exu_n2914));
AND2X1 exu_U14950(.A(shft_rshift4_b1[8]), .B(exu_n16223), .Y(exu_n27382));
INVX1 exu_U14951(.A(exu_n27382), .Y(exu_n2915));
AND2X1 exu_U14952(.A(shft_rshift4_b1[10]), .B(exu_n16227), .Y(exu_n27384));
INVX1 exu_U14953(.A(exu_n27384), .Y(exu_n2916));
AND2X1 exu_U14954(.A(shft_rshift4_b1[7]), .B(exu_n16223), .Y(exu_n27388));
INVX1 exu_U14955(.A(exu_n27388), .Y(exu_n2917));
AND2X1 exu_U14956(.A(shft_rshift4_b1[9]), .B(exu_n15402), .Y(exu_n27390));
INVX1 exu_U14957(.A(exu_n27390), .Y(exu_n2918));
AND2X1 exu_U14958(.A(shft_rshift4_b1[6]), .B(exu_n16224), .Y(exu_n27394));
INVX1 exu_U14959(.A(exu_n27394), .Y(exu_n2919));
AND2X1 exu_U14960(.A(shft_rshift4_b1[8]), .B(exu_n15402), .Y(exu_n27396));
INVX1 exu_U14961(.A(exu_n27396), .Y(exu_n2920));
AND2X1 exu_U14962(.A(shft_rshift4_b1[63]), .B(exu_n16224), .Y(exu_n27400));
INVX1 exu_U14963(.A(exu_n27400), .Y(exu_n2921));
AND2X1 exu_U14964(.A(shft_rshift4_b1[62]), .B(exu_n16224), .Y(exu_n27403));
INVX1 exu_U14965(.A(exu_n27403), .Y(exu_n2922));
AND2X1 exu_U14966(.A(exu_n16191), .B(exu_n15402), .Y(exu_n27405));
INVX1 exu_U14967(.A(exu_n27405), .Y(exu_n2923));
AND2X1 exu_U14968(.A(shft_rshift4_b1[61]), .B(exu_n16224), .Y(exu_n27409));
INVX1 exu_U14969(.A(exu_n27409), .Y(exu_n2924));
AND2X1 exu_U14970(.A(shft_rshift4_b1[63]), .B(exu_n15402), .Y(exu_n27411));
INVX1 exu_U14971(.A(exu_n27411), .Y(exu_n2925));
AND2X1 exu_U14972(.A(shft_rshift4_b1[60]), .B(exu_n16224), .Y(exu_n27414));
INVX1 exu_U14973(.A(exu_n27414), .Y(exu_n2926));
AND2X1 exu_U14974(.A(shft_rshift4_b1[62]), .B(exu_n16227), .Y(exu_n27416));
INVX1 exu_U14975(.A(exu_n27416), .Y(exu_n2927));
AND2X1 exu_U14976(.A(shft_rshift4_b1[5]), .B(exu_n16224), .Y(exu_n27420));
INVX1 exu_U14977(.A(exu_n27420), .Y(exu_n2928));
AND2X1 exu_U14978(.A(shft_rshift4_b1[7]), .B(exu_n16227), .Y(exu_n27422));
INVX1 exu_U14979(.A(exu_n27422), .Y(exu_n2929));
AND2X1 exu_U14980(.A(shft_rshift4_b1[59]), .B(exu_n16224), .Y(exu_n27426));
INVX1 exu_U14981(.A(exu_n27426), .Y(exu_n2930));
AND2X1 exu_U14982(.A(shft_rshift4_b1[61]), .B(exu_n15402), .Y(exu_n27428));
INVX1 exu_U14983(.A(exu_n27428), .Y(exu_n2931));
AND2X1 exu_U14984(.A(shft_rshift4_b1[58]), .B(exu_n16224), .Y(exu_n27432));
INVX1 exu_U14985(.A(exu_n27432), .Y(exu_n2932));
AND2X1 exu_U14986(.A(shft_rshift4_b1[60]), .B(exu_n15402), .Y(exu_n27434));
INVX1 exu_U14987(.A(exu_n27434), .Y(exu_n2933));
AND2X1 exu_U14988(.A(shft_rshift4_b1[57]), .B(exu_n16223), .Y(exu_n27438));
INVX1 exu_U14989(.A(exu_n27438), .Y(exu_n2934));
AND2X1 exu_U14990(.A(shft_rshift4_b1[59]), .B(exu_n16227), .Y(exu_n27440));
INVX1 exu_U14991(.A(exu_n27440), .Y(exu_n2935));
AND2X1 exu_U14992(.A(shft_rshift4_b1[56]), .B(exu_n16224), .Y(exu_n27444));
INVX1 exu_U14993(.A(exu_n27444), .Y(exu_n2936));
AND2X1 exu_U14994(.A(shft_rshift4_b1[58]), .B(exu_n15402), .Y(exu_n27446));
INVX1 exu_U14995(.A(exu_n27446), .Y(exu_n2937));
AND2X1 exu_U14996(.A(shft_rshift4_b1[55]), .B(exu_n16223), .Y(exu_n27450));
INVX1 exu_U14997(.A(exu_n27450), .Y(exu_n2938));
AND2X1 exu_U14998(.A(shft_rshift4_b1[57]), .B(exu_n16227), .Y(exu_n27452));
INVX1 exu_U14999(.A(exu_n27452), .Y(exu_n2939));
AND2X1 exu_U15000(.A(shft_rshift4_b1[54]), .B(exu_n16224), .Y(exu_n27456));
INVX1 exu_U15001(.A(exu_n27456), .Y(exu_n2940));
AND2X1 exu_U15002(.A(shft_rshift4_b1[56]), .B(exu_n16227), .Y(exu_n27458));
INVX1 exu_U15003(.A(exu_n27458), .Y(exu_n2941));
AND2X1 exu_U15004(.A(shft_rshift4_b1[53]), .B(exu_n16223), .Y(exu_n27462));
INVX1 exu_U15005(.A(exu_n27462), .Y(exu_n2942));
AND2X1 exu_U15006(.A(shft_rshift4_b1[55]), .B(exu_n16227), .Y(exu_n27464));
INVX1 exu_U15007(.A(exu_n27464), .Y(exu_n2943));
AND2X1 exu_U15008(.A(shft_rshift4_b1[52]), .B(exu_n16223), .Y(exu_n27468));
INVX1 exu_U15009(.A(exu_n27468), .Y(exu_n2944));
AND2X1 exu_U15010(.A(shft_rshift4_b1[54]), .B(exu_n16227), .Y(exu_n27470));
INVX1 exu_U15011(.A(exu_n27470), .Y(exu_n2945));
AND2X1 exu_U15012(.A(shft_rshift4_b1[51]), .B(exu_n16223), .Y(exu_n27474));
INVX1 exu_U15013(.A(exu_n27474), .Y(exu_n2946));
AND2X1 exu_U15014(.A(shft_rshift4_b1[53]), .B(exu_n15402), .Y(exu_n27476));
INVX1 exu_U15015(.A(exu_n27476), .Y(exu_n2947));
AND2X1 exu_U15016(.A(shft_rshift4_b1[50]), .B(exu_n16223), .Y(exu_n27480));
INVX1 exu_U15017(.A(exu_n27480), .Y(exu_n2948));
AND2X1 exu_U15018(.A(shft_rshift4_b1[52]), .B(exu_n16227), .Y(exu_n27482));
INVX1 exu_U15019(.A(exu_n27482), .Y(exu_n2949));
AND2X1 exu_U15020(.A(shft_rshift4_b1[4]), .B(exu_n16223), .Y(exu_n27486));
INVX1 exu_U15021(.A(exu_n27486), .Y(exu_n2950));
AND2X1 exu_U15022(.A(shft_rshift4_b1[6]), .B(exu_n15402), .Y(exu_n27488));
INVX1 exu_U15023(.A(exu_n27488), .Y(exu_n2951));
AND2X1 exu_U15024(.A(shft_rshift4_b1[49]), .B(exu_n16224), .Y(exu_n27492));
INVX1 exu_U15025(.A(exu_n27492), .Y(exu_n2952));
AND2X1 exu_U15026(.A(shft_rshift4_b1[51]), .B(exu_n15402), .Y(exu_n27494));
INVX1 exu_U15027(.A(exu_n27494), .Y(exu_n2953));
AND2X1 exu_U15028(.A(shft_rshift4_b1[48]), .B(exu_n16223), .Y(exu_n27498));
INVX1 exu_U15029(.A(exu_n27498), .Y(exu_n2954));
AND2X1 exu_U15030(.A(shft_rshift4_b1[50]), .B(exu_n16227), .Y(exu_n27500));
INVX1 exu_U15031(.A(exu_n27500), .Y(exu_n2955));
AND2X1 exu_U15032(.A(shft_rshift4_b1[47]), .B(exu_n16224), .Y(exu_n27504));
INVX1 exu_U15033(.A(exu_n27504), .Y(exu_n2956));
AND2X1 exu_U15034(.A(shft_rshift4_b1[49]), .B(exu_n16227), .Y(exu_n27506));
INVX1 exu_U15035(.A(exu_n27506), .Y(exu_n2957));
AND2X1 exu_U15036(.A(shft_rshift4_b1[46]), .B(exu_n16223), .Y(exu_n27510));
INVX1 exu_U15037(.A(exu_n27510), .Y(exu_n2958));
AND2X1 exu_U15038(.A(shft_rshift4_b1[48]), .B(exu_n15402), .Y(exu_n27512));
INVX1 exu_U15039(.A(exu_n27512), .Y(exu_n2959));
AND2X1 exu_U15040(.A(shft_rshift4_b1[45]), .B(exu_n16224), .Y(exu_n27516));
INVX1 exu_U15041(.A(exu_n27516), .Y(exu_n2960));
AND2X1 exu_U15042(.A(shft_rshift4_b1[47]), .B(exu_n16227), .Y(exu_n27518));
INVX1 exu_U15043(.A(exu_n27518), .Y(exu_n2961));
AND2X1 exu_U15044(.A(shft_rshift4_b1[44]), .B(exu_n16224), .Y(exu_n27522));
INVX1 exu_U15045(.A(exu_n27522), .Y(exu_n2962));
AND2X1 exu_U15046(.A(shft_rshift4_b1[46]), .B(exu_n16227), .Y(exu_n27524));
INVX1 exu_U15047(.A(exu_n27524), .Y(exu_n2963));
AND2X1 exu_U15048(.A(shft_rshift4_b1[43]), .B(exu_n16223), .Y(exu_n27528));
INVX1 exu_U15049(.A(exu_n27528), .Y(exu_n2964));
AND2X1 exu_U15050(.A(shft_rshift4_b1[45]), .B(exu_n15402), .Y(exu_n27530));
INVX1 exu_U15051(.A(exu_n27530), .Y(exu_n2965));
AND2X1 exu_U15052(.A(shft_rshift4_b1[42]), .B(exu_n16223), .Y(exu_n27534));
INVX1 exu_U15053(.A(exu_n27534), .Y(exu_n2966));
AND2X1 exu_U15054(.A(shft_rshift4_b1[44]), .B(exu_n16227), .Y(exu_n27536));
INVX1 exu_U15055(.A(exu_n27536), .Y(exu_n2967));
AND2X1 exu_U15056(.A(shft_rshift4_b1[41]), .B(exu_n16223), .Y(exu_n27540));
INVX1 exu_U15057(.A(exu_n27540), .Y(exu_n2968));
AND2X1 exu_U15058(.A(shft_rshift4_b1[43]), .B(exu_n16227), .Y(exu_n27542));
INVX1 exu_U15059(.A(exu_n27542), .Y(exu_n2969));
AND2X1 exu_U15060(.A(shft_rshift4_b1[40]), .B(exu_n16224), .Y(exu_n27546));
INVX1 exu_U15061(.A(exu_n27546), .Y(exu_n2970));
AND2X1 exu_U15062(.A(shft_rshift4_b1[42]), .B(exu_n16227), .Y(exu_n27548));
INVX1 exu_U15063(.A(exu_n27548), .Y(exu_n2971));
AND2X1 exu_U15064(.A(shft_rshift4_b1[3]), .B(exu_n16223), .Y(exu_n27552));
INVX1 exu_U15065(.A(exu_n27552), .Y(exu_n2972));
AND2X1 exu_U15066(.A(shft_rshift4_b1[5]), .B(exu_n16227), .Y(exu_n27554));
INVX1 exu_U15067(.A(exu_n27554), .Y(exu_n2973));
AND2X1 exu_U15068(.A(shft_rshift4_b1[39]), .B(exu_n16223), .Y(exu_n27558));
INVX1 exu_U15069(.A(exu_n27558), .Y(exu_n2974));
AND2X1 exu_U15070(.A(shft_rshift4_b1[41]), .B(exu_n16227), .Y(exu_n27560));
INVX1 exu_U15071(.A(exu_n27560), .Y(exu_n2975));
AND2X1 exu_U15072(.A(shft_rshift4_b1[38]), .B(exu_n16224), .Y(exu_n27564));
INVX1 exu_U15073(.A(exu_n27564), .Y(exu_n2976));
AND2X1 exu_U15074(.A(shft_rshift4_b1[40]), .B(exu_n16227), .Y(exu_n27566));
INVX1 exu_U15075(.A(exu_n27566), .Y(exu_n2977));
AND2X1 exu_U15076(.A(shft_rshift4_b1[37]), .B(exu_n16224), .Y(exu_n27570));
INVX1 exu_U15077(.A(exu_n27570), .Y(exu_n2978));
AND2X1 exu_U15078(.A(shft_rshift4_b1[39]), .B(exu_n16227), .Y(exu_n27572));
INVX1 exu_U15079(.A(exu_n27572), .Y(exu_n2979));
AND2X1 exu_U15080(.A(shft_rshift4_b1[36]), .B(exu_n16224), .Y(exu_n27576));
INVX1 exu_U15081(.A(exu_n27576), .Y(exu_n2980));
AND2X1 exu_U15082(.A(shft_rshift4_b1[38]), .B(exu_n16227), .Y(exu_n27578));
INVX1 exu_U15083(.A(exu_n27578), .Y(exu_n2981));
AND2X1 exu_U15084(.A(shft_rshift4_b1[35]), .B(exu_n16223), .Y(exu_n27582));
INVX1 exu_U15085(.A(exu_n27582), .Y(exu_n2982));
AND2X1 exu_U15086(.A(shft_rshift4_b1[37]), .B(exu_n16227), .Y(exu_n27584));
INVX1 exu_U15087(.A(exu_n27584), .Y(exu_n2983));
AND2X1 exu_U15088(.A(shft_rshift4_b1[34]), .B(exu_n16223), .Y(exu_n27588));
INVX1 exu_U15089(.A(exu_n27588), .Y(exu_n2984));
AND2X1 exu_U15090(.A(shft_rshift4_b1[36]), .B(exu_n16227), .Y(exu_n27590));
INVX1 exu_U15091(.A(exu_n27590), .Y(exu_n2985));
AND2X1 exu_U15092(.A(shft_rshift4_b1[33]), .B(exu_n16224), .Y(exu_n27594));
INVX1 exu_U15093(.A(exu_n27594), .Y(exu_n2986));
AND2X1 exu_U15094(.A(shft_rshift4_b1[35]), .B(exu_n16227), .Y(exu_n27596));
INVX1 exu_U15095(.A(exu_n27596), .Y(exu_n2987));
AND2X1 exu_U15096(.A(shft_rshift4_b1[32]), .B(exu_n16223), .Y(exu_n27600));
INVX1 exu_U15097(.A(exu_n27600), .Y(exu_n2988));
AND2X1 exu_U15098(.A(shft_rshift4_b1[34]), .B(exu_n16227), .Y(exu_n27602));
INVX1 exu_U15099(.A(exu_n27602), .Y(exu_n2989));
AND2X1 exu_U15100(.A(shft_rshift4_b1[31]), .B(exu_n16224), .Y(exu_n27606));
INVX1 exu_U15101(.A(exu_n27606), .Y(exu_n2990));
AND2X1 exu_U15102(.A(shft_rshift4_b1[33]), .B(exu_n16227), .Y(exu_n27608));
INVX1 exu_U15103(.A(exu_n27608), .Y(exu_n2991));
AND2X1 exu_U15104(.A(shft_rshift4_b1[30]), .B(exu_n16223), .Y(exu_n27612));
INVX1 exu_U15105(.A(exu_n27612), .Y(exu_n2992));
AND2X1 exu_U15106(.A(shft_rshift4_b1[32]), .B(exu_n16227), .Y(exu_n27614));
INVX1 exu_U15107(.A(exu_n27614), .Y(exu_n2993));
AND2X1 exu_U15108(.A(shft_rshift4_b1[2]), .B(exu_n16224), .Y(exu_n27618));
INVX1 exu_U15109(.A(exu_n27618), .Y(exu_n2994));
AND2X1 exu_U15110(.A(shft_rshift4_b1[4]), .B(exu_n15402), .Y(exu_n27620));
INVX1 exu_U15111(.A(exu_n27620), .Y(exu_n2995));
AND2X1 exu_U15112(.A(shft_rshift4_b1[29]), .B(exu_n16224), .Y(exu_n27624));
INVX1 exu_U15113(.A(exu_n27624), .Y(exu_n2996));
AND2X1 exu_U15114(.A(shft_rshift4_b1[31]), .B(exu_n16227), .Y(exu_n27626));
INVX1 exu_U15115(.A(exu_n27626), .Y(exu_n2997));
AND2X1 exu_U15116(.A(shft_rshift4_b1[28]), .B(exu_n16224), .Y(exu_n27630));
INVX1 exu_U15117(.A(exu_n27630), .Y(exu_n2998));
AND2X1 exu_U15118(.A(shft_rshift4_b1[30]), .B(exu_n15402), .Y(exu_n27632));
INVX1 exu_U15119(.A(exu_n27632), .Y(exu_n2999));
AND2X1 exu_U15120(.A(shft_rshift4_b1[27]), .B(exu_n16224), .Y(exu_n27636));
INVX1 exu_U15121(.A(exu_n27636), .Y(exu_n3000));
AND2X1 exu_U15122(.A(shft_rshift4_b1[29]), .B(exu_n16227), .Y(exu_n27638));
INVX1 exu_U15123(.A(exu_n27638), .Y(exu_n3001));
AND2X1 exu_U15124(.A(shft_rshift4_b1[26]), .B(exu_n16223), .Y(exu_n27642));
INVX1 exu_U15125(.A(exu_n27642), .Y(exu_n3002));
AND2X1 exu_U15126(.A(shft_rshift4_b1[28]), .B(exu_n15402), .Y(exu_n27644));
INVX1 exu_U15127(.A(exu_n27644), .Y(exu_n3003));
AND2X1 exu_U15128(.A(shft_rshift4_b1[25]), .B(exu_n16224), .Y(exu_n27648));
INVX1 exu_U15129(.A(exu_n27648), .Y(exu_n3004));
AND2X1 exu_U15130(.A(shft_rshift4_b1[27]), .B(exu_n15402), .Y(exu_n27650));
INVX1 exu_U15131(.A(exu_n27650), .Y(exu_n3005));
AND2X1 exu_U15132(.A(shft_rshift4_b1[24]), .B(exu_n16223), .Y(exu_n27654));
INVX1 exu_U15133(.A(exu_n27654), .Y(exu_n3006));
AND2X1 exu_U15134(.A(shft_rshift4_b1[26]), .B(exu_n16227), .Y(exu_n27656));
INVX1 exu_U15135(.A(exu_n27656), .Y(exu_n3007));
AND2X1 exu_U15136(.A(shft_rshift4_b1[23]), .B(exu_n16224), .Y(exu_n27660));
INVX1 exu_U15137(.A(exu_n27660), .Y(exu_n3008));
AND2X1 exu_U15138(.A(shft_rshift4_b1[25]), .B(exu_n16227), .Y(exu_n27662));
INVX1 exu_U15139(.A(exu_n27662), .Y(exu_n3009));
AND2X1 exu_U15140(.A(shft_rshift4_b1[22]), .B(exu_n16223), .Y(exu_n27666));
INVX1 exu_U15141(.A(exu_n27666), .Y(exu_n3010));
AND2X1 exu_U15142(.A(shft_rshift4_b1[24]), .B(exu_n15402), .Y(exu_n27668));
INVX1 exu_U15143(.A(exu_n27668), .Y(exu_n3011));
AND2X1 exu_U15144(.A(shft_rshift4_b1[21]), .B(exu_n16223), .Y(exu_n27672));
INVX1 exu_U15145(.A(exu_n27672), .Y(exu_n3012));
AND2X1 exu_U15146(.A(shft_rshift4_b1[23]), .B(exu_n16227), .Y(exu_n27674));
INVX1 exu_U15147(.A(exu_n27674), .Y(exu_n3013));
AND2X1 exu_U15148(.A(shft_rshift4_b1[20]), .B(exu_n16224), .Y(exu_n27678));
INVX1 exu_U15149(.A(exu_n27678), .Y(exu_n3014));
AND2X1 exu_U15150(.A(shft_rshift4_b1[22]), .B(exu_n15402), .Y(exu_n27680));
INVX1 exu_U15151(.A(exu_n27680), .Y(exu_n3015));
AND2X1 exu_U15152(.A(shft_rshift4_b1[1]), .B(exu_n16223), .Y(exu_n27684));
INVX1 exu_U15153(.A(exu_n27684), .Y(exu_n3016));
AND2X1 exu_U15154(.A(shft_rshift4_b1[3]), .B(exu_n15402), .Y(exu_n27686));
INVX1 exu_U15155(.A(exu_n27686), .Y(exu_n3017));
AND2X1 exu_U15156(.A(shft_rshift4_b1[19]), .B(exu_n16224), .Y(exu_n27690));
INVX1 exu_U15157(.A(exu_n27690), .Y(exu_n3018));
AND2X1 exu_U15158(.A(shft_rshift4_b1[21]), .B(exu_n16227), .Y(exu_n27692));
INVX1 exu_U15159(.A(exu_n27692), .Y(exu_n3019));
AND2X1 exu_U15160(.A(shft_rshift4_b1[18]), .B(exu_n16224), .Y(exu_n27696));
INVX1 exu_U15161(.A(exu_n27696), .Y(exu_n3020));
AND2X1 exu_U15162(.A(shft_rshift4_b1[20]), .B(exu_n15402), .Y(exu_n27698));
INVX1 exu_U15163(.A(exu_n27698), .Y(exu_n3021));
AND2X1 exu_U15164(.A(shft_rshift4_b1[17]), .B(exu_n16224), .Y(exu_n27702));
INVX1 exu_U15165(.A(exu_n27702), .Y(exu_n3022));
AND2X1 exu_U15166(.A(shft_rshift4_b1[19]), .B(exu_n15402), .Y(exu_n27704));
INVX1 exu_U15167(.A(exu_n27704), .Y(exu_n3023));
AND2X1 exu_U15168(.A(shft_rshift4_b1[16]), .B(exu_n16223), .Y(exu_n27708));
INVX1 exu_U15169(.A(exu_n27708), .Y(exu_n3024));
AND2X1 exu_U15170(.A(shft_rshift4_b1[18]), .B(exu_n15402), .Y(exu_n27710));
INVX1 exu_U15171(.A(exu_n27710), .Y(exu_n3025));
AND2X1 exu_U15172(.A(shft_rshift4_b1[15]), .B(exu_n16224), .Y(exu_n27714));
INVX1 exu_U15173(.A(exu_n27714), .Y(exu_n3026));
AND2X1 exu_U15174(.A(shft_rshift4_b1[17]), .B(exu_n15402), .Y(exu_n27716));
INVX1 exu_U15175(.A(exu_n27716), .Y(exu_n3027));
AND2X1 exu_U15176(.A(shft_rshift4_b1[14]), .B(exu_n16223), .Y(exu_n27720));
INVX1 exu_U15177(.A(exu_n27720), .Y(exu_n3028));
AND2X1 exu_U15178(.A(shft_rshift4_b1[16]), .B(exu_n15402), .Y(exu_n27722));
INVX1 exu_U15179(.A(exu_n27722), .Y(exu_n3029));
AND2X1 exu_U15180(.A(shft_rshift4_b1[13]), .B(exu_n16224), .Y(exu_n27726));
INVX1 exu_U15181(.A(exu_n27726), .Y(exu_n3030));
AND2X1 exu_U15182(.A(shft_rshift4_b1[15]), .B(exu_n15402), .Y(exu_n27728));
INVX1 exu_U15183(.A(exu_n27728), .Y(exu_n3031));
AND2X1 exu_U15184(.A(shft_rshift4_b1[12]), .B(exu_n16224), .Y(exu_n27732));
INVX1 exu_U15185(.A(exu_n27732), .Y(exu_n3032));
AND2X1 exu_U15186(.A(shft_rshift4_b1[14]), .B(exu_n16227), .Y(exu_n27734));
INVX1 exu_U15187(.A(exu_n27734), .Y(exu_n3033));
AND2X1 exu_U15188(.A(shft_rshift4_b1[11]), .B(exu_n16224), .Y(exu_n27738));
INVX1 exu_U15189(.A(exu_n27738), .Y(exu_n3034));
AND2X1 exu_U15190(.A(shft_rshift4_b1[13]), .B(exu_n15402), .Y(exu_n27740));
INVX1 exu_U15191(.A(exu_n27740), .Y(exu_n3035));
AND2X1 exu_U15192(.A(shft_rshift4_b1[10]), .B(exu_n16223), .Y(exu_n27744));
INVX1 exu_U15193(.A(exu_n27744), .Y(exu_n3036));
AND2X1 exu_U15194(.A(shft_rshift4_b1[12]), .B(exu_n16227), .Y(exu_n27746));
INVX1 exu_U15195(.A(exu_n27746), .Y(exu_n3037));
AND2X1 exu_U15196(.A(shft_rshift4_b1[0]), .B(exu_n16224), .Y(exu_n27750));
INVX1 exu_U15197(.A(exu_n27750), .Y(exu_n3038));
AND2X1 exu_U15198(.A(shft_rshift4_b1[2]), .B(exu_n16227), .Y(exu_n27752));
INVX1 exu_U15199(.A(exu_n27752), .Y(exu_n3039));
AND2X1 exu_U15200(.A(shft_shifter_input_b1[63]), .B(shft_shift16_e[0]), .Y(exu_n27760));
INVX1 exu_U15201(.A(exu_n27760), .Y(exu_n3040));
AND2X1 exu_U15202(.A(shft_rshifterinput_b1[31]), .B(exu_n16145), .Y(exu_n27762));
INVX1 exu_U15203(.A(exu_n27762), .Y(exu_n3041));
AND2X1 exu_U15204(.A(shft_shifter_input_b1[62]), .B(exu_n16148), .Y(exu_n27766));
INVX1 exu_U15205(.A(exu_n27766), .Y(exu_n3042));
AND2X1 exu_U15206(.A(shft_rshifterinput_b1[30]), .B(exu_n16145), .Y(exu_n27768));
INVX1 exu_U15207(.A(exu_n27768), .Y(exu_n3043));
AND2X1 exu_U15208(.A(shft_shifter_input_b1[61]), .B(exu_n16148), .Y(exu_n27772));
INVX1 exu_U15209(.A(exu_n27772), .Y(exu_n3044));
AND2X1 exu_U15210(.A(shft_rshifterinput_b1[29]), .B(exu_n16145), .Y(exu_n27774));
INVX1 exu_U15211(.A(exu_n27774), .Y(exu_n3045));
AND2X1 exu_U15212(.A(shft_shifter_input_b1[60]), .B(exu_n16148), .Y(exu_n27778));
INVX1 exu_U15213(.A(exu_n27778), .Y(exu_n3046));
AND2X1 exu_U15214(.A(shft_rshifterinput_b1[28]), .B(exu_n16145), .Y(exu_n27780));
INVX1 exu_U15215(.A(exu_n27780), .Y(exu_n3047));
AND2X1 exu_U15216(.A(shft_shifter_input_b1[59]), .B(shft_shift16_e[0]), .Y(exu_n27785));
INVX1 exu_U15217(.A(exu_n27785), .Y(exu_n3048));
AND2X1 exu_U15218(.A(shft_rshifterinput_b1[27]), .B(exu_n16145), .Y(exu_n27787));
INVX1 exu_U15219(.A(exu_n27787), .Y(exu_n3049));
AND2X1 exu_U15220(.A(shft_shifter_input_b1[58]), .B(exu_n16148), .Y(exu_n27791));
INVX1 exu_U15221(.A(exu_n27791), .Y(exu_n3050));
AND2X1 exu_U15222(.A(shft_rshifterinput_b1[26]), .B(exu_n16145), .Y(exu_n27793));
INVX1 exu_U15223(.A(exu_n27793), .Y(exu_n3051));
AND2X1 exu_U15224(.A(shft_shifter_input_b1[57]), .B(shft_shift16_e[0]), .Y(exu_n27797));
INVX1 exu_U15225(.A(exu_n27797), .Y(exu_n3052));
AND2X1 exu_U15226(.A(shft_rshifterinput_b1[25]), .B(exu_n16145), .Y(exu_n27799));
INVX1 exu_U15227(.A(exu_n27799), .Y(exu_n3053));
AND2X1 exu_U15228(.A(shft_shifter_input_b1[56]), .B(shft_shift16_e[0]), .Y(exu_n27803));
INVX1 exu_U15229(.A(exu_n27803), .Y(exu_n3054));
AND2X1 exu_U15230(.A(shft_rshifterinput_b1[24]), .B(exu_n16145), .Y(exu_n27805));
INVX1 exu_U15231(.A(exu_n27805), .Y(exu_n3055));
AND2X1 exu_U15232(.A(shft_shifter_input_b1[55]), .B(shft_shift16_e[0]), .Y(exu_n27809));
INVX1 exu_U15233(.A(exu_n27809), .Y(exu_n3056));
AND2X1 exu_U15234(.A(shft_rshifterinput_b1[23]), .B(exu_n16145), .Y(exu_n27811));
INVX1 exu_U15235(.A(exu_n27811), .Y(exu_n3057));
AND2X1 exu_U15236(.A(shft_shifter_input_b1[54]), .B(shft_shift16_e[0]), .Y(exu_n27815));
INVX1 exu_U15237(.A(exu_n27815), .Y(exu_n3058));
AND2X1 exu_U15238(.A(shft_rshifterinput_b1[22]), .B(exu_n16145), .Y(exu_n27817));
INVX1 exu_U15239(.A(exu_n27817), .Y(exu_n3059));
AND2X1 exu_U15240(.A(shft_shifter_input_b1[53]), .B(shft_shift16_e[0]), .Y(exu_n27821));
INVX1 exu_U15241(.A(exu_n27821), .Y(exu_n3060));
AND2X1 exu_U15242(.A(shft_rshifterinput_b1[21]), .B(exu_n16145), .Y(exu_n27823));
INVX1 exu_U15243(.A(exu_n27823), .Y(exu_n3061));
AND2X1 exu_U15244(.A(shft_shifter_input_b1[52]), .B(shft_shift16_e[0]), .Y(exu_n27827));
INVX1 exu_U15245(.A(exu_n27827), .Y(exu_n3062));
AND2X1 exu_U15246(.A(shft_rshifterinput_b1[20]), .B(exu_n16145), .Y(exu_n27829));
INVX1 exu_U15247(.A(exu_n27829), .Y(exu_n3063));
AND2X1 exu_U15248(.A(shft_shifter_input_b1[51]), .B(shft_shift16_e[0]), .Y(exu_n27833));
INVX1 exu_U15249(.A(exu_n27833), .Y(exu_n3064));
AND2X1 exu_U15250(.A(shft_rshifterinput_b1[19]), .B(exu_n16145), .Y(exu_n27835));
INVX1 exu_U15251(.A(exu_n27835), .Y(exu_n3065));
AND2X1 exu_U15252(.A(shft_shifter_input_b1[50]), .B(shft_shift16_e[0]), .Y(exu_n27839));
INVX1 exu_U15253(.A(exu_n27839), .Y(exu_n3066));
AND2X1 exu_U15254(.A(shft_rshifterinput_b1[18]), .B(exu_n16145), .Y(exu_n27841));
INVX1 exu_U15255(.A(exu_n27841), .Y(exu_n3067));
AND2X1 exu_U15256(.A(shft_shifter_input_b1[49]), .B(shft_shift16_e[0]), .Y(exu_n27846));
INVX1 exu_U15257(.A(exu_n27846), .Y(exu_n3068));
AND2X1 exu_U15258(.A(shft_rshifterinput_b1[17]), .B(exu_n16145), .Y(exu_n27848));
INVX1 exu_U15259(.A(exu_n27848), .Y(exu_n3069));
AND2X1 exu_U15260(.A(shft_shifter_input_b1[48]), .B(shft_shift16_e[0]), .Y(exu_n27852));
INVX1 exu_U15261(.A(exu_n27852), .Y(exu_n3070));
AND2X1 exu_U15262(.A(shft_rshifterinput_b1[16]), .B(exu_n16145), .Y(exu_n27854));
INVX1 exu_U15263(.A(exu_n27854), .Y(exu_n3071));
AND2X1 exu_U15264(.A(shft_shifter_input_b1[47]), .B(exu_n16148), .Y(exu_n27857));
INVX1 exu_U15265(.A(exu_n27857), .Y(exu_n3072));
AND2X1 exu_U15266(.A(shft_shifter_input_b1[46]), .B(exu_n16148), .Y(exu_n27861));
INVX1 exu_U15267(.A(exu_n27861), .Y(exu_n3073));
AND2X1 exu_U15268(.A(shft_shifter_input_b1[45]), .B(exu_n16148), .Y(exu_n27865));
INVX1 exu_U15269(.A(exu_n27865), .Y(exu_n3074));
AND2X1 exu_U15270(.A(shft_shifter_input_b1[44]), .B(exu_n16148), .Y(exu_n27869));
INVX1 exu_U15271(.A(exu_n27869), .Y(exu_n3075));
AND2X1 exu_U15272(.A(shft_shifter_input_b1[43]), .B(exu_n16148), .Y(exu_n27873));
INVX1 exu_U15273(.A(exu_n27873), .Y(exu_n3076));
AND2X1 exu_U15274(.A(shft_shifter_input_b1[42]), .B(exu_n16148), .Y(exu_n27877));
INVX1 exu_U15275(.A(exu_n27877), .Y(exu_n3077));
AND2X1 exu_U15276(.A(shft_shifter_input_b1[41]), .B(exu_n16148), .Y(exu_n27881));
INVX1 exu_U15277(.A(exu_n27881), .Y(exu_n3078));
AND2X1 exu_U15278(.A(shft_shifter_input_b1[40]), .B(exu_n16148), .Y(exu_n27885));
INVX1 exu_U15279(.A(exu_n27885), .Y(exu_n3079));
AND2X1 exu_U15280(.A(shft_shifter_input_b1[39]), .B(exu_n16148), .Y(exu_n27890));
INVX1 exu_U15281(.A(exu_n27890), .Y(exu_n3080));
AND2X1 exu_U15282(.A(shft_shifter_input_b1[38]), .B(exu_n16148), .Y(exu_n27894));
INVX1 exu_U15283(.A(exu_n27894), .Y(exu_n3081));
AND2X1 exu_U15284(.A(shft_shifter_input_b1[37]), .B(exu_n16148), .Y(exu_n27898));
INVX1 exu_U15285(.A(exu_n27898), .Y(exu_n3082));
AND2X1 exu_U15286(.A(shft_shifter_input_b1[36]), .B(exu_n16148), .Y(exu_n27902));
INVX1 exu_U15287(.A(exu_n27902), .Y(exu_n3083));
AND2X1 exu_U15288(.A(shft_shifter_input_b1[35]), .B(exu_n16148), .Y(exu_n27906));
INVX1 exu_U15289(.A(exu_n27906), .Y(exu_n3084));
AND2X1 exu_U15290(.A(shft_shifter_input_b1[34]), .B(exu_n16148), .Y(exu_n27910));
INVX1 exu_U15291(.A(exu_n27910), .Y(exu_n3085));
AND2X1 exu_U15292(.A(shft_shifter_input_b1[33]), .B(exu_n16148), .Y(exu_n27914));
INVX1 exu_U15293(.A(exu_n27914), .Y(exu_n3086));
AND2X1 exu_U15294(.A(shft_shifter_input_b1[32]), .B(exu_n16148), .Y(exu_n27918));
INVX1 exu_U15295(.A(exu_n27918), .Y(exu_n3087));
AND2X1 exu_U15296(.A(shft_rshifterinput_b1[31]), .B(exu_n16148), .Y(exu_n27922));
INVX1 exu_U15297(.A(exu_n27922), .Y(exu_n3088));
AND2X1 exu_U15298(.A(shft_rshifterinput_b1[30]), .B(shft_shift16_e[0]), .Y(exu_n27925));
INVX1 exu_U15299(.A(exu_n27925), .Y(exu_n3089));
AND2X1 exu_U15300(.A(shft_rshifterinput_b1[29]), .B(exu_n16148), .Y(exu_n27929));
INVX1 exu_U15301(.A(exu_n27929), .Y(exu_n3090));
AND2X1 exu_U15302(.A(shft_rshifterinput_b1[28]), .B(shft_shift16_e[0]), .Y(exu_n27932));
INVX1 exu_U15303(.A(exu_n27932), .Y(exu_n3091));
AND2X1 exu_U15304(.A(shft_rshifterinput_b1[27]), .B(exu_n16148), .Y(exu_n27935));
INVX1 exu_U15305(.A(exu_n27935), .Y(exu_n3092));
AND2X1 exu_U15306(.A(shft_rshifterinput_b1[26]), .B(shft_shift16_e[0]), .Y(exu_n27938));
INVX1 exu_U15307(.A(exu_n27938), .Y(exu_n3093));
AND2X1 exu_U15308(.A(shft_rshifterinput_b1[25]), .B(exu_n16148), .Y(exu_n27941));
INVX1 exu_U15309(.A(exu_n27941), .Y(exu_n3094));
AND2X1 exu_U15310(.A(shft_rshifterinput_b1[24]), .B(shft_shift16_e[0]), .Y(exu_n27944));
INVX1 exu_U15311(.A(exu_n27944), .Y(exu_n3095));
AND2X1 exu_U15312(.A(shft_rshifterinput_b1[23]), .B(exu_n16148), .Y(exu_n27947));
INVX1 exu_U15313(.A(exu_n27947), .Y(exu_n3096));
AND2X1 exu_U15314(.A(shft_rshifterinput_b1[22]), .B(shft_shift16_e[0]), .Y(exu_n27950));
INVX1 exu_U15315(.A(exu_n27950), .Y(exu_n3097));
AND2X1 exu_U15316(.A(shft_rshifterinput_b1[21]), .B(exu_n16148), .Y(exu_n27953));
INVX1 exu_U15317(.A(exu_n27953), .Y(exu_n3098));
AND2X1 exu_U15318(.A(shft_rshifterinput_b1[20]), .B(shft_shift16_e[0]), .Y(exu_n27956));
INVX1 exu_U15319(.A(exu_n27956), .Y(exu_n3099));
AND2X1 exu_U15320(.A(shft_rshifterinput_b1[19]), .B(exu_n16148), .Y(exu_n27960));
INVX1 exu_U15321(.A(exu_n27960), .Y(exu_n3100));
AND2X1 exu_U15322(.A(shft_rshifterinput_b1[18]), .B(shft_shift16_e[0]), .Y(exu_n27963));
INVX1 exu_U15323(.A(exu_n27963), .Y(exu_n3101));
AND2X1 exu_U15324(.A(shft_rshifterinput_b1[17]), .B(shft_shift16_e[0]), .Y(exu_n27966));
INVX1 exu_U15325(.A(exu_n27966), .Y(exu_n3102));
AND2X1 exu_U15326(.A(shft_rshifterinput_b1[16]), .B(shft_shift16_e[0]), .Y(exu_n27969));
INVX1 exu_U15327(.A(exu_n27969), .Y(exu_n3103));
AND2X1 exu_U15328(.A(exu_n15401), .B(exu_n27754), .Y(exu_n27979));
INVX1 exu_U15329(.A(exu_n27979), .Y(exu_n3104));
AND2X1 exu_U15330(.A(exu_n27755), .B(exu_n15401), .Y(exu_n27983));
INVX1 exu_U15331(.A(exu_n27983), .Y(exu_n3105));
AND2X1 exu_U15332(.A(exu_n27756), .B(exu_n16230), .Y(exu_n27987));
INVX1 exu_U15333(.A(exu_n27987), .Y(exu_n3106));
AND2X1 exu_U15334(.A(exu_n27757), .B(exu_n15401), .Y(exu_n27990));
INVX1 exu_U15335(.A(exu_n27990), .Y(exu_n3107));
AND2X1 exu_U15336(.A(shft_lshift16_b1[63]), .B(exu_n15401), .Y(exu_n27994));
INVX1 exu_U15337(.A(exu_n27994), .Y(exu_n3108));
AND2X1 exu_U15338(.A(shft_lshift16_b1[55]), .B(exu_n16233), .Y(exu_n27996));
INVX1 exu_U15339(.A(exu_n27996), .Y(exu_n3109));
AND2X1 exu_U15340(.A(shft_lshift16_b1[62]), .B(exu_n16230), .Y(exu_n28000));
INVX1 exu_U15341(.A(exu_n28000), .Y(exu_n3110));
AND2X1 exu_U15342(.A(shft_lshift16_b1[54]), .B(exu_n16232), .Y(exu_n28002));
INVX1 exu_U15343(.A(exu_n28002), .Y(exu_n3111));
AND2X1 exu_U15344(.A(shft_lshift16_b1[61]), .B(exu_n15401), .Y(exu_n28006));
INVX1 exu_U15345(.A(exu_n28006), .Y(exu_n3112));
AND2X1 exu_U15346(.A(shft_lshift16_b1[53]), .B(exu_n16233), .Y(exu_n28008));
INVX1 exu_U15347(.A(exu_n28008), .Y(exu_n3113));
AND2X1 exu_U15348(.A(shft_lshift16_b1[60]), .B(exu_n16230), .Y(exu_n28012));
INVX1 exu_U15349(.A(exu_n28012), .Y(exu_n3114));
AND2X1 exu_U15350(.A(shft_lshift16_b1[52]), .B(exu_n16232), .Y(exu_n28014));
INVX1 exu_U15351(.A(exu_n28014), .Y(exu_n3115));
AND2X1 exu_U15352(.A(exu_n27782), .B(exu_n16230), .Y(exu_n28017));
INVX1 exu_U15353(.A(exu_n28017), .Y(exu_n3116));
AND2X1 exu_U15354(.A(shft_lshift16_b1[59]), .B(exu_n15401), .Y(exu_n28021));
INVX1 exu_U15355(.A(exu_n28021), .Y(exu_n3117));
AND2X1 exu_U15356(.A(shft_lshift16_b1[51]), .B(exu_n16233), .Y(exu_n28023));
INVX1 exu_U15357(.A(exu_n28023), .Y(exu_n3118));
AND2X1 exu_U15358(.A(shft_lshift16_b1[58]), .B(exu_n15401), .Y(exu_n28027));
INVX1 exu_U15359(.A(exu_n28027), .Y(exu_n3119));
AND2X1 exu_U15360(.A(shft_lshift16_b1[50]), .B(exu_n16233), .Y(exu_n28029));
INVX1 exu_U15361(.A(exu_n28029), .Y(exu_n3120));
AND2X1 exu_U15362(.A(shft_lshift16_b1[57]), .B(exu_n15401), .Y(exu_n28033));
INVX1 exu_U15363(.A(exu_n28033), .Y(exu_n3121));
AND2X1 exu_U15364(.A(shft_lshift16_b1[49]), .B(exu_n16233), .Y(exu_n28035));
INVX1 exu_U15365(.A(exu_n28035), .Y(exu_n3122));
AND2X1 exu_U15366(.A(shft_lshift16_b1[56]), .B(exu_n15401), .Y(exu_n28039));
INVX1 exu_U15367(.A(exu_n28039), .Y(exu_n3123));
AND2X1 exu_U15368(.A(shft_lshift16_b1[48]), .B(exu_n16233), .Y(exu_n28041));
INVX1 exu_U15369(.A(exu_n28041), .Y(exu_n3124));
AND2X1 exu_U15370(.A(shft_lshift16_b1[55]), .B(exu_n15401), .Y(exu_n28045));
INVX1 exu_U15371(.A(exu_n28045), .Y(exu_n3125));
AND2X1 exu_U15372(.A(shft_lshift16_b1[47]), .B(exu_n16233), .Y(exu_n28047));
INVX1 exu_U15373(.A(exu_n28047), .Y(exu_n3126));
AND2X1 exu_U15374(.A(shft_lshift16_b1[54]), .B(exu_n16230), .Y(exu_n28051));
INVX1 exu_U15375(.A(exu_n28051), .Y(exu_n3127));
AND2X1 exu_U15376(.A(shft_lshift16_b1[46]), .B(exu_n16232), .Y(exu_n28053));
INVX1 exu_U15377(.A(exu_n28053), .Y(exu_n3128));
AND2X1 exu_U15378(.A(shft_lshift16_b1[53]), .B(exu_n15401), .Y(exu_n28057));
INVX1 exu_U15379(.A(exu_n28057), .Y(exu_n3129));
AND2X1 exu_U15380(.A(shft_lshift16_b1[45]), .B(exu_n16232), .Y(exu_n28059));
INVX1 exu_U15381(.A(exu_n28059), .Y(exu_n3130));
AND2X1 exu_U15382(.A(shft_lshift16_b1[52]), .B(exu_n16230), .Y(exu_n28063));
INVX1 exu_U15383(.A(exu_n28063), .Y(exu_n3131));
AND2X1 exu_U15384(.A(shft_lshift16_b1[44]), .B(exu_n16233), .Y(exu_n28065));
INVX1 exu_U15385(.A(exu_n28065), .Y(exu_n3132));
AND2X1 exu_U15386(.A(shft_lshift16_b1[51]), .B(exu_n15401), .Y(exu_n28069));
INVX1 exu_U15387(.A(exu_n28069), .Y(exu_n3133));
AND2X1 exu_U15388(.A(shft_lshift16_b1[43]), .B(exu_n16233), .Y(exu_n28071));
INVX1 exu_U15389(.A(exu_n28071), .Y(exu_n3134));
AND2X1 exu_U15390(.A(shft_lshift16_b1[50]), .B(exu_n15401), .Y(exu_n28075));
INVX1 exu_U15391(.A(exu_n28075), .Y(exu_n3135));
AND2X1 exu_U15392(.A(shft_lshift16_b1[42]), .B(exu_n16233), .Y(exu_n28077));
INVX1 exu_U15393(.A(exu_n28077), .Y(exu_n3136));
AND2X1 exu_U15394(.A(exu_n27843), .B(exu_n16230), .Y(exu_n28080));
INVX1 exu_U15395(.A(exu_n28080), .Y(exu_n3137));
AND2X1 exu_U15396(.A(shft_lshift16_b1[49]), .B(exu_n16230), .Y(exu_n28084));
INVX1 exu_U15397(.A(exu_n28084), .Y(exu_n3138));
AND2X1 exu_U15398(.A(shft_lshift16_b1[41]), .B(exu_n16233), .Y(exu_n28086));
INVX1 exu_U15399(.A(exu_n28086), .Y(exu_n3139));
AND2X1 exu_U15400(.A(shft_lshift16_b1[48]), .B(exu_n16230), .Y(exu_n28090));
INVX1 exu_U15401(.A(exu_n28090), .Y(exu_n3140));
AND2X1 exu_U15402(.A(shft_lshift16_b1[40]), .B(exu_n16233), .Y(exu_n28092));
INVX1 exu_U15403(.A(exu_n28092), .Y(exu_n3141));
AND2X1 exu_U15404(.A(shft_lshift16_b1[47]), .B(exu_n15401), .Y(exu_n28096));
INVX1 exu_U15405(.A(exu_n28096), .Y(exu_n3142));
AND2X1 exu_U15406(.A(shft_lshift16_b1[39]), .B(exu_n16232), .Y(exu_n28098));
INVX1 exu_U15407(.A(exu_n28098), .Y(exu_n3143));
AND2X1 exu_U15408(.A(shft_lshift16_b1[46]), .B(exu_n16230), .Y(exu_n28102));
INVX1 exu_U15409(.A(exu_n28102), .Y(exu_n3144));
AND2X1 exu_U15410(.A(shft_lshift16_b1[38]), .B(exu_n16232), .Y(exu_n28104));
INVX1 exu_U15411(.A(exu_n28104), .Y(exu_n3145));
AND2X1 exu_U15412(.A(shft_lshift16_b1[45]), .B(exu_n16230), .Y(exu_n28108));
INVX1 exu_U15413(.A(exu_n28108), .Y(exu_n3146));
AND2X1 exu_U15414(.A(shft_lshift16_b1[37]), .B(exu_n16232), .Y(exu_n28110));
INVX1 exu_U15415(.A(exu_n28110), .Y(exu_n3147));
AND2X1 exu_U15416(.A(shft_lshift16_b1[44]), .B(exu_n16230), .Y(exu_n28114));
INVX1 exu_U15417(.A(exu_n28114), .Y(exu_n3148));
AND2X1 exu_U15418(.A(shft_lshift16_b1[36]), .B(exu_n16233), .Y(exu_n28116));
INVX1 exu_U15419(.A(exu_n28116), .Y(exu_n3149));
AND2X1 exu_U15420(.A(shft_lshift16_b1[43]), .B(exu_n15401), .Y(exu_n28120));
INVX1 exu_U15421(.A(exu_n28120), .Y(exu_n3150));
AND2X1 exu_U15422(.A(shft_lshift16_b1[35]), .B(exu_n16232), .Y(exu_n28122));
INVX1 exu_U15423(.A(exu_n28122), .Y(exu_n3151));
AND2X1 exu_U15424(.A(shft_lshift16_b1[42]), .B(exu_n15401), .Y(exu_n28126));
INVX1 exu_U15425(.A(exu_n28126), .Y(exu_n3152));
AND2X1 exu_U15426(.A(shft_lshift16_b1[34]), .B(exu_n16232), .Y(exu_n28128));
INVX1 exu_U15427(.A(exu_n28128), .Y(exu_n3153));
AND2X1 exu_U15428(.A(shft_lshift16_b1[41]), .B(exu_n16230), .Y(exu_n28132));
INVX1 exu_U15429(.A(exu_n28132), .Y(exu_n3154));
AND2X1 exu_U15430(.A(shft_lshift16_b1[33]), .B(exu_n16233), .Y(exu_n28134));
INVX1 exu_U15431(.A(exu_n28134), .Y(exu_n3155));
AND2X1 exu_U15432(.A(shft_lshift16_b1[40]), .B(exu_n15401), .Y(exu_n28138));
INVX1 exu_U15433(.A(exu_n28138), .Y(exu_n3156));
AND2X1 exu_U15434(.A(shft_lshift16_b1[32]), .B(exu_n16232), .Y(exu_n28140));
INVX1 exu_U15435(.A(exu_n28140), .Y(exu_n3157));
AND2X1 exu_U15436(.A(shft_lshift16_b1[39]), .B(exu_n16230), .Y(exu_n28145));
INVX1 exu_U15437(.A(exu_n28145), .Y(exu_n3158));
AND2X1 exu_U15438(.A(exu_n15703), .B(exu_n16233), .Y(exu_n28147));
INVX1 exu_U15439(.A(exu_n28147), .Y(exu_n3159));
AND2X1 exu_U15440(.A(shft_lshift16_b1[38]), .B(exu_n15401), .Y(exu_n28151));
INVX1 exu_U15441(.A(exu_n28151), .Y(exu_n3160));
AND2X1 exu_U15442(.A(exu_n15704), .B(exu_n16233), .Y(exu_n28153));
INVX1 exu_U15443(.A(exu_n28153), .Y(exu_n3161));
AND2X1 exu_U15444(.A(shft_lshift16_b1[37]), .B(exu_n15401), .Y(exu_n28157));
INVX1 exu_U15445(.A(exu_n28157), .Y(exu_n3162));
AND2X1 exu_U15446(.A(exu_n15705), .B(exu_n16232), .Y(exu_n28159));
INVX1 exu_U15447(.A(exu_n28159), .Y(exu_n3163));
AND2X1 exu_U15448(.A(shft_lshift16_b1[36]), .B(exu_n16230), .Y(exu_n28163));
INVX1 exu_U15449(.A(exu_n28163), .Y(exu_n3164));
AND2X1 exu_U15450(.A(exu_n15706), .B(exu_n16232), .Y(exu_n28165));
INVX1 exu_U15451(.A(exu_n28165), .Y(exu_n3165));
AND2X1 exu_U15452(.A(shft_lshift16_b1[35]), .B(exu_n15401), .Y(exu_n28169));
INVX1 exu_U15453(.A(exu_n28169), .Y(exu_n3166));
AND2X1 exu_U15454(.A(exu_n15707), .B(exu_n16232), .Y(exu_n28171));
INVX1 exu_U15455(.A(exu_n28171), .Y(exu_n3167));
AND2X1 exu_U15456(.A(shft_lshift16_b1[34]), .B(exu_n15401), .Y(exu_n28175));
INVX1 exu_U15457(.A(exu_n28175), .Y(exu_n3168));
AND2X1 exu_U15458(.A(exu_n15708), .B(exu_n16233), .Y(exu_n28177));
INVX1 exu_U15459(.A(exu_n28177), .Y(exu_n3169));
AND2X1 exu_U15460(.A(shft_lshift16_b1[33]), .B(exu_n16230), .Y(exu_n28181));
INVX1 exu_U15461(.A(exu_n28181), .Y(exu_n3170));
AND2X1 exu_U15462(.A(exu_n15709), .B(exu_n16232), .Y(exu_n28183));
INVX1 exu_U15463(.A(exu_n28183), .Y(exu_n3171));
AND2X1 exu_U15464(.A(shft_lshift16_b1[32]), .B(exu_n15401), .Y(exu_n28187));
INVX1 exu_U15465(.A(exu_n28187), .Y(exu_n3172));
AND2X1 exu_U15466(.A(exu_n15710), .B(exu_n16232), .Y(exu_n28189));
INVX1 exu_U15467(.A(exu_n28189), .Y(exu_n3173));
AND2X1 exu_U15468(.A(exu_n15703), .B(exu_n15401), .Y(exu_n28193));
INVX1 exu_U15469(.A(exu_n28193), .Y(exu_n3174));
AND2X1 exu_U15470(.A(exu_n15711), .B(exu_n16232), .Y(exu_n28195));
INVX1 exu_U15471(.A(exu_n28195), .Y(exu_n3175));
AND2X1 exu_U15472(.A(exu_n15704), .B(exu_n16230), .Y(exu_n28199));
INVX1 exu_U15473(.A(exu_n28199), .Y(exu_n3176));
AND2X1 exu_U15474(.A(exu_n15712), .B(exu_n16233), .Y(exu_n28201));
INVX1 exu_U15475(.A(exu_n28201), .Y(exu_n3177));
AND2X1 exu_U15476(.A(exu_n15705), .B(exu_n16230), .Y(exu_n28206));
INVX1 exu_U15477(.A(exu_n28206), .Y(exu_n3178));
AND2X1 exu_U15478(.A(exu_n15713), .B(exu_n16233), .Y(exu_n28208));
INVX1 exu_U15479(.A(exu_n28208), .Y(exu_n3179));
AND2X1 exu_U15480(.A(exu_n15706), .B(exu_n15401), .Y(exu_n28212));
INVX1 exu_U15481(.A(exu_n28212), .Y(exu_n3180));
AND2X1 exu_U15482(.A(exu_n15714), .B(exu_n16232), .Y(exu_n28214));
INVX1 exu_U15483(.A(exu_n28214), .Y(exu_n3181));
AND2X1 exu_U15484(.A(exu_n15707), .B(exu_n16230), .Y(exu_n28218));
INVX1 exu_U15485(.A(exu_n28218), .Y(exu_n3182));
AND2X1 exu_U15486(.A(exu_n15715), .B(exu_n16233), .Y(exu_n28220));
INVX1 exu_U15487(.A(exu_n28220), .Y(exu_n3183));
AND2X1 exu_U15488(.A(exu_n15708), .B(exu_n15401), .Y(exu_n28224));
INVX1 exu_U15489(.A(exu_n28224), .Y(exu_n3184));
AND2X1 exu_U15490(.A(exu_n15716), .B(exu_n16232), .Y(exu_n28226));
INVX1 exu_U15491(.A(exu_n28226), .Y(exu_n3185));
AND2X1 exu_U15492(.A(exu_n15709), .B(exu_n16230), .Y(exu_n28230));
INVX1 exu_U15493(.A(exu_n28230), .Y(exu_n3186));
AND2X1 exu_U15494(.A(exu_n15717), .B(exu_n16233), .Y(exu_n28232));
INVX1 exu_U15495(.A(exu_n28232), .Y(exu_n3187));
AND2X1 exu_U15496(.A(exu_n15710), .B(exu_n15401), .Y(exu_n28236));
INVX1 exu_U15497(.A(exu_n28236), .Y(exu_n3188));
AND2X1 exu_U15498(.A(exu_n15718), .B(exu_n16233), .Y(exu_n28238));
INVX1 exu_U15499(.A(exu_n28238), .Y(exu_n3189));
AND2X1 exu_U15500(.A(exu_n15711), .B(exu_n16230), .Y(exu_n28242));
INVX1 exu_U15501(.A(exu_n28242), .Y(exu_n3190));
AND2X1 exu_U15502(.A(exu_n27971), .B(exu_n16232), .Y(exu_n28244));
INVX1 exu_U15503(.A(exu_n28244), .Y(exu_n3191));
AND2X1 exu_U15504(.A(exu_n15712), .B(exu_n16230), .Y(exu_n28248));
INVX1 exu_U15505(.A(exu_n28248), .Y(exu_n3192));
AND2X1 exu_U15506(.A(exu_n27972), .B(exu_n16232), .Y(exu_n28250));
INVX1 exu_U15507(.A(exu_n28250), .Y(exu_n3193));
AND2X1 exu_U15508(.A(exu_n15713), .B(exu_n16230), .Y(exu_n28254));
INVX1 exu_U15509(.A(exu_n28254), .Y(exu_n3194));
AND2X1 exu_U15510(.A(exu_n27973), .B(exu_n16232), .Y(exu_n28256));
INVX1 exu_U15511(.A(exu_n28256), .Y(exu_n3195));
AND2X1 exu_U15512(.A(exu_n15714), .B(exu_n15401), .Y(exu_n28260));
INVX1 exu_U15513(.A(exu_n28260), .Y(exu_n3196));
AND2X1 exu_U15514(.A(exu_n27974), .B(exu_n16233), .Y(exu_n28262));
INVX1 exu_U15515(.A(exu_n28262), .Y(exu_n3197));
AND2X1 exu_U15516(.A(exu_n15715), .B(exu_n15401), .Y(exu_n28267));
INVX1 exu_U15517(.A(exu_n28267), .Y(exu_n3198));
AND2X1 exu_U15518(.A(exu_n27975), .B(exu_n16232), .Y(exu_n28269));
INVX1 exu_U15519(.A(exu_n28269), .Y(exu_n3199));
AND2X1 exu_U15520(.A(exu_n15716), .B(exu_n16230), .Y(exu_n28273));
INVX1 exu_U15521(.A(exu_n28273), .Y(exu_n3200));
AND2X1 exu_U15522(.A(exu_n27976), .B(exu_n16233), .Y(exu_n28275));
INVX1 exu_U15523(.A(exu_n28275), .Y(exu_n3201));
AND2X1 exu_U15524(.A(exu_n15717), .B(exu_n15401), .Y(exu_n28279));
INVX1 exu_U15525(.A(exu_n28279), .Y(exu_n3202));
AND2X1 exu_U15526(.A(exu_n27754), .B(exu_n16232), .Y(exu_n28281));
INVX1 exu_U15527(.A(exu_n28281), .Y(exu_n3203));
AND2X1 exu_U15528(.A(exu_n15718), .B(exu_n16230), .Y(exu_n28285));
INVX1 exu_U15529(.A(exu_n28285), .Y(exu_n3204));
AND2X1 exu_U15530(.A(exu_n27755), .B(exu_n16233), .Y(exu_n28287));
INVX1 exu_U15531(.A(exu_n28287), .Y(exu_n3205));
AND2X1 exu_U15532(.A(exu_n27971), .B(exu_n15401), .Y(exu_n28291));
INVX1 exu_U15533(.A(exu_n28291), .Y(exu_n3206));
AND2X1 exu_U15534(.A(exu_n27756), .B(exu_n16233), .Y(exu_n28293));
INVX1 exu_U15535(.A(exu_n28293), .Y(exu_n3207));
AND2X1 exu_U15536(.A(exu_n27972), .B(exu_n15401), .Y(exu_n28297));
INVX1 exu_U15537(.A(exu_n28297), .Y(exu_n3208));
AND2X1 exu_U15538(.A(exu_n27757), .B(exu_n16233), .Y(exu_n28299));
INVX1 exu_U15539(.A(exu_n28299), .Y(exu_n3209));
AND2X1 exu_U15540(.A(exu_n27973), .B(exu_n16230), .Y(exu_n28303));
INVX1 exu_U15541(.A(exu_n28303), .Y(exu_n3210));
AND2X1 exu_U15542(.A(exu_n27782), .B(exu_n16232), .Y(exu_n28305));
INVX1 exu_U15543(.A(exu_n28305), .Y(exu_n3211));
AND2X1 exu_U15544(.A(exu_n27974), .B(exu_n16230), .Y(exu_n28309));
INVX1 exu_U15545(.A(exu_n28309), .Y(exu_n3212));
AND2X1 exu_U15546(.A(exu_n27843), .B(exu_n16233), .Y(exu_n28311));
INVX1 exu_U15547(.A(exu_n28311), .Y(exu_n3213));
AND2X1 exu_U15548(.A(exu_n27975), .B(exu_n15401), .Y(exu_n28314));
INVX1 exu_U15549(.A(exu_n28314), .Y(exu_n3214));
AND2X1 exu_U15550(.A(exu_n27976), .B(exu_n15401), .Y(exu_n28318));
INVX1 exu_U15551(.A(exu_n28318), .Y(exu_n3215));
AND2X1 exu_U15552(.A(exu_n16224), .B(shft_lshift4_b1[9]), .Y(exu_n28324));
INVX1 exu_U15553(.A(exu_n28324), .Y(exu_n3216));
AND2X1 exu_U15554(.A(exu_n15402), .B(exu_n15693), .Y(exu_n28326));
INVX1 exu_U15555(.A(exu_n28326), .Y(exu_n3217));
AND2X1 exu_U15556(.A(shft_lshift4_b1[8]), .B(exu_n16224), .Y(exu_n28330));
INVX1 exu_U15557(.A(exu_n28330), .Y(exu_n3218));
AND2X1 exu_U15558(.A(exu_n15695), .B(exu_n15402), .Y(exu_n28332));
INVX1 exu_U15559(.A(exu_n28332), .Y(exu_n3219));
AND2X1 exu_U15560(.A(exu_n15693), .B(exu_n16224), .Y(exu_n28336));
INVX1 exu_U15561(.A(exu_n28336), .Y(exu_n3220));
AND2X1 exu_U15562(.A(exu_n15719), .B(exu_n16227), .Y(exu_n28338));
INVX1 exu_U15563(.A(exu_n28338), .Y(exu_n3221));
AND2X1 exu_U15564(.A(exu_n15695), .B(exu_n16224), .Y(exu_n28342));
INVX1 exu_U15565(.A(exu_n28342), .Y(exu_n3222));
AND2X1 exu_U15566(.A(exu_n15720), .B(exu_n15402), .Y(exu_n28344));
INVX1 exu_U15567(.A(exu_n28344), .Y(exu_n3223));
AND2X1 exu_U15568(.A(shft_lshift4_b1[63]), .B(exu_n16223), .Y(exu_n28348));
INVX1 exu_U15569(.A(exu_n28348), .Y(exu_n3224));
AND2X1 exu_U15570(.A(shft_lshift4_b1[61]), .B(exu_n16227), .Y(exu_n28350));
INVX1 exu_U15571(.A(exu_n28350), .Y(exu_n3225));
AND2X1 exu_U15572(.A(shft_lshift4_b1[62]), .B(exu_n16223), .Y(exu_n28354));
INVX1 exu_U15573(.A(exu_n28354), .Y(exu_n3226));
AND2X1 exu_U15574(.A(shft_lshift4_b1[60]), .B(exu_n15402), .Y(exu_n28356));
INVX1 exu_U15575(.A(exu_n28356), .Y(exu_n3227));
AND2X1 exu_U15576(.A(shft_lshift4_b1[61]), .B(exu_n16224), .Y(exu_n28360));
INVX1 exu_U15577(.A(exu_n28360), .Y(exu_n3228));
AND2X1 exu_U15578(.A(shft_lshift4_b1[59]), .B(exu_n15402), .Y(exu_n28362));
INVX1 exu_U15579(.A(exu_n28362), .Y(exu_n3229));
AND2X1 exu_U15580(.A(shft_lshift4_b1[60]), .B(exu_n16224), .Y(exu_n28366));
INVX1 exu_U15581(.A(exu_n28366), .Y(exu_n3230));
AND2X1 exu_U15582(.A(shft_lshift4_b1[58]), .B(exu_n15402), .Y(exu_n28368));
INVX1 exu_U15583(.A(exu_n28368), .Y(exu_n3231));
AND2X1 exu_U15584(.A(exu_n15719), .B(exu_n16223), .Y(exu_n28372));
INVX1 exu_U15585(.A(exu_n28372), .Y(exu_n3232));
AND2X1 exu_U15586(.A(exu_n28142), .B(exu_n16227), .Y(exu_n28374));
INVX1 exu_U15587(.A(exu_n28374), .Y(exu_n3233));
AND2X1 exu_U15588(.A(shft_lshift4_b1[59]), .B(exu_n16224), .Y(exu_n28378));
INVX1 exu_U15589(.A(exu_n28378), .Y(exu_n3234));
AND2X1 exu_U15590(.A(shft_lshift4_b1[57]), .B(exu_n15402), .Y(exu_n28380));
INVX1 exu_U15591(.A(exu_n28380), .Y(exu_n3235));
AND2X1 exu_U15592(.A(shft_lshift4_b1[58]), .B(exu_n16223), .Y(exu_n28384));
INVX1 exu_U15593(.A(exu_n28384), .Y(exu_n3236));
AND2X1 exu_U15594(.A(shft_lshift4_b1[56]), .B(exu_n15402), .Y(exu_n28386));
INVX1 exu_U15595(.A(exu_n28386), .Y(exu_n3237));
AND2X1 exu_U15596(.A(shft_lshift4_b1[57]), .B(exu_n16224), .Y(exu_n28390));
INVX1 exu_U15597(.A(exu_n28390), .Y(exu_n3238));
AND2X1 exu_U15598(.A(shft_lshift4_b1[55]), .B(exu_n15402), .Y(exu_n28392));
INVX1 exu_U15599(.A(exu_n28392), .Y(exu_n3239));
AND2X1 exu_U15600(.A(shft_lshift4_b1[56]), .B(exu_n16224), .Y(exu_n28396));
INVX1 exu_U15601(.A(exu_n28396), .Y(exu_n3240));
AND2X1 exu_U15602(.A(shft_lshift4_b1[54]), .B(exu_n15402), .Y(exu_n28398));
INVX1 exu_U15603(.A(exu_n28398), .Y(exu_n3241));
AND2X1 exu_U15604(.A(shft_lshift4_b1[55]), .B(exu_n16223), .Y(exu_n28402));
INVX1 exu_U15605(.A(exu_n28402), .Y(exu_n3242));
AND2X1 exu_U15606(.A(shft_lshift4_b1[53]), .B(exu_n15402), .Y(exu_n28404));
INVX1 exu_U15607(.A(exu_n28404), .Y(exu_n3243));
AND2X1 exu_U15608(.A(shft_lshift4_b1[54]), .B(exu_n16223), .Y(exu_n28408));
INVX1 exu_U15609(.A(exu_n28408), .Y(exu_n3244));
AND2X1 exu_U15610(.A(shft_lshift4_b1[52]), .B(exu_n16227), .Y(exu_n28410));
INVX1 exu_U15611(.A(exu_n28410), .Y(exu_n3245));
AND2X1 exu_U15612(.A(shft_lshift4_b1[53]), .B(exu_n16224), .Y(exu_n28414));
INVX1 exu_U15613(.A(exu_n28414), .Y(exu_n3246));
AND2X1 exu_U15614(.A(shft_lshift4_b1[51]), .B(exu_n16227), .Y(exu_n28416));
INVX1 exu_U15615(.A(exu_n28416), .Y(exu_n3247));
AND2X1 exu_U15616(.A(shft_lshift4_b1[52]), .B(exu_n16224), .Y(exu_n28420));
INVX1 exu_U15617(.A(exu_n28420), .Y(exu_n3248));
AND2X1 exu_U15618(.A(shft_lshift4_b1[50]), .B(exu_n15402), .Y(exu_n28422));
INVX1 exu_U15619(.A(exu_n28422), .Y(exu_n3249));
AND2X1 exu_U15620(.A(shft_lshift4_b1[51]), .B(exu_n16223), .Y(exu_n28426));
INVX1 exu_U15621(.A(exu_n28426), .Y(exu_n3250));
AND2X1 exu_U15622(.A(shft_lshift4_b1[49]), .B(exu_n16227), .Y(exu_n28428));
INVX1 exu_U15623(.A(exu_n28428), .Y(exu_n3251));
AND2X1 exu_U15624(.A(shft_lshift4_b1[50]), .B(exu_n16223), .Y(exu_n28432));
INVX1 exu_U15625(.A(exu_n28432), .Y(exu_n3252));
AND2X1 exu_U15626(.A(shft_lshift4_b1[48]), .B(exu_n15402), .Y(exu_n28434));
INVX1 exu_U15627(.A(exu_n28434), .Y(exu_n3253));
AND2X1 exu_U15628(.A(exu_n15720), .B(exu_n16224), .Y(exu_n28438));
INVX1 exu_U15629(.A(exu_n28438), .Y(exu_n3254));
AND2X1 exu_U15630(.A(exu_n28203), .B(exu_n16227), .Y(exu_n28440));
INVX1 exu_U15631(.A(exu_n28440), .Y(exu_n3255));
AND2X1 exu_U15632(.A(shft_lshift4_b1[49]), .B(exu_n16224), .Y(exu_n28444));
INVX1 exu_U15633(.A(exu_n28444), .Y(exu_n3256));
AND2X1 exu_U15634(.A(shft_lshift4_b1[47]), .B(exu_n15402), .Y(exu_n28446));
INVX1 exu_U15635(.A(exu_n28446), .Y(exu_n3257));
AND2X1 exu_U15636(.A(shft_lshift4_b1[48]), .B(exu_n16223), .Y(exu_n28450));
INVX1 exu_U15637(.A(exu_n28450), .Y(exu_n3258));
AND2X1 exu_U15638(.A(shft_lshift4_b1[46]), .B(exu_n15402), .Y(exu_n28452));
INVX1 exu_U15639(.A(exu_n28452), .Y(exu_n3259));
AND2X1 exu_U15640(.A(shft_lshift4_b1[47]), .B(exu_n16224), .Y(exu_n28456));
INVX1 exu_U15641(.A(exu_n28456), .Y(exu_n3260));
AND2X1 exu_U15642(.A(shft_lshift4_b1[45]), .B(exu_n15402), .Y(exu_n28458));
INVX1 exu_U15643(.A(exu_n28458), .Y(exu_n3261));
AND2X1 exu_U15644(.A(shft_lshift4_b1[46]), .B(exu_n16223), .Y(exu_n28462));
INVX1 exu_U15645(.A(exu_n28462), .Y(exu_n3262));
AND2X1 exu_U15646(.A(shft_lshift4_b1[44]), .B(exu_n16227), .Y(exu_n28464));
INVX1 exu_U15647(.A(exu_n28464), .Y(exu_n3263));
AND2X1 exu_U15648(.A(shft_lshift4_b1[45]), .B(exu_n16223), .Y(exu_n28468));
INVX1 exu_U15649(.A(exu_n28468), .Y(exu_n3264));
AND2X1 exu_U15650(.A(shft_lshift4_b1[43]), .B(exu_n16227), .Y(exu_n28470));
INVX1 exu_U15651(.A(exu_n28470), .Y(exu_n3265));
AND2X1 exu_U15652(.A(shft_lshift4_b1[44]), .B(exu_n16224), .Y(exu_n28474));
INVX1 exu_U15653(.A(exu_n28474), .Y(exu_n3266));
AND2X1 exu_U15654(.A(shft_lshift4_b1[42]), .B(exu_n16227), .Y(exu_n28476));
INVX1 exu_U15655(.A(exu_n28476), .Y(exu_n3267));
AND2X1 exu_U15656(.A(shft_lshift4_b1[43]), .B(exu_n16224), .Y(exu_n28480));
INVX1 exu_U15657(.A(exu_n28480), .Y(exu_n3268));
AND2X1 exu_U15658(.A(shft_lshift4_b1[41]), .B(exu_n15402), .Y(exu_n28482));
INVX1 exu_U15659(.A(exu_n28482), .Y(exu_n3269));
AND2X1 exu_U15660(.A(shft_lshift4_b1[42]), .B(exu_n16223), .Y(exu_n28486));
INVX1 exu_U15661(.A(exu_n28486), .Y(exu_n3270));
AND2X1 exu_U15662(.A(shft_lshift4_b1[40]), .B(exu_n15402), .Y(exu_n28488));
INVX1 exu_U15663(.A(exu_n28488), .Y(exu_n3271));
AND2X1 exu_U15664(.A(shft_lshift4_b1[41]), .B(exu_n16224), .Y(exu_n28492));
INVX1 exu_U15665(.A(exu_n28492), .Y(exu_n3272));
AND2X1 exu_U15666(.A(shft_lshift4_b1[39]), .B(exu_n16227), .Y(exu_n28494));
INVX1 exu_U15667(.A(exu_n28494), .Y(exu_n3273));
AND2X1 exu_U15668(.A(shft_lshift4_b1[40]), .B(exu_n16224), .Y(exu_n28498));
INVX1 exu_U15669(.A(exu_n28498), .Y(exu_n3274));
AND2X1 exu_U15670(.A(shft_lshift4_b1[38]), .B(exu_n16227), .Y(exu_n28500));
INVX1 exu_U15671(.A(exu_n28500), .Y(exu_n3275));
AND2X1 exu_U15672(.A(exu_n28142), .B(exu_n16223), .Y(exu_n28504));
INVX1 exu_U15673(.A(exu_n28504), .Y(exu_n3276));
AND2X1 exu_U15674(.A(exu_n28264), .B(exu_n15402), .Y(exu_n28506));
INVX1 exu_U15675(.A(exu_n28506), .Y(exu_n3277));
AND2X1 exu_U15676(.A(shft_lshift4_b1[39]), .B(exu_n16224), .Y(exu_n28510));
INVX1 exu_U15677(.A(exu_n28510), .Y(exu_n3278));
AND2X1 exu_U15678(.A(shft_lshift4_b1[37]), .B(exu_n15402), .Y(exu_n28512));
INVX1 exu_U15679(.A(exu_n28512), .Y(exu_n3279));
AND2X1 exu_U15680(.A(shft_lshift4_b1[38]), .B(exu_n16224), .Y(exu_n28516));
INVX1 exu_U15681(.A(exu_n28516), .Y(exu_n3280));
AND2X1 exu_U15682(.A(shft_lshift4_b1[36]), .B(exu_n15402), .Y(exu_n28518));
INVX1 exu_U15683(.A(exu_n28518), .Y(exu_n3281));
AND2X1 exu_U15684(.A(shft_lshift4_b1[37]), .B(exu_n16224), .Y(exu_n28522));
INVX1 exu_U15685(.A(exu_n28522), .Y(exu_n3282));
AND2X1 exu_U15686(.A(shft_lshift4_b1[35]), .B(exu_n15402), .Y(exu_n28524));
INVX1 exu_U15687(.A(exu_n28524), .Y(exu_n3283));
AND2X1 exu_U15688(.A(shft_lshift4_b1[36]), .B(exu_n16224), .Y(exu_n28528));
INVX1 exu_U15689(.A(exu_n28528), .Y(exu_n3284));
AND2X1 exu_U15690(.A(shft_lshift4_b1[34]), .B(exu_n15402), .Y(exu_n28530));
INVX1 exu_U15691(.A(exu_n28530), .Y(exu_n3285));
AND2X1 exu_U15692(.A(shft_lshift4_b1[35]), .B(exu_n16223), .Y(exu_n28534));
INVX1 exu_U15693(.A(exu_n28534), .Y(exu_n3286));
AND2X1 exu_U15694(.A(shft_lshift4_b1[33]), .B(exu_n15402), .Y(exu_n28536));
INVX1 exu_U15695(.A(exu_n28536), .Y(exu_n3287));
AND2X1 exu_U15696(.A(shft_lshift4_b1[34]), .B(exu_n16223), .Y(exu_n28540));
INVX1 exu_U15697(.A(exu_n28540), .Y(exu_n3288));
AND2X1 exu_U15698(.A(shft_lshift4_b1[32]), .B(exu_n15402), .Y(exu_n28542));
INVX1 exu_U15699(.A(exu_n28542), .Y(exu_n3289));
AND2X1 exu_U15700(.A(shft_lshift4_b1[33]), .B(exu_n16224), .Y(exu_n28546));
INVX1 exu_U15701(.A(exu_n28546), .Y(exu_n3290));
AND2X1 exu_U15702(.A(shft_lshift4_b1[31]), .B(exu_n16227), .Y(exu_n28548));
INVX1 exu_U15703(.A(exu_n28548), .Y(exu_n3291));
AND2X1 exu_U15704(.A(shft_lshift4_b1[32]), .B(exu_n16223), .Y(exu_n28552));
INVX1 exu_U15705(.A(exu_n28552), .Y(exu_n3292));
AND2X1 exu_U15706(.A(shft_lshift4_b1[30]), .B(exu_n15402), .Y(exu_n28554));
INVX1 exu_U15707(.A(exu_n28554), .Y(exu_n3293));
AND2X1 exu_U15708(.A(shft_lshift4_b1[31]), .B(exu_n16223), .Y(exu_n28558));
INVX1 exu_U15709(.A(exu_n28558), .Y(exu_n3294));
AND2X1 exu_U15710(.A(shft_lshift4_b1[29]), .B(exu_n16227), .Y(exu_n28560));
INVX1 exu_U15711(.A(exu_n28560), .Y(exu_n3295));
AND2X1 exu_U15712(.A(shft_lshift4_b1[30]), .B(exu_n16224), .Y(exu_n28564));
INVX1 exu_U15713(.A(exu_n28564), .Y(exu_n3296));
AND2X1 exu_U15714(.A(shft_lshift4_b1[28]), .B(exu_n16227), .Y(exu_n28566));
INVX1 exu_U15715(.A(exu_n28566), .Y(exu_n3297));
AND2X1 exu_U15716(.A(exu_n28203), .B(exu_n16223), .Y(exu_n28569));
INVX1 exu_U15717(.A(exu_n28569), .Y(exu_n3298));
AND2X1 exu_U15718(.A(shft_lshift4_b1[29]), .B(exu_n16224), .Y(exu_n28574));
INVX1 exu_U15719(.A(exu_n28574), .Y(exu_n3299));
AND2X1 exu_U15720(.A(shft_lshift4_b1[27]), .B(exu_n16227), .Y(exu_n28576));
INVX1 exu_U15721(.A(exu_n28576), .Y(exu_n3300));
AND2X1 exu_U15722(.A(shft_lshift4_b1[28]), .B(exu_n16224), .Y(exu_n28580));
INVX1 exu_U15723(.A(exu_n28580), .Y(exu_n3301));
AND2X1 exu_U15724(.A(shft_lshift4_b1[26]), .B(exu_n16227), .Y(exu_n28582));
INVX1 exu_U15725(.A(exu_n28582), .Y(exu_n3302));
AND2X1 exu_U15726(.A(shft_lshift4_b1[27]), .B(exu_n16224), .Y(exu_n28586));
INVX1 exu_U15727(.A(exu_n28586), .Y(exu_n3303));
AND2X1 exu_U15728(.A(shft_lshift4_b1[25]), .B(exu_n15402), .Y(exu_n28588));
INVX1 exu_U15729(.A(exu_n28588), .Y(exu_n3304));
AND2X1 exu_U15730(.A(shft_lshift4_b1[26]), .B(exu_n16223), .Y(exu_n28592));
INVX1 exu_U15731(.A(exu_n28592), .Y(exu_n3305));
AND2X1 exu_U15732(.A(shft_lshift4_b1[24]), .B(exu_n15402), .Y(exu_n28594));
INVX1 exu_U15733(.A(exu_n28594), .Y(exu_n3306));
AND2X1 exu_U15734(.A(shft_lshift4_b1[25]), .B(exu_n16223), .Y(exu_n28598));
INVX1 exu_U15735(.A(exu_n28598), .Y(exu_n3307));
AND2X1 exu_U15736(.A(shft_lshift4_b1[23]), .B(exu_n16227), .Y(exu_n28600));
INVX1 exu_U15737(.A(exu_n28600), .Y(exu_n3308));
AND2X1 exu_U15738(.A(shft_lshift4_b1[24]), .B(exu_n16223), .Y(exu_n28604));
INVX1 exu_U15739(.A(exu_n28604), .Y(exu_n3309));
AND2X1 exu_U15740(.A(shft_lshift4_b1[22]), .B(exu_n16227), .Y(exu_n28606));
INVX1 exu_U15741(.A(exu_n28606), .Y(exu_n3310));
AND2X1 exu_U15742(.A(shft_lshift4_b1[23]), .B(exu_n16224), .Y(exu_n28610));
INVX1 exu_U15743(.A(exu_n28610), .Y(exu_n3311));
AND2X1 exu_U15744(.A(shft_lshift4_b1[21]), .B(exu_n15402), .Y(exu_n28612));
INVX1 exu_U15745(.A(exu_n28612), .Y(exu_n3312));
AND2X1 exu_U15746(.A(shft_lshift4_b1[22]), .B(exu_n16223), .Y(exu_n28616));
INVX1 exu_U15747(.A(exu_n28616), .Y(exu_n3313));
AND2X1 exu_U15748(.A(shft_lshift4_b1[20]), .B(exu_n15402), .Y(exu_n28618));
INVX1 exu_U15749(.A(exu_n28618), .Y(exu_n3314));
AND2X1 exu_U15750(.A(shft_lshift4_b1[21]), .B(exu_n16223), .Y(exu_n28622));
INVX1 exu_U15751(.A(exu_n28622), .Y(exu_n3315));
AND2X1 exu_U15752(.A(shft_lshift4_b1[19]), .B(exu_n16227), .Y(exu_n28624));
INVX1 exu_U15753(.A(exu_n28624), .Y(exu_n3316));
AND2X1 exu_U15754(.A(shft_lshift4_b1[20]), .B(exu_n16223), .Y(exu_n28628));
INVX1 exu_U15755(.A(exu_n28628), .Y(exu_n3317));
AND2X1 exu_U15756(.A(shft_lshift4_b1[18]), .B(exu_n15402), .Y(exu_n28630));
INVX1 exu_U15757(.A(exu_n28630), .Y(exu_n3318));
AND2X1 exu_U15758(.A(shft_lshift4_b1[19]), .B(exu_n16223), .Y(exu_n28637));
INVX1 exu_U15759(.A(exu_n28637), .Y(exu_n3319));
AND2X1 exu_U15760(.A(shft_lshift4_b1[17]), .B(exu_n16227), .Y(exu_n28639));
INVX1 exu_U15761(.A(exu_n28639), .Y(exu_n3320));
AND2X1 exu_U15762(.A(shft_lshift4_b1[18]), .B(exu_n16223), .Y(exu_n28643));
INVX1 exu_U15763(.A(exu_n28643), .Y(exu_n3321));
AND2X1 exu_U15764(.A(shft_lshift4_b1[16]), .B(exu_n16227), .Y(exu_n28645));
INVX1 exu_U15765(.A(exu_n28645), .Y(exu_n3322));
AND2X1 exu_U15766(.A(shft_lshift4_b1[17]), .B(exu_n16223), .Y(exu_n28649));
INVX1 exu_U15767(.A(exu_n28649), .Y(exu_n3323));
AND2X1 exu_U15768(.A(shft_lshift4_b1[15]), .B(exu_n15402), .Y(exu_n28651));
INVX1 exu_U15769(.A(exu_n28651), .Y(exu_n3324));
AND2X1 exu_U15770(.A(shft_lshift4_b1[16]), .B(exu_n16223), .Y(exu_n28655));
INVX1 exu_U15771(.A(exu_n28655), .Y(exu_n3325));
AND2X1 exu_U15772(.A(shft_lshift4_b1[14]), .B(exu_n16227), .Y(exu_n28657));
INVX1 exu_U15773(.A(exu_n28657), .Y(exu_n3326));
AND2X1 exu_U15774(.A(shft_lshift4_b1[15]), .B(exu_n16223), .Y(exu_n28661));
INVX1 exu_U15775(.A(exu_n28661), .Y(exu_n3327));
AND2X1 exu_U15776(.A(shft_lshift4_b1[13]), .B(exu_n15402), .Y(exu_n28663));
INVX1 exu_U15777(.A(exu_n28663), .Y(exu_n3328));
AND2X1 exu_U15778(.A(shft_lshift4_b1[14]), .B(exu_n16223), .Y(exu_n28667));
INVX1 exu_U15779(.A(exu_n28667), .Y(exu_n3329));
AND2X1 exu_U15780(.A(shft_lshift4_b1[12]), .B(exu_n15402), .Y(exu_n28669));
INVX1 exu_U15781(.A(exu_n28669), .Y(exu_n3330));
AND2X1 exu_U15782(.A(shft_lshift4_b1[13]), .B(exu_n16223), .Y(exu_n28673));
INVX1 exu_U15783(.A(exu_n28673), .Y(exu_n3331));
AND2X1 exu_U15784(.A(shft_lshift4_b1[11]), .B(exu_n16227), .Y(exu_n28675));
INVX1 exu_U15785(.A(exu_n28675), .Y(exu_n3332));
AND2X1 exu_U15786(.A(shft_lshift4_b1[12]), .B(exu_n16223), .Y(exu_n28679));
INVX1 exu_U15787(.A(exu_n28679), .Y(exu_n3333));
AND2X1 exu_U15788(.A(shft_lshift4_b1[10]), .B(exu_n16227), .Y(exu_n28681));
INVX1 exu_U15789(.A(exu_n28681), .Y(exu_n3334));
AND2X1 exu_U15790(.A(shft_lshift4_b1[11]), .B(exu_n16223), .Y(exu_n28685));
INVX1 exu_U15791(.A(exu_n28685), .Y(exu_n3335));
AND2X1 exu_U15792(.A(shft_lshift4_b1[9]), .B(exu_n15402), .Y(exu_n28687));
INVX1 exu_U15793(.A(exu_n28687), .Y(exu_n3336));
AND2X1 exu_U15794(.A(shft_lshift4_b1[10]), .B(exu_n16223), .Y(exu_n28691));
INVX1 exu_U15795(.A(exu_n28691), .Y(exu_n3337));
AND2X1 exu_U15796(.A(shft_lshift4_b1[8]), .B(exu_n16227), .Y(exu_n28693));
INVX1 exu_U15797(.A(exu_n28693), .Y(exu_n3338));
AND2X1 exu_U15798(.A(exu_n16248), .B(div_neg32[9]), .Y(exu_n28698));
INVX1 exu_U15799(.A(exu_n28698), .Y(exu_n3339));
AND2X1 exu_U15800(.A(exu_n16247), .B(exu_n10695), .Y(exu_n28700));
INVX1 exu_U15801(.A(exu_n28700), .Y(exu_n3340));
AND2X1 exu_U15802(.A(div_neg32[8]), .B(exu_n16248), .Y(exu_n28704));
INVX1 exu_U15803(.A(exu_n28704), .Y(exu_n3341));
AND2X1 exu_U15804(.A(exu_n11861), .B(exu_n16247), .Y(exu_n28706));
INVX1 exu_U15805(.A(exu_n28706), .Y(exu_n3342));
AND2X1 exu_U15806(.A(div_neg32[7]), .B(ecl_div_sel_neg32), .Y(exu_n28710));
INVX1 exu_U15807(.A(exu_n28710), .Y(exu_n3343));
AND2X1 exu_U15808(.A(exu_n11862), .B(exu_n16247), .Y(exu_n28712));
INVX1 exu_U15809(.A(exu_n28712), .Y(exu_n3344));
AND2X1 exu_U15810(.A(div_neg32[6]), .B(ecl_div_sel_neg32), .Y(exu_n28716));
INVX1 exu_U15811(.A(exu_n28716), .Y(exu_n3345));
AND2X1 exu_U15812(.A(exu_n11863), .B(exu_n16247), .Y(exu_n28718));
INVX1 exu_U15813(.A(exu_n28718), .Y(exu_n3346));
AND2X1 exu_U15814(.A(div_neg32[5]), .B(exu_n16248), .Y(exu_n28726));
INVX1 exu_U15815(.A(exu_n28726), .Y(exu_n3347));
AND2X1 exu_U15816(.A(exu_n11864), .B(exu_n16247), .Y(exu_n28728));
INVX1 exu_U15817(.A(exu_n28728), .Y(exu_n3348));
AND2X1 exu_U15818(.A(div_neg32[4]), .B(ecl_div_sel_neg32), .Y(exu_n28742));
INVX1 exu_U15819(.A(exu_n28742), .Y(exu_n3349));
AND2X1 exu_U15820(.A(exu_n11865), .B(exu_n16247), .Y(exu_n28744));
INVX1 exu_U15821(.A(exu_n28744), .Y(exu_n3350));
AND2X1 exu_U15822(.A(div_neg32[3]), .B(ecl_div_sel_neg32), .Y(exu_n28758));
INVX1 exu_U15823(.A(exu_n28758), .Y(exu_n3351));
AND2X1 exu_U15824(.A(exu_n11866), .B(exu_n16247), .Y(exu_n28760));
INVX1 exu_U15825(.A(exu_n28760), .Y(exu_n3352));
AND2X1 exu_U15826(.A(exu_n11867), .B(exu_n16247), .Y(exu_n28771));
INVX1 exu_U15827(.A(exu_n28771), .Y(exu_n3353));
AND2X1 exu_U15828(.A(div_neg32[30]), .B(exu_n16248), .Y(exu_n28775));
INVX1 exu_U15829(.A(exu_n28775), .Y(exu_n3354));
AND2X1 exu_U15830(.A(exu_n11868), .B(exu_n16247), .Y(exu_n28777));
INVX1 exu_U15831(.A(exu_n28777), .Y(exu_n3355));
AND2X1 exu_U15832(.A(div_neg32[2]), .B(ecl_div_sel_neg32), .Y(exu_n28781));
INVX1 exu_U15833(.A(exu_n28781), .Y(exu_n3356));
AND2X1 exu_U15834(.A(exu_n11869), .B(exu_n16247), .Y(exu_n28783));
INVX1 exu_U15835(.A(exu_n28783), .Y(exu_n3357));
AND2X1 exu_U15836(.A(div_neg32[29]), .B(ecl_div_sel_neg32), .Y(exu_n28787));
INVX1 exu_U15837(.A(exu_n28787), .Y(exu_n3358));
AND2X1 exu_U15838(.A(exu_n11870), .B(exu_n16247), .Y(exu_n28789));
INVX1 exu_U15839(.A(exu_n28789), .Y(exu_n3359));
AND2X1 exu_U15840(.A(div_neg32[28]), .B(exu_n16248), .Y(exu_n28793));
INVX1 exu_U15841(.A(exu_n28793), .Y(exu_n3360));
AND2X1 exu_U15842(.A(exu_n11871), .B(exu_n16247), .Y(exu_n28795));
INVX1 exu_U15843(.A(exu_n28795), .Y(exu_n3361));
AND2X1 exu_U15844(.A(div_neg32[27]), .B(ecl_div_sel_neg32), .Y(exu_n28799));
INVX1 exu_U15845(.A(exu_n28799), .Y(exu_n3362));
AND2X1 exu_U15846(.A(exu_n11872), .B(exu_n16247), .Y(exu_n28801));
INVX1 exu_U15847(.A(exu_n28801), .Y(exu_n3363));
AND2X1 exu_U15848(.A(div_neg32[26]), .B(ecl_div_sel_neg32), .Y(exu_n28805));
INVX1 exu_U15849(.A(exu_n28805), .Y(exu_n3364));
AND2X1 exu_U15850(.A(exu_n11873), .B(exu_n16247), .Y(exu_n28807));
INVX1 exu_U15851(.A(exu_n28807), .Y(exu_n3365));
AND2X1 exu_U15852(.A(div_neg32[25]), .B(exu_n16248), .Y(exu_n28811));
INVX1 exu_U15853(.A(exu_n28811), .Y(exu_n3366));
AND2X1 exu_U15854(.A(exu_n11874), .B(exu_n16247), .Y(exu_n28813));
INVX1 exu_U15855(.A(exu_n28813), .Y(exu_n3367));
AND2X1 exu_U15856(.A(div_neg32[24]), .B(exu_n16248), .Y(exu_n28817));
INVX1 exu_U15857(.A(exu_n28817), .Y(exu_n3368));
AND2X1 exu_U15858(.A(exu_n11875), .B(exu_n16247), .Y(exu_n28819));
INVX1 exu_U15859(.A(exu_n28819), .Y(exu_n3369));
AND2X1 exu_U15860(.A(div_neg32[23]), .B(exu_n16248), .Y(exu_n28823));
INVX1 exu_U15861(.A(exu_n28823), .Y(exu_n3370));
AND2X1 exu_U15862(.A(exu_n11876), .B(exu_n16247), .Y(exu_n28825));
INVX1 exu_U15863(.A(exu_n28825), .Y(exu_n3371));
AND2X1 exu_U15864(.A(div_neg32[22]), .B(exu_n16248), .Y(exu_n28829));
INVX1 exu_U15865(.A(exu_n28829), .Y(exu_n3372));
AND2X1 exu_U15866(.A(exu_n11877), .B(exu_n16247), .Y(exu_n28831));
INVX1 exu_U15867(.A(exu_n28831), .Y(exu_n3373));
AND2X1 exu_U15868(.A(div_neg32[21]), .B(exu_n16248), .Y(exu_n28835));
INVX1 exu_U15869(.A(exu_n28835), .Y(exu_n3374));
AND2X1 exu_U15870(.A(exu_n11878), .B(exu_n16247), .Y(exu_n28837));
INVX1 exu_U15871(.A(exu_n28837), .Y(exu_n3375));
AND2X1 exu_U15872(.A(div_neg32[20]), .B(exu_n16248), .Y(exu_n28841));
INVX1 exu_U15873(.A(exu_n28841), .Y(exu_n3376));
AND2X1 exu_U15874(.A(exu_n11879), .B(exu_n16247), .Y(exu_n28843));
INVX1 exu_U15875(.A(exu_n28843), .Y(exu_n3377));
AND2X1 exu_U15876(.A(div_neg32[1]), .B(exu_n16248), .Y(exu_n28847));
INVX1 exu_U15877(.A(exu_n28847), .Y(exu_n3378));
AND2X1 exu_U15878(.A(exu_n11880), .B(exu_n16247), .Y(exu_n28849));
INVX1 exu_U15879(.A(exu_n28849), .Y(exu_n3379));
AND2X1 exu_U15880(.A(div_neg32[19]), .B(exu_n16248), .Y(exu_n28853));
INVX1 exu_U15881(.A(exu_n28853), .Y(exu_n3380));
AND2X1 exu_U15882(.A(exu_n11881), .B(exu_n16247), .Y(exu_n28855));
INVX1 exu_U15883(.A(exu_n28855), .Y(exu_n3381));
AND2X1 exu_U15884(.A(div_neg32[18]), .B(exu_n16248), .Y(exu_n28859));
INVX1 exu_U15885(.A(exu_n28859), .Y(exu_n3382));
AND2X1 exu_U15886(.A(exu_n11882), .B(exu_n16247), .Y(exu_n28861));
INVX1 exu_U15887(.A(exu_n28861), .Y(exu_n3383));
AND2X1 exu_U15888(.A(div_neg32[17]), .B(exu_n16248), .Y(exu_n28865));
INVX1 exu_U15889(.A(exu_n28865), .Y(exu_n3384));
AND2X1 exu_U15890(.A(exu_n11883), .B(exu_n16247), .Y(exu_n28867));
INVX1 exu_U15891(.A(exu_n28867), .Y(exu_n3385));
AND2X1 exu_U15892(.A(div_neg32[16]), .B(exu_n16248), .Y(exu_n28871));
INVX1 exu_U15893(.A(exu_n28871), .Y(exu_n3386));
AND2X1 exu_U15894(.A(exu_n11884), .B(exu_n16247), .Y(exu_n28873));
INVX1 exu_U15895(.A(exu_n28873), .Y(exu_n3387));
AND2X1 exu_U15896(.A(div_neg32[15]), .B(exu_n16248), .Y(exu_n28877));
INVX1 exu_U15897(.A(exu_n28877), .Y(exu_n3388));
AND2X1 exu_U15898(.A(exu_n11885), .B(exu_n16247), .Y(exu_n28879));
INVX1 exu_U15899(.A(exu_n28879), .Y(exu_n3389));
AND2X1 exu_U15900(.A(div_neg32[14]), .B(exu_n16248), .Y(exu_n28883));
INVX1 exu_U15901(.A(exu_n28883), .Y(exu_n3390));
AND2X1 exu_U15902(.A(exu_n11886), .B(exu_n16247), .Y(exu_n28885));
INVX1 exu_U15903(.A(exu_n28885), .Y(exu_n3391));
AND2X1 exu_U15904(.A(div_neg32[13]), .B(exu_n16248), .Y(exu_n28889));
INVX1 exu_U15905(.A(exu_n28889), .Y(exu_n3392));
AND2X1 exu_U15906(.A(exu_n11887), .B(exu_n16247), .Y(exu_n28891));
INVX1 exu_U15907(.A(exu_n28891), .Y(exu_n3393));
AND2X1 exu_U15908(.A(div_neg32[12]), .B(exu_n16248), .Y(exu_n28895));
INVX1 exu_U15909(.A(exu_n28895), .Y(exu_n3394));
AND2X1 exu_U15910(.A(exu_n11888), .B(exu_n16247), .Y(exu_n28897));
INVX1 exu_U15911(.A(exu_n28897), .Y(exu_n3395));
AND2X1 exu_U15912(.A(div_neg32[11]), .B(exu_n16248), .Y(exu_n28901));
INVX1 exu_U15913(.A(exu_n28901), .Y(exu_n3396));
AND2X1 exu_U15914(.A(exu_n11889), .B(exu_n16247), .Y(exu_n28903));
INVX1 exu_U15915(.A(exu_n28903), .Y(exu_n3397));
AND2X1 exu_U15916(.A(div_neg32[10]), .B(ecl_div_sel_neg32), .Y(exu_n28907));
INVX1 exu_U15917(.A(exu_n28907), .Y(exu_n3398));
AND2X1 exu_U15918(.A(exu_n11890), .B(exu_n16247), .Y(exu_n28909));
INVX1 exu_U15919(.A(exu_n28909), .Y(exu_n3399));
AND2X1 exu_U15920(.A(div_neg32[0]), .B(exu_n16248), .Y(exu_n28913));
INVX1 exu_U15921(.A(exu_n28913), .Y(exu_n3400));
AND2X1 exu_U15922(.A(exu_n11891), .B(exu_n16247), .Y(exu_n28915));
INVX1 exu_U15923(.A(exu_n28915), .Y(exu_n3401));
AND2X1 exu_U15924(.A(exu_n16237), .B(div_input_data_e[73]), .Y(exu_n28919));
INVX1 exu_U15925(.A(exu_n28919), .Y(exu_n3402));
AND2X1 exu_U15926(.A(exu_n16239), .B(alu_logic_result_or[9]), .Y(exu_n28921));
INVX1 exu_U15927(.A(exu_n28921), .Y(exu_n3403));
AND2X1 exu_U15928(.A(div_input_data_e[72]), .B(exu_n16237), .Y(exu_n28925));
INVX1 exu_U15929(.A(exu_n28925), .Y(exu_n3404));
AND2X1 exu_U15930(.A(alu_logic_result_or[8]), .B(exu_n16239), .Y(exu_n28927));
INVX1 exu_U15931(.A(exu_n28927), .Y(exu_n3405));
AND2X1 exu_U15932(.A(div_input_data_e[71]), .B(exu_n16237), .Y(exu_n28931));
INVX1 exu_U15933(.A(exu_n28931), .Y(exu_n3406));
AND2X1 exu_U15934(.A(alu_logic_result_or[7]), .B(exu_n16239), .Y(exu_n28933));
INVX1 exu_U15935(.A(exu_n28933), .Y(exu_n3407));
AND2X1 exu_U15936(.A(div_input_data_e[70]), .B(exu_n16237), .Y(exu_n28937));
INVX1 exu_U15937(.A(exu_n28937), .Y(exu_n3408));
AND2X1 exu_U15938(.A(alu_logic_result_or[6]), .B(exu_n16239), .Y(exu_n28939));
INVX1 exu_U15939(.A(exu_n28939), .Y(exu_n3409));
AND2X1 exu_U15940(.A(exu_n11618), .B(exu_n16237), .Y(exu_n28943));
INVX1 exu_U15941(.A(exu_n28943), .Y(exu_n3410));
AND2X1 exu_U15942(.A(alu_logic_result_or[63]), .B(exu_n16239), .Y(exu_n28945));
INVX1 exu_U15943(.A(exu_n28945), .Y(exu_n3411));
AND2X1 exu_U15944(.A(exu_n11619), .B(exu_n16237), .Y(exu_n28949));
INVX1 exu_U15945(.A(exu_n28949), .Y(exu_n3412));
AND2X1 exu_U15946(.A(alu_logic_result_or[62]), .B(exu_n16239), .Y(exu_n28951));
INVX1 exu_U15947(.A(exu_n28951), .Y(exu_n3413));
AND2X1 exu_U15948(.A(exu_n11620), .B(exu_n16237), .Y(exu_n28955));
INVX1 exu_U15949(.A(exu_n28955), .Y(exu_n3414));
AND2X1 exu_U15950(.A(alu_logic_result_or[61]), .B(exu_n16239), .Y(exu_n28957));
INVX1 exu_U15951(.A(exu_n28957), .Y(exu_n3415));
AND2X1 exu_U15952(.A(exu_n11621), .B(exu_n16237), .Y(exu_n28961));
INVX1 exu_U15953(.A(exu_n28961), .Y(exu_n3416));
AND2X1 exu_U15954(.A(alu_logic_result_or[60]), .B(exu_n16239), .Y(exu_n28963));
INVX1 exu_U15955(.A(exu_n28963), .Y(exu_n3417));
AND2X1 exu_U15956(.A(div_input_data_e[69]), .B(exu_n16237), .Y(exu_n28967));
INVX1 exu_U15957(.A(exu_n28967), .Y(exu_n3418));
AND2X1 exu_U15958(.A(alu_logic_result_or[5]), .B(exu_n16239), .Y(exu_n28969));
INVX1 exu_U15959(.A(exu_n28969), .Y(exu_n3419));
AND2X1 exu_U15960(.A(exu_n11622), .B(exu_n16237), .Y(exu_n28973));
INVX1 exu_U15961(.A(exu_n28973), .Y(exu_n3420));
AND2X1 exu_U15962(.A(alu_logic_result_or[59]), .B(exu_n16239), .Y(exu_n28975));
INVX1 exu_U15963(.A(exu_n28975), .Y(exu_n3421));
AND2X1 exu_U15964(.A(exu_n11623), .B(exu_n16237), .Y(exu_n28979));
INVX1 exu_U15965(.A(exu_n28979), .Y(exu_n3422));
AND2X1 exu_U15966(.A(alu_logic_result_or[58]), .B(exu_n16239), .Y(exu_n28981));
INVX1 exu_U15967(.A(exu_n28981), .Y(exu_n3423));
AND2X1 exu_U15968(.A(exu_n11624), .B(exu_n16237), .Y(exu_n28985));
INVX1 exu_U15969(.A(exu_n28985), .Y(exu_n3424));
AND2X1 exu_U15970(.A(alu_logic_result_or[57]), .B(exu_n16239), .Y(exu_n28987));
INVX1 exu_U15971(.A(exu_n28987), .Y(exu_n3425));
AND2X1 exu_U15972(.A(exu_n11625), .B(exu_n16237), .Y(exu_n28991));
INVX1 exu_U15973(.A(exu_n28991), .Y(exu_n3426));
AND2X1 exu_U15974(.A(alu_logic_result_or[56]), .B(exu_n16239), .Y(exu_n28993));
INVX1 exu_U15975(.A(exu_n28993), .Y(exu_n3427));
AND2X1 exu_U15976(.A(exu_n11626), .B(exu_n16237), .Y(exu_n28997));
INVX1 exu_U15977(.A(exu_n28997), .Y(exu_n3428));
AND2X1 exu_U15978(.A(alu_logic_result_or[55]), .B(exu_n16239), .Y(exu_n28999));
INVX1 exu_U15979(.A(exu_n28999), .Y(exu_n3429));
AND2X1 exu_U15980(.A(exu_n11627), .B(exu_n16237), .Y(exu_n29003));
INVX1 exu_U15981(.A(exu_n29003), .Y(exu_n3430));
AND2X1 exu_U15982(.A(alu_logic_result_or[54]), .B(exu_n16239), .Y(exu_n29005));
INVX1 exu_U15983(.A(exu_n29005), .Y(exu_n3431));
AND2X1 exu_U15984(.A(exu_n11628), .B(exu_n16237), .Y(exu_n29009));
INVX1 exu_U15985(.A(exu_n29009), .Y(exu_n3432));
AND2X1 exu_U15986(.A(alu_logic_result_or[53]), .B(exu_n16239), .Y(exu_n29011));
INVX1 exu_U15987(.A(exu_n29011), .Y(exu_n3433));
AND2X1 exu_U15988(.A(exu_n11629), .B(exu_n16237), .Y(exu_n29015));
INVX1 exu_U15989(.A(exu_n29015), .Y(exu_n3434));
AND2X1 exu_U15990(.A(alu_logic_result_or[52]), .B(exu_n16239), .Y(exu_n29017));
INVX1 exu_U15991(.A(exu_n29017), .Y(exu_n3435));
AND2X1 exu_U15992(.A(exu_n11630), .B(exu_n16237), .Y(exu_n29021));
INVX1 exu_U15993(.A(exu_n29021), .Y(exu_n3436));
AND2X1 exu_U15994(.A(alu_logic_result_or[51]), .B(exu_n16239), .Y(exu_n29023));
INVX1 exu_U15995(.A(exu_n29023), .Y(exu_n3437));
AND2X1 exu_U15996(.A(exu_n11631), .B(exu_n16237), .Y(exu_n29027));
INVX1 exu_U15997(.A(exu_n29027), .Y(exu_n3438));
AND2X1 exu_U15998(.A(alu_logic_result_or[50]), .B(exu_n16239), .Y(exu_n29029));
INVX1 exu_U15999(.A(exu_n29029), .Y(exu_n3439));
AND2X1 exu_U16000(.A(div_input_data_e[68]), .B(exu_n16237), .Y(exu_n29033));
INVX1 exu_U16001(.A(exu_n29033), .Y(exu_n3440));
AND2X1 exu_U16002(.A(alu_logic_result_or[4]), .B(exu_n16239), .Y(exu_n29035));
INVX1 exu_U16003(.A(exu_n29035), .Y(exu_n3441));
AND2X1 exu_U16004(.A(exu_n11632), .B(exu_n16237), .Y(exu_n29039));
INVX1 exu_U16005(.A(exu_n29039), .Y(exu_n3442));
AND2X1 exu_U16006(.A(alu_logic_result_or[49]), .B(exu_n16239), .Y(exu_n29041));
INVX1 exu_U16007(.A(exu_n29041), .Y(exu_n3443));
AND2X1 exu_U16008(.A(exu_n11633), .B(exu_n16237), .Y(exu_n29045));
INVX1 exu_U16009(.A(exu_n29045), .Y(exu_n3444));
AND2X1 exu_U16010(.A(alu_logic_result_or[48]), .B(exu_n16239), .Y(exu_n29047));
INVX1 exu_U16011(.A(exu_n29047), .Y(exu_n3445));
AND2X1 exu_U16012(.A(exu_n11634), .B(exu_n16237), .Y(exu_n29051));
INVX1 exu_U16013(.A(exu_n29051), .Y(exu_n3446));
AND2X1 exu_U16014(.A(alu_logic_result_or[47]), .B(exu_n16239), .Y(exu_n29053));
INVX1 exu_U16015(.A(exu_n29053), .Y(exu_n3447));
AND2X1 exu_U16016(.A(exu_n11635), .B(exu_n16237), .Y(exu_n29057));
INVX1 exu_U16017(.A(exu_n29057), .Y(exu_n3448));
AND2X1 exu_U16018(.A(alu_logic_result_or[46]), .B(exu_n16239), .Y(exu_n29059));
INVX1 exu_U16019(.A(exu_n29059), .Y(exu_n3449));
AND2X1 exu_U16020(.A(exu_n11636), .B(exu_n16237), .Y(exu_n29063));
INVX1 exu_U16021(.A(exu_n29063), .Y(exu_n3450));
AND2X1 exu_U16022(.A(alu_logic_result_or[45]), .B(exu_n16239), .Y(exu_n29065));
INVX1 exu_U16023(.A(exu_n29065), .Y(exu_n3451));
AND2X1 exu_U16024(.A(exu_n11637), .B(exu_n16237), .Y(exu_n29069));
INVX1 exu_U16025(.A(exu_n29069), .Y(exu_n3452));
AND2X1 exu_U16026(.A(alu_logic_result_or[44]), .B(exu_n16239), .Y(exu_n29071));
INVX1 exu_U16027(.A(exu_n29071), .Y(exu_n3453));
AND2X1 exu_U16028(.A(exu_n11638), .B(exu_n16237), .Y(exu_n29075));
INVX1 exu_U16029(.A(exu_n29075), .Y(exu_n3454));
AND2X1 exu_U16030(.A(alu_logic_result_or[43]), .B(exu_n16239), .Y(exu_n29077));
INVX1 exu_U16031(.A(exu_n29077), .Y(exu_n3455));
AND2X1 exu_U16032(.A(exu_n11639), .B(exu_n16237), .Y(exu_n29081));
INVX1 exu_U16033(.A(exu_n29081), .Y(exu_n3456));
AND2X1 exu_U16034(.A(alu_logic_result_or[42]), .B(exu_n16239), .Y(exu_n29083));
INVX1 exu_U16035(.A(exu_n29083), .Y(exu_n3457));
AND2X1 exu_U16036(.A(exu_n11640), .B(exu_n16237), .Y(exu_n29087));
INVX1 exu_U16037(.A(exu_n29087), .Y(exu_n3458));
AND2X1 exu_U16038(.A(alu_logic_result_or[41]), .B(exu_n16239), .Y(exu_n29089));
INVX1 exu_U16039(.A(exu_n29089), .Y(exu_n3459));
AND2X1 exu_U16040(.A(exu_n11641), .B(exu_n16237), .Y(exu_n29093));
INVX1 exu_U16041(.A(exu_n29093), .Y(exu_n3460));
AND2X1 exu_U16042(.A(alu_logic_result_or[40]), .B(exu_n16239), .Y(exu_n29095));
INVX1 exu_U16043(.A(exu_n29095), .Y(exu_n3461));
AND2X1 exu_U16044(.A(div_input_data_e[67]), .B(exu_n16237), .Y(exu_n29099));
INVX1 exu_U16045(.A(exu_n29099), .Y(exu_n3462));
AND2X1 exu_U16046(.A(alu_logic_result_or[3]), .B(exu_n16239), .Y(exu_n29101));
INVX1 exu_U16047(.A(exu_n29101), .Y(exu_n3463));
AND2X1 exu_U16048(.A(exu_n11642), .B(exu_n16237), .Y(exu_n29105));
INVX1 exu_U16049(.A(exu_n29105), .Y(exu_n3464));
AND2X1 exu_U16050(.A(alu_logic_result_or[39]), .B(exu_n16239), .Y(exu_n29107));
INVX1 exu_U16051(.A(exu_n29107), .Y(exu_n3465));
AND2X1 exu_U16052(.A(exu_n11643), .B(exu_n16237), .Y(exu_n29111));
INVX1 exu_U16053(.A(exu_n29111), .Y(exu_n3466));
AND2X1 exu_U16054(.A(alu_logic_result_or[38]), .B(exu_n16239), .Y(exu_n29113));
INVX1 exu_U16055(.A(exu_n29113), .Y(exu_n3467));
AND2X1 exu_U16056(.A(exu_n11644), .B(exu_n16237), .Y(exu_n29117));
INVX1 exu_U16057(.A(exu_n29117), .Y(exu_n3468));
AND2X1 exu_U16058(.A(alu_logic_result_or[37]), .B(exu_n16239), .Y(exu_n29119));
INVX1 exu_U16059(.A(exu_n29119), .Y(exu_n3469));
AND2X1 exu_U16060(.A(exu_n11645), .B(exu_n16237), .Y(exu_n29123));
INVX1 exu_U16061(.A(exu_n29123), .Y(exu_n3470));
AND2X1 exu_U16062(.A(alu_logic_result_or[36]), .B(exu_n16239), .Y(exu_n29125));
INVX1 exu_U16063(.A(exu_n29125), .Y(exu_n3471));
AND2X1 exu_U16064(.A(exu_n11646), .B(exu_n16237), .Y(exu_n29129));
INVX1 exu_U16065(.A(exu_n29129), .Y(exu_n3472));
AND2X1 exu_U16066(.A(alu_logic_result_or[35]), .B(exu_n16239), .Y(exu_n29131));
INVX1 exu_U16067(.A(exu_n29131), .Y(exu_n3473));
AND2X1 exu_U16068(.A(exu_n11647), .B(exu_n16237), .Y(exu_n29135));
INVX1 exu_U16069(.A(exu_n29135), .Y(exu_n3474));
AND2X1 exu_U16070(.A(alu_logic_result_or[34]), .B(exu_n16239), .Y(exu_n29137));
INVX1 exu_U16071(.A(exu_n29137), .Y(exu_n3475));
AND2X1 exu_U16072(.A(exu_n11648), .B(exu_n16237), .Y(exu_n29141));
INVX1 exu_U16073(.A(exu_n29141), .Y(exu_n3476));
AND2X1 exu_U16074(.A(alu_logic_result_or[33]), .B(exu_n16239), .Y(exu_n29143));
INVX1 exu_U16075(.A(exu_n29143), .Y(exu_n3477));
AND2X1 exu_U16076(.A(exu_n11649), .B(exu_n16237), .Y(exu_n29147));
INVX1 exu_U16077(.A(exu_n29147), .Y(exu_n3478));
AND2X1 exu_U16078(.A(alu_logic_result_or[32]), .B(exu_n16239), .Y(exu_n29149));
INVX1 exu_U16079(.A(exu_n29149), .Y(exu_n3479));
AND2X1 exu_U16080(.A(div_input_data_e[95]), .B(exu_n16237), .Y(exu_n29153));
INVX1 exu_U16081(.A(exu_n29153), .Y(exu_n3480));
AND2X1 exu_U16082(.A(alu_logic_result_or[31]), .B(exu_n16239), .Y(exu_n29155));
INVX1 exu_U16083(.A(exu_n29155), .Y(exu_n3481));
AND2X1 exu_U16084(.A(div_input_data_e[94]), .B(exu_n16237), .Y(exu_n29159));
INVX1 exu_U16085(.A(exu_n29159), .Y(exu_n3482));
AND2X1 exu_U16086(.A(alu_logic_result_or[30]), .B(exu_n16239), .Y(exu_n29161));
INVX1 exu_U16087(.A(exu_n29161), .Y(exu_n3483));
AND2X1 exu_U16088(.A(div_input_data_e[66]), .B(exu_n16237), .Y(exu_n29165));
INVX1 exu_U16089(.A(exu_n29165), .Y(exu_n3484));
AND2X1 exu_U16090(.A(alu_logic_result_or[2]), .B(exu_n16239), .Y(exu_n29167));
INVX1 exu_U16091(.A(exu_n29167), .Y(exu_n3485));
AND2X1 exu_U16092(.A(div_input_data_e[93]), .B(exu_n16237), .Y(exu_n29171));
INVX1 exu_U16093(.A(exu_n29171), .Y(exu_n3486));
AND2X1 exu_U16094(.A(alu_logic_result_or[29]), .B(exu_n16239), .Y(exu_n29173));
INVX1 exu_U16095(.A(exu_n29173), .Y(exu_n3487));
AND2X1 exu_U16096(.A(div_input_data_e[92]), .B(exu_n16237), .Y(exu_n29177));
INVX1 exu_U16097(.A(exu_n29177), .Y(exu_n3488));
AND2X1 exu_U16098(.A(alu_logic_result_or[28]), .B(exu_n16239), .Y(exu_n29179));
INVX1 exu_U16099(.A(exu_n29179), .Y(exu_n3489));
AND2X1 exu_U16100(.A(div_input_data_e[91]), .B(exu_n16237), .Y(exu_n29183));
INVX1 exu_U16101(.A(exu_n29183), .Y(exu_n3490));
AND2X1 exu_U16102(.A(alu_logic_result_or[27]), .B(exu_n16239), .Y(exu_n29185));
INVX1 exu_U16103(.A(exu_n29185), .Y(exu_n3491));
AND2X1 exu_U16104(.A(div_input_data_e[90]), .B(exu_n16237), .Y(exu_n29189));
INVX1 exu_U16105(.A(exu_n29189), .Y(exu_n3492));
AND2X1 exu_U16106(.A(alu_logic_result_or[26]), .B(exu_n16239), .Y(exu_n29191));
INVX1 exu_U16107(.A(exu_n29191), .Y(exu_n3493));
AND2X1 exu_U16108(.A(div_input_data_e[89]), .B(exu_n16237), .Y(exu_n29195));
INVX1 exu_U16109(.A(exu_n29195), .Y(exu_n3494));
AND2X1 exu_U16110(.A(alu_logic_result_or[25]), .B(exu_n16239), .Y(exu_n29197));
INVX1 exu_U16111(.A(exu_n29197), .Y(exu_n3495));
AND2X1 exu_U16112(.A(div_input_data_e[88]), .B(exu_n16237), .Y(exu_n29201));
INVX1 exu_U16113(.A(exu_n29201), .Y(exu_n3496));
AND2X1 exu_U16114(.A(alu_logic_result_or[24]), .B(exu_n16239), .Y(exu_n29203));
INVX1 exu_U16115(.A(exu_n29203), .Y(exu_n3497));
AND2X1 exu_U16116(.A(div_input_data_e[87]), .B(exu_n16237), .Y(exu_n29207));
INVX1 exu_U16117(.A(exu_n29207), .Y(exu_n3498));
AND2X1 exu_U16118(.A(alu_logic_result_or[23]), .B(exu_n16239), .Y(exu_n29209));
INVX1 exu_U16119(.A(exu_n29209), .Y(exu_n3499));
AND2X1 exu_U16120(.A(div_input_data_e[86]), .B(exu_n16237), .Y(exu_n29213));
INVX1 exu_U16121(.A(exu_n29213), .Y(exu_n3500));
AND2X1 exu_U16122(.A(alu_logic_result_or[22]), .B(exu_n16239), .Y(exu_n29215));
INVX1 exu_U16123(.A(exu_n29215), .Y(exu_n3501));
AND2X1 exu_U16124(.A(div_input_data_e[85]), .B(exu_n16237), .Y(exu_n29219));
INVX1 exu_U16125(.A(exu_n29219), .Y(exu_n3502));
AND2X1 exu_U16126(.A(alu_logic_result_or[21]), .B(exu_n16239), .Y(exu_n29221));
INVX1 exu_U16127(.A(exu_n29221), .Y(exu_n3503));
AND2X1 exu_U16128(.A(div_input_data_e[84]), .B(exu_n16237), .Y(exu_n29225));
INVX1 exu_U16129(.A(exu_n29225), .Y(exu_n3504));
AND2X1 exu_U16130(.A(alu_logic_result_or[20]), .B(exu_n16239), .Y(exu_n29227));
INVX1 exu_U16131(.A(exu_n29227), .Y(exu_n3505));
AND2X1 exu_U16132(.A(div_input_data_e[65]), .B(exu_n16237), .Y(exu_n29231));
INVX1 exu_U16133(.A(exu_n29231), .Y(exu_n3506));
AND2X1 exu_U16134(.A(alu_logic_result_or[1]), .B(exu_n16239), .Y(exu_n29233));
INVX1 exu_U16135(.A(exu_n29233), .Y(exu_n3507));
AND2X1 exu_U16136(.A(div_input_data_e[83]), .B(exu_n16237), .Y(exu_n29237));
INVX1 exu_U16137(.A(exu_n29237), .Y(exu_n3508));
AND2X1 exu_U16138(.A(alu_logic_result_or[19]), .B(exu_n16239), .Y(exu_n29239));
INVX1 exu_U16139(.A(exu_n29239), .Y(exu_n3509));
AND2X1 exu_U16140(.A(div_input_data_e[82]), .B(exu_n16237), .Y(exu_n29243));
INVX1 exu_U16141(.A(exu_n29243), .Y(exu_n3510));
AND2X1 exu_U16142(.A(alu_logic_result_or[18]), .B(exu_n16239), .Y(exu_n29245));
INVX1 exu_U16143(.A(exu_n29245), .Y(exu_n3511));
AND2X1 exu_U16144(.A(div_input_data_e[81]), .B(exu_n16237), .Y(exu_n29249));
INVX1 exu_U16145(.A(exu_n29249), .Y(exu_n3512));
AND2X1 exu_U16146(.A(alu_logic_result_or[17]), .B(exu_n16239), .Y(exu_n29251));
INVX1 exu_U16147(.A(exu_n29251), .Y(exu_n3513));
AND2X1 exu_U16148(.A(div_input_data_e[80]), .B(exu_n16237), .Y(exu_n29255));
INVX1 exu_U16149(.A(exu_n29255), .Y(exu_n3514));
AND2X1 exu_U16150(.A(alu_logic_result_or[16]), .B(exu_n16239), .Y(exu_n29257));
INVX1 exu_U16151(.A(exu_n29257), .Y(exu_n3515));
AND2X1 exu_U16152(.A(div_input_data_e[79]), .B(exu_n16237), .Y(exu_n29261));
INVX1 exu_U16153(.A(exu_n29261), .Y(exu_n3516));
AND2X1 exu_U16154(.A(alu_logic_result_or[15]), .B(exu_n16239), .Y(exu_n29263));
INVX1 exu_U16155(.A(exu_n29263), .Y(exu_n3517));
AND2X1 exu_U16156(.A(div_input_data_e[78]), .B(exu_n16237), .Y(exu_n29267));
INVX1 exu_U16157(.A(exu_n29267), .Y(exu_n3518));
AND2X1 exu_U16158(.A(alu_logic_result_or[14]), .B(exu_n16239), .Y(exu_n29269));
INVX1 exu_U16159(.A(exu_n29269), .Y(exu_n3519));
AND2X1 exu_U16160(.A(div_input_data_e[77]), .B(exu_n16237), .Y(exu_n29273));
INVX1 exu_U16161(.A(exu_n29273), .Y(exu_n3520));
AND2X1 exu_U16162(.A(alu_logic_result_or[13]), .B(exu_n16239), .Y(exu_n29275));
INVX1 exu_U16163(.A(exu_n29275), .Y(exu_n3521));
AND2X1 exu_U16164(.A(div_input_data_e[76]), .B(exu_n16237), .Y(exu_n29279));
INVX1 exu_U16165(.A(exu_n29279), .Y(exu_n3522));
AND2X1 exu_U16166(.A(alu_logic_result_or[12]), .B(exu_n16239), .Y(exu_n29281));
INVX1 exu_U16167(.A(exu_n29281), .Y(exu_n3523));
AND2X1 exu_U16168(.A(div_input_data_e[75]), .B(exu_n16237), .Y(exu_n29285));
INVX1 exu_U16169(.A(exu_n29285), .Y(exu_n3524));
AND2X1 exu_U16170(.A(alu_logic_result_or[11]), .B(exu_n16239), .Y(exu_n29287));
INVX1 exu_U16171(.A(exu_n29287), .Y(exu_n3525));
AND2X1 exu_U16172(.A(div_input_data_e[74]), .B(exu_n16237), .Y(exu_n29291));
INVX1 exu_U16173(.A(exu_n29291), .Y(exu_n3526));
AND2X1 exu_U16174(.A(alu_logic_result_or[10]), .B(exu_n16239), .Y(exu_n29293));
INVX1 exu_U16175(.A(exu_n29293), .Y(exu_n3527));
AND2X1 exu_U16176(.A(div_input_data_e[64]), .B(exu_n16237), .Y(exu_n29297));
INVX1 exu_U16177(.A(exu_n29297), .Y(exu_n3528));
AND2X1 exu_U16178(.A(alu_logic_result_or[0]), .B(exu_n16239), .Y(exu_n29299));
INVX1 exu_U16179(.A(exu_n29299), .Y(exu_n3529));
AND2X1 exu_U16180(.A(exu_n11059), .B(exu_n10065), .Y(bypass_restore_rd_data_next[9]));
INVX1 exu_U16181(.A(bypass_restore_rd_data_next[9]), .Y(exu_n3530));
AND2X1 exu_U16182(.A(exu_n11060), .B(exu_n10066), .Y(bypass_restore_rd_data_next[8]));
INVX1 exu_U16183(.A(bypass_restore_rd_data_next[8]), .Y(exu_n3531));
AND2X1 exu_U16184(.A(exu_n11061), .B(exu_n10067), .Y(bypass_restore_rd_data_next[7]));
INVX1 exu_U16185(.A(bypass_restore_rd_data_next[7]), .Y(exu_n3532));
AND2X1 exu_U16186(.A(exu_n11062), .B(exu_n10068), .Y(bypass_restore_rd_data_next[6]));
INVX1 exu_U16187(.A(bypass_restore_rd_data_next[6]), .Y(exu_n3533));
AND2X1 exu_U16188(.A(exu_n11063), .B(exu_n10069), .Y(bypass_restore_rd_data_next[63]));
INVX1 exu_U16189(.A(bypass_restore_rd_data_next[63]), .Y(exu_n3534));
AND2X1 exu_U16190(.A(exu_n11064), .B(exu_n10070), .Y(bypass_restore_rd_data_next[62]));
INVX1 exu_U16191(.A(bypass_restore_rd_data_next[62]), .Y(exu_n3535));
AND2X1 exu_U16192(.A(exu_n11065), .B(exu_n10071), .Y(bypass_restore_rd_data_next[61]));
INVX1 exu_U16193(.A(bypass_restore_rd_data_next[61]), .Y(exu_n3536));
AND2X1 exu_U16194(.A(exu_n11066), .B(exu_n10072), .Y(bypass_restore_rd_data_next[60]));
INVX1 exu_U16195(.A(bypass_restore_rd_data_next[60]), .Y(exu_n3537));
AND2X1 exu_U16196(.A(exu_n11067), .B(exu_n10073), .Y(bypass_restore_rd_data_next[5]));
INVX1 exu_U16197(.A(bypass_restore_rd_data_next[5]), .Y(exu_n3538));
AND2X1 exu_U16198(.A(exu_n11068), .B(exu_n10074), .Y(bypass_restore_rd_data_next[59]));
INVX1 exu_U16199(.A(bypass_restore_rd_data_next[59]), .Y(exu_n3539));
AND2X1 exu_U16200(.A(exu_n11069), .B(exu_n10075), .Y(bypass_restore_rd_data_next[58]));
INVX1 exu_U16201(.A(bypass_restore_rd_data_next[58]), .Y(exu_n3540));
AND2X1 exu_U16202(.A(exu_n11070), .B(exu_n10076), .Y(bypass_restore_rd_data_next[57]));
INVX1 exu_U16203(.A(bypass_restore_rd_data_next[57]), .Y(exu_n3541));
AND2X1 exu_U16204(.A(exu_n11071), .B(exu_n10077), .Y(bypass_restore_rd_data_next[56]));
INVX1 exu_U16205(.A(bypass_restore_rd_data_next[56]), .Y(exu_n3542));
AND2X1 exu_U16206(.A(exu_n11072), .B(exu_n10078), .Y(bypass_restore_rd_data_next[55]));
INVX1 exu_U16207(.A(bypass_restore_rd_data_next[55]), .Y(exu_n3543));
AND2X1 exu_U16208(.A(exu_n11073), .B(exu_n10079), .Y(bypass_restore_rd_data_next[54]));
INVX1 exu_U16209(.A(bypass_restore_rd_data_next[54]), .Y(exu_n3544));
AND2X1 exu_U16210(.A(exu_n11074), .B(exu_n10080), .Y(bypass_restore_rd_data_next[53]));
INVX1 exu_U16211(.A(bypass_restore_rd_data_next[53]), .Y(exu_n3545));
AND2X1 exu_U16212(.A(exu_n11075), .B(exu_n10081), .Y(bypass_restore_rd_data_next[52]));
INVX1 exu_U16213(.A(bypass_restore_rd_data_next[52]), .Y(exu_n3546));
AND2X1 exu_U16214(.A(exu_n11076), .B(exu_n10082), .Y(bypass_restore_rd_data_next[51]));
INVX1 exu_U16215(.A(bypass_restore_rd_data_next[51]), .Y(exu_n3547));
AND2X1 exu_U16216(.A(exu_n11077), .B(exu_n10083), .Y(bypass_restore_rd_data_next[50]));
INVX1 exu_U16217(.A(bypass_restore_rd_data_next[50]), .Y(exu_n3548));
AND2X1 exu_U16218(.A(exu_n11078), .B(exu_n10084), .Y(bypass_restore_rd_data_next[4]));
INVX1 exu_U16219(.A(bypass_restore_rd_data_next[4]), .Y(exu_n3549));
AND2X1 exu_U16220(.A(exu_n11079), .B(exu_n10085), .Y(bypass_restore_rd_data_next[49]));
INVX1 exu_U16221(.A(bypass_restore_rd_data_next[49]), .Y(exu_n3550));
AND2X1 exu_U16222(.A(exu_n11080), .B(exu_n10086), .Y(bypass_restore_rd_data_next[48]));
INVX1 exu_U16223(.A(bypass_restore_rd_data_next[48]), .Y(exu_n3551));
AND2X1 exu_U16224(.A(exu_n11081), .B(exu_n10087), .Y(bypass_restore_rd_data_next[47]));
INVX1 exu_U16225(.A(bypass_restore_rd_data_next[47]), .Y(exu_n3552));
AND2X1 exu_U16226(.A(exu_n11082), .B(exu_n10088), .Y(bypass_restore_rd_data_next[46]));
INVX1 exu_U16227(.A(bypass_restore_rd_data_next[46]), .Y(exu_n3553));
AND2X1 exu_U16228(.A(exu_n11083), .B(exu_n10089), .Y(bypass_restore_rd_data_next[45]));
INVX1 exu_U16229(.A(bypass_restore_rd_data_next[45]), .Y(exu_n3554));
AND2X1 exu_U16230(.A(exu_n11084), .B(exu_n10090), .Y(bypass_restore_rd_data_next[44]));
INVX1 exu_U16231(.A(bypass_restore_rd_data_next[44]), .Y(exu_n3555));
AND2X1 exu_U16232(.A(exu_n11085), .B(exu_n10091), .Y(bypass_restore_rd_data_next[43]));
INVX1 exu_U16233(.A(bypass_restore_rd_data_next[43]), .Y(exu_n3556));
AND2X1 exu_U16234(.A(exu_n11086), .B(exu_n10092), .Y(bypass_restore_rd_data_next[42]));
INVX1 exu_U16235(.A(bypass_restore_rd_data_next[42]), .Y(exu_n3557));
AND2X1 exu_U16236(.A(exu_n11087), .B(exu_n10093), .Y(bypass_restore_rd_data_next[41]));
INVX1 exu_U16237(.A(bypass_restore_rd_data_next[41]), .Y(exu_n3558));
AND2X1 exu_U16238(.A(exu_n11088), .B(exu_n10094), .Y(bypass_restore_rd_data_next[40]));
INVX1 exu_U16239(.A(bypass_restore_rd_data_next[40]), .Y(exu_n3559));
AND2X1 exu_U16240(.A(exu_n11089), .B(exu_n10095), .Y(bypass_restore_rd_data_next[3]));
INVX1 exu_U16241(.A(bypass_restore_rd_data_next[3]), .Y(exu_n3560));
AND2X1 exu_U16242(.A(exu_n11090), .B(exu_n10096), .Y(bypass_restore_rd_data_next[39]));
INVX1 exu_U16243(.A(bypass_restore_rd_data_next[39]), .Y(exu_n3561));
AND2X1 exu_U16244(.A(exu_n11091), .B(exu_n10097), .Y(bypass_restore_rd_data_next[38]));
INVX1 exu_U16245(.A(bypass_restore_rd_data_next[38]), .Y(exu_n3562));
AND2X1 exu_U16246(.A(exu_n11092), .B(exu_n10098), .Y(bypass_restore_rd_data_next[37]));
INVX1 exu_U16247(.A(bypass_restore_rd_data_next[37]), .Y(exu_n3563));
AND2X1 exu_U16248(.A(exu_n11093), .B(exu_n10099), .Y(bypass_restore_rd_data_next[36]));
INVX1 exu_U16249(.A(bypass_restore_rd_data_next[36]), .Y(exu_n3564));
AND2X1 exu_U16250(.A(exu_n11094), .B(exu_n10100), .Y(bypass_restore_rd_data_next[35]));
INVX1 exu_U16251(.A(bypass_restore_rd_data_next[35]), .Y(exu_n3565));
AND2X1 exu_U16252(.A(exu_n11095), .B(exu_n10101), .Y(bypass_restore_rd_data_next[34]));
INVX1 exu_U16253(.A(bypass_restore_rd_data_next[34]), .Y(exu_n3566));
AND2X1 exu_U16254(.A(exu_n11096), .B(exu_n10102), .Y(bypass_restore_rd_data_next[33]));
INVX1 exu_U16255(.A(bypass_restore_rd_data_next[33]), .Y(exu_n3567));
AND2X1 exu_U16256(.A(exu_n11097), .B(exu_n10103), .Y(bypass_restore_rd_data_next[32]));
INVX1 exu_U16257(.A(bypass_restore_rd_data_next[32]), .Y(exu_n3568));
AND2X1 exu_U16258(.A(exu_n11098), .B(exu_n10104), .Y(bypass_restore_rd_data_next[31]));
INVX1 exu_U16259(.A(bypass_restore_rd_data_next[31]), .Y(exu_n3569));
AND2X1 exu_U16260(.A(exu_n11099), .B(exu_n10105), .Y(bypass_restore_rd_data_next[30]));
INVX1 exu_U16261(.A(bypass_restore_rd_data_next[30]), .Y(exu_n3570));
AND2X1 exu_U16262(.A(exu_n11100), .B(exu_n10106), .Y(bypass_restore_rd_data_next[2]));
INVX1 exu_U16263(.A(bypass_restore_rd_data_next[2]), .Y(exu_n3571));
AND2X1 exu_U16264(.A(exu_n11101), .B(exu_n10107), .Y(bypass_restore_rd_data_next[29]));
INVX1 exu_U16265(.A(bypass_restore_rd_data_next[29]), .Y(exu_n3572));
AND2X1 exu_U16266(.A(exu_n11102), .B(exu_n10108), .Y(bypass_restore_rd_data_next[28]));
INVX1 exu_U16267(.A(bypass_restore_rd_data_next[28]), .Y(exu_n3573));
AND2X1 exu_U16268(.A(exu_n11103), .B(exu_n10109), .Y(bypass_restore_rd_data_next[27]));
INVX1 exu_U16269(.A(bypass_restore_rd_data_next[27]), .Y(exu_n3574));
AND2X1 exu_U16270(.A(exu_n11104), .B(exu_n10110), .Y(bypass_restore_rd_data_next[26]));
INVX1 exu_U16271(.A(bypass_restore_rd_data_next[26]), .Y(exu_n3575));
AND2X1 exu_U16272(.A(exu_n11105), .B(exu_n10111), .Y(bypass_restore_rd_data_next[25]));
INVX1 exu_U16273(.A(bypass_restore_rd_data_next[25]), .Y(exu_n3576));
AND2X1 exu_U16274(.A(exu_n11106), .B(exu_n10112), .Y(bypass_restore_rd_data_next[24]));
INVX1 exu_U16275(.A(bypass_restore_rd_data_next[24]), .Y(exu_n3577));
AND2X1 exu_U16276(.A(exu_n11107), .B(exu_n10113), .Y(bypass_restore_rd_data_next[23]));
INVX1 exu_U16277(.A(bypass_restore_rd_data_next[23]), .Y(exu_n3578));
AND2X1 exu_U16278(.A(exu_n11108), .B(exu_n10114), .Y(bypass_restore_rd_data_next[22]));
INVX1 exu_U16279(.A(bypass_restore_rd_data_next[22]), .Y(exu_n3579));
AND2X1 exu_U16280(.A(exu_n11109), .B(exu_n10115), .Y(bypass_restore_rd_data_next[21]));
INVX1 exu_U16281(.A(bypass_restore_rd_data_next[21]), .Y(exu_n3580));
AND2X1 exu_U16282(.A(exu_n11110), .B(exu_n10116), .Y(bypass_restore_rd_data_next[20]));
INVX1 exu_U16283(.A(bypass_restore_rd_data_next[20]), .Y(exu_n3581));
AND2X1 exu_U16284(.A(exu_n11111), .B(exu_n10117), .Y(bypass_restore_rd_data_next[1]));
INVX1 exu_U16285(.A(bypass_restore_rd_data_next[1]), .Y(exu_n3582));
AND2X1 exu_U16286(.A(exu_n11112), .B(exu_n10118), .Y(bypass_restore_rd_data_next[19]));
INVX1 exu_U16287(.A(bypass_restore_rd_data_next[19]), .Y(exu_n3583));
AND2X1 exu_U16288(.A(exu_n11113), .B(exu_n10119), .Y(bypass_restore_rd_data_next[18]));
INVX1 exu_U16289(.A(bypass_restore_rd_data_next[18]), .Y(exu_n3584));
AND2X1 exu_U16290(.A(exu_n11114), .B(exu_n10120), .Y(bypass_restore_rd_data_next[17]));
INVX1 exu_U16291(.A(bypass_restore_rd_data_next[17]), .Y(exu_n3585));
AND2X1 exu_U16292(.A(exu_n11115), .B(exu_n10121), .Y(bypass_restore_rd_data_next[16]));
INVX1 exu_U16293(.A(bypass_restore_rd_data_next[16]), .Y(exu_n3586));
AND2X1 exu_U16294(.A(exu_n11116), .B(exu_n10122), .Y(bypass_restore_rd_data_next[15]));
INVX1 exu_U16295(.A(bypass_restore_rd_data_next[15]), .Y(exu_n3587));
AND2X1 exu_U16296(.A(exu_n11117), .B(exu_n10123), .Y(bypass_restore_rd_data_next[14]));
INVX1 exu_U16297(.A(bypass_restore_rd_data_next[14]), .Y(exu_n3588));
AND2X1 exu_U16298(.A(exu_n11118), .B(exu_n10124), .Y(bypass_restore_rd_data_next[13]));
INVX1 exu_U16299(.A(bypass_restore_rd_data_next[13]), .Y(exu_n3589));
AND2X1 exu_U16300(.A(exu_n11119), .B(exu_n10125), .Y(bypass_restore_rd_data_next[12]));
INVX1 exu_U16301(.A(bypass_restore_rd_data_next[12]), .Y(exu_n3590));
AND2X1 exu_U16302(.A(exu_n11120), .B(exu_n10126), .Y(bypass_restore_rd_data_next[11]));
INVX1 exu_U16303(.A(bypass_restore_rd_data_next[11]), .Y(exu_n3591));
AND2X1 exu_U16304(.A(exu_n11121), .B(exu_n10127), .Y(bypass_restore_rd_data_next[10]));
INVX1 exu_U16305(.A(bypass_restore_rd_data_next[10]), .Y(exu_n3592));
AND2X1 exu_U16306(.A(exu_n11122), .B(exu_n10128), .Y(bypass_restore_rd_data_next[0]));
INVX1 exu_U16307(.A(bypass_restore_rd_data_next[0]), .Y(exu_n3593));
AND2X1 exu_U16308(.A(exu_n16162), .B(bypass_rs3h_data_e[9]), .Y(exu_n30401));
INVX1 exu_U16309(.A(exu_n30401), .Y(exu_n3594));
AND2X1 exu_U16310(.A(bypass_rs3h_data_e[8]), .B(exu_n16165), .Y(exu_n30403));
INVX1 exu_U16311(.A(exu_n30403), .Y(exu_n3595));
AND2X1 exu_U16312(.A(bypass_rs3h_data_e[7]), .B(exu_n16165), .Y(exu_n30405));
INVX1 exu_U16313(.A(exu_n30405), .Y(exu_n3596));
AND2X1 exu_U16314(.A(bypass_rs3h_data_e[6]), .B(exu_n16165), .Y(exu_n30407));
INVX1 exu_U16315(.A(exu_n30407), .Y(exu_n3597));
AND2X1 exu_U16316(.A(bypass_rs3h_data_e[5]), .B(exu_n16165), .Y(exu_n30413));
INVX1 exu_U16317(.A(exu_n30413), .Y(exu_n3598));
AND2X1 exu_U16318(.A(bypass_rs3h_data_e[4]), .B(exu_n16164), .Y(exu_n30425));
INVX1 exu_U16319(.A(exu_n30425), .Y(exu_n3599));
AND2X1 exu_U16320(.A(bypass_rs3h_data_e[3]), .B(exu_n16164), .Y(exu_n30437));
INVX1 exu_U16321(.A(exu_n30437), .Y(exu_n3600));
AND2X1 exu_U16322(.A(bypass_rs3h_data_e[31]), .B(exu_n16164), .Y(exu_n30447));
INVX1 exu_U16323(.A(exu_n30447), .Y(exu_n3601));
AND2X1 exu_U16324(.A(bypass_rs3h_data_e[30]), .B(exu_n16164), .Y(exu_n30449));
INVX1 exu_U16325(.A(exu_n30449), .Y(exu_n3602));
AND2X1 exu_U16326(.A(bypass_rs3h_data_e[2]), .B(exu_n16165), .Y(exu_n30451));
INVX1 exu_U16327(.A(exu_n30451), .Y(exu_n3603));
AND2X1 exu_U16328(.A(bypass_rs3h_data_e[29]), .B(exu_n16164), .Y(exu_n30453));
INVX1 exu_U16329(.A(exu_n30453), .Y(exu_n3604));
AND2X1 exu_U16330(.A(bypass_rs3h_data_e[28]), .B(exu_n16164), .Y(exu_n30455));
INVX1 exu_U16331(.A(exu_n30455), .Y(exu_n3605));
AND2X1 exu_U16332(.A(bypass_rs3h_data_e[27]), .B(exu_n16164), .Y(exu_n30457));
INVX1 exu_U16333(.A(exu_n30457), .Y(exu_n3606));
AND2X1 exu_U16334(.A(bypass_rs3h_data_e[26]), .B(exu_n16164), .Y(exu_n30459));
INVX1 exu_U16335(.A(exu_n30459), .Y(exu_n3607));
AND2X1 exu_U16336(.A(bypass_rs3h_data_e[25]), .B(exu_n16164), .Y(exu_n30461));
INVX1 exu_U16337(.A(exu_n30461), .Y(exu_n3608));
AND2X1 exu_U16338(.A(bypass_rs3h_data_e[24]), .B(ecl_std_e), .Y(exu_n30463));
INVX1 exu_U16339(.A(exu_n30463), .Y(exu_n3609));
AND2X1 exu_U16340(.A(bypass_rs3h_data_e[23]), .B(exu_n16164), .Y(exu_n30465));
INVX1 exu_U16341(.A(exu_n30465), .Y(exu_n3610));
AND2X1 exu_U16342(.A(bypass_rs3h_data_e[22]), .B(exu_n16164), .Y(exu_n30467));
INVX1 exu_U16343(.A(exu_n30467), .Y(exu_n3611));
AND2X1 exu_U16344(.A(bypass_rs3h_data_e[21]), .B(exu_n16164), .Y(exu_n30469));
INVX1 exu_U16345(.A(exu_n30469), .Y(exu_n3612));
AND2X1 exu_U16346(.A(bypass_rs3h_data_e[20]), .B(exu_n16164), .Y(exu_n30471));
INVX1 exu_U16347(.A(exu_n30471), .Y(exu_n3613));
AND2X1 exu_U16348(.A(bypass_rs3h_data_e[1]), .B(exu_n16164), .Y(exu_n30473));
INVX1 exu_U16349(.A(exu_n30473), .Y(exu_n3614));
AND2X1 exu_U16350(.A(bypass_rs3h_data_e[19]), .B(exu_n16163), .Y(exu_n30475));
INVX1 exu_U16351(.A(exu_n30475), .Y(exu_n3615));
AND2X1 exu_U16352(.A(bypass_rs3h_data_e[18]), .B(exu_n16163), .Y(exu_n30477));
INVX1 exu_U16353(.A(exu_n30477), .Y(exu_n3616));
AND2X1 exu_U16354(.A(bypass_rs3h_data_e[17]), .B(exu_n16163), .Y(exu_n30479));
INVX1 exu_U16355(.A(exu_n30479), .Y(exu_n3617));
AND2X1 exu_U16356(.A(bypass_rs3h_data_e[16]), .B(exu_n16163), .Y(exu_n30481));
INVX1 exu_U16357(.A(exu_n30481), .Y(exu_n3618));
AND2X1 exu_U16358(.A(bypass_rs3h_data_e[15]), .B(exu_n16163), .Y(exu_n30483));
INVX1 exu_U16359(.A(exu_n30483), .Y(exu_n3619));
AND2X1 exu_U16360(.A(bypass_rs3h_data_e[14]), .B(exu_n16163), .Y(exu_n30485));
INVX1 exu_U16361(.A(exu_n30485), .Y(exu_n3620));
AND2X1 exu_U16362(.A(bypass_rs3h_data_e[13]), .B(exu_n16163), .Y(exu_n30487));
INVX1 exu_U16363(.A(exu_n30487), .Y(exu_n3621));
AND2X1 exu_U16364(.A(bypass_rs3h_data_e[12]), .B(exu_n16163), .Y(exu_n30489));
INVX1 exu_U16365(.A(exu_n30489), .Y(exu_n3622));
AND2X1 exu_U16366(.A(bypass_rs3h_data_e[11]), .B(exu_n16164), .Y(exu_n30491));
INVX1 exu_U16367(.A(exu_n30491), .Y(exu_n3623));
AND2X1 exu_U16368(.A(bypass_rs3h_data_e[10]), .B(exu_n16163), .Y(exu_n30493));
INVX1 exu_U16369(.A(exu_n30493), .Y(exu_n3624));
AND2X1 exu_U16370(.A(bypass_rs3h_data_e[0]), .B(exu_n16164), .Y(exu_n30495));
INVX1 exu_U16371(.A(exu_n30495), .Y(exu_n3625));
AND2X1 exu_U16372(.A(alu_logic_rs1_data_bf1[63]), .B(ecl_alu_casa_e), .Y(exu_n30505));
INVX1 exu_U16373(.A(exu_n30505), .Y(exu_n3626));
AND2X1 exu_U16374(.A(alu_logic_rs1_data_bf1[62]), .B(ecl_alu_casa_e), .Y(exu_n30507));
INVX1 exu_U16375(.A(exu_n30507), .Y(exu_n3627));
AND2X1 exu_U16376(.A(alu_logic_rs1_data_bf1[61]), .B(ecl_alu_casa_e), .Y(exu_n30509));
INVX1 exu_U16377(.A(exu_n30509), .Y(exu_n3628));
AND2X1 exu_U16378(.A(alu_logic_rs1_data_bf1[60]), .B(ecl_alu_casa_e), .Y(exu_n30511));
INVX1 exu_U16379(.A(exu_n30511), .Y(exu_n3629));
AND2X1 exu_U16380(.A(alu_logic_rs1_data_bf1[59]), .B(ecl_alu_casa_e), .Y(exu_n30515));
INVX1 exu_U16381(.A(exu_n30515), .Y(exu_n3630));
AND2X1 exu_U16382(.A(alu_logic_rs1_data_bf1[58]), .B(ecl_alu_casa_e), .Y(exu_n30517));
INVX1 exu_U16383(.A(exu_n30517), .Y(exu_n3631));
AND2X1 exu_U16384(.A(alu_logic_rs1_data_bf1[57]), .B(ecl_alu_casa_e), .Y(exu_n30519));
INVX1 exu_U16385(.A(exu_n30519), .Y(exu_n3632));
AND2X1 exu_U16386(.A(alu_logic_rs1_data_bf1[56]), .B(ecl_alu_casa_e), .Y(exu_n30521));
INVX1 exu_U16387(.A(exu_n30521), .Y(exu_n3633));
AND2X1 exu_U16388(.A(alu_logic_rs1_data_bf1[55]), .B(ecl_alu_casa_e), .Y(exu_n30523));
INVX1 exu_U16389(.A(exu_n30523), .Y(exu_n3634));
AND2X1 exu_U16390(.A(alu_logic_rs1_data_bf1[54]), .B(ecl_alu_casa_e), .Y(exu_n30525));
INVX1 exu_U16391(.A(exu_n30525), .Y(exu_n3635));
AND2X1 exu_U16392(.A(alu_logic_rs1_data_bf1[53]), .B(ecl_alu_casa_e), .Y(exu_n30527));
INVX1 exu_U16393(.A(exu_n30527), .Y(exu_n3636));
AND2X1 exu_U16394(.A(alu_logic_rs1_data_bf1[52]), .B(ecl_alu_casa_e), .Y(exu_n30529));
INVX1 exu_U16395(.A(exu_n30529), .Y(exu_n3637));
AND2X1 exu_U16396(.A(alu_logic_rs1_data_bf1[51]), .B(ecl_alu_casa_e), .Y(exu_n30531));
INVX1 exu_U16397(.A(exu_n30531), .Y(exu_n3638));
AND2X1 exu_U16398(.A(alu_logic_rs1_data_bf1[50]), .B(ecl_alu_casa_e), .Y(exu_n30533));
INVX1 exu_U16399(.A(exu_n30533), .Y(exu_n3639));
AND2X1 exu_U16400(.A(alu_logic_rs1_data_bf1[49]), .B(ecl_alu_casa_e), .Y(exu_n30537));
INVX1 exu_U16401(.A(exu_n30537), .Y(exu_n3640));
AND2X1 exu_U16402(.A(alu_logic_rs1_data_bf1[48]), .B(ecl_alu_casa_e), .Y(exu_n30539));
INVX1 exu_U16403(.A(exu_n30539), .Y(exu_n3641));
AND2X1 exu_U16404(.A(alu_logic_rs1_data_bf1[47]), .B(ecl_alu_casa_e), .Y(exu_n30541));
INVX1 exu_U16405(.A(exu_n30541), .Y(exu_n3642));
AND2X1 exu_U16406(.A(exu_n16155), .B(alu_spr_out[9]), .Y(exu_n30625));
INVX1 exu_U16407(.A(exu_n30625), .Y(exu_n3643));
AND2X1 exu_U16408(.A(alu_spr_out[8]), .B(exu_n16155), .Y(exu_n30627));
INVX1 exu_U16409(.A(exu_n30627), .Y(exu_n3644));
AND2X1 exu_U16410(.A(alu_spr_out[7]), .B(exu_n16158), .Y(exu_n30629));
INVX1 exu_U16411(.A(exu_n30629), .Y(exu_n3645));
AND2X1 exu_U16412(.A(alu_spr_out[6]), .B(ecl_sel_sum_e), .Y(exu_n30631));
INVX1 exu_U16413(.A(exu_n30631), .Y(exu_n3646));
AND2X1 exu_U16414(.A(alu_spr_out[63]), .B(exu_n16155), .Y(exu_n30633));
INVX1 exu_U16415(.A(exu_n30633), .Y(exu_n3647));
AND2X1 exu_U16416(.A(alu_spr_out[62]), .B(exu_n16157), .Y(exu_n30635));
INVX1 exu_U16417(.A(exu_n30635), .Y(exu_n3648));
AND2X1 exu_U16418(.A(alu_spr_out[61]), .B(exu_n16158), .Y(exu_n30637));
INVX1 exu_U16419(.A(exu_n30637), .Y(exu_n3649));
AND2X1 exu_U16420(.A(alu_spr_out[60]), .B(exu_n16157), .Y(exu_n30639));
INVX1 exu_U16421(.A(exu_n30639), .Y(exu_n3650));
AND2X1 exu_U16422(.A(alu_spr_out[5]), .B(ecl_sel_sum_e), .Y(exu_n30641));
INVX1 exu_U16423(.A(exu_n30641), .Y(exu_n3651));
AND2X1 exu_U16424(.A(alu_spr_out[59]), .B(exu_n16157), .Y(exu_n30643));
INVX1 exu_U16425(.A(exu_n30643), .Y(exu_n3652));
AND2X1 exu_U16426(.A(alu_spr_out[58]), .B(ecl_sel_sum_e), .Y(exu_n30645));
INVX1 exu_U16427(.A(exu_n30645), .Y(exu_n3653));
AND2X1 exu_U16428(.A(alu_spr_out[57]), .B(exu_n16155), .Y(exu_n30647));
INVX1 exu_U16429(.A(exu_n30647), .Y(exu_n3654));
AND2X1 exu_U16430(.A(alu_spr_out[56]), .B(exu_n16157), .Y(exu_n30649));
INVX1 exu_U16431(.A(exu_n30649), .Y(exu_n3655));
AND2X1 exu_U16432(.A(alu_spr_out[55]), .B(exu_n16158), .Y(exu_n30651));
INVX1 exu_U16433(.A(exu_n30651), .Y(exu_n3656));
AND2X1 exu_U16434(.A(alu_spr_out[54]), .B(exu_n16158), .Y(exu_n30653));
INVX1 exu_U16435(.A(exu_n30653), .Y(exu_n3657));
AND2X1 exu_U16436(.A(alu_spr_out[53]), .B(ecl_sel_sum_e), .Y(exu_n30655));
INVX1 exu_U16437(.A(exu_n30655), .Y(exu_n3658));
AND2X1 exu_U16438(.A(alu_spr_out[52]), .B(ecl_sel_sum_e), .Y(exu_n30657));
INVX1 exu_U16439(.A(exu_n30657), .Y(exu_n3659));
AND2X1 exu_U16440(.A(alu_spr_out[51]), .B(ecl_sel_sum_e), .Y(exu_n30659));
INVX1 exu_U16441(.A(exu_n30659), .Y(exu_n3660));
AND2X1 exu_U16442(.A(alu_spr_out[50]), .B(exu_n16157), .Y(exu_n30661));
INVX1 exu_U16443(.A(exu_n30661), .Y(exu_n3661));
AND2X1 exu_U16444(.A(alu_spr_out[4]), .B(ecl_sel_sum_e), .Y(exu_n30663));
INVX1 exu_U16445(.A(exu_n30663), .Y(exu_n3662));
AND2X1 exu_U16446(.A(alu_spr_out[49]), .B(exu_n16155), .Y(exu_n30665));
INVX1 exu_U16447(.A(exu_n30665), .Y(exu_n3663));
AND2X1 exu_U16448(.A(alu_spr_out[48]), .B(exu_n16157), .Y(exu_n30667));
INVX1 exu_U16449(.A(exu_n30667), .Y(exu_n3664));
AND2X1 exu_U16450(.A(alu_spr_out[47]), .B(exu_n16158), .Y(exu_n30669));
INVX1 exu_U16451(.A(exu_n30669), .Y(exu_n3665));
AND2X1 exu_U16452(.A(alu_spr_out[46]), .B(exu_n16155), .Y(exu_n30671));
INVX1 exu_U16453(.A(exu_n30671), .Y(exu_n3666));
AND2X1 exu_U16454(.A(alu_spr_out[45]), .B(exu_n16155), .Y(exu_n30673));
INVX1 exu_U16455(.A(exu_n30673), .Y(exu_n3667));
AND2X1 exu_U16456(.A(alu_spr_out[44]), .B(exu_n16155), .Y(exu_n30675));
INVX1 exu_U16457(.A(exu_n30675), .Y(exu_n3668));
AND2X1 exu_U16458(.A(alu_spr_out[43]), .B(exu_n16158), .Y(exu_n30677));
INVX1 exu_U16459(.A(exu_n30677), .Y(exu_n3669));
AND2X1 exu_U16460(.A(alu_spr_out[42]), .B(ecl_sel_sum_e), .Y(exu_n30679));
INVX1 exu_U16461(.A(exu_n30679), .Y(exu_n3670));
AND2X1 exu_U16462(.A(alu_spr_out[41]), .B(exu_n16155), .Y(exu_n30681));
INVX1 exu_U16463(.A(exu_n30681), .Y(exu_n3671));
AND2X1 exu_U16464(.A(alu_spr_out[40]), .B(exu_n16157), .Y(exu_n30683));
INVX1 exu_U16465(.A(exu_n30683), .Y(exu_n3672));
AND2X1 exu_U16466(.A(alu_spr_out[3]), .B(exu_n16157), .Y(exu_n30685));
INVX1 exu_U16467(.A(exu_n30685), .Y(exu_n3673));
AND2X1 exu_U16468(.A(alu_spr_out[39]), .B(exu_n16157), .Y(exu_n30687));
INVX1 exu_U16469(.A(exu_n30687), .Y(exu_n3674));
AND2X1 exu_U16470(.A(alu_spr_out[38]), .B(exu_n16157), .Y(exu_n30689));
INVX1 exu_U16471(.A(exu_n30689), .Y(exu_n3675));
AND2X1 exu_U16472(.A(alu_spr_out[37]), .B(exu_n16157), .Y(exu_n30691));
INVX1 exu_U16473(.A(exu_n30691), .Y(exu_n3676));
AND2X1 exu_U16474(.A(alu_spr_out[36]), .B(exu_n16157), .Y(exu_n30693));
INVX1 exu_U16475(.A(exu_n30693), .Y(exu_n3677));
AND2X1 exu_U16476(.A(alu_spr_out[35]), .B(exu_n16157), .Y(exu_n30695));
INVX1 exu_U16477(.A(exu_n30695), .Y(exu_n3678));
AND2X1 exu_U16478(.A(alu_spr_out[34]), .B(exu_n16157), .Y(exu_n30697));
INVX1 exu_U16479(.A(exu_n30697), .Y(exu_n3679));
AND2X1 exu_U16480(.A(alu_spr_out[33]), .B(exu_n16157), .Y(exu_n30699));
INVX1 exu_U16481(.A(exu_n30699), .Y(exu_n3680));
AND2X1 exu_U16482(.A(alu_spr_out[32]), .B(exu_n16157), .Y(exu_n30701));
INVX1 exu_U16483(.A(exu_n30701), .Y(exu_n3681));
AND2X1 exu_U16484(.A(alu_spr_out[31]), .B(exu_n16157), .Y(exu_n30703));
INVX1 exu_U16485(.A(exu_n30703), .Y(exu_n3682));
AND2X1 exu_U16486(.A(alu_spr_out[30]), .B(exu_n16157), .Y(exu_n30705));
INVX1 exu_U16487(.A(exu_n30705), .Y(exu_n3683));
AND2X1 exu_U16488(.A(alu_spr_out[2]), .B(exu_n16157), .Y(exu_n30707));
INVX1 exu_U16489(.A(exu_n30707), .Y(exu_n3684));
AND2X1 exu_U16490(.A(alu_spr_out[29]), .B(exu_n16157), .Y(exu_n30709));
INVX1 exu_U16491(.A(exu_n30709), .Y(exu_n3685));
AND2X1 exu_U16492(.A(alu_spr_out[28]), .B(exu_n16158), .Y(exu_n30711));
INVX1 exu_U16493(.A(exu_n30711), .Y(exu_n3686));
AND2X1 exu_U16494(.A(alu_spr_out[27]), .B(exu_n16158), .Y(exu_n30713));
INVX1 exu_U16495(.A(exu_n30713), .Y(exu_n3687));
AND2X1 exu_U16496(.A(alu_spr_out[26]), .B(exu_n16158), .Y(exu_n30715));
INVX1 exu_U16497(.A(exu_n30715), .Y(exu_n3688));
AND2X1 exu_U16498(.A(alu_spr_out[25]), .B(exu_n16158), .Y(exu_n30717));
INVX1 exu_U16499(.A(exu_n30717), .Y(exu_n3689));
AND2X1 exu_U16500(.A(alu_spr_out[24]), .B(exu_n16158), .Y(exu_n30719));
INVX1 exu_U16501(.A(exu_n30719), .Y(exu_n3690));
AND2X1 exu_U16502(.A(alu_spr_out[23]), .B(exu_n16158), .Y(exu_n30721));
INVX1 exu_U16503(.A(exu_n30721), .Y(exu_n3691));
AND2X1 exu_U16504(.A(alu_spr_out[22]), .B(exu_n16158), .Y(exu_n30723));
INVX1 exu_U16505(.A(exu_n30723), .Y(exu_n3692));
AND2X1 exu_U16506(.A(alu_spr_out[21]), .B(exu_n16158), .Y(exu_n30725));
INVX1 exu_U16507(.A(exu_n30725), .Y(exu_n3693));
AND2X1 exu_U16508(.A(alu_spr_out[20]), .B(exu_n16158), .Y(exu_n30727));
INVX1 exu_U16509(.A(exu_n30727), .Y(exu_n3694));
AND2X1 exu_U16510(.A(alu_spr_out[1]), .B(exu_n16158), .Y(exu_n30729));
INVX1 exu_U16511(.A(exu_n30729), .Y(exu_n3695));
AND2X1 exu_U16512(.A(alu_spr_out[19]), .B(exu_n16158), .Y(exu_n30731));
INVX1 exu_U16513(.A(exu_n30731), .Y(exu_n3696));
AND2X1 exu_U16514(.A(alu_spr_out[18]), .B(exu_n16158), .Y(exu_n30733));
INVX1 exu_U16515(.A(exu_n30733), .Y(exu_n3697));
AND2X1 exu_U16516(.A(alu_spr_out[17]), .B(exu_n16158), .Y(exu_n30735));
INVX1 exu_U16517(.A(exu_n30735), .Y(exu_n3698));
AND2X1 exu_U16518(.A(alu_spr_out[16]), .B(exu_n16158), .Y(exu_n30737));
INVX1 exu_U16519(.A(exu_n30737), .Y(exu_n3699));
AND2X1 exu_U16520(.A(alu_spr_out[15]), .B(ecl_sel_sum_e), .Y(exu_n30739));
INVX1 exu_U16521(.A(exu_n30739), .Y(exu_n3700));
AND2X1 exu_U16522(.A(alu_spr_out[14]), .B(ecl_sel_sum_e), .Y(exu_n30741));
INVX1 exu_U16523(.A(exu_n30741), .Y(exu_n3701));
AND2X1 exu_U16524(.A(alu_spr_out[13]), .B(ecl_sel_sum_e), .Y(exu_n30743));
INVX1 exu_U16525(.A(exu_n30743), .Y(exu_n3702));
AND2X1 exu_U16526(.A(alu_spr_out[12]), .B(ecl_sel_sum_e), .Y(exu_n30745));
INVX1 exu_U16527(.A(exu_n30745), .Y(exu_n3703));
AND2X1 exu_U16528(.A(alu_spr_out[11]), .B(ecl_sel_sum_e), .Y(exu_n30747));
INVX1 exu_U16529(.A(exu_n30747), .Y(exu_n3704));
AND2X1 exu_U16530(.A(alu_spr_out[10]), .B(ecl_sel_sum_e), .Y(exu_n30749));
INVX1 exu_U16531(.A(exu_n30749), .Y(exu_n3705));
AND2X1 exu_U16532(.A(alu_spr_out[0]), .B(exu_n16155), .Y(exu_n30751));
INVX1 exu_U16533(.A(exu_n30751), .Y(exu_n3706));
AND2X1 exu_U16534(.A(exu_n16194), .B(div_curr_q[9]), .Y(exu_n30946));
INVX1 exu_U16535(.A(exu_n30946), .Y(exu_n3707));
AND2X1 exu_U16536(.A(div_curr_q[8]), .B(exu_n16195), .Y(exu_n30947));
INVX1 exu_U16537(.A(exu_n30947), .Y(exu_n3708));
AND2X1 exu_U16538(.A(div_curr_q[7]), .B(exu_n16195), .Y(exu_n30949));
INVX1 exu_U16539(.A(exu_n30949), .Y(exu_n3709));
AND2X1 exu_U16540(.A(div_curr_q[6]), .B(exu_n16193), .Y(exu_n30951));
INVX1 exu_U16541(.A(exu_n30951), .Y(exu_n3710));
AND2X1 exu_U16542(.A(div_ecl_d_msb), .B(ecl_div_sel_div), .Y(exu_n30953));
INVX1 exu_U16543(.A(exu_n30953), .Y(exu_n3711));
AND2X1 exu_U16544(.A(div_curr_q[62]), .B(exu_n16194), .Y(exu_n30955));
INVX1 exu_U16545(.A(exu_n30955), .Y(exu_n3712));
AND2X1 exu_U16546(.A(div_curr_q[61]), .B(exu_n16197), .Y(exu_n30957));
INVX1 exu_U16547(.A(exu_n30957), .Y(exu_n3713));
AND2X1 exu_U16548(.A(div_curr_q[60]), .B(exu_n16194), .Y(exu_n30959));
INVX1 exu_U16549(.A(exu_n30959), .Y(exu_n3714));
AND2X1 exu_U16550(.A(div_curr_q[5]), .B(exu_n16197), .Y(exu_n30961));
INVX1 exu_U16551(.A(exu_n30961), .Y(exu_n3715));
AND2X1 exu_U16552(.A(div_curr_q[59]), .B(exu_n16197), .Y(exu_n30963));
INVX1 exu_U16553(.A(exu_n30963), .Y(exu_n3716));
AND2X1 exu_U16554(.A(div_curr_q[58]), .B(exu_n16195), .Y(exu_n30965));
INVX1 exu_U16555(.A(exu_n30965), .Y(exu_n3717));
AND2X1 exu_U16556(.A(div_curr_q[57]), .B(exu_n16193), .Y(exu_n30967));
INVX1 exu_U16557(.A(exu_n30967), .Y(exu_n3718));
AND2X1 exu_U16558(.A(div_curr_q[56]), .B(ecl_div_sel_div), .Y(exu_n30969));
INVX1 exu_U16559(.A(exu_n30969), .Y(exu_n3719));
AND2X1 exu_U16560(.A(div_curr_q[55]), .B(exu_n16197), .Y(exu_n30971));
INVX1 exu_U16561(.A(exu_n30971), .Y(exu_n3720));
AND2X1 exu_U16562(.A(div_curr_q[54]), .B(exu_n16194), .Y(exu_n30973));
INVX1 exu_U16563(.A(exu_n30973), .Y(exu_n3721));
AND2X1 exu_U16564(.A(div_curr_q[53]), .B(exu_n16197), .Y(exu_n30975));
INVX1 exu_U16565(.A(exu_n30975), .Y(exu_n3722));
AND2X1 exu_U16566(.A(div_curr_q[52]), .B(ecl_div_sel_div), .Y(exu_n30977));
INVX1 exu_U16567(.A(exu_n30977), .Y(exu_n3723));
AND2X1 exu_U16568(.A(div_curr_q[51]), .B(exu_n16195), .Y(exu_n30979));
INVX1 exu_U16569(.A(exu_n30979), .Y(exu_n3724));
AND2X1 exu_U16570(.A(div_curr_q[50]), .B(exu_n16193), .Y(exu_n30981));
INVX1 exu_U16571(.A(exu_n30981), .Y(exu_n3725));
AND2X1 exu_U16572(.A(div_curr_q[4]), .B(exu_n16193), .Y(exu_n30983));
INVX1 exu_U16573(.A(exu_n30983), .Y(exu_n3726));
AND2X1 exu_U16574(.A(div_curr_q[49]), .B(ecl_div_sel_div), .Y(exu_n30985));
INVX1 exu_U16575(.A(exu_n30985), .Y(exu_n3727));
AND2X1 exu_U16576(.A(div_curr_q[48]), .B(exu_n16195), .Y(exu_n30987));
INVX1 exu_U16577(.A(exu_n30987), .Y(exu_n3728));
AND2X1 exu_U16578(.A(div_curr_q[47]), .B(exu_n16193), .Y(exu_n30989));
INVX1 exu_U16579(.A(exu_n30989), .Y(exu_n3729));
AND2X1 exu_U16580(.A(div_curr_q[46]), .B(exu_n16195), .Y(exu_n30991));
INVX1 exu_U16581(.A(exu_n30991), .Y(exu_n3730));
AND2X1 exu_U16582(.A(div_curr_q[45]), .B(ecl_div_sel_div), .Y(exu_n30993));
INVX1 exu_U16583(.A(exu_n30993), .Y(exu_n3731));
AND2X1 exu_U16584(.A(div_curr_q[44]), .B(exu_n16194), .Y(exu_n30995));
INVX1 exu_U16585(.A(exu_n30995), .Y(exu_n3732));
AND2X1 exu_U16586(.A(div_curr_q[43]), .B(exu_n16194), .Y(exu_n30997));
INVX1 exu_U16587(.A(exu_n30997), .Y(exu_n3733));
AND2X1 exu_U16588(.A(div_curr_q[42]), .B(exu_n16197), .Y(exu_n30999));
INVX1 exu_U16589(.A(exu_n30999), .Y(exu_n3734));
AND2X1 exu_U16590(.A(div_curr_q[41]), .B(ecl_div_sel_div), .Y(exu_n31001));
INVX1 exu_U16591(.A(exu_n31001), .Y(exu_n3735));
AND2X1 exu_U16592(.A(div_curr_q[40]), .B(exu_n16197), .Y(exu_n31003));
INVX1 exu_U16593(.A(exu_n31003), .Y(exu_n3736));
AND2X1 exu_U16594(.A(div_curr_q[3]), .B(exu_n16197), .Y(exu_n31005));
INVX1 exu_U16595(.A(exu_n31005), .Y(exu_n3737));
AND2X1 exu_U16596(.A(div_curr_q[39]), .B(exu_n16195), .Y(exu_n31007));
INVX1 exu_U16597(.A(exu_n31007), .Y(exu_n3738));
AND2X1 exu_U16598(.A(div_curr_q[38]), .B(ecl_div_sel_div), .Y(exu_n31009));
INVX1 exu_U16599(.A(exu_n31009), .Y(exu_n3739));
AND2X1 exu_U16600(.A(div_curr_q[37]), .B(exu_n16193), .Y(exu_n31011));
INVX1 exu_U16601(.A(exu_n31011), .Y(exu_n3740));
AND2X1 exu_U16602(.A(div_curr_q[36]), .B(exu_n16193), .Y(exu_n31013));
INVX1 exu_U16603(.A(exu_n31013), .Y(exu_n3741));
AND2X1 exu_U16604(.A(div_curr_q[35]), .B(exu_n16193), .Y(exu_n31015));
INVX1 exu_U16605(.A(exu_n31015), .Y(exu_n3742));
AND2X1 exu_U16606(.A(div_curr_q[34]), .B(exu_n16193), .Y(exu_n31017));
INVX1 exu_U16607(.A(exu_n31017), .Y(exu_n3743));
AND2X1 exu_U16608(.A(div_curr_q[33]), .B(exu_n16194), .Y(exu_n31019));
INVX1 exu_U16609(.A(exu_n31019), .Y(exu_n3744));
AND2X1 exu_U16610(.A(div_curr_q[32]), .B(exu_n16193), .Y(exu_n31021));
INVX1 exu_U16611(.A(exu_n31021), .Y(exu_n3745));
AND2X1 exu_U16612(.A(div_curr_q[31]), .B(exu_n16195), .Y(exu_n31023));
INVX1 exu_U16613(.A(exu_n31023), .Y(exu_n3746));
AND2X1 exu_U16614(.A(div_curr_q[30]), .B(ecl_div_sel_div), .Y(exu_n31025));
INVX1 exu_U16615(.A(exu_n31025), .Y(exu_n3747));
AND2X1 exu_U16616(.A(div_curr_q[2]), .B(exu_n16197), .Y(exu_n31027));
INVX1 exu_U16617(.A(exu_n31027), .Y(exu_n3748));
AND2X1 exu_U16618(.A(div_curr_q[29]), .B(exu_n16194), .Y(exu_n31029));
INVX1 exu_U16619(.A(exu_n31029), .Y(exu_n3749));
AND2X1 exu_U16620(.A(div_curr_q[28]), .B(exu_n16193), .Y(exu_n31031));
INVX1 exu_U16621(.A(exu_n31031), .Y(exu_n3750));
AND2X1 exu_U16622(.A(div_curr_q[27]), .B(exu_n16194), .Y(exu_n31033));
INVX1 exu_U16623(.A(exu_n31033), .Y(exu_n3751));
AND2X1 exu_U16624(.A(div_curr_q[26]), .B(exu_n16197), .Y(exu_n31035));
INVX1 exu_U16625(.A(exu_n31035), .Y(exu_n3752));
AND2X1 exu_U16626(.A(div_curr_q[25]), .B(exu_n16193), .Y(exu_n31037));
INVX1 exu_U16627(.A(exu_n31037), .Y(exu_n3753));
AND2X1 exu_U16628(.A(div_curr_q[24]), .B(ecl_div_sel_div), .Y(exu_n31039));
INVX1 exu_U16629(.A(exu_n31039), .Y(exu_n3754));
AND2X1 exu_U16630(.A(div_curr_q[23]), .B(exu_n16193), .Y(exu_n31041));
INVX1 exu_U16631(.A(exu_n31041), .Y(exu_n3755));
AND2X1 exu_U16632(.A(div_curr_q[22]), .B(exu_n16195), .Y(exu_n31043));
INVX1 exu_U16633(.A(exu_n31043), .Y(exu_n3756));
AND2X1 exu_U16634(.A(div_curr_q[21]), .B(exu_n16193), .Y(exu_n31045));
INVX1 exu_U16635(.A(exu_n31045), .Y(exu_n3757));
AND2X1 exu_U16636(.A(div_curr_q[20]), .B(exu_n16195), .Y(exu_n31047));
INVX1 exu_U16637(.A(exu_n31047), .Y(exu_n3758));
AND2X1 exu_U16638(.A(div_curr_q[1]), .B(exu_n16193), .Y(exu_n31049));
INVX1 exu_U16639(.A(exu_n31049), .Y(exu_n3759));
AND2X1 exu_U16640(.A(div_curr_q[19]), .B(exu_n16195), .Y(exu_n31051));
INVX1 exu_U16641(.A(exu_n31051), .Y(exu_n3760));
AND2X1 exu_U16642(.A(div_curr_q[18]), .B(exu_n16193), .Y(exu_n31053));
INVX1 exu_U16643(.A(exu_n31053), .Y(exu_n3761));
AND2X1 exu_U16644(.A(div_curr_q[17]), .B(ecl_div_sel_div), .Y(exu_n31055));
INVX1 exu_U16645(.A(exu_n31055), .Y(exu_n3762));
AND2X1 exu_U16646(.A(div_curr_q[16]), .B(exu_n16194), .Y(exu_n31057));
INVX1 exu_U16647(.A(exu_n31057), .Y(exu_n3763));
AND2X1 exu_U16648(.A(div_curr_q[15]), .B(exu_n16195), .Y(exu_n31059));
INVX1 exu_U16649(.A(exu_n31059), .Y(exu_n3764));
AND2X1 exu_U16650(.A(div_curr_q[14]), .B(exu_n16193), .Y(exu_n31061));
INVX1 exu_U16651(.A(exu_n31061), .Y(exu_n3765));
AND2X1 exu_U16652(.A(div_curr_q[13]), .B(ecl_div_sel_div), .Y(exu_n31063));
INVX1 exu_U16653(.A(exu_n31063), .Y(exu_n3766));
AND2X1 exu_U16654(.A(div_curr_q[12]), .B(exu_n16197), .Y(exu_n31065));
INVX1 exu_U16655(.A(exu_n31065), .Y(exu_n3767));
AND2X1 exu_U16656(.A(div_curr_q[11]), .B(exu_n16197), .Y(exu_n31067));
INVX1 exu_U16657(.A(exu_n31067), .Y(exu_n3768));
AND2X1 exu_U16658(.A(div_curr_q[10]), .B(exu_n16197), .Y(exu_n31069));
INVX1 exu_U16659(.A(exu_n31069), .Y(exu_n3769));
AND2X1 exu_U16660(.A(div_curr_q[0]), .B(exu_n16197), .Y(exu_n31071));
INVX1 exu_U16661(.A(exu_n31071), .Y(exu_n3770));
AND2X1 exu_U16662(.A(ecl_div_last_cycle), .B(div_d[8]), .Y(exu_n31073));
INVX1 exu_U16663(.A(exu_n31073), .Y(exu_n3771));
AND2X1 exu_U16664(.A(div_d[7]), .B(ecl_div_last_cycle), .Y(exu_n31075));
INVX1 exu_U16665(.A(exu_n31075), .Y(exu_n3772));
AND2X1 exu_U16666(.A(div_d[6]), .B(ecl_div_last_cycle), .Y(exu_n31077));
INVX1 exu_U16667(.A(exu_n31077), .Y(exu_n3773));
AND2X1 exu_U16668(.A(div_d[5]), .B(ecl_div_last_cycle), .Y(exu_n31079));
INVX1 exu_U16669(.A(exu_n31079), .Y(exu_n3774));
AND2X1 exu_U16670(.A(div_ecl_d_62), .B(ecl_div_last_cycle), .Y(exu_n31081));
INVX1 exu_U16671(.A(exu_n31081), .Y(exu_n3775));
AND2X1 exu_U16672(.A(div_d[61]), .B(ecl_div_last_cycle), .Y(exu_n31083));
INVX1 exu_U16673(.A(exu_n31083), .Y(exu_n3776));
AND2X1 exu_U16674(.A(div_d[60]), .B(ecl_div_last_cycle), .Y(exu_n31085));
INVX1 exu_U16675(.A(exu_n31085), .Y(exu_n3777));
AND2X1 exu_U16676(.A(div_d[59]), .B(ecl_div_last_cycle), .Y(exu_n31087));
INVX1 exu_U16677(.A(exu_n31087), .Y(exu_n3778));
AND2X1 exu_U16678(.A(div_d[4]), .B(ecl_div_last_cycle), .Y(exu_n31089));
INVX1 exu_U16679(.A(exu_n31089), .Y(exu_n3779));
AND2X1 exu_U16680(.A(div_d[58]), .B(ecl_div_last_cycle), .Y(exu_n31091));
INVX1 exu_U16681(.A(exu_n31091), .Y(exu_n3780));
AND2X1 exu_U16682(.A(div_d[57]), .B(ecl_div_last_cycle), .Y(exu_n31093));
INVX1 exu_U16683(.A(exu_n31093), .Y(exu_n3781));
AND2X1 exu_U16684(.A(div_d[56]), .B(ecl_div_last_cycle), .Y(exu_n31095));
INVX1 exu_U16685(.A(exu_n31095), .Y(exu_n3782));
AND2X1 exu_U16686(.A(div_d[55]), .B(ecl_div_last_cycle), .Y(exu_n31097));
INVX1 exu_U16687(.A(exu_n31097), .Y(exu_n3783));
AND2X1 exu_U16688(.A(div_d[54]), .B(ecl_div_last_cycle), .Y(exu_n31099));
INVX1 exu_U16689(.A(exu_n31099), .Y(exu_n3784));
AND2X1 exu_U16690(.A(div_d[53]), .B(ecl_div_last_cycle), .Y(exu_n31101));
INVX1 exu_U16691(.A(exu_n31101), .Y(exu_n3785));
AND2X1 exu_U16692(.A(div_d[52]), .B(ecl_div_last_cycle), .Y(exu_n31103));
INVX1 exu_U16693(.A(exu_n31103), .Y(exu_n3786));
AND2X1 exu_U16694(.A(div_d[51]), .B(ecl_div_last_cycle), .Y(exu_n31105));
INVX1 exu_U16695(.A(exu_n31105), .Y(exu_n3787));
AND2X1 exu_U16696(.A(div_d[50]), .B(ecl_div_last_cycle), .Y(exu_n31107));
INVX1 exu_U16697(.A(exu_n31107), .Y(exu_n3788));
AND2X1 exu_U16698(.A(div_d[49]), .B(ecl_div_last_cycle), .Y(exu_n31109));
INVX1 exu_U16699(.A(exu_n31109), .Y(exu_n3789));
AND2X1 exu_U16700(.A(div_d[3]), .B(ecl_div_last_cycle), .Y(exu_n31111));
INVX1 exu_U16701(.A(exu_n31111), .Y(exu_n3790));
AND2X1 exu_U16702(.A(div_d[48]), .B(ecl_div_last_cycle), .Y(exu_n31113));
INVX1 exu_U16703(.A(exu_n31113), .Y(exu_n3791));
AND2X1 exu_U16704(.A(div_d[47]), .B(ecl_div_last_cycle), .Y(exu_n31115));
INVX1 exu_U16705(.A(exu_n31115), .Y(exu_n3792));
AND2X1 exu_U16706(.A(div_d[46]), .B(ecl_div_last_cycle), .Y(exu_n31117));
INVX1 exu_U16707(.A(exu_n31117), .Y(exu_n3793));
AND2X1 exu_U16708(.A(div_d[45]), .B(ecl_div_last_cycle), .Y(exu_n31119));
INVX1 exu_U16709(.A(exu_n31119), .Y(exu_n3794));
AND2X1 exu_U16710(.A(div_d[44]), .B(ecl_div_last_cycle), .Y(exu_n31121));
INVX1 exu_U16711(.A(exu_n31121), .Y(exu_n3795));
AND2X1 exu_U16712(.A(div_d[43]), .B(ecl_div_last_cycle), .Y(exu_n31123));
INVX1 exu_U16713(.A(exu_n31123), .Y(exu_n3796));
AND2X1 exu_U16714(.A(div_d[42]), .B(ecl_div_last_cycle), .Y(exu_n31125));
INVX1 exu_U16715(.A(exu_n31125), .Y(exu_n3797));
AND2X1 exu_U16716(.A(div_d[41]), .B(ecl_div_last_cycle), .Y(exu_n31127));
INVX1 exu_U16717(.A(exu_n31127), .Y(exu_n3798));
AND2X1 exu_U16718(.A(div_d[40]), .B(ecl_div_last_cycle), .Y(exu_n31129));
INVX1 exu_U16719(.A(exu_n31129), .Y(exu_n3799));
AND2X1 exu_U16720(.A(div_d[39]), .B(ecl_div_last_cycle), .Y(exu_n31131));
INVX1 exu_U16721(.A(exu_n31131), .Y(exu_n3800));
AND2X1 exu_U16722(.A(div_d[2]), .B(ecl_div_last_cycle), .Y(exu_n31133));
INVX1 exu_U16723(.A(exu_n31133), .Y(exu_n3801));
AND2X1 exu_U16724(.A(div_d[38]), .B(ecl_div_last_cycle), .Y(exu_n31135));
INVX1 exu_U16725(.A(exu_n31135), .Y(exu_n3802));
AND2X1 exu_U16726(.A(div_d[37]), .B(ecl_div_last_cycle), .Y(exu_n31137));
INVX1 exu_U16727(.A(exu_n31137), .Y(exu_n3803));
AND2X1 exu_U16728(.A(div_d[36]), .B(ecl_div_last_cycle), .Y(exu_n31139));
INVX1 exu_U16729(.A(exu_n31139), .Y(exu_n3804));
AND2X1 exu_U16730(.A(div_d[35]), .B(ecl_div_last_cycle), .Y(exu_n31141));
INVX1 exu_U16731(.A(exu_n31141), .Y(exu_n3805));
AND2X1 exu_U16732(.A(div_d[34]), .B(ecl_div_last_cycle), .Y(exu_n31143));
INVX1 exu_U16733(.A(exu_n31143), .Y(exu_n3806));
AND2X1 exu_U16734(.A(div_d[33]), .B(ecl_div_last_cycle), .Y(exu_n31145));
INVX1 exu_U16735(.A(exu_n31145), .Y(exu_n3807));
AND2X1 exu_U16736(.A(div_d[32]), .B(ecl_div_last_cycle), .Y(exu_n31147));
INVX1 exu_U16737(.A(exu_n31147), .Y(exu_n3808));
AND2X1 exu_U16738(.A(div_d[31]), .B(ecl_div_last_cycle), .Y(exu_n31149));
INVX1 exu_U16739(.A(exu_n31149), .Y(exu_n3809));
AND2X1 exu_U16740(.A(div_d[30]), .B(ecl_div_last_cycle), .Y(exu_n31151));
INVX1 exu_U16741(.A(exu_n31151), .Y(exu_n3810));
AND2X1 exu_U16742(.A(div_d[29]), .B(ecl_div_last_cycle), .Y(exu_n31153));
INVX1 exu_U16743(.A(exu_n31153), .Y(exu_n3811));
AND2X1 exu_U16744(.A(div_d[1]), .B(ecl_div_last_cycle), .Y(exu_n31155));
INVX1 exu_U16745(.A(exu_n31155), .Y(exu_n3812));
AND2X1 exu_U16746(.A(div_d[28]), .B(ecl_div_last_cycle), .Y(exu_n31157));
INVX1 exu_U16747(.A(exu_n31157), .Y(exu_n3813));
AND2X1 exu_U16748(.A(div_d[27]), .B(ecl_div_last_cycle), .Y(exu_n31159));
INVX1 exu_U16749(.A(exu_n31159), .Y(exu_n3814));
AND2X1 exu_U16750(.A(div_d[26]), .B(ecl_div_last_cycle), .Y(exu_n31161));
INVX1 exu_U16751(.A(exu_n31161), .Y(exu_n3815));
AND2X1 exu_U16752(.A(div_d[25]), .B(ecl_div_last_cycle), .Y(exu_n31163));
INVX1 exu_U16753(.A(exu_n31163), .Y(exu_n3816));
AND2X1 exu_U16754(.A(div_d[24]), .B(ecl_div_last_cycle), .Y(exu_n31165));
INVX1 exu_U16755(.A(exu_n31165), .Y(exu_n3817));
AND2X1 exu_U16756(.A(div_d[23]), .B(ecl_div_last_cycle), .Y(exu_n31167));
INVX1 exu_U16757(.A(exu_n31167), .Y(exu_n3818));
AND2X1 exu_U16758(.A(div_d[22]), .B(ecl_div_last_cycle), .Y(exu_n31169));
INVX1 exu_U16759(.A(exu_n31169), .Y(exu_n3819));
AND2X1 exu_U16760(.A(div_d[21]), .B(ecl_div_last_cycle), .Y(exu_n31171));
INVX1 exu_U16761(.A(exu_n31171), .Y(exu_n3820));
AND2X1 exu_U16762(.A(div_d[20]), .B(ecl_div_last_cycle), .Y(exu_n31173));
INVX1 exu_U16763(.A(exu_n31173), .Y(exu_n3821));
AND2X1 exu_U16764(.A(div_d[19]), .B(ecl_div_last_cycle), .Y(exu_n31175));
INVX1 exu_U16765(.A(exu_n31175), .Y(exu_n3822));
AND2X1 exu_U16766(.A(div_d[0]), .B(ecl_div_last_cycle), .Y(exu_n31177));
INVX1 exu_U16767(.A(exu_n31177), .Y(exu_n3823));
AND2X1 exu_U16768(.A(div_d[18]), .B(ecl_div_last_cycle), .Y(exu_n31179));
INVX1 exu_U16769(.A(exu_n31179), .Y(exu_n3824));
AND2X1 exu_U16770(.A(div_d[17]), .B(ecl_div_last_cycle), .Y(exu_n31181));
INVX1 exu_U16771(.A(exu_n31181), .Y(exu_n3825));
AND2X1 exu_U16772(.A(div_d[16]), .B(ecl_div_last_cycle), .Y(exu_n31183));
INVX1 exu_U16773(.A(exu_n31183), .Y(exu_n3826));
AND2X1 exu_U16774(.A(div_d[15]), .B(ecl_div_last_cycle), .Y(exu_n31185));
INVX1 exu_U16775(.A(exu_n31185), .Y(exu_n3827));
AND2X1 exu_U16776(.A(div_d[14]), .B(ecl_div_last_cycle), .Y(exu_n31187));
INVX1 exu_U16777(.A(exu_n31187), .Y(exu_n3828));
AND2X1 exu_U16778(.A(div_d[13]), .B(ecl_div_last_cycle), .Y(exu_n31189));
INVX1 exu_U16779(.A(exu_n31189), .Y(exu_n3829));
AND2X1 exu_U16780(.A(div_d[12]), .B(ecl_div_last_cycle), .Y(exu_n31191));
INVX1 exu_U16781(.A(exu_n31191), .Y(exu_n3830));
AND2X1 exu_U16782(.A(div_d[11]), .B(ecl_div_last_cycle), .Y(exu_n31193));
INVX1 exu_U16783(.A(exu_n31193), .Y(exu_n3831));
AND2X1 exu_U16784(.A(div_d[10]), .B(ecl_div_last_cycle), .Y(exu_n31195));
INVX1 exu_U16785(.A(exu_n31195), .Y(exu_n3832));
AND2X1 exu_U16786(.A(div_d[9]), .B(ecl_div_last_cycle), .Y(exu_n31197));
INVX1 exu_U16787(.A(exu_n31197), .Y(exu_n3833));
AND2X1 exu_U16788(.A(ecl_div_newq), .B(ecl_div_last_cycle), .Y(exu_n31199));
INVX1 exu_U16789(.A(exu_n31199), .Y(exu_n3834));
AND2X1 exu_U16790(.A(ecl_div_ld_inputs), .B(div_xin[9]), .Y(exu_n31201));
INVX1 exu_U16791(.A(exu_n31201), .Y(exu_n3835));
AND2X1 exu_U16792(.A(div_xin[8]), .B(ecl_div_ld_inputs), .Y(exu_n31203));
INVX1 exu_U16793(.A(exu_n31203), .Y(exu_n3836));
AND2X1 exu_U16794(.A(div_xin[7]), .B(exu_n16204), .Y(exu_n31205));
INVX1 exu_U16795(.A(exu_n31205), .Y(exu_n3837));
AND2X1 exu_U16796(.A(div_xin[6]), .B(exu_n16203), .Y(exu_n31207));
INVX1 exu_U16797(.A(exu_n31207), .Y(exu_n3838));
AND2X1 exu_U16798(.A(exu_n15492), .B(exu_n16204), .Y(exu_n31209));
INVX1 exu_U16799(.A(exu_n31209), .Y(exu_n3839));
AND2X1 exu_U16800(.A(exu_n15247), .B(ecl_div_ld_inputs), .Y(exu_n31211));
INVX1 exu_U16801(.A(exu_n31211), .Y(exu_n3840));
AND2X1 exu_U16802(.A(exu_n15249), .B(exu_n16204), .Y(exu_n31213));
INVX1 exu_U16803(.A(exu_n31213), .Y(exu_n3841));
AND2X1 exu_U16804(.A(exu_n15250), .B(exu_n16203), .Y(exu_n31215));
INVX1 exu_U16805(.A(exu_n31215), .Y(exu_n3842));
AND2X1 exu_U16806(.A(div_xin[5]), .B(exu_n16204), .Y(exu_n31217));
INVX1 exu_U16807(.A(exu_n31217), .Y(exu_n3843));
AND2X1 exu_U16808(.A(exu_n15251), .B(ecl_div_ld_inputs), .Y(exu_n31219));
INVX1 exu_U16809(.A(exu_n31219), .Y(exu_n3844));
AND2X1 exu_U16810(.A(exu_n15252), .B(exu_n16209), .Y(exu_n31221));
INVX1 exu_U16811(.A(exu_n31221), .Y(exu_n3845));
AND2X1 exu_U16812(.A(exu_n15253), .B(exu_n16210), .Y(exu_n31223));
INVX1 exu_U16813(.A(exu_n31223), .Y(exu_n3846));
AND2X1 exu_U16814(.A(exu_n15254), .B(exu_n16207), .Y(exu_n31225));
INVX1 exu_U16815(.A(exu_n31225), .Y(exu_n3847));
AND2X1 exu_U16816(.A(exu_n15255), .B(exu_n16208), .Y(exu_n31227));
INVX1 exu_U16817(.A(exu_n31227), .Y(exu_n3848));
AND2X1 exu_U16818(.A(exu_n15256), .B(exu_n16211), .Y(exu_n31229));
INVX1 exu_U16819(.A(exu_n31229), .Y(exu_n3849));
AND2X1 exu_U16820(.A(exu_n15257), .B(exu_n16212), .Y(exu_n31231));
INVX1 exu_U16821(.A(exu_n31231), .Y(exu_n3850));
AND2X1 exu_U16822(.A(exu_n15258), .B(exu_n16214), .Y(exu_n31233));
INVX1 exu_U16823(.A(exu_n31233), .Y(exu_n3851));
AND2X1 exu_U16824(.A(exu_n15260), .B(ecl_div_ld_inputs), .Y(exu_n31235));
INVX1 exu_U16825(.A(exu_n31235), .Y(exu_n3852));
AND2X1 exu_U16826(.A(exu_n15261), .B(exu_n16203), .Y(exu_n31237));
INVX1 exu_U16827(.A(exu_n31237), .Y(exu_n3853));
AND2X1 exu_U16828(.A(div_xin[4]), .B(exu_n16213), .Y(exu_n31239));
INVX1 exu_U16829(.A(exu_n31239), .Y(exu_n3854));
AND2X1 exu_U16830(.A(exu_n15262), .B(exu_n16204), .Y(exu_n31241));
INVX1 exu_U16831(.A(exu_n31241), .Y(exu_n3855));
AND2X1 exu_U16832(.A(exu_n15263), .B(exu_n16209), .Y(exu_n31243));
INVX1 exu_U16833(.A(exu_n31243), .Y(exu_n3856));
AND2X1 exu_U16834(.A(exu_n15264), .B(exu_n16210), .Y(exu_n31245));
INVX1 exu_U16835(.A(exu_n31245), .Y(exu_n3857));
AND2X1 exu_U16836(.A(exu_n15265), .B(exu_n16207), .Y(exu_n31247));
INVX1 exu_U16837(.A(exu_n31247), .Y(exu_n3858));
AND2X1 exu_U16838(.A(exu_n15266), .B(exu_n16203), .Y(exu_n31249));
INVX1 exu_U16839(.A(exu_n31249), .Y(exu_n3859));
AND2X1 exu_U16840(.A(exu_n15267), .B(exu_n16213), .Y(exu_n31251));
INVX1 exu_U16841(.A(exu_n31251), .Y(exu_n3860));
AND2X1 exu_U16842(.A(exu_n15268), .B(exu_n16204), .Y(exu_n31253));
INVX1 exu_U16843(.A(exu_n31253), .Y(exu_n3861));
AND2X1 exu_U16844(.A(exu_n15269), .B(exu_n16207), .Y(exu_n31255));
INVX1 exu_U16845(.A(exu_n31255), .Y(exu_n3862));
AND2X1 exu_U16846(.A(exu_n15240), .B(ecl_div_ld_inputs), .Y(exu_n31257));
INVX1 exu_U16847(.A(exu_n31257), .Y(exu_n3863));
AND2X1 exu_U16848(.A(exu_n15241), .B(exu_n16203), .Y(exu_n31259));
INVX1 exu_U16849(.A(exu_n31259), .Y(exu_n3864));
AND2X1 exu_U16850(.A(div_xin[3]), .B(exu_n16213), .Y(exu_n31261));
INVX1 exu_U16851(.A(exu_n31261), .Y(exu_n3865));
AND2X1 exu_U16852(.A(exu_n15242), .B(exu_n16204), .Y(exu_n31263));
INVX1 exu_U16853(.A(exu_n31263), .Y(exu_n3866));
AND2X1 exu_U16854(.A(exu_n15243), .B(exu_n16207), .Y(exu_n31265));
INVX1 exu_U16855(.A(exu_n31265), .Y(exu_n3867));
AND2X1 exu_U16856(.A(exu_n15244), .B(exu_n16214), .Y(exu_n31267));
INVX1 exu_U16857(.A(exu_n31267), .Y(exu_n3868));
AND2X1 exu_U16858(.A(exu_n15245), .B(ecl_div_ld_inputs), .Y(exu_n31269));
INVX1 exu_U16859(.A(exu_n31269), .Y(exu_n3869));
AND2X1 exu_U16860(.A(exu_n15246), .B(exu_n16203), .Y(exu_n31271));
INVX1 exu_U16861(.A(exu_n31271), .Y(exu_n3870));
AND2X1 exu_U16862(.A(exu_n15248), .B(exu_n16213), .Y(exu_n31273));
INVX1 exu_U16863(.A(exu_n31273), .Y(exu_n3871));
AND2X1 exu_U16864(.A(exu_n15259), .B(exu_n16204), .Y(exu_n31275));
INVX1 exu_U16865(.A(exu_n31275), .Y(exu_n3872));
AND2X1 exu_U16866(.A(exu_n15270), .B(exu_n16213), .Y(exu_n31277));
INVX1 exu_U16867(.A(exu_n31277), .Y(exu_n3873));
AND2X1 exu_U16868(.A(div_xin[31]), .B(exu_n16204), .Y(exu_n31279));
INVX1 exu_U16869(.A(exu_n31279), .Y(exu_n3874));
AND2X1 exu_U16870(.A(div_xin[30]), .B(exu_n16207), .Y(exu_n31281));
INVX1 exu_U16871(.A(exu_n31281), .Y(exu_n3875));
AND2X1 exu_U16872(.A(div_xin[2]), .B(ecl_div_ld_inputs), .Y(exu_n31283));
INVX1 exu_U16873(.A(exu_n31283), .Y(exu_n3876));
AND2X1 exu_U16874(.A(div_xin[29]), .B(exu_n16203), .Y(exu_n31285));
INVX1 exu_U16875(.A(exu_n31285), .Y(exu_n3877));
AND2X1 exu_U16876(.A(div_xin[28]), .B(exu_n16213), .Y(exu_n31287));
INVX1 exu_U16877(.A(exu_n31287), .Y(exu_n3878));
AND2X1 exu_U16878(.A(div_xin[27]), .B(exu_n16204), .Y(exu_n31289));
INVX1 exu_U16879(.A(exu_n31289), .Y(exu_n3879));
AND2X1 exu_U16880(.A(div_xin[26]), .B(exu_n16207), .Y(exu_n31291));
INVX1 exu_U16881(.A(exu_n31291), .Y(exu_n3880));
AND2X1 exu_U16882(.A(div_xin[25]), .B(ecl_div_ld_inputs), .Y(exu_n31293));
INVX1 exu_U16883(.A(exu_n31293), .Y(exu_n3881));
AND2X1 exu_U16884(.A(div_xin[24]), .B(exu_n16203), .Y(exu_n31295));
INVX1 exu_U16885(.A(exu_n31295), .Y(exu_n3882));
AND2X1 exu_U16886(.A(div_xin[23]), .B(exu_n16213), .Y(exu_n31297));
INVX1 exu_U16887(.A(exu_n31297), .Y(exu_n3883));
AND2X1 exu_U16888(.A(div_xin[22]), .B(exu_n16204), .Y(exu_n31299));
INVX1 exu_U16889(.A(exu_n31299), .Y(exu_n3884));
AND2X1 exu_U16890(.A(div_xin[21]), .B(exu_n16207), .Y(exu_n31301));
INVX1 exu_U16891(.A(exu_n31301), .Y(exu_n3885));
AND2X1 exu_U16892(.A(div_xin[20]), .B(ecl_div_ld_inputs), .Y(exu_n31303));
INVX1 exu_U16893(.A(exu_n31303), .Y(exu_n3886));
AND2X1 exu_U16894(.A(div_xin[1]), .B(exu_n16214), .Y(exu_n31305));
INVX1 exu_U16895(.A(exu_n31305), .Y(exu_n3887));
AND2X1 exu_U16896(.A(div_xin[19]), .B(exu_n16214), .Y(exu_n31307));
INVX1 exu_U16897(.A(exu_n31307), .Y(exu_n3888));
AND2X1 exu_U16898(.A(div_xin[18]), .B(exu_n16214), .Y(exu_n31309));
INVX1 exu_U16899(.A(exu_n31309), .Y(exu_n3889));
AND2X1 exu_U16900(.A(div_xin[17]), .B(exu_n16214), .Y(exu_n31311));
INVX1 exu_U16901(.A(exu_n31311), .Y(exu_n3890));
AND2X1 exu_U16902(.A(div_xin[16]), .B(exu_n16214), .Y(exu_n31313));
INVX1 exu_U16903(.A(exu_n31313), .Y(exu_n3891));
AND2X1 exu_U16904(.A(div_xin[15]), .B(exu_n16214), .Y(exu_n31315));
INVX1 exu_U16905(.A(exu_n31315), .Y(exu_n3892));
AND2X1 exu_U16906(.A(div_xin[14]), .B(exu_n16214), .Y(exu_n31317));
INVX1 exu_U16907(.A(exu_n31317), .Y(exu_n3893));
AND2X1 exu_U16908(.A(div_xin[13]), .B(exu_n16214), .Y(exu_n31319));
INVX1 exu_U16909(.A(exu_n31319), .Y(exu_n3894));
AND2X1 exu_U16910(.A(div_xin[12]), .B(exu_n16214), .Y(exu_n31321));
INVX1 exu_U16911(.A(exu_n31321), .Y(exu_n3895));
AND2X1 exu_U16912(.A(div_xin[11]), .B(exu_n16214), .Y(exu_n31323));
INVX1 exu_U16913(.A(exu_n31323), .Y(exu_n3896));
AND2X1 exu_U16914(.A(div_xin[10]), .B(exu_n16214), .Y(exu_n31325));
INVX1 exu_U16915(.A(exu_n31325), .Y(exu_n3897));
AND2X1 exu_U16916(.A(div_xin[0]), .B(exu_n16214), .Y(exu_n31327));
INVX1 exu_U16917(.A(exu_n31327), .Y(exu_n3898));
AND2X1 exu_U16918(.A(exu_n11488), .B(exu_n10244), .Y(div_mul_result_next[9]));
INVX1 exu_U16919(.A(div_mul_result_next[9]), .Y(exu_n3899));
AND2X1 exu_U16920(.A(exu_n11489), .B(exu_n10245), .Y(div_mul_result_next[8]));
INVX1 exu_U16921(.A(div_mul_result_next[8]), .Y(exu_n3900));
AND2X1 exu_U16922(.A(exu_n11490), .B(exu_n10246), .Y(div_mul_result_next[7]));
INVX1 exu_U16923(.A(div_mul_result_next[7]), .Y(exu_n3901));
AND2X1 exu_U16924(.A(exu_n11491), .B(exu_n10247), .Y(div_mul_result_next[6]));
INVX1 exu_U16925(.A(div_mul_result_next[6]), .Y(exu_n3902));
AND2X1 exu_U16926(.A(exu_n11492), .B(exu_n10248), .Y(div_mul_result_next[63]));
INVX1 exu_U16927(.A(div_mul_result_next[63]), .Y(exu_n3903));
AND2X1 exu_U16928(.A(exu_n11493), .B(exu_n10249), .Y(div_mul_result_next[62]));
INVX1 exu_U16929(.A(div_mul_result_next[62]), .Y(exu_n3904));
AND2X1 exu_U16930(.A(exu_n11494), .B(exu_n10250), .Y(div_mul_result_next[61]));
INVX1 exu_U16931(.A(div_mul_result_next[61]), .Y(exu_n3905));
AND2X1 exu_U16932(.A(exu_n11495), .B(exu_n10251), .Y(div_mul_result_next[60]));
INVX1 exu_U16933(.A(div_mul_result_next[60]), .Y(exu_n3906));
AND2X1 exu_U16934(.A(exu_n11496), .B(exu_n10252), .Y(div_mul_result_next[5]));
INVX1 exu_U16935(.A(div_mul_result_next[5]), .Y(exu_n3907));
AND2X1 exu_U16936(.A(exu_n11497), .B(exu_n10253), .Y(div_mul_result_next[59]));
INVX1 exu_U16937(.A(div_mul_result_next[59]), .Y(exu_n3908));
AND2X1 exu_U16938(.A(exu_n11498), .B(exu_n10254), .Y(div_mul_result_next[58]));
INVX1 exu_U16939(.A(div_mul_result_next[58]), .Y(exu_n3909));
AND2X1 exu_U16940(.A(exu_n11499), .B(exu_n10255), .Y(div_mul_result_next[57]));
INVX1 exu_U16941(.A(div_mul_result_next[57]), .Y(exu_n3910));
AND2X1 exu_U16942(.A(exu_n11500), .B(exu_n10256), .Y(div_mul_result_next[56]));
INVX1 exu_U16943(.A(div_mul_result_next[56]), .Y(exu_n3911));
AND2X1 exu_U16944(.A(exu_n11501), .B(exu_n10257), .Y(div_mul_result_next[55]));
INVX1 exu_U16945(.A(div_mul_result_next[55]), .Y(exu_n3912));
AND2X1 exu_U16946(.A(exu_n11502), .B(exu_n10258), .Y(div_mul_result_next[54]));
INVX1 exu_U16947(.A(div_mul_result_next[54]), .Y(exu_n3913));
AND2X1 exu_U16948(.A(exu_n11503), .B(exu_n10259), .Y(div_mul_result_next[53]));
INVX1 exu_U16949(.A(div_mul_result_next[53]), .Y(exu_n3914));
AND2X1 exu_U16950(.A(exu_n11504), .B(exu_n10260), .Y(div_mul_result_next[52]));
INVX1 exu_U16951(.A(div_mul_result_next[52]), .Y(exu_n3915));
AND2X1 exu_U16952(.A(exu_n11505), .B(exu_n10261), .Y(div_mul_result_next[51]));
INVX1 exu_U16953(.A(div_mul_result_next[51]), .Y(exu_n3916));
AND2X1 exu_U16954(.A(exu_n11506), .B(exu_n10262), .Y(div_mul_result_next[50]));
INVX1 exu_U16955(.A(div_mul_result_next[50]), .Y(exu_n3917));
AND2X1 exu_U16956(.A(exu_n11507), .B(exu_n10263), .Y(div_mul_result_next[4]));
INVX1 exu_U16957(.A(div_mul_result_next[4]), .Y(exu_n3918));
AND2X1 exu_U16958(.A(exu_n11508), .B(exu_n10264), .Y(div_mul_result_next[49]));
INVX1 exu_U16959(.A(div_mul_result_next[49]), .Y(exu_n3919));
AND2X1 exu_U16960(.A(exu_n11509), .B(exu_n10265), .Y(div_mul_result_next[48]));
INVX1 exu_U16961(.A(div_mul_result_next[48]), .Y(exu_n3920));
AND2X1 exu_U16962(.A(exu_n11510), .B(exu_n10266), .Y(div_mul_result_next[47]));
INVX1 exu_U16963(.A(div_mul_result_next[47]), .Y(exu_n3921));
AND2X1 exu_U16964(.A(exu_n11511), .B(exu_n10267), .Y(div_mul_result_next[46]));
INVX1 exu_U16965(.A(div_mul_result_next[46]), .Y(exu_n3922));
AND2X1 exu_U16966(.A(exu_n11512), .B(exu_n10268), .Y(div_mul_result_next[45]));
INVX1 exu_U16967(.A(div_mul_result_next[45]), .Y(exu_n3923));
AND2X1 exu_U16968(.A(exu_n11513), .B(exu_n10269), .Y(div_mul_result_next[44]));
INVX1 exu_U16969(.A(div_mul_result_next[44]), .Y(exu_n3924));
AND2X1 exu_U16970(.A(exu_n11514), .B(exu_n10270), .Y(div_mul_result_next[43]));
INVX1 exu_U16971(.A(div_mul_result_next[43]), .Y(exu_n3925));
AND2X1 exu_U16972(.A(exu_n11515), .B(exu_n10271), .Y(div_mul_result_next[42]));
INVX1 exu_U16973(.A(div_mul_result_next[42]), .Y(exu_n3926));
AND2X1 exu_U16974(.A(exu_n11516), .B(exu_n10272), .Y(div_mul_result_next[41]));
INVX1 exu_U16975(.A(div_mul_result_next[41]), .Y(exu_n3927));
AND2X1 exu_U16976(.A(exu_n11517), .B(exu_n10273), .Y(div_mul_result_next[40]));
INVX1 exu_U16977(.A(div_mul_result_next[40]), .Y(exu_n3928));
AND2X1 exu_U16978(.A(exu_n11518), .B(exu_n10274), .Y(div_mul_result_next[3]));
INVX1 exu_U16979(.A(div_mul_result_next[3]), .Y(exu_n3929));
AND2X1 exu_U16980(.A(exu_n11519), .B(exu_n10275), .Y(div_mul_result_next[39]));
INVX1 exu_U16981(.A(div_mul_result_next[39]), .Y(exu_n3930));
AND2X1 exu_U16982(.A(exu_n11520), .B(exu_n10276), .Y(div_mul_result_next[38]));
INVX1 exu_U16983(.A(div_mul_result_next[38]), .Y(exu_n3931));
AND2X1 exu_U16984(.A(exu_n11521), .B(exu_n10277), .Y(div_mul_result_next[37]));
INVX1 exu_U16985(.A(div_mul_result_next[37]), .Y(exu_n3932));
AND2X1 exu_U16986(.A(exu_n11522), .B(exu_n10278), .Y(div_mul_result_next[36]));
INVX1 exu_U16987(.A(div_mul_result_next[36]), .Y(exu_n3933));
AND2X1 exu_U16988(.A(exu_n11523), .B(exu_n10279), .Y(div_mul_result_next[35]));
INVX1 exu_U16989(.A(div_mul_result_next[35]), .Y(exu_n3934));
AND2X1 exu_U16990(.A(exu_n11524), .B(exu_n10280), .Y(div_mul_result_next[34]));
INVX1 exu_U16991(.A(div_mul_result_next[34]), .Y(exu_n3935));
AND2X1 exu_U16992(.A(exu_n11525), .B(exu_n10281), .Y(div_mul_result_next[33]));
INVX1 exu_U16993(.A(div_mul_result_next[33]), .Y(exu_n3936));
AND2X1 exu_U16994(.A(exu_n11526), .B(exu_n10282), .Y(div_mul_result_next[32]));
INVX1 exu_U16995(.A(div_mul_result_next[32]), .Y(exu_n3937));
AND2X1 exu_U16996(.A(exu_n11527), .B(exu_n10283), .Y(div_mul_result_next[31]));
INVX1 exu_U16997(.A(div_mul_result_next[31]), .Y(exu_n3938));
AND2X1 exu_U16998(.A(exu_n11528), .B(exu_n10284), .Y(div_mul_result_next[30]));
INVX1 exu_U16999(.A(div_mul_result_next[30]), .Y(exu_n3939));
AND2X1 exu_U17000(.A(exu_n11529), .B(exu_n10285), .Y(div_mul_result_next[2]));
INVX1 exu_U17001(.A(div_mul_result_next[2]), .Y(exu_n3940));
AND2X1 exu_U17002(.A(exu_n11530), .B(exu_n10286), .Y(div_mul_result_next[29]));
INVX1 exu_U17003(.A(div_mul_result_next[29]), .Y(exu_n3941));
AND2X1 exu_U17004(.A(exu_n11531), .B(exu_n10287), .Y(div_mul_result_next[28]));
INVX1 exu_U17005(.A(div_mul_result_next[28]), .Y(exu_n3942));
AND2X1 exu_U17006(.A(exu_n11532), .B(exu_n10288), .Y(div_mul_result_next[27]));
INVX1 exu_U17007(.A(div_mul_result_next[27]), .Y(exu_n3943));
AND2X1 exu_U17008(.A(exu_n11533), .B(exu_n10289), .Y(div_mul_result_next[26]));
INVX1 exu_U17009(.A(div_mul_result_next[26]), .Y(exu_n3944));
AND2X1 exu_U17010(.A(exu_n11534), .B(exu_n10290), .Y(div_mul_result_next[25]));
INVX1 exu_U17011(.A(div_mul_result_next[25]), .Y(exu_n3945));
AND2X1 exu_U17012(.A(exu_n11535), .B(exu_n10291), .Y(div_mul_result_next[24]));
INVX1 exu_U17013(.A(div_mul_result_next[24]), .Y(exu_n3946));
AND2X1 exu_U17014(.A(exu_n11536), .B(exu_n10292), .Y(div_mul_result_next[23]));
INVX1 exu_U17015(.A(div_mul_result_next[23]), .Y(exu_n3947));
AND2X1 exu_U17016(.A(exu_n11537), .B(exu_n10293), .Y(div_mul_result_next[22]));
INVX1 exu_U17017(.A(div_mul_result_next[22]), .Y(exu_n3948));
AND2X1 exu_U17018(.A(exu_n11538), .B(exu_n10294), .Y(div_mul_result_next[21]));
INVX1 exu_U17019(.A(div_mul_result_next[21]), .Y(exu_n3949));
AND2X1 exu_U17020(.A(exu_n11539), .B(exu_n10295), .Y(div_mul_result_next[20]));
INVX1 exu_U17021(.A(div_mul_result_next[20]), .Y(exu_n3950));
AND2X1 exu_U17022(.A(exu_n11540), .B(exu_n10296), .Y(div_mul_result_next[1]));
INVX1 exu_U17023(.A(div_mul_result_next[1]), .Y(exu_n3951));
AND2X1 exu_U17024(.A(exu_n11541), .B(exu_n10297), .Y(div_mul_result_next[19]));
INVX1 exu_U17025(.A(div_mul_result_next[19]), .Y(exu_n3952));
AND2X1 exu_U17026(.A(exu_n11542), .B(exu_n10298), .Y(div_mul_result_next[18]));
INVX1 exu_U17027(.A(div_mul_result_next[18]), .Y(exu_n3953));
AND2X1 exu_U17028(.A(exu_n11543), .B(exu_n10299), .Y(div_mul_result_next[17]));
INVX1 exu_U17029(.A(div_mul_result_next[17]), .Y(exu_n3954));
AND2X1 exu_U17030(.A(exu_n11544), .B(exu_n10300), .Y(div_mul_result_next[16]));
INVX1 exu_U17031(.A(div_mul_result_next[16]), .Y(exu_n3955));
AND2X1 exu_U17032(.A(exu_n11545), .B(exu_n10301), .Y(div_mul_result_next[15]));
INVX1 exu_U17033(.A(div_mul_result_next[15]), .Y(exu_n3956));
AND2X1 exu_U17034(.A(exu_n11546), .B(exu_n10302), .Y(div_mul_result_next[14]));
INVX1 exu_U17035(.A(div_mul_result_next[14]), .Y(exu_n3957));
AND2X1 exu_U17036(.A(exu_n11547), .B(exu_n10303), .Y(div_mul_result_next[13]));
INVX1 exu_U17037(.A(div_mul_result_next[13]), .Y(exu_n3958));
AND2X1 exu_U17038(.A(exu_n11548), .B(exu_n10304), .Y(div_mul_result_next[12]));
INVX1 exu_U17039(.A(div_mul_result_next[12]), .Y(exu_n3959));
AND2X1 exu_U17040(.A(exu_n11549), .B(exu_n10305), .Y(div_mul_result_next[11]));
INVX1 exu_U17041(.A(div_mul_result_next[11]), .Y(exu_n3960));
AND2X1 exu_U17042(.A(exu_n11550), .B(exu_n10306), .Y(div_mul_result_next[10]));
INVX1 exu_U17043(.A(div_mul_result_next[10]), .Y(exu_n3961));
AND2X1 exu_U17044(.A(exu_n11551), .B(exu_n10307), .Y(div_mul_result_next[0]));
INVX1 exu_U17045(.A(div_mul_result_next[0]), .Y(exu_n3962));
AND2X1 exu_U17046(.A(ecl_writeback_n129), .B(ecl_writeback_restore_tid[1]), .Y(exu_n31459));
INVX1 exu_U17047(.A(exu_n31459), .Y(exu_n3963));
AND2X1 exu_U17048(.A(ecl_writeback_ecl_sel_div_g), .B(ecl_mdqctl_wb_divthr_g[1]), .Y(exu_n31461));
INVX1 exu_U17049(.A(exu_n31461), .Y(exu_n3964));
AND2X1 exu_U17050(.A(ecl_writeback_restore_tid[0]), .B(exu_n15988), .Y(exu_n31465));
INVX1 exu_U17051(.A(exu_n31465), .Y(exu_n3965));
AND2X1 exu_U17052(.A(ecl_mdqctl_wb_divthr_g[0]), .B(ecl_writeback_ecl_sel_div_g), .Y(exu_n31467));
INVX1 exu_U17053(.A(exu_n31467), .Y(exu_n3966));
AND2X1 exu_U17054(.A(rml_cwp_swap_next_state[0]), .B(rml_cwp_swap_slot0_state_valid[0]), .Y(exu_n31470));
INVX1 exu_U17055(.A(exu_n31470), .Y(exu_n3967));
AND2X1 exu_U17056(.A(exu_n11611), .B(rml_cwp_swap_slot1_state_valid[0]), .Y(exu_n31475));
INVX1 exu_U17057(.A(exu_n31475), .Y(exu_n3968));
AND2X1 exu_U17058(.A(exu_n11610), .B(rml_cwp_swap_slot2_state_valid[0]), .Y(exu_n31480));
INVX1 exu_U17059(.A(exu_n31480), .Y(exu_n3969));
AND2X1 exu_U17060(.A(exu_n11609), .B(rml_cwp_swap_slot3_state_valid[0]), .Y(exu_n31485));
INVX1 exu_U17061(.A(exu_n31485), .Y(exu_n3970));
OR2X1 exu_U17062(.A(byp_alu_rcc_data_e[18]), .B(byp_alu_rcc_data_e[17]), .Y(exu_n31622));
INVX1 exu_U17063(.A(exu_n31622), .Y(exu_n3971));
OR2X1 exu_U17064(.A(byp_alu_rcc_data_e[21]), .B(byp_alu_rcc_data_e[20]), .Y(exu_n31624));
INVX1 exu_U17065(.A(exu_n31624), .Y(exu_n3972));
OR2X1 exu_U17066(.A(exu_n12040), .B(exu_n14928), .Y(exu_n31618));
INVX1 exu_U17067(.A(exu_n31618), .Y(exu_n3973));
OR2X1 exu_U17068(.A(byp_alu_rcc_data_e[10]), .B(byp_alu_rcc_data_e[0]), .Y(exu_n31628));
INVX1 exu_U17069(.A(exu_n31628), .Y(exu_n3974));
OR2X1 exu_U17070(.A(byp_alu_rcc_data_e[14]), .B(byp_alu_rcc_data_e[13]), .Y(exu_n31630));
INVX1 exu_U17071(.A(exu_n31630), .Y(exu_n3975));
OR2X1 exu_U17072(.A(byp_alu_rcc_data_e[3]), .B(byp_alu_rcc_data_e[31]), .Y(exu_n31636));
INVX1 exu_U17073(.A(exu_n31636), .Y(exu_n3976));
OR2X1 exu_U17074(.A(byp_alu_rcc_data_e[7]), .B(byp_alu_rcc_data_e[6]), .Y(exu_n31638));
INVX1 exu_U17075(.A(exu_n31638), .Y(exu_n3977));
OR2X1 exu_U17076(.A(exu_n12042), .B(exu_n14930), .Y(exu_n31632));
INVX1 exu_U17077(.A(exu_n31632), .Y(exu_n3978));
OR2X1 exu_U17078(.A(byp_alu_rcc_data_e[25]), .B(byp_alu_rcc_data_e[24]), .Y(exu_n31642));
INVX1 exu_U17079(.A(exu_n31642), .Y(exu_n3979));
OR2X1 exu_U17080(.A(byp_alu_rcc_data_e[29]), .B(byp_alu_rcc_data_e[28]), .Y(exu_n31644));
INVX1 exu_U17081(.A(exu_n31644), .Y(exu_n3980));
OR2X1 exu_U17082(.A(byp_alu_rcc_data_e[50]), .B(byp_alu_rcc_data_e[49]), .Y(exu_n31652));
INVX1 exu_U17083(.A(exu_n31652), .Y(exu_n3981));
OR2X1 exu_U17084(.A(byp_alu_rcc_data_e[53]), .B(byp_alu_rcc_data_e[52]), .Y(exu_n31654));
INVX1 exu_U17085(.A(exu_n31654), .Y(exu_n3982));
OR2X1 exu_U17086(.A(exu_n12044), .B(exu_n14932), .Y(exu_n31648));
INVX1 exu_U17087(.A(exu_n31648), .Y(exu_n3983));
OR2X1 exu_U17088(.A(byp_alu_rcc_data_e[42]), .B(byp_alu_rcc_data_e[32]), .Y(exu_n31658));
INVX1 exu_U17089(.A(exu_n31658), .Y(exu_n3984));
OR2X1 exu_U17090(.A(byp_alu_rcc_data_e[46]), .B(byp_alu_rcc_data_e[45]), .Y(exu_n31660));
INVX1 exu_U17091(.A(exu_n31660), .Y(exu_n3985));
OR2X1 exu_U17092(.A(byp_alu_rcc_data_e[35]), .B(exu_ifu_regn_e), .Y(exu_n31666));
INVX1 exu_U17093(.A(exu_n31666), .Y(exu_n3986));
OR2X1 exu_U17094(.A(byp_alu_rcc_data_e[39]), .B(byp_alu_rcc_data_e[38]), .Y(exu_n31668));
INVX1 exu_U17095(.A(exu_n31668), .Y(exu_n3987));
OR2X1 exu_U17096(.A(exu_n12046), .B(exu_n14934), .Y(exu_n31662));
INVX1 exu_U17097(.A(exu_n31662), .Y(exu_n3988));
OR2X1 exu_U17098(.A(byp_alu_rcc_data_e[57]), .B(byp_alu_rcc_data_e[56]), .Y(exu_n31672));
INVX1 exu_U17099(.A(exu_n31672), .Y(exu_n3989));
OR2X1 exu_U17100(.A(byp_alu_rcc_data_e[61]), .B(byp_alu_rcc_data_e[60]), .Y(exu_n31674));
INVX1 exu_U17101(.A(exu_n31674), .Y(exu_n3990));
OR2X1 exu_U17102(.A(div_u32eql_inxor[18]), .B(div_u32eql_inxor[17]), .Y(exu_n31682));
INVX1 exu_U17103(.A(exu_n31682), .Y(exu_n3991));
OR2X1 exu_U17104(.A(div_u32eql_inxor[21]), .B(div_u32eql_inxor[20]), .Y(exu_n31684));
INVX1 exu_U17105(.A(exu_n31684), .Y(exu_n3992));
OR2X1 exu_U17106(.A(exu_n12048), .B(exu_n14936), .Y(exu_n31678));
INVX1 exu_U17107(.A(exu_n31678), .Y(exu_n3993));
OR2X1 exu_U17108(.A(div_u32eql_inxor[14]), .B(div_u32eql_inxor[13]), .Y(exu_n31689));
INVX1 exu_U17109(.A(exu_n31689), .Y(exu_n3994));
OR2X1 exu_U17110(.A(div_u32eql_inxor[3]), .B(div_u32eql_inxor[31]), .Y(exu_n31695));
INVX1 exu_U17111(.A(exu_n31695), .Y(exu_n3995));
OR2X1 exu_U17112(.A(div_u32eql_inxor[7]), .B(div_u32eql_inxor[6]), .Y(exu_n31697));
INVX1 exu_U17113(.A(exu_n31697), .Y(exu_n3996));
OR2X1 exu_U17114(.A(exu_n12050), .B(exu_n14938), .Y(exu_n31691));
INVX1 exu_U17115(.A(exu_n31691), .Y(exu_n3997));
OR2X1 exu_U17116(.A(div_u32eql_inxor[25]), .B(div_u32eql_inxor[24]), .Y(exu_n31701));
INVX1 exu_U17117(.A(exu_n31701), .Y(exu_n3998));
OR2X1 exu_U17118(.A(div_u32eql_inxor[29]), .B(div_u32eql_inxor[28]), .Y(exu_n31703));
INVX1 exu_U17119(.A(exu_n31703), .Y(exu_n3999));
AND2X1 exu_U17120(.A(rml_cwp_swap_sel[3]), .B(rml_cwp_swap_slot3_data[9]), .Y(rml_cwp_cwp_output_mux_n3));
INVX1 exu_U17121(.A(rml_cwp_cwp_output_mux_n3), .Y(exu_n4000));
AND2X1 exu_U17122(.A(rml_cwp_swap_sel[1]), .B(rml_cwp_swap_slot1_data[9]), .Y(rml_cwp_cwp_output_mux_n5));
INVX1 exu_U17123(.A(rml_cwp_cwp_output_mux_n5), .Y(exu_n4001));
AND2X1 exu_U17124(.A(rml_cwp_swap_slot3_data[8]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n9));
INVX1 exu_U17125(.A(rml_cwp_cwp_output_mux_n9), .Y(exu_n4002));
AND2X1 exu_U17126(.A(rml_cwp_swap_slot1_data[8]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n11));
INVX1 exu_U17127(.A(rml_cwp_cwp_output_mux_n11), .Y(exu_n4003));
AND2X1 exu_U17128(.A(rml_cwp_swap_slot3_data[7]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n15));
INVX1 exu_U17129(.A(rml_cwp_cwp_output_mux_n15), .Y(exu_n4004));
AND2X1 exu_U17130(.A(rml_cwp_swap_slot1_data[7]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n17));
INVX1 exu_U17131(.A(rml_cwp_cwp_output_mux_n17), .Y(exu_n4005));
AND2X1 exu_U17132(.A(rml_cwp_swap_slot3_data[6]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n21));
INVX1 exu_U17133(.A(rml_cwp_cwp_output_mux_n21), .Y(exu_n4006));
AND2X1 exu_U17134(.A(rml_cwp_swap_slot1_data[6]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n23));
INVX1 exu_U17135(.A(rml_cwp_cwp_output_mux_n23), .Y(exu_n4007));
AND2X1 exu_U17136(.A(rml_cwp_swap_slot3_data[5]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n27));
INVX1 exu_U17137(.A(rml_cwp_cwp_output_mux_n27), .Y(exu_n4008));
AND2X1 exu_U17138(.A(rml_cwp_swap_slot1_data[5]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n29));
INVX1 exu_U17139(.A(rml_cwp_cwp_output_mux_n29), .Y(exu_n4009));
AND2X1 exu_U17140(.A(rml_cwp_swap_slot3_data[4]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n33));
INVX1 exu_U17141(.A(rml_cwp_cwp_output_mux_n33), .Y(exu_n4010));
AND2X1 exu_U17142(.A(rml_cwp_swap_slot1_data[4]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n35));
INVX1 exu_U17143(.A(rml_cwp_cwp_output_mux_n35), .Y(exu_n4011));
AND2X1 exu_U17144(.A(rml_cwp_swap_slot3_data[3]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n39));
INVX1 exu_U17145(.A(rml_cwp_cwp_output_mux_n39), .Y(exu_n4012));
AND2X1 exu_U17146(.A(rml_cwp_swap_slot1_data[3]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n41));
INVX1 exu_U17147(.A(rml_cwp_cwp_output_mux_n41), .Y(exu_n4013));
AND2X1 exu_U17148(.A(rml_cwp_swap_slot3_data[2]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n45));
INVX1 exu_U17149(.A(rml_cwp_cwp_output_mux_n45), .Y(exu_n4014));
AND2X1 exu_U17150(.A(rml_cwp_swap_slot1_data[2]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n47));
INVX1 exu_U17151(.A(rml_cwp_cwp_output_mux_n47), .Y(exu_n4015));
AND2X1 exu_U17152(.A(rml_cwp_swap_slot3_data[1]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n51));
INVX1 exu_U17153(.A(rml_cwp_cwp_output_mux_n51), .Y(exu_n4016));
AND2X1 exu_U17154(.A(rml_cwp_swap_slot1_data[1]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n53));
INVX1 exu_U17155(.A(rml_cwp_cwp_output_mux_n53), .Y(exu_n4017));
AND2X1 exu_U17156(.A(rml_cwp_swap_slot3_state[1]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n57));
INVX1 exu_U17157(.A(rml_cwp_cwp_output_mux_n57), .Y(exu_n4018));
AND2X1 exu_U17158(.A(rml_cwp_swap_slot1_state[1]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n59));
INVX1 exu_U17159(.A(rml_cwp_cwp_output_mux_n59), .Y(exu_n4019));
AND2X1 exu_U17160(.A(rml_cwp_swap_slot3_state_valid[0]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n63));
INVX1 exu_U17161(.A(rml_cwp_cwp_output_mux_n63), .Y(exu_n4020));
AND2X1 exu_U17162(.A(rml_cwp_swap_slot1_state_valid[0]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n65));
INVX1 exu_U17163(.A(rml_cwp_cwp_output_mux_n65), .Y(exu_n4021));
AND2X1 exu_U17164(.A(rml_cwp_swap_slot3_data[12]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n69));
INVX1 exu_U17165(.A(rml_cwp_cwp_output_mux_n69), .Y(exu_n4022));
AND2X1 exu_U17166(.A(rml_cwp_swap_slot1_data[12]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n71));
INVX1 exu_U17167(.A(rml_cwp_cwp_output_mux_n71), .Y(exu_n4023));
AND2X1 exu_U17168(.A(rml_cwp_swap_slot3_data[11]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n75));
INVX1 exu_U17169(.A(rml_cwp_cwp_output_mux_n75), .Y(exu_n4024));
AND2X1 exu_U17170(.A(rml_cwp_swap_slot1_data[11]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n77));
INVX1 exu_U17171(.A(rml_cwp_cwp_output_mux_n77), .Y(exu_n4025));
AND2X1 exu_U17172(.A(rml_cwp_swap_slot3_data[10]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n81));
INVX1 exu_U17173(.A(rml_cwp_cwp_output_mux_n81), .Y(exu_n4026));
AND2X1 exu_U17174(.A(rml_cwp_swap_slot1_data[10]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n83));
INVX1 exu_U17175(.A(rml_cwp_cwp_output_mux_n83), .Y(exu_n4027));
AND2X1 exu_U17176(.A(rml_cwp_swap_slot3_data[0]), .B(rml_cwp_swap_sel[3]), .Y(rml_cwp_cwp_output_mux_n87));
INVX1 exu_U17177(.A(rml_cwp_cwp_output_mux_n87), .Y(exu_n4028));
AND2X1 exu_U17178(.A(rml_cwp_swap_slot1_data[0]), .B(rml_cwp_swap_sel[1]), .Y(rml_cwp_cwp_output_mux_n89));
INVX1 exu_U17179(.A(rml_cwp_cwp_output_mux_n89), .Y(exu_n4029));
AND2X1 exu_U17180(.A(exu_n11552), .B(exu_n10308), .Y(rml_cwp_cwp_output_queue_next_pv[3]));
INVX1 exu_U17181(.A(rml_cwp_cwp_output_queue_next_pv[3]), .Y(exu_n4030));
AND2X1 exu_U17182(.A(exu_n11553), .B(exu_n10309), .Y(rml_cwp_cwp_output_queue_next_pv[2]));
INVX1 exu_U17183(.A(rml_cwp_cwp_output_queue_next_pv[2]), .Y(exu_n4031));
AND2X1 exu_U17184(.A(exu_n11554), .B(exu_n10310), .Y(rml_cwp_cwp_output_queue_next_pv[1]));
INVX1 exu_U17185(.A(rml_cwp_cwp_output_queue_next_pv[1]), .Y(exu_n4032));
AND2X1 exu_U17186(.A(exu_n11555), .B(exu_n10311), .Y(rml_cwp_cwp_output_queue_next_pv[0]));
INVX1 exu_U17187(.A(rml_cwp_cwp_output_queue_next_pv[0]), .Y(exu_n4033));
AND2X1 exu_U17188(.A(rml_cwp_cwp_output_queue_pv[3]), .B(rml_cwp_swap_req_vec[0]), .Y(rml_cwp_cwp_output_queue_n33));
INVX1 exu_U17189(.A(rml_cwp_cwp_output_queue_n33), .Y(exu_n4034));
AND2X1 exu_U17190(.A(exu_n11559), .B(exu_n10317), .Y(rml_cwp_next_slot0_data[9]));
INVX1 exu_U17191(.A(rml_cwp_next_slot0_data[9]), .Y(exu_n4035));
AND2X1 exu_U17192(.A(exu_n11560), .B(exu_n10318), .Y(rml_cwp_next_slot0_data[8]));
INVX1 exu_U17193(.A(rml_cwp_next_slot0_data[8]), .Y(exu_n4036));
AND2X1 exu_U17194(.A(exu_n16393), .B(exu_n10319), .Y(rml_cwp_next_slot0_data[7]));
INVX1 exu_U17195(.A(rml_cwp_next_slot0_data[7]), .Y(exu_n4037));
AND2X1 exu_U17196(.A(exu_n11561), .B(exu_n10320), .Y(rml_cwp_next_slot0_data[6]));
INVX1 exu_U17197(.A(rml_cwp_next_slot0_data[6]), .Y(exu_n4038));
AND2X1 exu_U17198(.A(rml_cwp_slot0_data_mux_n17), .B(exu_n10321), .Y(rml_cwp_next_slot0_data[5]));
INVX1 exu_U17199(.A(rml_cwp_next_slot0_data[5]), .Y(exu_n4039));
AND2X1 exu_U17200(.A(rml_cwp_tlu_exu_cwp_w[2]), .B(rml_cwp_swap_sel_tlu[0]), .Y(rml_cwp_slot0_data_mux_n19));
INVX1 exu_U17201(.A(rml_cwp_slot0_data_mux_n19), .Y(exu_n4040));
AND2X1 exu_U17202(.A(rml_cwp_slot0_data_mux_n21), .B(exu_n10322), .Y(rml_cwp_next_slot0_data[4]));
INVX1 exu_U17203(.A(rml_cwp_next_slot0_data[4]), .Y(exu_n4041));
AND2X1 exu_U17204(.A(rml_cwp_tlu_exu_cwp_w[1]), .B(rml_cwp_swap_sel_tlu[0]), .Y(rml_cwp_slot0_data_mux_n23));
INVX1 exu_U17205(.A(rml_cwp_slot0_data_mux_n23), .Y(exu_n4042));
AND2X1 exu_U17206(.A(rml_cwp_slot0_data_mux_n25), .B(exu_n10323), .Y(rml_cwp_next_slot0_data[3]));
INVX1 exu_U17207(.A(rml_cwp_next_slot0_data[3]), .Y(exu_n4043));
AND2X1 exu_U17208(.A(rml_cwp_tlu_exu_cwp_w[0]), .B(rml_cwp_swap_sel_tlu[0]), .Y(rml_cwp_slot0_data_mux_n27));
INVX1 exu_U17209(.A(rml_cwp_slot0_data_mux_n27), .Y(exu_n4044));
AND2X1 exu_U17210(.A(rml_cwp_slot0_data_mux_n29), .B(exu_n10324), .Y(rml_cwp_next_slot0_data[2]));
INVX1 exu_U17211(.A(rml_cwp_next_slot0_data[2]), .Y(exu_n4045));
AND2X1 exu_U17212(.A(rml_cwp_old_cwp_w[2]), .B(rml_cwp_swap_sel_tlu[0]), .Y(rml_cwp_slot0_data_mux_n31));
INVX1 exu_U17213(.A(rml_cwp_slot0_data_mux_n31), .Y(exu_n4046));
AND2X1 exu_U17214(.A(rml_cwp_slot0_data_mux_n33), .B(exu_n10325), .Y(rml_cwp_next_slot0_data[1]));
INVX1 exu_U17215(.A(rml_cwp_next_slot0_data[1]), .Y(exu_n4047));
AND2X1 exu_U17216(.A(rml_cwp_old_cwp_w[1]), .B(rml_cwp_swap_sel_tlu[0]), .Y(rml_cwp_slot0_data_mux_n35));
INVX1 exu_U17217(.A(rml_cwp_slot0_data_mux_n35), .Y(exu_n4048));
AND2X1 exu_U17218(.A(exu_n11562), .B(exu_n10326), .Y(rml_cwp_next_slot0_data[12]));
INVX1 exu_U17219(.A(rml_cwp_next_slot0_data[12]), .Y(exu_n4049));
AND2X1 exu_U17220(.A(exu_n11563), .B(exu_n10327), .Y(rml_cwp_next_slot0_data[11]));
INVX1 exu_U17221(.A(rml_cwp_next_slot0_data[11]), .Y(exu_n4050));
AND2X1 exu_U17222(.A(exu_n11564), .B(exu_n10328), .Y(rml_cwp_next_slot0_data[10]));
INVX1 exu_U17223(.A(rml_cwp_next_slot0_data[10]), .Y(exu_n4051));
AND2X1 exu_U17224(.A(rml_cwp_slot0_data_mux_n49), .B(exu_n10329), .Y(rml_cwp_next_slot0_data[0]));
INVX1 exu_U17225(.A(rml_cwp_next_slot0_data[0]), .Y(exu_n4052));
AND2X1 exu_U17226(.A(rml_cwp_old_cwp_w[0]), .B(rml_cwp_swap_sel_tlu[0]), .Y(rml_cwp_slot0_data_mux_n51));
INVX1 exu_U17227(.A(rml_cwp_slot0_data_mux_n51), .Y(exu_n4053));
AND2X1 exu_U17228(.A(exu_n11565), .B(exu_n10330), .Y(ecl_mdqctl_div_data_next[0]));
INVX1 exu_U17229(.A(ecl_mdqctl_div_data_next[0]), .Y(exu_n4054));
AND2X1 exu_U17230(.A(exu_n11566), .B(exu_n10331), .Y(ecl_mdqctl_div_data_next[1]));
INVX1 exu_U17231(.A(ecl_mdqctl_div_data_next[1]), .Y(exu_n4055));
AND2X1 exu_U17232(.A(exu_n11567), .B(exu_n10332), .Y(ecl_mdqctl_div_data_next[2]));
INVX1 exu_U17233(.A(ecl_mdqctl_div_data_next[2]), .Y(exu_n4056));
AND2X1 exu_U17234(.A(exu_n11568), .B(exu_n10333), .Y(ecl_mdqctl_div_data_next[3]));
INVX1 exu_U17235(.A(ecl_mdqctl_div_data_next[3]), .Y(exu_n4057));
AND2X1 exu_U17236(.A(exu_n11569), .B(exu_n10334), .Y(ecl_mdqctl_div_data_next[4]));
INVX1 exu_U17237(.A(ecl_mdqctl_div_data_next[4]), .Y(exu_n4058));
AND2X1 exu_U17238(.A(exu_n11570), .B(exu_n10335), .Y(ecl_mdqctl_div_data_next[5]));
INVX1 exu_U17239(.A(ecl_mdqctl_div_data_next[5]), .Y(exu_n4059));
AND2X1 exu_U17240(.A(exu_n11571), .B(exu_n10336), .Y(ecl_mdqctl_div_data_next[6]));
INVX1 exu_U17241(.A(ecl_mdqctl_div_data_next[6]), .Y(exu_n4060));
AND2X1 exu_U17242(.A(exu_n11572), .B(exu_n10337), .Y(ecl_mdqctl_div_data_next[7]));
INVX1 exu_U17243(.A(ecl_mdqctl_div_data_next[7]), .Y(exu_n4061));
AND2X1 exu_U17244(.A(exu_n11573), .B(exu_n10338), .Y(ecl_mdqctl_div_data_next[8]));
INVX1 exu_U17245(.A(ecl_mdqctl_div_data_next[8]), .Y(exu_n4062));
AND2X1 exu_U17246(.A(exu_n11574), .B(exu_n10339), .Y(ecl_mdqctl_div_data_next[9]));
INVX1 exu_U17247(.A(ecl_mdqctl_div_data_next[9]), .Y(exu_n4063));
AND2X1 exu_U17248(.A(exu_n11575), .B(exu_n10340), .Y(ecl_mdqctl_div_data_next[10]));
INVX1 exu_U17249(.A(ecl_mdqctl_div_data_next[10]), .Y(exu_n4064));
AND2X1 exu_U17250(.A(exu_n16387), .B(exu_n10341), .Y(ecl_mdqctl_div_data_next[11]));
INVX1 exu_U17251(.A(ecl_mdqctl_div_data_next[11]), .Y(exu_n4065));
AND2X1 exu_U17252(.A(exu_n11577), .B(exu_n10343), .Y(ecl_divcntl_q_next));
INVX1 exu_U17253(.A(ecl_divcntl_q_next), .Y(exu_n4066));
OR2X1 exu_U17254(.A(exu_n16438), .B(ecl_divcntl_cnt6_n9), .Y(ecl_divcntl_cnt6_next_cntr[5]));
INVX1 exu_U17255(.A(ecl_divcntl_cnt6_next_cntr[5]), .Y(exu_n4067));
AND2X1 exu_U17256(.A(exu_n11578), .B(ecl_divcntl_cnt6_n15), .Y(ecl_divcntl_cnt6_next_cntr[4]));
INVX1 exu_U17257(.A(ecl_divcntl_cnt6_next_cntr[4]), .Y(exu_n4068));
AND2X1 exu_U17258(.A(exu_n11579), .B(ecl_divcntl_cnt6_n22), .Y(ecl_divcntl_cnt6_next_cntr[3]));
INVX1 exu_U17259(.A(ecl_divcntl_cnt6_next_cntr[3]), .Y(exu_n4069));
AND2X1 exu_U17260(.A(exu_n11580), .B(exu_n10345), .Y(ecl_divcntl_cnt6_next_cntr[2]));
INVX1 exu_U17261(.A(ecl_divcntl_cnt6_next_cntr[2]), .Y(exu_n4070));
OR2X1 exu_U17262(.A(exu_n16438), .B(exu_n16621), .Y(ecl_divcntl_cnt6_n29));
INVX1 exu_U17263(.A(ecl_divcntl_cnt6_n29), .Y(exu_n4071));
OR2X1 exu_U17264(.A(ecl_byplog_rs1_w_comp7_n9), .B(exu_n14941), .Y(ecl_byplog_rs1_w_comp7_n1));
INVX1 exu_U17265(.A(ecl_byplog_rs1_w_comp7_n1), .Y(exu_n4072));
AND2X1 exu_U17266(.A(ecl_ecc_log_rs2_m), .B(ecl_eccctl_rs2_ce_m), .Y(ecl_eccctl_ecc_synd7_mux_n3));
INVX1 exu_U17267(.A(ecl_eccctl_ecc_synd7_mux_n3), .Y(exu_n4073));
AND2X1 exu_U17268(.A(ecl_ecc_sel_rs2_m_l), .B(ecl_ifu_exu_rs2_m[4]), .Y(ecl_eccctl_ecc_rd_mux_n3));
INVX1 exu_U17269(.A(ecl_eccctl_ecc_rd_mux_n3), .Y(exu_n4074));
AND2X1 exu_U17270(.A(ecl_ifu_exu_rs2_m[3]), .B(ecl_ecc_sel_rs2_m_l), .Y(ecl_eccctl_ecc_rd_mux_n7));
INVX1 exu_U17271(.A(ecl_eccctl_ecc_rd_mux_n7), .Y(exu_n4075));
AND2X1 exu_U17272(.A(ecl_ifu_exu_rs2_m[2]), .B(exu_n15974), .Y(ecl_eccctl_ecc_rd_mux_n11));
INVX1 exu_U17273(.A(ecl_eccctl_ecc_rd_mux_n11), .Y(exu_n4076));
AND2X1 exu_U17274(.A(ecl_ifu_exu_rs2_m[1]), .B(ecl_ecc_sel_rs2_m_l), .Y(ecl_eccctl_ecc_rd_mux_n15));
INVX1 exu_U17275(.A(ecl_eccctl_ecc_rd_mux_n15), .Y(exu_n4077));
AND2X1 exu_U17276(.A(ecl_ifu_exu_rs2_m[0]), .B(ecl_ecc_sel_rs2_m_l), .Y(ecl_eccctl_ecc_rd_mux_n19));
INVX1 exu_U17277(.A(ecl_eccctl_ecc_rd_mux_n19), .Y(exu_n4078));
AND2X1 exu_U17278(.A(ecl_writeback_n70), .B(rml_ecl_otherwin_d[2]), .Y(ecl_writeback_rdpr_mux1_n3));
INVX1 exu_U17279(.A(ecl_writeback_rdpr_mux1_n3), .Y(exu_n4079));
AND2X1 exu_U17280(.A(exu_n15432), .B(rml_ecl_cleanwin_d[2]), .Y(ecl_writeback_rdpr_mux1_n5));
INVX1 exu_U17281(.A(ecl_writeback_rdpr_mux1_n5), .Y(exu_n4080));
AND2X1 exu_U17282(.A(rml_ecl_otherwin_d[1]), .B(ecl_writeback_n70), .Y(ecl_writeback_rdpr_mux1_n9));
INVX1 exu_U17283(.A(ecl_writeback_rdpr_mux1_n9), .Y(exu_n4081));
AND2X1 exu_U17284(.A(rml_ecl_cleanwin_d[1]), .B(exu_n15432), .Y(ecl_writeback_rdpr_mux1_n11));
INVX1 exu_U17285(.A(ecl_writeback_rdpr_mux1_n11), .Y(exu_n4082));
AND2X1 exu_U17286(.A(rml_ecl_otherwin_d[0]), .B(ecl_writeback_n70), .Y(ecl_writeback_rdpr_mux1_n15));
INVX1 exu_U17287(.A(ecl_writeback_rdpr_mux1_n15), .Y(exu_n4083));
AND2X1 exu_U17288(.A(rml_ecl_cleanwin_d[0]), .B(exu_n15432), .Y(ecl_writeback_rdpr_mux1_n17));
INVX1 exu_U17289(.A(ecl_writeback_rdpr_mux1_n17), .Y(exu_n4084));
AND2X1 exu_U17290(.A(exu_n11592), .B(exu_n10356), .Y(ecl_writeback_setcc_g));
INVX1 exu_U17291(.A(ecl_writeback_setcc_g), .Y(exu_n4085));
AND2X1 exu_U17292(.A(exu_n15988), .B(ecl_writeback_restore_rd[4]), .Y(ecl_writeback_rd_g_mux_n3));
INVX1 exu_U17293(.A(ecl_writeback_rd_g_mux_n3), .Y(exu_n4086));
AND2X1 exu_U17294(.A(ecl_writeback_ecl_sel_div_g), .B(ecl_mdqctl_wb_divrd_g[4]), .Y(ecl_writeback_rd_g_mux_n5));
INVX1 exu_U17295(.A(ecl_writeback_rd_g_mux_n5), .Y(exu_n4087));
AND2X1 exu_U17296(.A(ecl_writeback_restore_rd[3]), .B(ecl_writeback_n129), .Y(ecl_writeback_rd_g_mux_n9));
INVX1 exu_U17297(.A(ecl_writeback_rd_g_mux_n9), .Y(exu_n4088));
AND2X1 exu_U17298(.A(ecl_mdqctl_wb_divrd_g[3]), .B(ecl_writeback_ecl_sel_div_g), .Y(ecl_writeback_rd_g_mux_n11));
INVX1 exu_U17299(.A(ecl_writeback_rd_g_mux_n11), .Y(exu_n4089));
AND2X1 exu_U17300(.A(ecl_writeback_restore_rd[2]), .B(exu_n15988), .Y(ecl_writeback_rd_g_mux_n15));
INVX1 exu_U17301(.A(ecl_writeback_rd_g_mux_n15), .Y(exu_n4090));
AND2X1 exu_U17302(.A(ecl_mdqctl_wb_divrd_g[2]), .B(ecl_writeback_ecl_sel_div_g), .Y(ecl_writeback_rd_g_mux_n17));
INVX1 exu_U17303(.A(ecl_writeback_rd_g_mux_n17), .Y(exu_n4091));
AND2X1 exu_U17304(.A(ecl_writeback_restore_rd[1]), .B(ecl_writeback_n129), .Y(ecl_writeback_rd_g_mux_n21));
INVX1 exu_U17305(.A(ecl_writeback_rd_g_mux_n21), .Y(exu_n4092));
AND2X1 exu_U17306(.A(ecl_mdqctl_wb_divrd_g[1]), .B(ecl_writeback_ecl_sel_div_g), .Y(ecl_writeback_rd_g_mux_n23));
INVX1 exu_U17307(.A(ecl_writeback_rd_g_mux_n23), .Y(exu_n4093));
AND2X1 exu_U17308(.A(ecl_writeback_restore_rd[0]), .B(ecl_writeback_n129), .Y(ecl_writeback_rd_g_mux_n27));
INVX1 exu_U17309(.A(ecl_writeback_rd_g_mux_n27), .Y(exu_n4094));
AND2X1 exu_U17310(.A(ecl_mdqctl_wb_divrd_g[0]), .B(ecl_writeback_ecl_sel_div_g), .Y(ecl_writeback_rd_g_mux_n29));
INVX1 exu_U17311(.A(ecl_writeback_rd_g_mux_n29), .Y(exu_n4095));
AND2X1 exu_U17312(.A(ecl_thr_d[3]), .B(exu_tlu_ccr3_w[7]), .Y(ecl_ccr_mux_ccr_out_n3));
INVX1 exu_U17313(.A(ecl_ccr_mux_ccr_out_n3), .Y(exu_n4096));
AND2X1 exu_U17314(.A(exu_n15934), .B(exu_tlu_ccr1_w[7]), .Y(ecl_ccr_mux_ccr_out_n5));
INVX1 exu_U17315(.A(ecl_ccr_mux_ccr_out_n5), .Y(exu_n4097));
AND2X1 exu_U17316(.A(exu_tlu_ccr3_w[6]), .B(ecl_thr_d[3]), .Y(ecl_ccr_mux_ccr_out_n9));
INVX1 exu_U17317(.A(ecl_ccr_mux_ccr_out_n9), .Y(exu_n4098));
AND2X1 exu_U17318(.A(exu_tlu_ccr1_w[6]), .B(exu_n15934), .Y(ecl_ccr_mux_ccr_out_n11));
INVX1 exu_U17319(.A(ecl_ccr_mux_ccr_out_n11), .Y(exu_n4099));
AND2X1 exu_U17320(.A(exu_tlu_ccr3_w[5]), .B(ecl_thr_d[3]), .Y(ecl_ccr_mux_ccr_out_n15));
INVX1 exu_U17321(.A(ecl_ccr_mux_ccr_out_n15), .Y(exu_n4100));
AND2X1 exu_U17322(.A(exu_tlu_ccr1_w[5]), .B(exu_n15934), .Y(ecl_ccr_mux_ccr_out_n17));
INVX1 exu_U17323(.A(ecl_ccr_mux_ccr_out_n17), .Y(exu_n4101));
AND2X1 exu_U17324(.A(exu_tlu_ccr3_w[4]), .B(ecl_thr_d[3]), .Y(ecl_ccr_mux_ccr_out_n21));
INVX1 exu_U17325(.A(ecl_ccr_mux_ccr_out_n21), .Y(exu_n4102));
AND2X1 exu_U17326(.A(exu_tlu_ccr1_w[4]), .B(exu_n15934), .Y(ecl_ccr_mux_ccr_out_n23));
INVX1 exu_U17327(.A(ecl_ccr_mux_ccr_out_n23), .Y(exu_n4103));
AND2X1 exu_U17328(.A(exu_tlu_ccr3_w[3]), .B(ecl_thr_d[3]), .Y(ecl_ccr_mux_ccr_out_n27));
INVX1 exu_U17329(.A(ecl_ccr_mux_ccr_out_n27), .Y(exu_n4104));
AND2X1 exu_U17330(.A(exu_tlu_ccr1_w[3]), .B(exu_n15934), .Y(ecl_ccr_mux_ccr_out_n29));
INVX1 exu_U17331(.A(ecl_ccr_mux_ccr_out_n29), .Y(exu_n4105));
AND2X1 exu_U17332(.A(exu_tlu_ccr3_w[2]), .B(ecl_thr_d[3]), .Y(ecl_ccr_mux_ccr_out_n33));
INVX1 exu_U17333(.A(ecl_ccr_mux_ccr_out_n33), .Y(exu_n4106));
AND2X1 exu_U17334(.A(exu_tlu_ccr1_w[2]), .B(exu_n15934), .Y(ecl_ccr_mux_ccr_out_n35));
INVX1 exu_U17335(.A(ecl_ccr_mux_ccr_out_n35), .Y(exu_n4107));
AND2X1 exu_U17336(.A(exu_tlu_ccr3_w[1]), .B(ecl_thr_d[3]), .Y(ecl_ccr_mux_ccr_out_n39));
INVX1 exu_U17337(.A(ecl_ccr_mux_ccr_out_n39), .Y(exu_n4108));
AND2X1 exu_U17338(.A(exu_tlu_ccr1_w[1]), .B(exu_n15934), .Y(ecl_ccr_mux_ccr_out_n41));
INVX1 exu_U17339(.A(ecl_ccr_mux_ccr_out_n41), .Y(exu_n4109));
AND2X1 exu_U17340(.A(exu_tlu_ccr3_w[0]), .B(ecl_thr_d[3]), .Y(ecl_ccr_mux_ccr_out_n45));
INVX1 exu_U17341(.A(ecl_ccr_mux_ccr_out_n45), .Y(exu_n4110));
AND2X1 exu_U17342(.A(exu_tlu_ccr1_w[0]), .B(exu_n15934), .Y(ecl_ccr_mux_ccr_out_n47));
INVX1 exu_U17343(.A(ecl_ccr_mux_ccr_out_n47), .Y(exu_n4111));
AND2X1 exu_U17344(.A(ecl_ccr_mux_ccrin0_n1), .B(exu_n10357), .Y(ecl_ccr_ccrin_thr0[7]));
INVX1 exu_U17345(.A(ecl_ccr_ccrin_thr0[7]), .Y(exu_n4112));
AND2X1 exu_U17346(.A(ecl_ccr_n19), .B(ecl_divcntl_ccr_cc_w2[7]), .Y(ecl_ccr_mux_ccrin0_n3));
INVX1 exu_U17347(.A(ecl_ccr_mux_ccrin0_n3), .Y(exu_n4113));
AND2X1 exu_U17348(.A(ecl_ccr_mux_ccrin0_n5), .B(exu_n10358), .Y(ecl_ccr_ccrin_thr0[6]));
INVX1 exu_U17349(.A(ecl_ccr_ccrin_thr0[6]), .Y(exu_n4114));
AND2X1 exu_U17350(.A(ecl_divcntl_ccr_cc_w2[6]), .B(ecl_ccr_n19), .Y(ecl_ccr_mux_ccrin0_n7));
INVX1 exu_U17351(.A(ecl_ccr_mux_ccrin0_n7), .Y(exu_n4115));
AND2X1 exu_U17352(.A(exu_n11593), .B(exu_n10359), .Y(ecl_ccr_ccrin_thr0[5]));
INVX1 exu_U17353(.A(ecl_ccr_ccrin_thr0[5]), .Y(exu_n4116));
AND2X1 exu_U17354(.A(exu_n11594), .B(exu_n10360), .Y(ecl_ccr_ccrin_thr0[4]));
INVX1 exu_U17355(.A(ecl_ccr_ccrin_thr0[4]), .Y(exu_n4117));
AND2X1 exu_U17356(.A(ecl_ccr_mux_ccrin0_n17), .B(exu_n10361), .Y(ecl_ccr_ccrin_thr0[3]));
INVX1 exu_U17357(.A(ecl_ccr_ccrin_thr0[3]), .Y(exu_n4118));
AND2X1 exu_U17358(.A(exu_n15736), .B(ecl_ccr_n19), .Y(ecl_ccr_mux_ccrin0_n19));
INVX1 exu_U17359(.A(ecl_ccr_mux_ccrin0_n19), .Y(exu_n4119));
AND2X1 exu_U17360(.A(ecl_ccr_mux_ccrin0_n21), .B(exu_n10362), .Y(ecl_ccr_ccrin_thr0[2]));
INVX1 exu_U17361(.A(ecl_ccr_ccrin_thr0[2]), .Y(exu_n4120));
AND2X1 exu_U17362(.A(exu_n15737), .B(ecl_ccr_n19), .Y(ecl_ccr_mux_ccrin0_n23));
INVX1 exu_U17363(.A(ecl_ccr_mux_ccrin0_n23), .Y(exu_n4121));
AND2X1 exu_U17364(.A(ecl_ccr_mux_ccrin0_n25), .B(exu_n10363), .Y(ecl_ccr_ccrin_thr0[1]));
INVX1 exu_U17365(.A(ecl_ccr_ccrin_thr0[1]), .Y(exu_n4122));
AND2X1 exu_U17366(.A(exu_n15738), .B(ecl_ccr_n19), .Y(ecl_ccr_mux_ccrin0_n27));
INVX1 exu_U17367(.A(ecl_ccr_mux_ccrin0_n27), .Y(exu_n4123));
AND2X1 exu_U17368(.A(ecl_ccr_mux_ccrin0_n29), .B(exu_n10364), .Y(ecl_ccr_ccrin_thr0[0]));
INVX1 exu_U17369(.A(ecl_ccr_ccrin_thr0[0]), .Y(exu_n4124));
AND2X1 exu_U17370(.A(ecl_divcntl_ccr_cc_w2[0]), .B(ecl_ccr_n19), .Y(ecl_ccr_mux_ccrin0_n31));
INVX1 exu_U17371(.A(ecl_ccr_mux_ccrin0_n31), .Y(exu_n4125));
AND2X1 exu_U17372(.A(exu_n11595), .B(exu_n10365), .Y(ecl_ccr_ccr_m[0]));
INVX1 exu_U17373(.A(ecl_ccr_ccr_m[0]), .Y(exu_n4126));
AND2X1 exu_U17374(.A(exu_n11596), .B(exu_n10366), .Y(ecl_ccr_ccr_m[1]));
INVX1 exu_U17375(.A(ecl_ccr_ccr_m[1]), .Y(exu_n4127));
AND2X1 exu_U17376(.A(exu_n11597), .B(exu_n10367), .Y(ecl_ccr_ccr_m[2]));
INVX1 exu_U17377(.A(ecl_ccr_ccr_m[2]), .Y(exu_n4128));
AND2X1 exu_U17378(.A(exu_n11598), .B(exu_n10368), .Y(ecl_ccr_ccr_m[3]));
INVX1 exu_U17379(.A(ecl_ccr_ccr_m[3]), .Y(exu_n4129));
AND2X1 exu_U17380(.A(exu_n11599), .B(exu_n10369), .Y(ecl_ccr_ccr_m[4]));
INVX1 exu_U17381(.A(ecl_ccr_ccr_m[4]), .Y(exu_n4130));
AND2X1 exu_U17382(.A(exu_n11600), .B(exu_n10370), .Y(ecl_ccr_ccr_m[5]));
INVX1 exu_U17383(.A(ecl_ccr_ccr_m[5]), .Y(exu_n4131));
AND2X1 exu_U17384(.A(exu_n11601), .B(exu_n10371), .Y(ecl_ccr_ccr_m[6]));
INVX1 exu_U17385(.A(ecl_ccr_ccr_m[6]), .Y(exu_n4132));
AND2X1 exu_U17386(.A(exu_n11602), .B(exu_n10372), .Y(ecl_ccr_ccr_m[7]));
INVX1 exu_U17387(.A(ecl_ccr_ccr_m[7]), .Y(exu_n4133));
AND2X1 exu_U17388(.A(exu_n11603), .B(exu_n10373), .Y(rml_agp_thr0_next[0]));
INVX1 exu_U17389(.A(rml_agp_thr0_next[0]), .Y(exu_n4134));
AND2X1 exu_U17390(.A(exu_n11604), .B(exu_n10374), .Y(rml_agp_thr0_next[1]));
INVX1 exu_U17391(.A(rml_agp_thr0_next[1]), .Y(exu_n4135));
AND2X1 exu_U17392(.A(rml_agp_thr[3]), .B(rml_agp_thr3[1]), .Y(rml_mux_agp_out1_n3));
INVX1 exu_U17393(.A(rml_mux_agp_out1_n3), .Y(exu_n4136));
AND2X1 exu_U17394(.A(exu_n15439), .B(rml_agp_thr1[1]), .Y(rml_mux_agp_out1_n5));
INVX1 exu_U17395(.A(rml_mux_agp_out1_n5), .Y(exu_n4137));
AND2X1 exu_U17396(.A(rml_agp_thr3[0]), .B(rml_agp_thr[3]), .Y(rml_mux_agp_out1_n9));
INVX1 exu_U17397(.A(rml_mux_agp_out1_n9), .Y(exu_n4138));
AND2X1 exu_U17398(.A(rml_agp_thr1[0]), .B(exu_n15439), .Y(rml_mux_agp_out1_n11));
INVX1 exu_U17399(.A(rml_mux_agp_out1_n11), .Y(exu_n4139));
AND2X1 exu_U17400(.A(exu_n11605), .B(exu_n10375), .Y(rml_next_cansave_e[0]));
INVX1 exu_U17401(.A(rml_next_cansave_e[0]), .Y(exu_n4140));
AND2X1 exu_U17402(.A(exu_n11606), .B(exu_n10376), .Y(rml_next_cansave_e[1]));
INVX1 exu_U17403(.A(rml_next_cansave_e[1]), .Y(exu_n4141));
AND2X1 exu_U17404(.A(exu_n11607), .B(exu_n10377), .Y(rml_next_cansave_e[2]));
INVX1 exu_U17405(.A(rml_next_cansave_e[2]), .Y(exu_n4142));
OR2X1 exu_U17406(.A(exu_n15766), .B(exu_n14942), .Y(rml_cwp_swap_done_next_cycle[3]));
INVX1 exu_U17407(.A(rml_cwp_swap_done_next_cycle[3]), .Y(exu_n4143));
OR2X1 exu_U17408(.A(exu_n15766), .B(exu_n14943), .Y(rml_cwp_swap_done_next_cycle[2]));
INVX1 exu_U17409(.A(rml_cwp_swap_done_next_cycle[2]), .Y(exu_n4144));
OR2X1 exu_U17410(.A(exu_n15766), .B(exu_n14944), .Y(rml_cwp_swap_done_next_cycle[1]));
INVX1 exu_U17411(.A(rml_cwp_swap_done_next_cycle[1]), .Y(exu_n4145));
OR2X1 exu_U17412(.A(exu_n15766), .B(exu_n14945), .Y(rml_cwp_swap_done_next_cycle[0]));
INVX1 exu_U17413(.A(rml_cwp_swap_done_next_cycle[0]), .Y(exu_n4146));
OR2X1 exu_U17414(.A(rml_cwp_swap_data[7]), .B(rml_cwp_swap_data[6]), .Y(rml_cwp_n52));
INVX1 exu_U17415(.A(rml_cwp_n52), .Y(exu_n4147));
OR2X1 exu_U17416(.A(exu_n15740), .B(rml_cwp_cwp_fastcmplt_w), .Y(rml_cwp_n90));
INVX1 exu_U17417(.A(rml_cwp_n90), .Y(exu_n4148));
OR2X1 exu_U17418(.A(exu_n15384), .B(rml_cwp_swap_data[7]), .Y(rml_cwp_n95));
INVX1 exu_U17419(.A(rml_cwp_n95), .Y(exu_n4149));
OR2X1 exu_U17420(.A(exu_n12052), .B(exu_n14946), .Y(rml_cwp_cwp_fastcmplt_m));
INVX1 exu_U17421(.A(rml_cwp_cwp_fastcmplt_m), .Y(exu_n4150));
OR2X1 exu_U17422(.A(ifu_exu_flushw_e), .B(exu_n15822), .Y(rml_cwp_n102));
INVX1 exu_U17423(.A(rml_cwp_n102), .Y(exu_n4151));
AND2X1 exu_U17424(.A(exu_n15822), .B(ecl_rml_xor_data_e[2]), .Y(rml_next_cwp_mux_n3));
INVX1 exu_U17425(.A(rml_next_cwp_mux_n3), .Y(exu_n4152));
AND2X1 exu_U17426(.A(ecl_rml_xor_data_e[1]), .B(exu_n15822), .Y(rml_next_cwp_mux_n7));
INVX1 exu_U17427(.A(rml_next_cwp_mux_n7), .Y(exu_n4153));
AND2X1 exu_U17428(.A(ecl_rml_xor_data_e[0]), .B(exu_n15822), .Y(rml_next_cwp_mux_n11));
INVX1 exu_U17429(.A(rml_next_cwp_mux_n11), .Y(exu_n4154));
AND2X1 exu_U17430(.A(rml_rml_ecl_cwp_e[1]), .B(rml_rml_ecl_cwp_e[0]), .Y(rml_cwp_inc_n4));
INVX1 exu_U17431(.A(rml_cwp_inc_n4), .Y(exu_n4155));
OR2X1 exu_U17432(.A(exu_n12053), .B(exu_n14947), .Y(rml_wtype_mux_n3));
INVX1 exu_U17433(.A(rml_wtype_mux_n3), .Y(exu_n4156));
OR2X1 exu_U17434(.A(exu_n12054), .B(exu_n14948), .Y(rml_wtype_mux_n4));
INVX1 exu_U17435(.A(rml_wtype_mux_n4), .Y(exu_n4157));
OR2X1 exu_U17436(.A(exu_n12055), .B(exu_n14949), .Y(rml_wtype_mux_n5));
INVX1 exu_U17437(.A(rml_wtype_mux_n5), .Y(exu_n4158));
AND2X1 exu_U17438(.A(div_d_mux_n1), .B(exu_n10385), .Y(div_dnext[9]));
INVX1 exu_U17439(.A(div_dnext[9]), .Y(exu_n4159));
AND2X1 exu_U17440(.A(ecl_div_sel_adder), .B(div_d[8]), .Y(div_d_mux_n3));
INVX1 exu_U17441(.A(div_d_mux_n3), .Y(exu_n4160));
AND2X1 exu_U17442(.A(div_d_mux_n5), .B(exu_n10777), .Y(div_dnext[99]));
INVX1 exu_U17443(.A(div_dnext[99]), .Y(exu_n4161));
AND2X1 exu_U17444(.A(div_adder_out[35]), .B(ecl_div_sel_adder), .Y(div_d_mux_n7));
INVX1 exu_U17445(.A(div_d_mux_n7), .Y(exu_n4162));
AND2X1 exu_U17446(.A(div_d_mux_n9), .B(exu_n10387), .Y(div_dnext[98]));
INVX1 exu_U17447(.A(div_dnext[98]), .Y(exu_n4163));
AND2X1 exu_U17448(.A(div_adder_out[34]), .B(ecl_div_sel_adder), .Y(div_d_mux_n11));
INVX1 exu_U17449(.A(div_d_mux_n11), .Y(exu_n4164));
AND2X1 exu_U17450(.A(div_d_mux_n13), .B(exu_n10387), .Y(div_dnext[97]));
INVX1 exu_U17451(.A(div_dnext[97]), .Y(exu_n4165));
AND2X1 exu_U17452(.A(div_adder_out[33]), .B(exu_n16250), .Y(div_d_mux_n15));
INVX1 exu_U17453(.A(div_d_mux_n15), .Y(exu_n4166));
AND2X1 exu_U17454(.A(div_d_mux_n17), .B(exu_n10389), .Y(div_dnext[96]));
INVX1 exu_U17455(.A(div_dnext[96]), .Y(exu_n4167));
AND2X1 exu_U17456(.A(div_adder_out[32]), .B(exu_n16250), .Y(div_d_mux_n19));
INVX1 exu_U17457(.A(div_d_mux_n19), .Y(exu_n4168));
AND2X1 exu_U17458(.A(div_d_mux_n21), .B(exu_n10391), .Y(div_dnext[95]));
INVX1 exu_U17459(.A(div_dnext[95]), .Y(exu_n4169));
AND2X1 exu_U17460(.A(div_ecl_adder_out_31), .B(ecl_div_sel_adder), .Y(div_d_mux_n23));
INVX1 exu_U17461(.A(div_d_mux_n23), .Y(exu_n4170));
AND2X1 exu_U17462(.A(div_d_mux_n25), .B(exu_n10392), .Y(div_dnext[94]));
INVX1 exu_U17463(.A(div_dnext[94]), .Y(exu_n4171));
AND2X1 exu_U17464(.A(div_adder_out_30), .B(exu_n16250), .Y(div_d_mux_n27));
INVX1 exu_U17465(.A(div_d_mux_n27), .Y(exu_n4172));
AND2X1 exu_U17466(.A(div_d_mux_n29), .B(exu_n10393), .Y(div_dnext[93]));
INVX1 exu_U17467(.A(div_dnext[93]), .Y(exu_n4173));
AND2X1 exu_U17468(.A(div_adder_out_29), .B(ecl_div_sel_adder), .Y(div_d_mux_n31));
INVX1 exu_U17469(.A(div_d_mux_n31), .Y(exu_n4174));
AND2X1 exu_U17470(.A(div_d_mux_n33), .B(exu_n10394), .Y(div_dnext[92]));
INVX1 exu_U17471(.A(div_dnext[92]), .Y(exu_n4175));
AND2X1 exu_U17472(.A(div_adder_out_28), .B(ecl_div_sel_adder), .Y(div_d_mux_n35));
INVX1 exu_U17473(.A(div_d_mux_n35), .Y(exu_n4176));
AND2X1 exu_U17474(.A(div_d_mux_n37), .B(exu_n10395), .Y(div_dnext[91]));
INVX1 exu_U17475(.A(div_dnext[91]), .Y(exu_n4177));
AND2X1 exu_U17476(.A(div_adder_out_27), .B(exu_n16250), .Y(div_d_mux_n39));
INVX1 exu_U17477(.A(div_d_mux_n39), .Y(exu_n4178));
AND2X1 exu_U17478(.A(div_d_mux_n41), .B(exu_n10396), .Y(div_dnext[90]));
INVX1 exu_U17479(.A(div_dnext[90]), .Y(exu_n4179));
AND2X1 exu_U17480(.A(div_adder_out_26), .B(exu_n16250), .Y(div_d_mux_n43));
INVX1 exu_U17481(.A(div_d_mux_n43), .Y(exu_n4180));
AND2X1 exu_U17482(.A(div_d_mux_n45), .B(exu_n10397), .Y(div_dnext[8]));
INVX1 exu_U17483(.A(div_dnext[8]), .Y(exu_n4181));
AND2X1 exu_U17484(.A(div_d[7]), .B(ecl_div_sel_adder), .Y(div_d_mux_n47));
INVX1 exu_U17485(.A(div_d_mux_n47), .Y(exu_n4182));
AND2X1 exu_U17486(.A(div_d_mux_n49), .B(exu_n10398), .Y(div_dnext[89]));
INVX1 exu_U17487(.A(div_dnext[89]), .Y(exu_n4183));
AND2X1 exu_U17488(.A(div_adder_out_25), .B(exu_n16250), .Y(div_d_mux_n51));
INVX1 exu_U17489(.A(div_d_mux_n51), .Y(exu_n4184));
AND2X1 exu_U17490(.A(div_d_mux_n53), .B(exu_n10399), .Y(div_dnext[88]));
INVX1 exu_U17491(.A(div_dnext[88]), .Y(exu_n4185));
AND2X1 exu_U17492(.A(div_adder_out_24), .B(ecl_div_sel_adder), .Y(div_d_mux_n55));
INVX1 exu_U17493(.A(div_d_mux_n55), .Y(exu_n4186));
AND2X1 exu_U17494(.A(div_d_mux_n57), .B(exu_n10400), .Y(div_dnext[87]));
INVX1 exu_U17495(.A(div_dnext[87]), .Y(exu_n4187));
AND2X1 exu_U17496(.A(div_adder_out_23), .B(exu_n16250), .Y(div_d_mux_n59));
INVX1 exu_U17497(.A(div_d_mux_n59), .Y(exu_n4188));
AND2X1 exu_U17498(.A(div_d_mux_n61), .B(exu_n10401), .Y(div_dnext[86]));
INVX1 exu_U17499(.A(div_dnext[86]), .Y(exu_n4189));
AND2X1 exu_U17500(.A(div_adder_out_22), .B(exu_n16250), .Y(div_d_mux_n63));
INVX1 exu_U17501(.A(div_d_mux_n63), .Y(exu_n4190));
AND2X1 exu_U17502(.A(div_d_mux_n65), .B(exu_n10402), .Y(div_dnext[85]));
INVX1 exu_U17503(.A(div_dnext[85]), .Y(exu_n4191));
AND2X1 exu_U17504(.A(div_adder_out_21), .B(exu_n16250), .Y(div_d_mux_n67));
INVX1 exu_U17505(.A(div_d_mux_n67), .Y(exu_n4192));
AND2X1 exu_U17506(.A(div_d_mux_n69), .B(exu_n10403), .Y(div_dnext[84]));
INVX1 exu_U17507(.A(div_dnext[84]), .Y(exu_n4193));
AND2X1 exu_U17508(.A(div_adder_out_20), .B(ecl_div_sel_adder), .Y(div_d_mux_n71));
INVX1 exu_U17509(.A(div_d_mux_n71), .Y(exu_n4194));
AND2X1 exu_U17510(.A(div_d_mux_n73), .B(exu_n10404), .Y(div_dnext[83]));
INVX1 exu_U17511(.A(div_dnext[83]), .Y(exu_n4195));
AND2X1 exu_U17512(.A(div_adder_out_19), .B(exu_n16250), .Y(div_d_mux_n75));
INVX1 exu_U17513(.A(div_d_mux_n75), .Y(exu_n4196));
AND2X1 exu_U17514(.A(div_d_mux_n77), .B(exu_n10405), .Y(div_dnext[82]));
INVX1 exu_U17515(.A(div_dnext[82]), .Y(exu_n4197));
AND2X1 exu_U17516(.A(div_adder_out_18), .B(exu_n16250), .Y(div_d_mux_n79));
INVX1 exu_U17517(.A(div_d_mux_n79), .Y(exu_n4198));
AND2X1 exu_U17518(.A(div_d_mux_n81), .B(exu_n10406), .Y(div_dnext[81]));
INVX1 exu_U17519(.A(div_dnext[81]), .Y(exu_n4199));
AND2X1 exu_U17520(.A(div_adder_out_17), .B(ecl_div_sel_adder), .Y(div_d_mux_n83));
INVX1 exu_U17521(.A(div_d_mux_n83), .Y(exu_n4200));
AND2X1 exu_U17522(.A(div_d_mux_n85), .B(exu_n10407), .Y(div_dnext[80]));
INVX1 exu_U17523(.A(div_dnext[80]), .Y(exu_n4201));
AND2X1 exu_U17524(.A(div_adder_out_16), .B(ecl_div_sel_adder), .Y(div_d_mux_n87));
INVX1 exu_U17525(.A(div_d_mux_n87), .Y(exu_n4202));
AND2X1 exu_U17526(.A(div_d_mux_n89), .B(exu_n10408), .Y(div_dnext[7]));
INVX1 exu_U17527(.A(div_dnext[7]), .Y(exu_n4203));
AND2X1 exu_U17528(.A(div_d[6]), .B(ecl_div_sel_adder), .Y(div_d_mux_n91));
INVX1 exu_U17529(.A(div_d_mux_n91), .Y(exu_n4204));
AND2X1 exu_U17530(.A(div_d_mux_n93), .B(exu_n10409), .Y(div_dnext[79]));
INVX1 exu_U17531(.A(div_dnext[79]), .Y(exu_n4205));
AND2X1 exu_U17532(.A(div_adder_out_15), .B(exu_n16250), .Y(div_d_mux_n95));
INVX1 exu_U17533(.A(div_d_mux_n95), .Y(exu_n4206));
AND2X1 exu_U17534(.A(div_d_mux_n97), .B(exu_n10410), .Y(div_dnext[78]));
INVX1 exu_U17535(.A(div_dnext[78]), .Y(exu_n4207));
AND2X1 exu_U17536(.A(div_adder_out_14), .B(exu_n16250), .Y(div_d_mux_n99));
INVX1 exu_U17537(.A(div_d_mux_n99), .Y(exu_n4208));
AND2X1 exu_U17538(.A(div_d_mux_n101), .B(exu_n10411), .Y(div_dnext[77]));
INVX1 exu_U17539(.A(div_dnext[77]), .Y(exu_n4209));
AND2X1 exu_U17540(.A(div_adder_out_13), .B(ecl_div_sel_adder), .Y(div_d_mux_n103));
INVX1 exu_U17541(.A(div_d_mux_n103), .Y(exu_n4210));
AND2X1 exu_U17542(.A(div_d_mux_n105), .B(exu_n10412), .Y(div_dnext[76]));
INVX1 exu_U17543(.A(div_dnext[76]), .Y(exu_n4211));
AND2X1 exu_U17544(.A(div_adder_out_12), .B(exu_n16250), .Y(div_d_mux_n107));
INVX1 exu_U17545(.A(div_d_mux_n107), .Y(exu_n4212));
AND2X1 exu_U17546(.A(div_d_mux_n109), .B(exu_n10413), .Y(div_dnext[75]));
INVX1 exu_U17547(.A(div_dnext[75]), .Y(exu_n4213));
AND2X1 exu_U17548(.A(div_adder_out_11), .B(exu_n16250), .Y(div_d_mux_n111));
INVX1 exu_U17549(.A(div_d_mux_n111), .Y(exu_n4214));
AND2X1 exu_U17550(.A(div_d_mux_n113), .B(exu_n10414), .Y(div_dnext[74]));
INVX1 exu_U17551(.A(div_dnext[74]), .Y(exu_n4215));
AND2X1 exu_U17552(.A(div_adder_out_10), .B(exu_n16250), .Y(div_d_mux_n115));
INVX1 exu_U17553(.A(div_d_mux_n115), .Y(exu_n4216));
AND2X1 exu_U17554(.A(div_d_mux_n117), .B(exu_n10415), .Y(div_dnext[73]));
INVX1 exu_U17555(.A(div_dnext[73]), .Y(exu_n4217));
AND2X1 exu_U17556(.A(div_adder_out_9), .B(exu_n16250), .Y(div_d_mux_n119));
INVX1 exu_U17557(.A(div_d_mux_n119), .Y(exu_n4218));
AND2X1 exu_U17558(.A(div_d_mux_n121), .B(exu_n10416), .Y(div_dnext[72]));
INVX1 exu_U17559(.A(div_dnext[72]), .Y(exu_n4219));
AND2X1 exu_U17560(.A(div_adder_out_8), .B(exu_n16250), .Y(div_d_mux_n123));
INVX1 exu_U17561(.A(div_d_mux_n123), .Y(exu_n4220));
AND2X1 exu_U17562(.A(div_d_mux_n125), .B(exu_n10417), .Y(div_dnext[71]));
INVX1 exu_U17563(.A(div_dnext[71]), .Y(exu_n4221));
AND2X1 exu_U17564(.A(div_adder_out_7), .B(exu_n16250), .Y(div_d_mux_n127));
INVX1 exu_U17565(.A(div_d_mux_n127), .Y(exu_n4222));
AND2X1 exu_U17566(.A(div_d_mux_n129), .B(exu_n10418), .Y(div_dnext[70]));
INVX1 exu_U17567(.A(div_dnext[70]), .Y(exu_n4223));
AND2X1 exu_U17568(.A(div_adder_out_6), .B(exu_n16250), .Y(div_d_mux_n131));
INVX1 exu_U17569(.A(div_d_mux_n131), .Y(exu_n4224));
AND2X1 exu_U17570(.A(div_d_mux_n133), .B(exu_n10419), .Y(div_dnext[6]));
INVX1 exu_U17571(.A(div_dnext[6]), .Y(exu_n4225));
AND2X1 exu_U17572(.A(div_d[5]), .B(exu_n16250), .Y(div_d_mux_n135));
INVX1 exu_U17573(.A(div_d_mux_n135), .Y(exu_n4226));
AND2X1 exu_U17574(.A(div_d_mux_n137), .B(exu_n10420), .Y(div_dnext[69]));
INVX1 exu_U17575(.A(div_dnext[69]), .Y(exu_n4227));
AND2X1 exu_U17576(.A(div_adder_out_5), .B(exu_n16250), .Y(div_d_mux_n139));
INVX1 exu_U17577(.A(div_d_mux_n139), .Y(exu_n4228));
AND2X1 exu_U17578(.A(div_d_mux_n141), .B(exu_n10421), .Y(div_dnext[68]));
INVX1 exu_U17579(.A(div_dnext[68]), .Y(exu_n4229));
AND2X1 exu_U17580(.A(div_adder_out_4), .B(exu_n16250), .Y(div_d_mux_n143));
INVX1 exu_U17581(.A(div_d_mux_n143), .Y(exu_n4230));
AND2X1 exu_U17582(.A(div_d_mux_n145), .B(exu_n10422), .Y(div_dnext[67]));
INVX1 exu_U17583(.A(div_dnext[67]), .Y(exu_n4231));
AND2X1 exu_U17584(.A(div_adder_out_3), .B(exu_n16250), .Y(div_d_mux_n147));
INVX1 exu_U17585(.A(div_d_mux_n147), .Y(exu_n4232));
AND2X1 exu_U17586(.A(div_d_mux_n149), .B(exu_n10423), .Y(div_dnext[66]));
INVX1 exu_U17587(.A(div_dnext[66]), .Y(exu_n4233));
AND2X1 exu_U17588(.A(div_adder_out_2), .B(exu_n16250), .Y(div_d_mux_n151));
INVX1 exu_U17589(.A(div_d_mux_n151), .Y(exu_n4234));
AND2X1 exu_U17590(.A(div_d_mux_n153), .B(exu_n10424), .Y(div_dnext[65]));
INVX1 exu_U17591(.A(div_dnext[65]), .Y(exu_n4235));
AND2X1 exu_U17592(.A(div_adder_out_1), .B(exu_n16250), .Y(div_d_mux_n155));
INVX1 exu_U17593(.A(div_d_mux_n155), .Y(exu_n4236));
AND2X1 exu_U17594(.A(div_d_mux_n157), .B(exu_n10425), .Y(div_dnext[64]));
INVX1 exu_U17595(.A(div_dnext[64]), .Y(exu_n4237));
AND2X1 exu_U17596(.A(div_adder_out_0), .B(exu_n16250), .Y(div_d_mux_n159));
INVX1 exu_U17597(.A(div_d_mux_n159), .Y(exu_n4238));
AND2X1 exu_U17598(.A(div_d_mux_n161), .B(exu_n10426), .Y(div_dnext[63]));
INVX1 exu_U17599(.A(div_dnext[63]), .Y(exu_n4239));
AND2X1 exu_U17600(.A(div_ecl_d_62), .B(exu_n16250), .Y(div_d_mux_n163));
INVX1 exu_U17601(.A(div_d_mux_n163), .Y(exu_n4240));
AND2X1 exu_U17602(.A(div_d_mux_n165), .B(exu_n10427), .Y(div_dnext[62]));
INVX1 exu_U17603(.A(div_dnext[62]), .Y(exu_n4241));
AND2X1 exu_U17604(.A(div_d[61]), .B(ecl_div_sel_adder), .Y(div_d_mux_n167));
INVX1 exu_U17605(.A(div_d_mux_n167), .Y(exu_n4242));
AND2X1 exu_U17606(.A(div_d_mux_n169), .B(exu_n10428), .Y(div_dnext[61]));
INVX1 exu_U17607(.A(div_dnext[61]), .Y(exu_n4243));
AND2X1 exu_U17608(.A(div_d[60]), .B(ecl_div_sel_adder), .Y(div_d_mux_n171));
INVX1 exu_U17609(.A(div_d_mux_n171), .Y(exu_n4244));
AND2X1 exu_U17610(.A(div_d_mux_n173), .B(exu_n10429), .Y(div_dnext[60]));
INVX1 exu_U17611(.A(div_dnext[60]), .Y(exu_n4245));
AND2X1 exu_U17612(.A(div_d[59]), .B(ecl_div_sel_adder), .Y(div_d_mux_n175));
INVX1 exu_U17613(.A(div_d_mux_n175), .Y(exu_n4246));
AND2X1 exu_U17614(.A(div_d_mux_n177), .B(exu_n10430), .Y(div_dnext[5]));
INVX1 exu_U17615(.A(div_dnext[5]), .Y(exu_n4247));
AND2X1 exu_U17616(.A(div_d[4]), .B(exu_n16250), .Y(div_d_mux_n179));
INVX1 exu_U17617(.A(div_d_mux_n179), .Y(exu_n4248));
AND2X1 exu_U17618(.A(div_d_mux_n181), .B(exu_n10431), .Y(div_dnext[59]));
INVX1 exu_U17619(.A(div_dnext[59]), .Y(exu_n4249));
AND2X1 exu_U17620(.A(div_d[58]), .B(ecl_div_sel_adder), .Y(div_d_mux_n183));
INVX1 exu_U17621(.A(div_d_mux_n183), .Y(exu_n4250));
AND2X1 exu_U17622(.A(div_d_mux_n185), .B(exu_n10432), .Y(div_dnext[58]));
INVX1 exu_U17623(.A(div_dnext[58]), .Y(exu_n4251));
AND2X1 exu_U17624(.A(div_d[57]), .B(exu_n16250), .Y(div_d_mux_n187));
INVX1 exu_U17625(.A(div_d_mux_n187), .Y(exu_n4252));
AND2X1 exu_U17626(.A(div_d_mux_n189), .B(exu_n10433), .Y(div_dnext[57]));
INVX1 exu_U17627(.A(div_dnext[57]), .Y(exu_n4253));
AND2X1 exu_U17628(.A(div_d[56]), .B(exu_n16250), .Y(div_d_mux_n191));
INVX1 exu_U17629(.A(div_d_mux_n191), .Y(exu_n4254));
AND2X1 exu_U17630(.A(div_d_mux_n193), .B(exu_n10434), .Y(div_dnext[56]));
INVX1 exu_U17631(.A(div_dnext[56]), .Y(exu_n4255));
AND2X1 exu_U17632(.A(div_d[55]), .B(exu_n16250), .Y(div_d_mux_n195));
INVX1 exu_U17633(.A(div_d_mux_n195), .Y(exu_n4256));
AND2X1 exu_U17634(.A(div_d_mux_n197), .B(exu_n10435), .Y(div_dnext[55]));
INVX1 exu_U17635(.A(div_dnext[55]), .Y(exu_n4257));
AND2X1 exu_U17636(.A(div_d[54]), .B(ecl_div_sel_adder), .Y(div_d_mux_n199));
INVX1 exu_U17637(.A(div_d_mux_n199), .Y(exu_n4258));
AND2X1 exu_U17638(.A(div_d_mux_n201), .B(exu_n10436), .Y(div_dnext[54]));
INVX1 exu_U17639(.A(div_dnext[54]), .Y(exu_n4259));
AND2X1 exu_U17640(.A(div_d[53]), .B(exu_n16250), .Y(div_d_mux_n203));
INVX1 exu_U17641(.A(div_d_mux_n203), .Y(exu_n4260));
AND2X1 exu_U17642(.A(div_d_mux_n205), .B(exu_n10437), .Y(div_dnext[53]));
INVX1 exu_U17643(.A(div_dnext[53]), .Y(exu_n4261));
AND2X1 exu_U17644(.A(div_d[52]), .B(ecl_div_sel_adder), .Y(div_d_mux_n207));
INVX1 exu_U17645(.A(div_d_mux_n207), .Y(exu_n4262));
AND2X1 exu_U17646(.A(div_d_mux_n209), .B(exu_n10438), .Y(div_dnext[52]));
INVX1 exu_U17647(.A(div_dnext[52]), .Y(exu_n4263));
AND2X1 exu_U17648(.A(div_d[51]), .B(exu_n16250), .Y(div_d_mux_n211));
INVX1 exu_U17649(.A(div_d_mux_n211), .Y(exu_n4264));
AND2X1 exu_U17650(.A(div_d_mux_n213), .B(exu_n10439), .Y(div_dnext[51]));
INVX1 exu_U17651(.A(div_dnext[51]), .Y(exu_n4265));
AND2X1 exu_U17652(.A(div_d[50]), .B(ecl_div_sel_adder), .Y(div_d_mux_n215));
INVX1 exu_U17653(.A(div_d_mux_n215), .Y(exu_n4266));
AND2X1 exu_U17654(.A(div_d_mux_n217), .B(exu_n10440), .Y(div_dnext[50]));
INVX1 exu_U17655(.A(div_dnext[50]), .Y(exu_n4267));
AND2X1 exu_U17656(.A(div_d[49]), .B(ecl_div_sel_adder), .Y(div_d_mux_n219));
INVX1 exu_U17657(.A(div_d_mux_n219), .Y(exu_n4268));
AND2X1 exu_U17658(.A(div_d_mux_n221), .B(exu_n10441), .Y(div_dnext[4]));
INVX1 exu_U17659(.A(div_dnext[4]), .Y(exu_n4269));
AND2X1 exu_U17660(.A(div_d[3]), .B(ecl_div_sel_adder), .Y(div_d_mux_n223));
INVX1 exu_U17661(.A(div_d_mux_n223), .Y(exu_n4270));
AND2X1 exu_U17662(.A(div_d_mux_n225), .B(exu_n10442), .Y(div_dnext[49]));
INVX1 exu_U17663(.A(div_dnext[49]), .Y(exu_n4271));
AND2X1 exu_U17664(.A(div_d[48]), .B(ecl_div_sel_adder), .Y(div_d_mux_n227));
INVX1 exu_U17665(.A(div_d_mux_n227), .Y(exu_n4272));
AND2X1 exu_U17666(.A(div_d_mux_n229), .B(exu_n10443), .Y(div_dnext[48]));
INVX1 exu_U17667(.A(div_dnext[48]), .Y(exu_n4273));
AND2X1 exu_U17668(.A(div_d[47]), .B(ecl_div_sel_adder), .Y(div_d_mux_n231));
INVX1 exu_U17669(.A(div_d_mux_n231), .Y(exu_n4274));
AND2X1 exu_U17670(.A(div_d_mux_n233), .B(exu_n10444), .Y(div_dnext[47]));
INVX1 exu_U17671(.A(div_dnext[47]), .Y(exu_n4275));
AND2X1 exu_U17672(.A(div_d[46]), .B(exu_n16250), .Y(div_d_mux_n235));
INVX1 exu_U17673(.A(div_d_mux_n235), .Y(exu_n4276));
AND2X1 exu_U17674(.A(div_d_mux_n237), .B(exu_n10445), .Y(div_dnext[46]));
INVX1 exu_U17675(.A(div_dnext[46]), .Y(exu_n4277));
AND2X1 exu_U17676(.A(div_d[45]), .B(ecl_div_sel_adder), .Y(div_d_mux_n239));
INVX1 exu_U17677(.A(div_d_mux_n239), .Y(exu_n4278));
AND2X1 exu_U17678(.A(div_d_mux_n241), .B(exu_n10446), .Y(div_dnext[45]));
INVX1 exu_U17679(.A(div_dnext[45]), .Y(exu_n4279));
AND2X1 exu_U17680(.A(div_d[44]), .B(exu_n16250), .Y(div_d_mux_n243));
INVX1 exu_U17681(.A(div_d_mux_n243), .Y(exu_n4280));
AND2X1 exu_U17682(.A(div_d_mux_n245), .B(exu_n10447), .Y(div_dnext[44]));
INVX1 exu_U17683(.A(div_dnext[44]), .Y(exu_n4281));
AND2X1 exu_U17684(.A(div_d[43]), .B(exu_n16250), .Y(div_d_mux_n247));
INVX1 exu_U17685(.A(div_d_mux_n247), .Y(exu_n4282));
AND2X1 exu_U17686(.A(div_d_mux_n249), .B(exu_n10448), .Y(div_dnext[43]));
INVX1 exu_U17687(.A(div_dnext[43]), .Y(exu_n4283));
AND2X1 exu_U17688(.A(div_d[42]), .B(ecl_div_sel_adder), .Y(div_d_mux_n251));
INVX1 exu_U17689(.A(div_d_mux_n251), .Y(exu_n4284));
AND2X1 exu_U17690(.A(div_d_mux_n253), .B(exu_n10449), .Y(div_dnext[42]));
INVX1 exu_U17691(.A(div_dnext[42]), .Y(exu_n4285));
AND2X1 exu_U17692(.A(div_d[41]), .B(exu_n16250), .Y(div_d_mux_n255));
INVX1 exu_U17693(.A(div_d_mux_n255), .Y(exu_n4286));
AND2X1 exu_U17694(.A(div_d_mux_n257), .B(exu_n10450), .Y(div_dnext[41]));
INVX1 exu_U17695(.A(div_dnext[41]), .Y(exu_n4287));
AND2X1 exu_U17696(.A(div_d[40]), .B(exu_n16250), .Y(div_d_mux_n259));
INVX1 exu_U17697(.A(div_d_mux_n259), .Y(exu_n4288));
AND2X1 exu_U17698(.A(div_d_mux_n261), .B(exu_n10451), .Y(div_dnext[40]));
INVX1 exu_U17699(.A(div_dnext[40]), .Y(exu_n4289));
AND2X1 exu_U17700(.A(div_d[39]), .B(ecl_div_sel_adder), .Y(div_d_mux_n263));
INVX1 exu_U17701(.A(div_d_mux_n263), .Y(exu_n4290));
AND2X1 exu_U17702(.A(div_d_mux_n265), .B(exu_n10452), .Y(div_dnext[3]));
INVX1 exu_U17703(.A(div_dnext[3]), .Y(exu_n4291));
AND2X1 exu_U17704(.A(div_d[2]), .B(exu_n16250), .Y(div_d_mux_n267));
INVX1 exu_U17705(.A(div_d_mux_n267), .Y(exu_n4292));
AND2X1 exu_U17706(.A(div_d_mux_n269), .B(exu_n10453), .Y(div_dnext[39]));
INVX1 exu_U17707(.A(div_dnext[39]), .Y(exu_n4293));
AND2X1 exu_U17708(.A(div_d[38]), .B(ecl_div_sel_adder), .Y(div_d_mux_n271));
INVX1 exu_U17709(.A(div_d_mux_n271), .Y(exu_n4294));
AND2X1 exu_U17710(.A(div_d_mux_n273), .B(exu_n10454), .Y(div_dnext[38]));
INVX1 exu_U17711(.A(div_dnext[38]), .Y(exu_n4295));
AND2X1 exu_U17712(.A(div_d[37]), .B(ecl_div_sel_adder), .Y(div_d_mux_n275));
INVX1 exu_U17713(.A(div_d_mux_n275), .Y(exu_n4296));
AND2X1 exu_U17714(.A(div_d_mux_n277), .B(exu_n10455), .Y(div_dnext[37]));
INVX1 exu_U17715(.A(div_dnext[37]), .Y(exu_n4297));
AND2X1 exu_U17716(.A(div_d[36]), .B(ecl_div_sel_adder), .Y(div_d_mux_n279));
INVX1 exu_U17717(.A(div_d_mux_n279), .Y(exu_n4298));
AND2X1 exu_U17718(.A(div_d_mux_n281), .B(exu_n10456), .Y(div_dnext[36]));
INVX1 exu_U17719(.A(div_dnext[36]), .Y(exu_n4299));
AND2X1 exu_U17720(.A(div_d[35]), .B(exu_n16250), .Y(div_d_mux_n283));
INVX1 exu_U17721(.A(div_d_mux_n283), .Y(exu_n4300));
AND2X1 exu_U17722(.A(div_d_mux_n285), .B(exu_n10457), .Y(div_dnext[35]));
INVX1 exu_U17723(.A(div_dnext[35]), .Y(exu_n4301));
AND2X1 exu_U17724(.A(div_d[34]), .B(exu_n16250), .Y(div_d_mux_n287));
INVX1 exu_U17725(.A(div_d_mux_n287), .Y(exu_n4302));
AND2X1 exu_U17726(.A(div_d_mux_n289), .B(exu_n10458), .Y(div_dnext[34]));
INVX1 exu_U17727(.A(div_dnext[34]), .Y(exu_n4303));
AND2X1 exu_U17728(.A(div_d[33]), .B(exu_n16250), .Y(div_d_mux_n291));
INVX1 exu_U17729(.A(div_d_mux_n291), .Y(exu_n4304));
AND2X1 exu_U17730(.A(div_d_mux_n293), .B(exu_n10459), .Y(div_dnext[33]));
INVX1 exu_U17731(.A(div_dnext[33]), .Y(exu_n4305));
AND2X1 exu_U17732(.A(div_d[32]), .B(ecl_div_sel_adder), .Y(div_d_mux_n295));
INVX1 exu_U17733(.A(div_d_mux_n295), .Y(exu_n4306));
AND2X1 exu_U17734(.A(div_d_mux_n297), .B(exu_n10460), .Y(div_dnext[32]));
INVX1 exu_U17735(.A(div_dnext[32]), .Y(exu_n4307));
AND2X1 exu_U17736(.A(div_d[31]), .B(exu_n16250), .Y(div_d_mux_n299));
INVX1 exu_U17737(.A(div_d_mux_n299), .Y(exu_n4308));
AND2X1 exu_U17738(.A(div_d_mux_n301), .B(exu_n10461), .Y(div_dnext[31]));
INVX1 exu_U17739(.A(div_dnext[31]), .Y(exu_n4309));
AND2X1 exu_U17740(.A(div_d[30]), .B(ecl_div_sel_adder), .Y(div_d_mux_n303));
INVX1 exu_U17741(.A(div_d_mux_n303), .Y(exu_n4310));
AND2X1 exu_U17742(.A(div_d_mux_n305), .B(exu_n10462), .Y(div_dnext[30]));
INVX1 exu_U17743(.A(div_dnext[30]), .Y(exu_n4311));
AND2X1 exu_U17744(.A(div_d[29]), .B(exu_n16250), .Y(div_d_mux_n307));
INVX1 exu_U17745(.A(div_d_mux_n307), .Y(exu_n4312));
AND2X1 exu_U17746(.A(div_d_mux_n309), .B(exu_n10463), .Y(div_dnext[2]));
INVX1 exu_U17747(.A(div_dnext[2]), .Y(exu_n4313));
AND2X1 exu_U17748(.A(div_d[1]), .B(exu_n16250), .Y(div_d_mux_n311));
INVX1 exu_U17749(.A(div_d_mux_n311), .Y(exu_n4314));
AND2X1 exu_U17750(.A(div_d_mux_n313), .B(exu_n10464), .Y(div_dnext[29]));
INVX1 exu_U17751(.A(div_dnext[29]), .Y(exu_n4315));
AND2X1 exu_U17752(.A(div_d[28]), .B(ecl_div_sel_adder), .Y(div_d_mux_n315));
INVX1 exu_U17753(.A(div_d_mux_n315), .Y(exu_n4316));
AND2X1 exu_U17754(.A(div_d_mux_n317), .B(exu_n10465), .Y(div_dnext[28]));
INVX1 exu_U17755(.A(div_dnext[28]), .Y(exu_n4317));
AND2X1 exu_U17756(.A(div_d[27]), .B(ecl_div_sel_adder), .Y(div_d_mux_n319));
INVX1 exu_U17757(.A(div_d_mux_n319), .Y(exu_n4318));
AND2X1 exu_U17758(.A(div_d_mux_n321), .B(exu_n10466), .Y(div_dnext[27]));
INVX1 exu_U17759(.A(div_dnext[27]), .Y(exu_n4319));
AND2X1 exu_U17760(.A(div_d[26]), .B(ecl_div_sel_adder), .Y(div_d_mux_n323));
INVX1 exu_U17761(.A(div_d_mux_n323), .Y(exu_n4320));
AND2X1 exu_U17762(.A(div_d_mux_n325), .B(exu_n10467), .Y(div_dnext[26]));
INVX1 exu_U17763(.A(div_dnext[26]), .Y(exu_n4321));
AND2X1 exu_U17764(.A(div_d[25]), .B(ecl_div_sel_adder), .Y(div_d_mux_n327));
INVX1 exu_U17765(.A(div_d_mux_n327), .Y(exu_n4322));
AND2X1 exu_U17766(.A(div_d_mux_n329), .B(exu_n10468), .Y(div_dnext[25]));
INVX1 exu_U17767(.A(div_dnext[25]), .Y(exu_n4323));
AND2X1 exu_U17768(.A(div_d[24]), .B(ecl_div_sel_adder), .Y(div_d_mux_n331));
INVX1 exu_U17769(.A(div_d_mux_n331), .Y(exu_n4324));
AND2X1 exu_U17770(.A(div_d_mux_n333), .B(exu_n10469), .Y(div_dnext[24]));
INVX1 exu_U17771(.A(div_dnext[24]), .Y(exu_n4325));
AND2X1 exu_U17772(.A(div_d[23]), .B(ecl_div_sel_adder), .Y(div_d_mux_n335));
INVX1 exu_U17773(.A(div_d_mux_n335), .Y(exu_n4326));
AND2X1 exu_U17774(.A(div_d_mux_n337), .B(exu_n10470), .Y(div_dnext[23]));
INVX1 exu_U17775(.A(div_dnext[23]), .Y(exu_n4327));
AND2X1 exu_U17776(.A(div_d[22]), .B(ecl_div_sel_adder), .Y(div_d_mux_n339));
INVX1 exu_U17777(.A(div_d_mux_n339), .Y(exu_n4328));
AND2X1 exu_U17778(.A(div_d_mux_n341), .B(exu_n10471), .Y(div_dnext[22]));
INVX1 exu_U17779(.A(div_dnext[22]), .Y(exu_n4329));
AND2X1 exu_U17780(.A(div_d[21]), .B(ecl_div_sel_adder), .Y(div_d_mux_n343));
INVX1 exu_U17781(.A(div_d_mux_n343), .Y(exu_n4330));
AND2X1 exu_U17782(.A(div_d_mux_n345), .B(exu_n10472), .Y(div_dnext[21]));
INVX1 exu_U17783(.A(div_dnext[21]), .Y(exu_n4331));
AND2X1 exu_U17784(.A(div_d[20]), .B(ecl_div_sel_adder), .Y(div_d_mux_n347));
INVX1 exu_U17785(.A(div_d_mux_n347), .Y(exu_n4332));
AND2X1 exu_U17786(.A(div_d_mux_n349), .B(exu_n10473), .Y(div_dnext[20]));
INVX1 exu_U17787(.A(div_dnext[20]), .Y(exu_n4333));
AND2X1 exu_U17788(.A(div_d[19]), .B(ecl_div_sel_adder), .Y(div_d_mux_n351));
INVX1 exu_U17789(.A(div_d_mux_n351), .Y(exu_n4334));
AND2X1 exu_U17790(.A(div_d_mux_n353), .B(exu_n10474), .Y(div_dnext[1]));
INVX1 exu_U17791(.A(div_dnext[1]), .Y(exu_n4335));
AND2X1 exu_U17792(.A(div_d[0]), .B(ecl_div_sel_adder), .Y(div_d_mux_n355));
INVX1 exu_U17793(.A(div_d_mux_n355), .Y(exu_n4336));
AND2X1 exu_U17794(.A(div_d_mux_n357), .B(exu_n10475), .Y(div_dnext[19]));
INVX1 exu_U17795(.A(div_dnext[19]), .Y(exu_n4337));
AND2X1 exu_U17796(.A(div_d[18]), .B(ecl_div_sel_adder), .Y(div_d_mux_n359));
INVX1 exu_U17797(.A(div_d_mux_n359), .Y(exu_n4338));
AND2X1 exu_U17798(.A(div_d_mux_n361), .B(exu_n10476), .Y(div_dnext[18]));
INVX1 exu_U17799(.A(div_dnext[18]), .Y(exu_n4339));
AND2X1 exu_U17800(.A(div_d[17]), .B(ecl_div_sel_adder), .Y(div_d_mux_n363));
INVX1 exu_U17801(.A(div_d_mux_n363), .Y(exu_n4340));
AND2X1 exu_U17802(.A(div_d_mux_n365), .B(exu_n10477), .Y(div_dnext[17]));
INVX1 exu_U17803(.A(div_dnext[17]), .Y(exu_n4341));
AND2X1 exu_U17804(.A(div_d[16]), .B(ecl_div_sel_adder), .Y(div_d_mux_n367));
INVX1 exu_U17805(.A(div_d_mux_n367), .Y(exu_n4342));
AND2X1 exu_U17806(.A(div_d_mux_n369), .B(exu_n10478), .Y(div_dnext[16]));
INVX1 exu_U17807(.A(div_dnext[16]), .Y(exu_n4343));
AND2X1 exu_U17808(.A(div_d[15]), .B(exu_n16250), .Y(div_d_mux_n371));
INVX1 exu_U17809(.A(div_d_mux_n371), .Y(exu_n4344));
AND2X1 exu_U17810(.A(div_d_mux_n373), .B(exu_n10479), .Y(div_dnext[15]));
INVX1 exu_U17811(.A(div_dnext[15]), .Y(exu_n4345));
AND2X1 exu_U17812(.A(div_d[14]), .B(ecl_div_sel_adder), .Y(div_d_mux_n375));
INVX1 exu_U17813(.A(div_d_mux_n375), .Y(exu_n4346));
AND2X1 exu_U17814(.A(div_d_mux_n377), .B(exu_n10480), .Y(div_dnext[14]));
INVX1 exu_U17815(.A(div_dnext[14]), .Y(exu_n4347));
AND2X1 exu_U17816(.A(div_d[13]), .B(exu_n16250), .Y(div_d_mux_n379));
INVX1 exu_U17817(.A(div_d_mux_n379), .Y(exu_n4348));
AND2X1 exu_U17818(.A(div_d_mux_n381), .B(exu_n10481), .Y(div_dnext[13]));
INVX1 exu_U17819(.A(div_dnext[13]), .Y(exu_n4349));
AND2X1 exu_U17820(.A(div_d[12]), .B(ecl_div_sel_adder), .Y(div_d_mux_n383));
INVX1 exu_U17821(.A(div_d_mux_n383), .Y(exu_n4350));
AND2X1 exu_U17822(.A(div_d_mux_n385), .B(exu_n10482), .Y(div_dnext[12]));
INVX1 exu_U17823(.A(div_dnext[12]), .Y(exu_n4351));
AND2X1 exu_U17824(.A(div_d[11]), .B(ecl_div_sel_adder), .Y(div_d_mux_n387));
INVX1 exu_U17825(.A(div_d_mux_n387), .Y(exu_n4352));
AND2X1 exu_U17826(.A(div_d_mux_n389), .B(exu_n10484), .Y(div_dnext[127]));
INVX1 exu_U17827(.A(div_dnext[127]), .Y(exu_n4353));
AND2X1 exu_U17828(.A(div_adder_out[63]), .B(exu_n16250), .Y(div_d_mux_n391));
INVX1 exu_U17829(.A(div_d_mux_n391), .Y(exu_n4354));
AND2X1 exu_U17830(.A(div_d_mux_n393), .B(exu_n10486), .Y(div_dnext[126]));
INVX1 exu_U17831(.A(div_dnext[126]), .Y(exu_n4355));
AND2X1 exu_U17832(.A(div_adder_out[62]), .B(exu_n16250), .Y(div_d_mux_n395));
INVX1 exu_U17833(.A(div_d_mux_n395), .Y(exu_n4356));
AND2X1 exu_U17834(.A(div_d_mux_n397), .B(exu_n10488), .Y(div_dnext[125]));
INVX1 exu_U17835(.A(div_dnext[125]), .Y(exu_n4357));
AND2X1 exu_U17836(.A(div_adder_out[61]), .B(ecl_div_sel_adder), .Y(div_d_mux_n399));
INVX1 exu_U17837(.A(div_d_mux_n399), .Y(exu_n4358));
AND2X1 exu_U17838(.A(div_d_mux_n401), .B(exu_n10490), .Y(div_dnext[124]));
INVX1 exu_U17839(.A(div_dnext[124]), .Y(exu_n4359));
AND2X1 exu_U17840(.A(div_adder_out[60]), .B(ecl_div_sel_adder), .Y(div_d_mux_n403));
INVX1 exu_U17841(.A(div_d_mux_n403), .Y(exu_n4360));
AND2X1 exu_U17842(.A(div_d_mux_n405), .B(exu_n10492), .Y(div_dnext[123]));
INVX1 exu_U17843(.A(div_dnext[123]), .Y(exu_n4361));
AND2X1 exu_U17844(.A(div_adder_out[59]), .B(exu_n16250), .Y(div_d_mux_n407));
INVX1 exu_U17845(.A(div_d_mux_n407), .Y(exu_n4362));
AND2X1 exu_U17846(.A(div_d_mux_n409), .B(exu_n10494), .Y(div_dnext[122]));
INVX1 exu_U17847(.A(div_dnext[122]), .Y(exu_n4363));
AND2X1 exu_U17848(.A(div_adder_out[58]), .B(exu_n16250), .Y(div_d_mux_n411));
INVX1 exu_U17849(.A(div_d_mux_n411), .Y(exu_n4364));
AND2X1 exu_U17850(.A(div_d_mux_n413), .B(exu_n10496), .Y(div_dnext[121]));
INVX1 exu_U17851(.A(div_dnext[121]), .Y(exu_n4365));
AND2X1 exu_U17852(.A(div_adder_out[57]), .B(ecl_div_sel_adder), .Y(div_d_mux_n415));
INVX1 exu_U17853(.A(div_d_mux_n415), .Y(exu_n4366));
AND2X1 exu_U17854(.A(div_d_mux_n417), .B(exu_n10498), .Y(div_dnext[120]));
INVX1 exu_U17855(.A(div_dnext[120]), .Y(exu_n4367));
AND2X1 exu_U17856(.A(div_adder_out[56]), .B(exu_n16250), .Y(div_d_mux_n419));
INVX1 exu_U17857(.A(div_d_mux_n419), .Y(exu_n4368));
AND2X1 exu_U17858(.A(div_d_mux_n421), .B(exu_n10499), .Y(div_dnext[11]));
INVX1 exu_U17859(.A(div_dnext[11]), .Y(exu_n4369));
AND2X1 exu_U17860(.A(div_d[10]), .B(exu_n16250), .Y(div_d_mux_n423));
INVX1 exu_U17861(.A(div_d_mux_n423), .Y(exu_n4370));
AND2X1 exu_U17862(.A(div_d_mux_n425), .B(exu_n10501), .Y(div_dnext[119]));
INVX1 exu_U17863(.A(div_dnext[119]), .Y(exu_n4371));
AND2X1 exu_U17864(.A(div_adder_out[55]), .B(exu_n16250), .Y(div_d_mux_n427));
INVX1 exu_U17865(.A(div_d_mux_n427), .Y(exu_n4372));
AND2X1 exu_U17866(.A(div_d_mux_n429), .B(exu_n10503), .Y(div_dnext[118]));
INVX1 exu_U17867(.A(div_dnext[118]), .Y(exu_n4373));
AND2X1 exu_U17868(.A(div_adder_out[54]), .B(exu_n16250), .Y(div_d_mux_n431));
INVX1 exu_U17869(.A(div_d_mux_n431), .Y(exu_n4374));
AND2X1 exu_U17870(.A(div_d_mux_n433), .B(exu_n10505), .Y(div_dnext[117]));
INVX1 exu_U17871(.A(div_dnext[117]), .Y(exu_n4375));
AND2X1 exu_U17872(.A(div_adder_out[53]), .B(exu_n16250), .Y(div_d_mux_n435));
INVX1 exu_U17873(.A(div_d_mux_n435), .Y(exu_n4376));
AND2X1 exu_U17874(.A(div_d_mux_n437), .B(exu_n10507), .Y(div_dnext[116]));
INVX1 exu_U17875(.A(div_dnext[116]), .Y(exu_n4377));
AND2X1 exu_U17876(.A(div_adder_out[52]), .B(exu_n16250), .Y(div_d_mux_n439));
INVX1 exu_U17877(.A(div_d_mux_n439), .Y(exu_n4378));
AND2X1 exu_U17878(.A(div_d_mux_n441), .B(exu_n10509), .Y(div_dnext[115]));
INVX1 exu_U17879(.A(div_dnext[115]), .Y(exu_n4379));
AND2X1 exu_U17880(.A(div_adder_out[51]), .B(exu_n16250), .Y(div_d_mux_n443));
INVX1 exu_U17881(.A(div_d_mux_n443), .Y(exu_n4380));
AND2X1 exu_U17882(.A(div_d_mux_n445), .B(exu_n10511), .Y(div_dnext[114]));
INVX1 exu_U17883(.A(div_dnext[114]), .Y(exu_n4381));
AND2X1 exu_U17884(.A(div_adder_out[50]), .B(exu_n16250), .Y(div_d_mux_n447));
INVX1 exu_U17885(.A(div_d_mux_n447), .Y(exu_n4382));
AND2X1 exu_U17886(.A(div_d_mux_n449), .B(exu_n10513), .Y(div_dnext[113]));
INVX1 exu_U17887(.A(div_dnext[113]), .Y(exu_n4383));
AND2X1 exu_U17888(.A(div_adder_out[49]), .B(exu_n16250), .Y(div_d_mux_n451));
INVX1 exu_U17889(.A(div_d_mux_n451), .Y(exu_n4384));
AND2X1 exu_U17890(.A(div_d_mux_n453), .B(exu_n10515), .Y(div_dnext[112]));
INVX1 exu_U17891(.A(div_dnext[112]), .Y(exu_n4385));
AND2X1 exu_U17892(.A(div_adder_out[48]), .B(exu_n16250), .Y(div_d_mux_n455));
INVX1 exu_U17893(.A(div_d_mux_n455), .Y(exu_n4386));
AND2X1 exu_U17894(.A(div_d_mux_n457), .B(exu_n10777), .Y(div_dnext[111]));
INVX1 exu_U17895(.A(div_dnext[111]), .Y(exu_n4387));
AND2X1 exu_U17896(.A(div_adder_out[47]), .B(exu_n16250), .Y(div_d_mux_n459));
INVX1 exu_U17897(.A(div_d_mux_n459), .Y(exu_n4388));
AND2X1 exu_U17898(.A(div_d_mux_n461), .B(exu_n10778), .Y(div_dnext[110]));
INVX1 exu_U17899(.A(div_dnext[110]), .Y(exu_n4389));
AND2X1 exu_U17900(.A(div_adder_out[46]), .B(exu_n16250), .Y(div_d_mux_n463));
INVX1 exu_U17901(.A(div_d_mux_n463), .Y(exu_n4390));
AND2X1 exu_U17902(.A(div_d_mux_n465), .B(exu_n10516), .Y(div_dnext[10]));
INVX1 exu_U17903(.A(div_dnext[10]), .Y(exu_n4391));
AND2X1 exu_U17904(.A(div_d[9]), .B(exu_n16250), .Y(div_d_mux_n467));
INVX1 exu_U17905(.A(div_d_mux_n467), .Y(exu_n4392));
AND2X1 exu_U17906(.A(div_d_mux_n469), .B(exu_n10777), .Y(div_dnext[109]));
INVX1 exu_U17907(.A(div_dnext[109]), .Y(exu_n4393));
AND2X1 exu_U17908(.A(div_adder_out[45]), .B(ecl_div_sel_adder), .Y(div_d_mux_n471));
INVX1 exu_U17909(.A(div_d_mux_n471), .Y(exu_n4394));
AND2X1 exu_U17910(.A(div_d_mux_n473), .B(exu_n10778), .Y(div_dnext[108]));
INVX1 exu_U17911(.A(div_dnext[108]), .Y(exu_n4395));
AND2X1 exu_U17912(.A(div_adder_out[44]), .B(exu_n16250), .Y(div_d_mux_n475));
INVX1 exu_U17913(.A(div_d_mux_n475), .Y(exu_n4396));
AND2X1 exu_U17914(.A(div_d_mux_n477), .B(exu_n10777), .Y(div_dnext[107]));
INVX1 exu_U17915(.A(div_dnext[107]), .Y(exu_n4397));
AND2X1 exu_U17916(.A(div_adder_out[43]), .B(ecl_div_sel_adder), .Y(div_d_mux_n479));
INVX1 exu_U17917(.A(div_d_mux_n479), .Y(exu_n4398));
AND2X1 exu_U17918(.A(div_d_mux_n481), .B(exu_n10778), .Y(div_dnext[106]));
INVX1 exu_U17919(.A(div_dnext[106]), .Y(exu_n4399));
AND2X1 exu_U17920(.A(div_adder_out[42]), .B(ecl_div_sel_adder), .Y(div_d_mux_n483));
INVX1 exu_U17921(.A(div_d_mux_n483), .Y(exu_n4400));
AND2X1 exu_U17922(.A(div_d_mux_n485), .B(exu_n10777), .Y(div_dnext[105]));
INVX1 exu_U17923(.A(div_dnext[105]), .Y(exu_n4401));
AND2X1 exu_U17924(.A(div_adder_out[41]), .B(exu_n16250), .Y(div_d_mux_n487));
INVX1 exu_U17925(.A(div_d_mux_n487), .Y(exu_n4402));
AND2X1 exu_U17926(.A(div_d_mux_n489), .B(exu_n10778), .Y(div_dnext[104]));
INVX1 exu_U17927(.A(div_dnext[104]), .Y(exu_n4403));
AND2X1 exu_U17928(.A(div_adder_out[40]), .B(exu_n16250), .Y(div_d_mux_n491));
INVX1 exu_U17929(.A(div_d_mux_n491), .Y(exu_n4404));
AND2X1 exu_U17930(.A(div_d_mux_n493), .B(exu_n10777), .Y(div_dnext[103]));
INVX1 exu_U17931(.A(div_dnext[103]), .Y(exu_n4405));
AND2X1 exu_U17932(.A(div_adder_out[39]), .B(ecl_div_sel_adder), .Y(div_d_mux_n495));
INVX1 exu_U17933(.A(div_d_mux_n495), .Y(exu_n4406));
AND2X1 exu_U17934(.A(div_d_mux_n497), .B(exu_n10778), .Y(div_dnext[102]));
INVX1 exu_U17935(.A(div_dnext[102]), .Y(exu_n4407));
AND2X1 exu_U17936(.A(div_adder_out[38]), .B(ecl_div_sel_adder), .Y(div_d_mux_n499));
INVX1 exu_U17937(.A(div_d_mux_n499), .Y(exu_n4408));
AND2X1 exu_U17938(.A(div_d_mux_n501), .B(exu_n10777), .Y(div_dnext[101]));
INVX1 exu_U17939(.A(div_dnext[101]), .Y(exu_n4409));
AND2X1 exu_U17940(.A(div_adder_out[37]), .B(exu_n16250), .Y(div_d_mux_n503));
INVX1 exu_U17941(.A(div_d_mux_n503), .Y(exu_n4410));
AND2X1 exu_U17942(.A(div_d_mux_n505), .B(exu_n10778), .Y(div_dnext[100]));
INVX1 exu_U17943(.A(div_dnext[100]), .Y(exu_n4411));
AND2X1 exu_U17944(.A(div_adder_out[36]), .B(exu_n16250), .Y(div_d_mux_n507));
INVX1 exu_U17945(.A(div_d_mux_n507), .Y(exu_n4412));
AND2X1 exu_U17946(.A(div_d_mux_n509), .B(exu_n10517), .Y(div_dnext[0]));
INVX1 exu_U17947(.A(div_dnext[0]), .Y(exu_n4413));
AND2X1 exu_U17948(.A(ecl_div_newq), .B(ecl_div_sel_adder), .Y(div_d_mux_n511));
INVX1 exu_U17949(.A(div_d_mux_n511), .Y(exu_n4414));
OR2X1 exu_U17950(.A(exu_n12002), .B(exu_n14890), .Y(div_low32or_n7));
INVX1 exu_U17951(.A(div_low32or_n7), .Y(exu_n4415));
OR2X1 exu_U17952(.A(exu_n12000), .B(exu_n14888), .Y(div_low32or_n9));
INVX1 exu_U17953(.A(div_low32or_n9), .Y(exu_n4416));
OR2X1 exu_U17954(.A(exu_n12057), .B(exu_n14951), .Y(div_low32or_n3));
INVX1 exu_U17955(.A(div_low32or_n3), .Y(exu_n4417));
OR2X1 exu_U17956(.A(exu_n12006), .B(exu_n14894), .Y(div_low32or_n13));
INVX1 exu_U17957(.A(div_low32or_n13), .Y(exu_n4418));
OR2X1 exu_U17958(.A(exu_n12004), .B(exu_n14892), .Y(div_low32or_n15));
INVX1 exu_U17959(.A(div_low32or_n15), .Y(exu_n4419));
OR2X1 exu_U17960(.A(exu_n11994), .B(exu_n15352), .Y(div_low32or_n21));
INVX1 exu_U17961(.A(div_low32or_n21), .Y(exu_n4420));
OR2X1 exu_U17962(.A(exu_n11992), .B(exu_n14881), .Y(div_low32or_n23));
INVX1 exu_U17963(.A(div_low32or_n23), .Y(exu_n4421));
OR2X1 exu_U17964(.A(exu_n12059), .B(exu_n14953), .Y(div_low32or_n17));
INVX1 exu_U17965(.A(div_low32or_n17), .Y(exu_n4422));
OR2X1 exu_U17966(.A(exu_n11998), .B(exu_n14886), .Y(div_low32or_n27));
INVX1 exu_U17967(.A(div_low32or_n27), .Y(exu_n4423));
OR2X1 exu_U17968(.A(exu_n11996), .B(exu_n14884), .Y(div_low32or_n29));
INVX1 exu_U17969(.A(div_low32or_n29), .Y(exu_n4424));
AND2X1 exu_U17970(.A(exu_n16154), .B(exu_n15350), .Y(shft_mux_rshift_extend_n2));
INVX1 exu_U17971(.A(shft_mux_rshift_extend_n2), .Y(exu_n4425));
INVX1 exu_U17972(.A(exu_n4428), .Y(exu_n4426));
INVX1 exu_U17973(.A(exu_n4426), .Y(exu_n4427));
AND2X1 exu_U17974(.A(ecl_shft_extend32bit_e_l), .B(exu_n16152), .Y(shft_mux_rshift_extend_n4));
INVX1 exu_U17975(.A(shft_mux_rshift_extend_n4), .Y(exu_n4428));
INVX1 exu_U17976(.A(exu_n4431), .Y(exu_n4429));
INVX1 exu_U17977(.A(exu_n4429), .Y(exu_n4430));
AND2X1 exu_U17978(.A(exu_n15984), .B(exu_n16152), .Y(shft_mux_rshift_extend_n6));
INVX1 exu_U17979(.A(shft_mux_rshift_extend_n6), .Y(exu_n4431));
INVX1 exu_U17980(.A(exu_n4434), .Y(exu_n4432));
INVX1 exu_U17981(.A(exu_n4432), .Y(exu_n4433));
AND2X1 exu_U17982(.A(ecl_shft_extend32bit_e_l), .B(exu_n16152), .Y(shft_mux_rshift_extend_n8));
INVX1 exu_U17983(.A(shft_mux_rshift_extend_n8), .Y(exu_n4434));
INVX1 exu_U17984(.A(exu_n4437), .Y(exu_n4435));
INVX1 exu_U17985(.A(exu_n4435), .Y(exu_n4436));
AND2X1 exu_U17986(.A(exu_n15350), .B(exu_n16152), .Y(shft_mux_rshift_extend_n10));
INVX1 exu_U17987(.A(shft_mux_rshift_extend_n10), .Y(exu_n4437));
INVX1 exu_U17988(.A(exu_n4440), .Y(exu_n4438));
INVX1 exu_U17989(.A(exu_n4438), .Y(exu_n4439));
AND2X1 exu_U17990(.A(ecl_shft_extend32bit_e_l), .B(exu_n16152), .Y(shft_mux_rshift_extend_n12));
INVX1 exu_U17991(.A(shft_mux_rshift_extend_n12), .Y(exu_n4440));
INVX1 exu_U17992(.A(exu_n4443), .Y(exu_n4441));
INVX1 exu_U17993(.A(exu_n4441), .Y(exu_n4442));
AND2X1 exu_U17994(.A(exu_n15350), .B(exu_n16152), .Y(shft_mux_rshift_extend_n14));
INVX1 exu_U17995(.A(shft_mux_rshift_extend_n14), .Y(exu_n4443));
INVX1 exu_U17996(.A(exu_n4446), .Y(exu_n4444));
INVX1 exu_U17997(.A(exu_n4444), .Y(exu_n4445));
AND2X1 exu_U17998(.A(exu_n15984), .B(exu_n16153), .Y(shft_mux_rshift_extend_n16));
INVX1 exu_U17999(.A(shft_mux_rshift_extend_n16), .Y(exu_n4446));
INVX1 exu_U18000(.A(exu_n4449), .Y(exu_n4447));
INVX1 exu_U18001(.A(exu_n4447), .Y(exu_n4448));
AND2X1 exu_U18002(.A(exu_n15983), .B(exu_n16152), .Y(shft_mux_rshift_extend_n18));
INVX1 exu_U18003(.A(shft_mux_rshift_extend_n18), .Y(exu_n4449));
INVX1 exu_U18004(.A(exu_n4452), .Y(exu_n4450));
INVX1 exu_U18005(.A(exu_n4450), .Y(exu_n4451));
AND2X1 exu_U18006(.A(ecl_shft_extend32bit_e_l), .B(exu_n16152), .Y(shft_mux_rshift_extend_n20));
INVX1 exu_U18007(.A(shft_mux_rshift_extend_n20), .Y(exu_n4452));
INVX1 exu_U18008(.A(exu_n4455), .Y(exu_n4453));
INVX1 exu_U18009(.A(exu_n4453), .Y(exu_n4454));
AND2X1 exu_U18010(.A(exu_n15983), .B(exu_n16152), .Y(shft_mux_rshift_extend_n22));
INVX1 exu_U18011(.A(shft_mux_rshift_extend_n22), .Y(exu_n4455));
AND2X1 exu_U18012(.A(exu_n15983), .B(exu_n16152), .Y(shft_mux_rshift_extend_n24));
INVX1 exu_U18013(.A(shft_mux_rshift_extend_n24), .Y(exu_n4456));
INVX1 exu_U18014(.A(exu_n4459), .Y(exu_n4457));
INVX1 exu_U18015(.A(exu_n4457), .Y(exu_n4458));
AND2X1 exu_U18016(.A(exu_n15983), .B(exu_n16152), .Y(shft_mux_rshift_extend_n30));
INVX1 exu_U18017(.A(shft_mux_rshift_extend_n30), .Y(exu_n4459));
INVX1 exu_U18018(.A(exu_n4462), .Y(exu_n4460));
INVX1 exu_U18019(.A(exu_n4460), .Y(exu_n4461));
AND2X1 exu_U18020(.A(exu_n15350), .B(exu_n16153), .Y(shft_mux_rshift_extend_n42));
INVX1 exu_U18021(.A(shft_mux_rshift_extend_n42), .Y(exu_n4462));
INVX1 exu_U18022(.A(exu_n4465), .Y(exu_n4463));
INVX1 exu_U18023(.A(exu_n4463), .Y(exu_n4464));
AND2X1 exu_U18024(.A(exu_n15984), .B(exu_n16153), .Y(shft_mux_rshift_extend_n52));
INVX1 exu_U18025(.A(shft_mux_rshift_extend_n52), .Y(exu_n4465));
INVX1 exu_U18026(.A(exu_n4468), .Y(exu_n4466));
INVX1 exu_U18027(.A(exu_n4466), .Y(exu_n4467));
AND2X1 exu_U18028(.A(exu_n15984), .B(exu_n16153), .Y(shft_mux_rshift_extend_n54));
INVX1 exu_U18029(.A(shft_mux_rshift_extend_n54), .Y(exu_n4468));
INVX1 exu_U18030(.A(exu_n4471), .Y(exu_n4469));
INVX1 exu_U18031(.A(exu_n4469), .Y(exu_n4470));
AND2X1 exu_U18032(.A(exu_n15984), .B(exu_n16153), .Y(shft_mux_rshift_extend_n56));
INVX1 exu_U18033(.A(shft_mux_rshift_extend_n56), .Y(exu_n4471));
INVX1 exu_U18034(.A(exu_n4474), .Y(exu_n4472));
INVX1 exu_U18035(.A(exu_n4472), .Y(exu_n4473));
AND2X1 exu_U18036(.A(exu_n15984), .B(exu_n16153), .Y(shft_mux_rshift_extend_n58));
INVX1 exu_U18037(.A(shft_mux_rshift_extend_n58), .Y(exu_n4474));
INVX1 exu_U18038(.A(exu_n4477), .Y(exu_n4475));
INVX1 exu_U18039(.A(exu_n4475), .Y(exu_n4476));
AND2X1 exu_U18040(.A(exu_n15984), .B(exu_n16153), .Y(shft_mux_rshift_extend_n60));
INVX1 exu_U18041(.A(shft_mux_rshift_extend_n60), .Y(exu_n4477));
INVX1 exu_U18042(.A(exu_n4480), .Y(exu_n4478));
INVX1 exu_U18043(.A(exu_n4478), .Y(exu_n4479));
AND2X1 exu_U18044(.A(exu_n15984), .B(exu_n16154), .Y(shft_mux_rshift_extend_n62));
INVX1 exu_U18045(.A(shft_mux_rshift_extend_n62), .Y(exu_n4480));
INVX1 exu_U18046(.A(exu_n4483), .Y(exu_n4481));
INVX1 exu_U18047(.A(exu_n4481), .Y(exu_n4482));
AND2X1 exu_U18048(.A(exu_n15983), .B(exu_n16152), .Y(shft_mux_rshift_extend_n64));
INVX1 exu_U18049(.A(shft_mux_rshift_extend_n64), .Y(exu_n4483));
OR2X1 exu_U18050(.A(exu_n12062), .B(exu_n14954), .Y(alu_ecl_mem_addr_invalid_e_l));
INVX1 exu_U18051(.A(alu_ecl_mem_addr_invalid_e_l), .Y(exu_n4484));
OR2X1 exu_U18052(.A(exu_n12061), .B(exu_n14956), .Y(alu_chk_mem_addr_n3));
INVX1 exu_U18053(.A(alu_chk_mem_addr_n3), .Y(exu_n4485));
OR2X1 exu_U18054(.A(exu_n12064), .B(exu_n14958), .Y(alu_chk_mem_addr_n17));
INVX1 exu_U18055(.A(alu_chk_mem_addr_n17), .Y(exu_n4486));
AND2X1 exu_U18056(.A(ecl_mdqctl_n13), .B(exu_n10518), .Y(ecl_mdqctl_n12));
INVX1 exu_U18057(.A(ecl_mdqctl_n12), .Y(exu_n4487));
AND2X1 exu_U18058(.A(exu_n15379), .B(ecl_mdqctl_n17), .Y(ecl_mdqctl_mul_ready_next));
INVX1 exu_U18059(.A(ecl_mdqctl_mul_ready_next), .Y(exu_n4488));
OR2X1 exu_U18060(.A(exu_n12065), .B(exu_n14959), .Y(ecl_mdqctl_mul_done_ack));
INVX1 exu_U18061(.A(ecl_mdqctl_mul_done_ack), .Y(exu_n4489));
AND2X1 exu_U18062(.A(exu_n11650), .B(exu_n10520), .Y(ecl_mdqctl_mul_data_next[9]));
INVX1 exu_U18063(.A(ecl_mdqctl_mul_data_next[9]), .Y(exu_n4490));
AND2X1 exu_U18064(.A(exu_n11651), .B(exu_n10521), .Y(ecl_mdqctl_mul_data_next[8]));
INVX1 exu_U18065(.A(ecl_mdqctl_mul_data_next[8]), .Y(exu_n4491));
AND2X1 exu_U18066(.A(exu_n11652), .B(exu_n10522), .Y(ecl_mdqctl_mul_data_next[7]));
INVX1 exu_U18067(.A(ecl_mdqctl_mul_data_next[7]), .Y(exu_n4492));
AND2X1 exu_U18068(.A(exu_n11653), .B(exu_n10523), .Y(ecl_mdqctl_mul_data_next[6]));
INVX1 exu_U18069(.A(ecl_mdqctl_mul_data_next[6]), .Y(exu_n4493));
AND2X1 exu_U18070(.A(exu_n11654), .B(exu_n10524), .Y(ecl_mdqctl_mul_data_next[5]));
INVX1 exu_U18071(.A(ecl_mdqctl_mul_data_next[5]), .Y(exu_n4494));
AND2X1 exu_U18072(.A(exu_n11655), .B(exu_n10525), .Y(ecl_mdqctl_mul_data_next[4]));
INVX1 exu_U18073(.A(ecl_mdqctl_mul_data_next[4]), .Y(exu_n4495));
AND2X1 exu_U18074(.A(exu_n11656), .B(exu_n10526), .Y(ecl_mdqctl_mul_data_next[3]));
INVX1 exu_U18075(.A(ecl_mdqctl_mul_data_next[3]), .Y(exu_n4496));
AND2X1 exu_U18076(.A(exu_n11657), .B(exu_n10527), .Y(ecl_mdqctl_mul_data_next[2]));
INVX1 exu_U18077(.A(ecl_mdqctl_mul_data_next[2]), .Y(exu_n4497));
AND2X1 exu_U18078(.A(exu_n11658), .B(exu_n10528), .Y(ecl_mdqctl_mul_data_next[1]));
INVX1 exu_U18079(.A(ecl_mdqctl_mul_data_next[1]), .Y(exu_n4498));
AND2X1 exu_U18080(.A(exu_n11659), .B(exu_n10529), .Y(ecl_mdqctl_mul_data_next[0]));
INVX1 exu_U18081(.A(ecl_mdqctl_mul_data_next[0]), .Y(exu_n4499));
OR2X1 exu_U18082(.A(exu_n12066), .B(exu_n14960), .Y(ecl_mdqctl_div_zero_e));
INVX1 exu_U18083(.A(ecl_mdqctl_div_zero_e), .Y(exu_n4500));
AND2X1 exu_U18084(.A(exu_n11663), .B(ecl_mdqctl_n61), .Y(ecl_mdqctl_n59));
INVX1 exu_U18085(.A(ecl_mdqctl_n59), .Y(exu_n4501));
OR2X1 exu_U18086(.A(exu_n16257), .B(ecl_divcntl_n24), .Y(ecl_divcntl_next_state[3]));
INVX1 exu_U18087(.A(ecl_divcntl_next_state[3]), .Y(exu_n4502));
OR2X1 exu_U18088(.A(ecl_divcntl_n24), .B(exu_n14961), .Y(ecl_divcntl_next_state[2]));
INVX1 exu_U18089(.A(ecl_divcntl_next_state[2]), .Y(exu_n4503));
AND2X1 exu_U18090(.A(ecl_divcntl_n35), .B(exu_n15815), .Y(ecl_divcntl_next_state[0]));
INVX1 exu_U18091(.A(ecl_divcntl_next_state[0]), .Y(exu_n4504));
AND2X1 exu_U18092(.A(ecl_divcntl_div_state_0), .B(exu_n16218), .Y(ecl_divcntl_n36));
INVX1 exu_U18093(.A(ecl_divcntl_n36), .Y(exu_n4505));
AND2X1 exu_U18094(.A(exu_n11667), .B(exu_n10531), .Y(ecl_divcntl_next_muls_v));
INVX1 exu_U18095(.A(ecl_divcntl_next_muls_v), .Y(exu_n4506));
AND2X1 exu_U18096(.A(exu_n11668), .B(exu_n10534), .Y(ecl_divcntl_next_muls_c));
INVX1 exu_U18097(.A(ecl_divcntl_next_muls_c), .Y(exu_n4507));
OR2X1 exu_U18098(.A(ecl_divcntl_n50), .B(exu_n16508), .Y(ecl_divcntl_last_cin_next));
INVX1 exu_U18099(.A(ecl_divcntl_last_cin_next), .Y(exu_n4508));
AND2X1 exu_U18100(.A(div_ecl_d_62), .B(exu_n15424), .Y(ecl_divcntl_n55));
INVX1 exu_U18101(.A(ecl_divcntl_n55), .Y(exu_n4509));
AND2X1 exu_U18102(.A(exu_n16257), .B(exu_n16438), .Y(ecl_divcntl_n62));
INVX1 exu_U18103(.A(ecl_divcntl_n62), .Y(exu_n4510));
AND2X1 exu_U18104(.A(ecl_divcntl_last_cin), .B(ecl_div_last_cycle), .Y(ecl_divcntl_n63));
INVX1 exu_U18105(.A(ecl_divcntl_n63), .Y(exu_n4511));
OR2X1 exu_U18106(.A(exu_n16508), .B(exu_n16252), .Y(ecl_divcntl_n77));
INVX1 exu_U18107(.A(ecl_divcntl_n77), .Y(exu_n4512));
OR2X1 exu_U18108(.A(exu_n16246), .B(exu_n15394), .Y(ecl_divcntl_n82));
INVX1 exu_U18109(.A(ecl_divcntl_n82), .Y(exu_n4513));
OR2X1 exu_U18110(.A(exu_n15221), .B(ecl_div_sel_64b), .Y(ecl_divcntl_n83));
INVX1 exu_U18111(.A(ecl_divcntl_n83), .Y(exu_n4514));
AND2X1 exu_U18112(.A(ecl_divcntl_n84), .B(ecl_divcntl_muls_v), .Y(ecl_divcntl_n81));
INVX1 exu_U18113(.A(ecl_divcntl_n81), .Y(exu_n4515));
AND2X1 exu_U18114(.A(ecl_byplog_rs2_n29), .B(exu_n10535), .Y(ecl_byplog_rs2_n16));
INVX1 exu_U18115(.A(ecl_byplog_rs2_n16), .Y(exu_n4516));
OR2X1 exu_U18116(.A(ifu_exu_useimm_d), .B(sehold), .Y(ecl_byplog_rs2_n47));
INVX1 exu_U18117(.A(ecl_byplog_rs2_n47), .Y(exu_n4517));
AND2X1 exu_U18118(.A(ecl_byplog_rs1_n20), .B(ecl_byplog_rs1_n19), .Y(ecl_byplog_rs1_n18));
INVX1 exu_U18119(.A(ecl_byplog_rs1_n18), .Y(exu_n4518));
OR2X1 exu_U18120(.A(ifu_exu_dbrinst_d), .B(sehold), .Y(ecl_byplog_rs1_n25));
INVX1 exu_U18121(.A(ecl_byplog_rs1_n25), .Y(exu_n4519));
OR2X1 exu_U18122(.A(ecl_ifu_exu_rs1_d[1]), .B(ecl_ifu_exu_rs1_d[0]), .Y(ecl_byplog_rs1_n39));
INVX1 exu_U18123(.A(ecl_byplog_rs1_n39), .Y(exu_n4520));
AND2X1 exu_U18124(.A(ecl_eccctl_n18), .B(exu_n10540), .Y(ecl_eccctl_flag_ecc_ue_e));
INVX1 exu_U18125(.A(ecl_eccctl_flag_ecc_ue_e), .Y(exu_n4521));
AND2X1 exu_U18126(.A(ifu_exu_disable_ce_e), .B(exu_n15373), .Y(ecl_eccctl_n20));
INVX1 exu_U18127(.A(ecl_eccctl_n20), .Y(exu_n4522));
OR2X1 exu_U18128(.A(ecl_eccctl_n21), .B(ifu_exu_disable_ce_e), .Y(ecl_eccctl_flag_ecc_ce_e));
INVX1 exu_U18129(.A(ecl_eccctl_flag_ecc_ce_e), .Y(exu_n4523));
AND2X1 exu_U18130(.A(exu_n16593), .B(exu_n10543), .Y(ecl_eccctl_n31));
INVX1 exu_U18131(.A(ecl_eccctl_n31), .Y(exu_n4524));
AND2X1 exu_U18132(.A(exu_n11676), .B(exu_n10544), .Y(ecl_writeback_wen_no_inst_vld_m));
INVX1 exu_U18133(.A(ecl_writeback_wen_no_inst_vld_m), .Y(exu_n4525));
OR2X1 exu_U18134(.A(exu_n12067), .B(exu_n14962), .Y(ecl_writeback_vld_restore_e));
INVX1 exu_U18135(.A(ecl_writeback_vld_restore_e), .Y(exu_n4526));
OR2X1 exu_U18136(.A(exu_n15030), .B(ecl_writeback_return_e), .Y(ecl_writeback_n61));
INVX1 exu_U18137(.A(ecl_writeback_n61), .Y(exu_n4527));
OR2X1 exu_U18138(.A(sehold), .B(rml_ecl_kill_m), .Y(ecl_writeback_n62));
INVX1 exu_U18139(.A(ecl_writeback_n62), .Y(exu_n4528));
OR2X1 exu_U18140(.A(exu_n12068), .B(exu_n14963), .Y(ecl_writeback_valid_e));
INVX1 exu_U18141(.A(ecl_writeback_valid_e), .Y(exu_n4529));
OR2X1 exu_U18142(.A(ecl_writeback_n50), .B(exu_n15238), .Y(ecl_writeback_restore_ready_next));
INVX1 exu_U18143(.A(ecl_writeback_restore_ready_next), .Y(exu_n4530));
AND2X1 exu_U18144(.A(ecl_writeback_n89), .B(exu_n10545), .Y(ecl_writeback_n88));
INVX1 exu_U18145(.A(ecl_writeback_n88), .Y(exu_n4531));
OR2X1 exu_U18146(.A(sehold), .B(exu_n16273), .Y(ecl_writeback_inst_vld_noflush_wen_m));
INVX1 exu_U18147(.A(ecl_writeback_inst_vld_noflush_wen_m), .Y(exu_n4532));
AND2X1 exu_U18148(.A(exu_n15921), .B(exu_n15687), .Y(ecl_writeback_n99));
INVX1 exu_U18149(.A(ecl_writeback_n99), .Y(exu_n4533));
AND2X1 exu_U18150(.A(exu_n15922), .B(exu_n15687), .Y(ecl_writeback_n107));
INVX1 exu_U18151(.A(ecl_writeback_n107), .Y(exu_n4534));
AND2X1 exu_U18152(.A(exu_n15923), .B(exu_n15687), .Y(ecl_writeback_n115));
INVX1 exu_U18153(.A(ecl_writeback_n115), .Y(exu_n4535));
AND2X1 exu_U18154(.A(ecl_mdqctl_wb_divthr_g[0]), .B(exu_n16193), .Y(ecl_writeback_n122));
INVX1 exu_U18155(.A(ecl_writeback_n122), .Y(exu_n4536));
AND2X1 exu_U18156(.A(ecl_mdqctl_wb_divthr_g[1]), .B(exu_n16195), .Y(ecl_writeback_n124));
INVX1 exu_U18157(.A(ecl_writeback_n124), .Y(exu_n4537));
AND2X1 exu_U18158(.A(exu_n15924), .B(exu_n15687), .Y(ecl_writeback_n126));
INVX1 exu_U18159(.A(ecl_writeback_n126), .Y(exu_n4538));
OR2X1 exu_U18160(.A(ecl_writeback_n131), .B(exu_n14971), .Y(ecl_rml_wstate_wen_w));
INVX1 exu_U18161(.A(ecl_rml_wstate_wen_w), .Y(exu_n4539));
OR2X1 exu_U18162(.A(ecl_writeback_sraddr_e[2]), .B(ecl_writeback_sraddr_e[1]), .Y(ecl_writeback_n138));
INVX1 exu_U18163(.A(ecl_writeback_n138), .Y(exu_n4540));
OR2X1 exu_U18164(.A(ecl_writeback_sraddr_w[6]), .B(ecl_writeback_sraddr_w[4]), .Y(ecl_writeback_n145));
INVX1 exu_U18165(.A(ecl_writeback_n145), .Y(exu_n4541));
AND2X1 exu_U18166(.A(exu_n11683), .B(exu_n10551), .Y(ecl_writeback_ecl_irf_wen_g));
INVX1 exu_U18167(.A(ecl_writeback_ecl_irf_wen_g), .Y(exu_n4542));
OR2X1 exu_U18168(.A(lsu_exu_ldst_miss_g2), .B(exu_n14973), .Y(ecl_writeback_n155));
INVX1 exu_U18169(.A(ecl_writeback_n155), .Y(exu_n4543));
AND2X1 exu_U18170(.A(ecl_writeback_n129), .B(exu_n15482), .Y(ecl_writeback_n160));
INVX1 exu_U18171(.A(ecl_writeback_n160), .Y(exu_n4544));
OR2X1 exu_U18172(.A(ecl_tid_w1[1]), .B(ecl_tid_w1[0]), .Y(ecl_writeback_n183));
INVX1 exu_U18173(.A(ecl_writeback_n183), .Y(exu_n4545));
OR2X1 exu_U18174(.A(ecl_mdqctl_wb_divthr_g[0]), .B(exu_n16507), .Y(ecl_writeback_n193));
INVX1 exu_U18175(.A(ecl_writeback_n193), .Y(exu_n4546));
OR2X1 exu_U18176(.A(ecl_mdqctl_wb_divthr_g[1]), .B(exu_n16506), .Y(ecl_writeback_n194));
INVX1 exu_U18177(.A(ecl_writeback_n194), .Y(exu_n4547));
OR2X1 exu_U18178(.A(ecl_mdqctl_wb_divthr_g[1]), .B(ecl_mdqctl_wb_divthr_g[0]), .Y(ecl_writeback_n195));
INVX1 exu_U18179(.A(ecl_writeback_n195), .Y(exu_n4548));
AND2X1 exu_U18180(.A(exu_n15765), .B(exu_n10554), .Y(ecl_writeback_n196));
INVX1 exu_U18181(.A(ecl_writeback_n196), .Y(exu_n4549));
OR2X1 exu_U18182(.A(ecl_writeback_wen_no_inst_vld_w), .B(ecl_writeback_wb_w), .Y(ecl_writeback_n200));
INVX1 exu_U18183(.A(ecl_writeback_n200), .Y(exu_n4550));
OR2X1 exu_U18184(.A(ecl_ccr_n25), .B(ecl_ccr_n26), .Y(ecl_ccr_n21));
INVX1 exu_U18185(.A(ecl_ccr_n21), .Y(exu_n4551));
AND2X1 exu_U18186(.A(ecl_rml_thr_w[3]), .B(exu_n15926), .Y(ecl_ccr_n27));
INVX1 exu_U18187(.A(ecl_ccr_n27), .Y(exu_n4552));
OR2X1 exu_U18188(.A(ecl_ccr_thr_w2[0]), .B(exu_n16584), .Y(ecl_ccr_n30));
INVX1 exu_U18189(.A(ecl_ccr_n30), .Y(exu_n4553));
AND2X1 exu_U18190(.A(ecl_rml_thr_w[2]), .B(exu_n15926), .Y(ecl_ccr_n29));
INVX1 exu_U18191(.A(ecl_ccr_n29), .Y(exu_n4554));
OR2X1 exu_U18192(.A(ecl_ccr_thr_w2[1]), .B(exu_n16584), .Y(ecl_ccr_n32));
INVX1 exu_U18193(.A(ecl_ccr_n32), .Y(exu_n4555));
AND2X1 exu_U18194(.A(exu_n15958), .B(exu_n15926), .Y(ecl_ccr_n31));
INVX1 exu_U18195(.A(ecl_ccr_n31), .Y(exu_n4556));
OR2X1 exu_U18196(.A(ecl_ccr_thr_w2[1]), .B(ecl_ccr_thr_w2[0]), .Y(ecl_ccr_n34));
INVX1 exu_U18197(.A(ecl_ccr_n34), .Y(exu_n4557));
AND2X1 exu_U18198(.A(exu_n15960), .B(exu_n15926), .Y(ecl_ccr_n33));
INVX1 exu_U18199(.A(ecl_ccr_n33), .Y(exu_n4558));
AND2X1 exu_U18200(.A(exu_n15338), .B(ecl_ccr_n40), .Y(ecl_ccr_n38));
INVX1 exu_U18201(.A(ecl_ccr_n38), .Y(exu_n4559));
AND2X1 exu_U18202(.A(ecl_alu_xcc_e[2]), .B(ecl_ccr_n40), .Y(ecl_ccr_n41));
INVX1 exu_U18203(.A(ecl_ccr_n41), .Y(exu_n4560));
AND2X1 exu_U18204(.A(ecl_adder_xcc[1]), .B(ecl_ccr_n40), .Y(ecl_ccr_n43));
INVX1 exu_U18205(.A(ecl_ccr_n43), .Y(exu_n4561));
AND2X1 exu_U18206(.A(ecl_adder_xcc[0]), .B(ecl_ccr_n40), .Y(ecl_ccr_n45));
INVX1 exu_U18207(.A(ecl_ccr_n45), .Y(exu_n4562));
AND2X1 exu_U18208(.A(exu_n15339), .B(ecl_ccr_n40), .Y(ecl_ccr_n47));
INVX1 exu_U18209(.A(ecl_ccr_n47), .Y(exu_n4563));
AND2X1 exu_U18210(.A(exu_n15426), .B(ecl_ccr_n40), .Y(ecl_ccr_n49));
INVX1 exu_U18211(.A(ecl_ccr_n49), .Y(exu_n4564));
AND2X1 exu_U18212(.A(ecl_adder_icc[1]), .B(ecl_ccr_n40), .Y(ecl_ccr_n51));
INVX1 exu_U18213(.A(ecl_ccr_n51), .Y(exu_n4565));
AND2X1 exu_U18214(.A(ecl_adder_icc[0]), .B(ecl_ccr_n40), .Y(ecl_ccr_n53));
INVX1 exu_U18215(.A(ecl_ccr_n53), .Y(exu_n4566));
AND2X1 exu_U18216(.A(exu_ifu_brpc_e[7]), .B(ifu_exu_tcc_e), .Y(ecl_ttype_mux_n7));
INVX1 exu_U18217(.A(ecl_ttype_mux_n7), .Y(exu_n4567));
AND2X1 exu_U18218(.A(exu_ifu_brpc_e[6]), .B(ifu_exu_tcc_e), .Y(ecl_ttype_mux_n11));
INVX1 exu_U18219(.A(ecl_ttype_mux_n11), .Y(exu_n4568));
AND2X1 exu_U18220(.A(ecl_ttype_mux_n13), .B(ecl_pick_not_aligned), .Y(ecl_early2_ttype_e[5]));
INVX1 exu_U18221(.A(ecl_early2_ttype_e[5]), .Y(exu_n4569));
AND2X1 exu_U18222(.A(exu_ifu_brpc_e[5]), .B(ifu_exu_tcc_e), .Y(ecl_ttype_mux_n15));
INVX1 exu_U18223(.A(ecl_ttype_mux_n15), .Y(exu_n4570));
AND2X1 exu_U18224(.A(ecl_ttype_mux_n17), .B(ecl_pick_not_aligned), .Y(ecl_early2_ttype_e[4]));
INVX1 exu_U18225(.A(ecl_early2_ttype_e[4]), .Y(exu_n4571));
AND2X1 exu_U18226(.A(exu_ifu_brpc_e[4]), .B(ifu_exu_tcc_e), .Y(ecl_ttype_mux_n19));
INVX1 exu_U18227(.A(ecl_ttype_mux_n19), .Y(exu_n4572));
AND2X1 exu_U18228(.A(exu_ifu_brpc_e[3]), .B(ifu_exu_tcc_e), .Y(ecl_ttype_mux_n23));
INVX1 exu_U18229(.A(ecl_ttype_mux_n23), .Y(exu_n4573));
AND2X1 exu_U18230(.A(ecl_ttype_mux_n25), .B(ecl_pick_not_aligned), .Y(ecl_early2_ttype_e[2]));
INVX1 exu_U18231(.A(ecl_early2_ttype_e[2]), .Y(exu_n4574));
AND2X1 exu_U18232(.A(exu_ifu_brpc_e[2]), .B(ifu_exu_tcc_e), .Y(ecl_ttype_mux_n27));
INVX1 exu_U18233(.A(ecl_ttype_mux_n27), .Y(exu_n4575));
AND2X1 exu_U18234(.A(exu_ifu_brpc_e[1]), .B(ifu_exu_tcc_e), .Y(ecl_ttype_mux_n31));
INVX1 exu_U18235(.A(ecl_ttype_mux_n31), .Y(exu_n4576));
AND2X1 exu_U18236(.A(exu_ifu_brpc_e[0]), .B(ifu_exu_tcc_e), .Y(ecl_ttype_mux_n35));
INVX1 exu_U18237(.A(ecl_ttype_mux_n35), .Y(exu_n4577));
AND2X1 exu_U18238(.A(ecl_thr_d[3]), .B(div_yreg_div_ecl_yreg_0[3]), .Y(ecl_yreg0_mux_n3));
INVX1 exu_U18239(.A(ecl_yreg0_mux_n3), .Y(exu_n4578));
AND2X1 exu_U18240(.A(exu_n15934), .B(div_yreg_div_ecl_yreg_0[1]), .Y(ecl_yreg0_mux_n5));
INVX1 exu_U18241(.A(ecl_yreg0_mux_n5), .Y(exu_n4579));
AND2X1 exu_U18242(.A(exu_n15974), .B(ecc_rs2_err_m[6]), .Y(ecc_syn_mux_n3));
INVX1 exu_U18243(.A(ecc_syn_mux_n3), .Y(exu_n4580));
AND2X1 exu_U18244(.A(ecc_rs2_err_m[5]), .B(exu_n15974), .Y(ecc_syn_mux_n7));
INVX1 exu_U18245(.A(ecc_syn_mux_n7), .Y(exu_n4581));
AND2X1 exu_U18246(.A(ecc_rs2_err_m[4]), .B(ecl_ecc_sel_rs2_m_l), .Y(ecc_syn_mux_n11));
INVX1 exu_U18247(.A(ecc_syn_mux_n11), .Y(exu_n4582));
AND2X1 exu_U18248(.A(ecc_rs2_err_m[3]), .B(exu_n15974), .Y(ecc_syn_mux_n15));
INVX1 exu_U18249(.A(ecc_syn_mux_n15), .Y(exu_n4583));
AND2X1 exu_U18250(.A(ecc_rs2_err_m[2]), .B(ecl_ecc_sel_rs2_m_l), .Y(ecc_syn_mux_n19));
INVX1 exu_U18251(.A(ecc_syn_mux_n19), .Y(exu_n4584));
AND2X1 exu_U18252(.A(ecc_rs2_err_m[1]), .B(exu_n15974), .Y(ecc_syn_mux_n23));
INVX1 exu_U18253(.A(ecc_syn_mux_n23), .Y(exu_n4585));
AND2X1 exu_U18254(.A(ecc_rs2_err_m[0]), .B(ecl_ecc_sel_rs2_m_l), .Y(ecc_syn_mux_n27));
INVX1 exu_U18255(.A(ecc_syn_mux_n27), .Y(exu_n4586));
AND2X1 exu_U18256(.A(exu_n11690), .B(ecc_chk_rs1_n6), .Y(ecc_chk_rs1_n3));
INVX1 exu_U18257(.A(ecc_chk_rs1_n3), .Y(exu_n4587));
OR2X1 exu_U18258(.A(ecc_rs1_err_e[4]), .B(ecc_rs1_err_e[3]), .Y(ecc_chk_rs1_n7));
INVX1 exu_U18259(.A(ecc_chk_rs1_n7), .Y(exu_n4588));
AND2X1 exu_U18260(.A(exu_n16285), .B(byp_irf_rd_data_w[9]), .Y(bypass_mux_rs3h_data_1_n5));
INVX1 exu_U18261(.A(bypass_mux_rs3h_data_1_n5), .Y(exu_n4589));
AND2X1 exu_U18262(.A(byp_irf_rd_data_w[8]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n11));
INVX1 exu_U18263(.A(bypass_mux_rs3h_data_1_n11), .Y(exu_n4590));
AND2X1 exu_U18264(.A(byp_irf_rd_data_w[7]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n17));
INVX1 exu_U18265(.A(bypass_mux_rs3h_data_1_n17), .Y(exu_n4591));
AND2X1 exu_U18266(.A(byp_irf_rd_data_w[6]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n23));
INVX1 exu_U18267(.A(bypass_mux_rs3h_data_1_n23), .Y(exu_n4592));
AND2X1 exu_U18268(.A(byp_irf_rd_data_w[5]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n29));
INVX1 exu_U18269(.A(bypass_mux_rs3h_data_1_n29), .Y(exu_n4593));
AND2X1 exu_U18270(.A(byp_irf_rd_data_w[4]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n35));
INVX1 exu_U18271(.A(bypass_mux_rs3h_data_1_n35), .Y(exu_n4594));
AND2X1 exu_U18272(.A(byp_irf_rd_data_w[3]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n41));
INVX1 exu_U18273(.A(bypass_mux_rs3h_data_1_n41), .Y(exu_n4595));
AND2X1 exu_U18274(.A(byp_irf_rd_data_w[31]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n47));
INVX1 exu_U18275(.A(bypass_mux_rs3h_data_1_n47), .Y(exu_n4596));
AND2X1 exu_U18276(.A(byp_irf_rd_data_w[30]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n53));
INVX1 exu_U18277(.A(bypass_mux_rs3h_data_1_n53), .Y(exu_n4597));
AND2X1 exu_U18278(.A(byp_irf_rd_data_w[2]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n59));
INVX1 exu_U18279(.A(bypass_mux_rs3h_data_1_n59), .Y(exu_n4598));
AND2X1 exu_U18280(.A(byp_irf_rd_data_w[29]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n65));
INVX1 exu_U18281(.A(bypass_mux_rs3h_data_1_n65), .Y(exu_n4599));
AND2X1 exu_U18282(.A(byp_irf_rd_data_w[28]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n71));
INVX1 exu_U18283(.A(bypass_mux_rs3h_data_1_n71), .Y(exu_n4600));
AND2X1 exu_U18284(.A(byp_irf_rd_data_w[27]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n77));
INVX1 exu_U18285(.A(bypass_mux_rs3h_data_1_n77), .Y(exu_n4601));
AND2X1 exu_U18286(.A(byp_irf_rd_data_w[26]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n83));
INVX1 exu_U18287(.A(bypass_mux_rs3h_data_1_n83), .Y(exu_n4602));
AND2X1 exu_U18288(.A(byp_irf_rd_data_w[25]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n89));
INVX1 exu_U18289(.A(bypass_mux_rs3h_data_1_n89), .Y(exu_n4603));
AND2X1 exu_U18290(.A(byp_irf_rd_data_w[24]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n95));
INVX1 exu_U18291(.A(bypass_mux_rs3h_data_1_n95), .Y(exu_n4604));
AND2X1 exu_U18292(.A(byp_irf_rd_data_w[23]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n101));
INVX1 exu_U18293(.A(bypass_mux_rs3h_data_1_n101), .Y(exu_n4605));
AND2X1 exu_U18294(.A(byp_irf_rd_data_w[22]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n107));
INVX1 exu_U18295(.A(bypass_mux_rs3h_data_1_n107), .Y(exu_n4606));
AND2X1 exu_U18296(.A(byp_irf_rd_data_w[21]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n113));
INVX1 exu_U18297(.A(bypass_mux_rs3h_data_1_n113), .Y(exu_n4607));
AND2X1 exu_U18298(.A(byp_irf_rd_data_w[20]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n119));
INVX1 exu_U18299(.A(bypass_mux_rs3h_data_1_n119), .Y(exu_n4608));
AND2X1 exu_U18300(.A(byp_irf_rd_data_w[1]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n125));
INVX1 exu_U18301(.A(bypass_mux_rs3h_data_1_n125), .Y(exu_n4609));
AND2X1 exu_U18302(.A(byp_irf_rd_data_w[19]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n131));
INVX1 exu_U18303(.A(bypass_mux_rs3h_data_1_n131), .Y(exu_n4610));
AND2X1 exu_U18304(.A(byp_irf_rd_data_w[18]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n137));
INVX1 exu_U18305(.A(bypass_mux_rs3h_data_1_n137), .Y(exu_n4611));
AND2X1 exu_U18306(.A(byp_irf_rd_data_w[17]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n143));
INVX1 exu_U18307(.A(bypass_mux_rs3h_data_1_n143), .Y(exu_n4612));
AND2X1 exu_U18308(.A(byp_irf_rd_data_w[16]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n149));
INVX1 exu_U18309(.A(bypass_mux_rs3h_data_1_n149), .Y(exu_n4613));
AND2X1 exu_U18310(.A(byp_irf_rd_data_w[15]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n155));
INVX1 exu_U18311(.A(bypass_mux_rs3h_data_1_n155), .Y(exu_n4614));
AND2X1 exu_U18312(.A(byp_irf_rd_data_w[14]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n161));
INVX1 exu_U18313(.A(bypass_mux_rs3h_data_1_n161), .Y(exu_n4615));
AND2X1 exu_U18314(.A(byp_irf_rd_data_w[13]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n167));
INVX1 exu_U18315(.A(bypass_mux_rs3h_data_1_n167), .Y(exu_n4616));
AND2X1 exu_U18316(.A(byp_irf_rd_data_w[12]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n173));
INVX1 exu_U18317(.A(bypass_mux_rs3h_data_1_n173), .Y(exu_n4617));
AND2X1 exu_U18318(.A(byp_irf_rd_data_w[11]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n179));
INVX1 exu_U18319(.A(bypass_mux_rs3h_data_1_n179), .Y(exu_n4618));
AND2X1 exu_U18320(.A(byp_irf_rd_data_w[10]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n185));
INVX1 exu_U18321(.A(bypass_mux_rs3h_data_1_n185), .Y(exu_n4619));
AND2X1 exu_U18322(.A(byp_irf_rd_data_w[0]), .B(exu_n16285), .Y(bypass_mux_rs3h_data_1_n191));
INVX1 exu_U18323(.A(bypass_mux_rs3h_data_1_n191), .Y(exu_n4620));
AND2X1 exu_U18324(.A(exu_n16275), .B(bypass_dfill_data_g2[9]), .Y(bypass_rs3h_w2_mux_n3));
INVX1 exu_U18325(.A(bypass_rs3h_w2_mux_n3), .Y(exu_n4621));
AND2X1 exu_U18326(.A(bypass_rs3h_w2_mux_n5), .B(exu_n10556), .Y(bypass_rs3h_data_w2[8]));
INVX1 exu_U18327(.A(bypass_rs3h_data_w2[8]), .Y(exu_n4622));
AND2X1 exu_U18328(.A(bypass_dfill_data_g2[8]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n7));
INVX1 exu_U18329(.A(bypass_rs3h_w2_mux_n7), .Y(exu_n4623));
AND2X1 exu_U18330(.A(bypass_rs3h_w2_mux_n9), .B(exu_n10557), .Y(bypass_rs3h_data_w2[7]));
INVX1 exu_U18331(.A(bypass_rs3h_data_w2[7]), .Y(exu_n4624));
AND2X1 exu_U18332(.A(bypass_dfill_data_g2[7]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n11));
INVX1 exu_U18333(.A(bypass_rs3h_w2_mux_n11), .Y(exu_n4625));
AND2X1 exu_U18334(.A(bypass_rs3h_w2_mux_n13), .B(exu_n10558), .Y(bypass_rs3h_data_w2[6]));
INVX1 exu_U18335(.A(bypass_rs3h_data_w2[6]), .Y(exu_n4626));
AND2X1 exu_U18336(.A(bypass_dfill_data_g2[6]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n15));
INVX1 exu_U18337(.A(bypass_rs3h_w2_mux_n15), .Y(exu_n4627));
AND2X1 exu_U18338(.A(bypass_rs3h_w2_mux_n17), .B(exu_n10559), .Y(bypass_rs3h_data_w2[5]));
INVX1 exu_U18339(.A(bypass_rs3h_data_w2[5]), .Y(exu_n4628));
AND2X1 exu_U18340(.A(bypass_dfill_data_g2[5]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n19));
INVX1 exu_U18341(.A(bypass_rs3h_w2_mux_n19), .Y(exu_n4629));
AND2X1 exu_U18342(.A(bypass_rs3h_w2_mux_n21), .B(exu_n10560), .Y(bypass_rs3h_data_w2[4]));
INVX1 exu_U18343(.A(bypass_rs3h_data_w2[4]), .Y(exu_n4630));
AND2X1 exu_U18344(.A(bypass_dfill_data_g2[4]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n23));
INVX1 exu_U18345(.A(bypass_rs3h_w2_mux_n23), .Y(exu_n4631));
AND2X1 exu_U18346(.A(bypass_rs3h_w2_mux_n25), .B(exu_n10561), .Y(bypass_rs3h_data_w2[3]));
INVX1 exu_U18347(.A(bypass_rs3h_data_w2[3]), .Y(exu_n4632));
AND2X1 exu_U18348(.A(bypass_dfill_data_g2[3]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n27));
INVX1 exu_U18349(.A(bypass_rs3h_w2_mux_n27), .Y(exu_n4633));
AND2X1 exu_U18350(.A(bypass_rs3h_w2_mux_n29), .B(exu_n10562), .Y(bypass_rs3h_data_w2[31]));
INVX1 exu_U18351(.A(bypass_rs3h_data_w2[31]), .Y(exu_n4634));
AND2X1 exu_U18352(.A(bypass_dfill_data_g2[31]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n31));
INVX1 exu_U18353(.A(bypass_rs3h_w2_mux_n31), .Y(exu_n4635));
AND2X1 exu_U18354(.A(bypass_rs3h_w2_mux_n33), .B(exu_n10563), .Y(bypass_rs3h_data_w2[30]));
INVX1 exu_U18355(.A(bypass_rs3h_data_w2[30]), .Y(exu_n4636));
AND2X1 exu_U18356(.A(bypass_dfill_data_g2[30]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n35));
INVX1 exu_U18357(.A(bypass_rs3h_w2_mux_n35), .Y(exu_n4637));
AND2X1 exu_U18358(.A(bypass_rs3h_w2_mux_n37), .B(exu_n10564), .Y(bypass_rs3h_data_w2[2]));
INVX1 exu_U18359(.A(bypass_rs3h_data_w2[2]), .Y(exu_n4638));
AND2X1 exu_U18360(.A(bypass_dfill_data_g2[2]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n39));
INVX1 exu_U18361(.A(bypass_rs3h_w2_mux_n39), .Y(exu_n4639));
AND2X1 exu_U18362(.A(bypass_rs3h_w2_mux_n41), .B(exu_n10565), .Y(bypass_rs3h_data_w2[29]));
INVX1 exu_U18363(.A(bypass_rs3h_data_w2[29]), .Y(exu_n4640));
AND2X1 exu_U18364(.A(bypass_dfill_data_g2[29]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n43));
INVX1 exu_U18365(.A(bypass_rs3h_w2_mux_n43), .Y(exu_n4641));
AND2X1 exu_U18366(.A(bypass_rs3h_w2_mux_n45), .B(exu_n10566), .Y(bypass_rs3h_data_w2[28]));
INVX1 exu_U18367(.A(bypass_rs3h_data_w2[28]), .Y(exu_n4642));
AND2X1 exu_U18368(.A(bypass_dfill_data_g2[28]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n47));
INVX1 exu_U18369(.A(bypass_rs3h_w2_mux_n47), .Y(exu_n4643));
AND2X1 exu_U18370(.A(bypass_rs3h_w2_mux_n49), .B(exu_n10567), .Y(bypass_rs3h_data_w2[27]));
INVX1 exu_U18371(.A(bypass_rs3h_data_w2[27]), .Y(exu_n4644));
AND2X1 exu_U18372(.A(bypass_dfill_data_g2[27]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n51));
INVX1 exu_U18373(.A(bypass_rs3h_w2_mux_n51), .Y(exu_n4645));
AND2X1 exu_U18374(.A(bypass_rs3h_w2_mux_n53), .B(exu_n10568), .Y(bypass_rs3h_data_w2[26]));
INVX1 exu_U18375(.A(bypass_rs3h_data_w2[26]), .Y(exu_n4646));
AND2X1 exu_U18376(.A(bypass_dfill_data_g2[26]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n55));
INVX1 exu_U18377(.A(bypass_rs3h_w2_mux_n55), .Y(exu_n4647));
AND2X1 exu_U18378(.A(bypass_rs3h_w2_mux_n57), .B(exu_n10569), .Y(bypass_rs3h_data_w2[25]));
INVX1 exu_U18379(.A(bypass_rs3h_data_w2[25]), .Y(exu_n4648));
AND2X1 exu_U18380(.A(bypass_dfill_data_g2[25]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n59));
INVX1 exu_U18381(.A(bypass_rs3h_w2_mux_n59), .Y(exu_n4649));
AND2X1 exu_U18382(.A(bypass_rs3h_w2_mux_n61), .B(exu_n10570), .Y(bypass_rs3h_data_w2[24]));
INVX1 exu_U18383(.A(bypass_rs3h_data_w2[24]), .Y(exu_n4650));
AND2X1 exu_U18384(.A(bypass_dfill_data_g2[24]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n63));
INVX1 exu_U18385(.A(bypass_rs3h_w2_mux_n63), .Y(exu_n4651));
AND2X1 exu_U18386(.A(bypass_rs3h_w2_mux_n65), .B(exu_n10571), .Y(bypass_rs3h_data_w2[23]));
INVX1 exu_U18387(.A(bypass_rs3h_data_w2[23]), .Y(exu_n4652));
AND2X1 exu_U18388(.A(bypass_dfill_data_g2[23]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n67));
INVX1 exu_U18389(.A(bypass_rs3h_w2_mux_n67), .Y(exu_n4653));
AND2X1 exu_U18390(.A(bypass_rs3h_w2_mux_n69), .B(exu_n10572), .Y(bypass_rs3h_data_w2[22]));
INVX1 exu_U18391(.A(bypass_rs3h_data_w2[22]), .Y(exu_n4654));
AND2X1 exu_U18392(.A(bypass_dfill_data_g2[22]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n71));
INVX1 exu_U18393(.A(bypass_rs3h_w2_mux_n71), .Y(exu_n4655));
AND2X1 exu_U18394(.A(bypass_rs3h_w2_mux_n73), .B(exu_n10573), .Y(bypass_rs3h_data_w2[21]));
INVX1 exu_U18395(.A(bypass_rs3h_data_w2[21]), .Y(exu_n4656));
AND2X1 exu_U18396(.A(bypass_dfill_data_g2[21]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n75));
INVX1 exu_U18397(.A(bypass_rs3h_w2_mux_n75), .Y(exu_n4657));
AND2X1 exu_U18398(.A(bypass_rs3h_w2_mux_n77), .B(exu_n10574), .Y(bypass_rs3h_data_w2[20]));
INVX1 exu_U18399(.A(bypass_rs3h_data_w2[20]), .Y(exu_n4658));
AND2X1 exu_U18400(.A(bypass_dfill_data_g2[20]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n79));
INVX1 exu_U18401(.A(bypass_rs3h_w2_mux_n79), .Y(exu_n4659));
AND2X1 exu_U18402(.A(bypass_rs3h_w2_mux_n81), .B(exu_n10575), .Y(bypass_rs3h_data_w2[1]));
INVX1 exu_U18403(.A(bypass_rs3h_data_w2[1]), .Y(exu_n4660));
AND2X1 exu_U18404(.A(bypass_dfill_data_g2[1]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n83));
INVX1 exu_U18405(.A(bypass_rs3h_w2_mux_n83), .Y(exu_n4661));
AND2X1 exu_U18406(.A(bypass_rs3h_w2_mux_n85), .B(exu_n10576), .Y(bypass_rs3h_data_w2[19]));
INVX1 exu_U18407(.A(bypass_rs3h_data_w2[19]), .Y(exu_n4662));
AND2X1 exu_U18408(.A(bypass_dfill_data_g2[19]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n87));
INVX1 exu_U18409(.A(bypass_rs3h_w2_mux_n87), .Y(exu_n4663));
AND2X1 exu_U18410(.A(bypass_rs3h_w2_mux_n89), .B(exu_n10577), .Y(bypass_rs3h_data_w2[18]));
INVX1 exu_U18411(.A(bypass_rs3h_data_w2[18]), .Y(exu_n4664));
AND2X1 exu_U18412(.A(bypass_dfill_data_g2[18]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n91));
INVX1 exu_U18413(.A(bypass_rs3h_w2_mux_n91), .Y(exu_n4665));
AND2X1 exu_U18414(.A(bypass_rs3h_w2_mux_n93), .B(exu_n10578), .Y(bypass_rs3h_data_w2[17]));
INVX1 exu_U18415(.A(bypass_rs3h_data_w2[17]), .Y(exu_n4666));
AND2X1 exu_U18416(.A(bypass_dfill_data_g2[17]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n95));
INVX1 exu_U18417(.A(bypass_rs3h_w2_mux_n95), .Y(exu_n4667));
AND2X1 exu_U18418(.A(bypass_rs3h_w2_mux_n97), .B(exu_n10579), .Y(bypass_rs3h_data_w2[16]));
INVX1 exu_U18419(.A(bypass_rs3h_data_w2[16]), .Y(exu_n4668));
AND2X1 exu_U18420(.A(bypass_dfill_data_g2[16]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n99));
INVX1 exu_U18421(.A(bypass_rs3h_w2_mux_n99), .Y(exu_n4669));
AND2X1 exu_U18422(.A(bypass_rs3h_w2_mux_n101), .B(exu_n10580), .Y(bypass_rs3h_data_w2[15]));
INVX1 exu_U18423(.A(bypass_rs3h_data_w2[15]), .Y(exu_n4670));
AND2X1 exu_U18424(.A(bypass_dfill_data_g2[15]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n103));
INVX1 exu_U18425(.A(bypass_rs3h_w2_mux_n103), .Y(exu_n4671));
AND2X1 exu_U18426(.A(bypass_rs3h_w2_mux_n105), .B(exu_n10581), .Y(bypass_rs3h_data_w2[14]));
INVX1 exu_U18427(.A(bypass_rs3h_data_w2[14]), .Y(exu_n4672));
AND2X1 exu_U18428(.A(bypass_dfill_data_g2[14]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n107));
INVX1 exu_U18429(.A(bypass_rs3h_w2_mux_n107), .Y(exu_n4673));
AND2X1 exu_U18430(.A(bypass_rs3h_w2_mux_n109), .B(exu_n10582), .Y(bypass_rs3h_data_w2[13]));
INVX1 exu_U18431(.A(bypass_rs3h_data_w2[13]), .Y(exu_n4674));
AND2X1 exu_U18432(.A(bypass_dfill_data_g2[13]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n111));
INVX1 exu_U18433(.A(bypass_rs3h_w2_mux_n111), .Y(exu_n4675));
AND2X1 exu_U18434(.A(bypass_rs3h_w2_mux_n113), .B(exu_n10583), .Y(bypass_rs3h_data_w2[12]));
INVX1 exu_U18435(.A(bypass_rs3h_data_w2[12]), .Y(exu_n4676));
AND2X1 exu_U18436(.A(bypass_dfill_data_g2[12]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n115));
INVX1 exu_U18437(.A(bypass_rs3h_w2_mux_n115), .Y(exu_n4677));
AND2X1 exu_U18438(.A(bypass_rs3h_w2_mux_n117), .B(exu_n10584), .Y(bypass_rs3h_data_w2[11]));
INVX1 exu_U18439(.A(bypass_rs3h_data_w2[11]), .Y(exu_n4678));
AND2X1 exu_U18440(.A(bypass_dfill_data_g2[11]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n119));
INVX1 exu_U18441(.A(bypass_rs3h_w2_mux_n119), .Y(exu_n4679));
AND2X1 exu_U18442(.A(bypass_rs3h_w2_mux_n121), .B(exu_n10585), .Y(bypass_rs3h_data_w2[10]));
INVX1 exu_U18443(.A(bypass_rs3h_data_w2[10]), .Y(exu_n4680));
AND2X1 exu_U18444(.A(bypass_dfill_data_g2[10]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n123));
INVX1 exu_U18445(.A(bypass_rs3h_w2_mux_n123), .Y(exu_n4681));
AND2X1 exu_U18446(.A(bypass_rs3h_w2_mux_n125), .B(exu_n10586), .Y(bypass_rs3h_data_w2[0]));
INVX1 exu_U18447(.A(bypass_rs3h_data_w2[0]), .Y(exu_n4682));
AND2X1 exu_U18448(.A(bypass_dfill_data_g2[0]), .B(exu_n16275), .Y(bypass_rs3h_w2_mux_n127));
INVX1 exu_U18449(.A(bypass_rs3h_w2_mux_n127), .Y(exu_n4683));
AND2X1 exu_U18450(.A(ecl_byp_sel_ffusr_m), .B(ffu_exu_rsr_data_m[9]), .Y(bypass_sr_out_mux_n3));
INVX1 exu_U18451(.A(bypass_sr_out_mux_n3), .Y(exu_n4684));
AND2X1 exu_U18452(.A(ffu_exu_rsr_data_m[8]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n7));
INVX1 exu_U18453(.A(bypass_sr_out_mux_n7), .Y(exu_n4685));
AND2X1 exu_U18454(.A(ffu_exu_rsr_data_m[7]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n11));
INVX1 exu_U18455(.A(bypass_sr_out_mux_n11), .Y(exu_n4686));
AND2X1 exu_U18456(.A(ffu_exu_rsr_data_m[6]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n15));
INVX1 exu_U18457(.A(bypass_sr_out_mux_n15), .Y(exu_n4687));
AND2X1 exu_U18458(.A(ffu_exu_rsr_data_m[63]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n19));
INVX1 exu_U18459(.A(bypass_sr_out_mux_n19), .Y(exu_n4688));
AND2X1 exu_U18460(.A(ffu_exu_rsr_data_m[62]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n23));
INVX1 exu_U18461(.A(bypass_sr_out_mux_n23), .Y(exu_n4689));
AND2X1 exu_U18462(.A(ffu_exu_rsr_data_m[61]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n27));
INVX1 exu_U18463(.A(bypass_sr_out_mux_n27), .Y(exu_n4690));
AND2X1 exu_U18464(.A(ffu_exu_rsr_data_m[60]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n31));
INVX1 exu_U18465(.A(bypass_sr_out_mux_n31), .Y(exu_n4691));
AND2X1 exu_U18466(.A(ffu_exu_rsr_data_m[5]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n35));
INVX1 exu_U18467(.A(bypass_sr_out_mux_n35), .Y(exu_n4692));
AND2X1 exu_U18468(.A(ffu_exu_rsr_data_m[59]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n39));
INVX1 exu_U18469(.A(bypass_sr_out_mux_n39), .Y(exu_n4693));
AND2X1 exu_U18470(.A(ffu_exu_rsr_data_m[58]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n43));
INVX1 exu_U18471(.A(bypass_sr_out_mux_n43), .Y(exu_n4694));
AND2X1 exu_U18472(.A(ffu_exu_rsr_data_m[57]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n47));
INVX1 exu_U18473(.A(bypass_sr_out_mux_n47), .Y(exu_n4695));
AND2X1 exu_U18474(.A(ffu_exu_rsr_data_m[56]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n51));
INVX1 exu_U18475(.A(bypass_sr_out_mux_n51), .Y(exu_n4696));
AND2X1 exu_U18476(.A(ffu_exu_rsr_data_m[55]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n55));
INVX1 exu_U18477(.A(bypass_sr_out_mux_n55), .Y(exu_n4697));
AND2X1 exu_U18478(.A(ffu_exu_rsr_data_m[54]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n59));
INVX1 exu_U18479(.A(bypass_sr_out_mux_n59), .Y(exu_n4698));
AND2X1 exu_U18480(.A(ffu_exu_rsr_data_m[53]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n63));
INVX1 exu_U18481(.A(bypass_sr_out_mux_n63), .Y(exu_n4699));
AND2X1 exu_U18482(.A(ffu_exu_rsr_data_m[52]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n67));
INVX1 exu_U18483(.A(bypass_sr_out_mux_n67), .Y(exu_n4700));
AND2X1 exu_U18484(.A(ffu_exu_rsr_data_m[51]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n71));
INVX1 exu_U18485(.A(bypass_sr_out_mux_n71), .Y(exu_n4701));
AND2X1 exu_U18486(.A(ffu_exu_rsr_data_m[50]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n75));
INVX1 exu_U18487(.A(bypass_sr_out_mux_n75), .Y(exu_n4702));
AND2X1 exu_U18488(.A(ffu_exu_rsr_data_m[4]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n79));
INVX1 exu_U18489(.A(bypass_sr_out_mux_n79), .Y(exu_n4703));
AND2X1 exu_U18490(.A(ffu_exu_rsr_data_m[49]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n83));
INVX1 exu_U18491(.A(bypass_sr_out_mux_n83), .Y(exu_n4704));
AND2X1 exu_U18492(.A(ffu_exu_rsr_data_m[48]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n87));
INVX1 exu_U18493(.A(bypass_sr_out_mux_n87), .Y(exu_n4705));
AND2X1 exu_U18494(.A(ffu_exu_rsr_data_m[47]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n91));
INVX1 exu_U18495(.A(bypass_sr_out_mux_n91), .Y(exu_n4706));
AND2X1 exu_U18496(.A(ffu_exu_rsr_data_m[46]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n95));
INVX1 exu_U18497(.A(bypass_sr_out_mux_n95), .Y(exu_n4707));
AND2X1 exu_U18498(.A(ffu_exu_rsr_data_m[45]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n99));
INVX1 exu_U18499(.A(bypass_sr_out_mux_n99), .Y(exu_n4708));
AND2X1 exu_U18500(.A(ffu_exu_rsr_data_m[44]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n103));
INVX1 exu_U18501(.A(bypass_sr_out_mux_n103), .Y(exu_n4709));
AND2X1 exu_U18502(.A(ffu_exu_rsr_data_m[43]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n107));
INVX1 exu_U18503(.A(bypass_sr_out_mux_n107), .Y(exu_n4710));
AND2X1 exu_U18504(.A(ffu_exu_rsr_data_m[42]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n111));
INVX1 exu_U18505(.A(bypass_sr_out_mux_n111), .Y(exu_n4711));
AND2X1 exu_U18506(.A(ffu_exu_rsr_data_m[41]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n115));
INVX1 exu_U18507(.A(bypass_sr_out_mux_n115), .Y(exu_n4712));
AND2X1 exu_U18508(.A(ffu_exu_rsr_data_m[40]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n119));
INVX1 exu_U18509(.A(bypass_sr_out_mux_n119), .Y(exu_n4713));
AND2X1 exu_U18510(.A(ffu_exu_rsr_data_m[3]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n123));
INVX1 exu_U18511(.A(bypass_sr_out_mux_n123), .Y(exu_n4714));
AND2X1 exu_U18512(.A(ffu_exu_rsr_data_m[39]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n127));
INVX1 exu_U18513(.A(bypass_sr_out_mux_n127), .Y(exu_n4715));
AND2X1 exu_U18514(.A(ffu_exu_rsr_data_m[38]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n131));
INVX1 exu_U18515(.A(bypass_sr_out_mux_n131), .Y(exu_n4716));
AND2X1 exu_U18516(.A(ffu_exu_rsr_data_m[37]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n135));
INVX1 exu_U18517(.A(bypass_sr_out_mux_n135), .Y(exu_n4717));
AND2X1 exu_U18518(.A(ffu_exu_rsr_data_m[36]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n139));
INVX1 exu_U18519(.A(bypass_sr_out_mux_n139), .Y(exu_n4718));
AND2X1 exu_U18520(.A(ffu_exu_rsr_data_m[35]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n143));
INVX1 exu_U18521(.A(bypass_sr_out_mux_n143), .Y(exu_n4719));
AND2X1 exu_U18522(.A(ffu_exu_rsr_data_m[34]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n147));
INVX1 exu_U18523(.A(bypass_sr_out_mux_n147), .Y(exu_n4720));
AND2X1 exu_U18524(.A(ffu_exu_rsr_data_m[33]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n151));
INVX1 exu_U18525(.A(bypass_sr_out_mux_n151), .Y(exu_n4721));
AND2X1 exu_U18526(.A(ffu_exu_rsr_data_m[32]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n155));
INVX1 exu_U18527(.A(bypass_sr_out_mux_n155), .Y(exu_n4722));
AND2X1 exu_U18528(.A(ffu_exu_rsr_data_m[31]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n159));
INVX1 exu_U18529(.A(bypass_sr_out_mux_n159), .Y(exu_n4723));
AND2X1 exu_U18530(.A(ffu_exu_rsr_data_m[30]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n163));
INVX1 exu_U18531(.A(bypass_sr_out_mux_n163), .Y(exu_n4724));
AND2X1 exu_U18532(.A(ffu_exu_rsr_data_m[2]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n167));
INVX1 exu_U18533(.A(bypass_sr_out_mux_n167), .Y(exu_n4725));
AND2X1 exu_U18534(.A(ffu_exu_rsr_data_m[29]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n171));
INVX1 exu_U18535(.A(bypass_sr_out_mux_n171), .Y(exu_n4726));
AND2X1 exu_U18536(.A(ffu_exu_rsr_data_m[28]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n175));
INVX1 exu_U18537(.A(bypass_sr_out_mux_n175), .Y(exu_n4727));
AND2X1 exu_U18538(.A(ffu_exu_rsr_data_m[27]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n179));
INVX1 exu_U18539(.A(bypass_sr_out_mux_n179), .Y(exu_n4728));
AND2X1 exu_U18540(.A(ffu_exu_rsr_data_m[26]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n183));
INVX1 exu_U18541(.A(bypass_sr_out_mux_n183), .Y(exu_n4729));
AND2X1 exu_U18542(.A(ffu_exu_rsr_data_m[25]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n187));
INVX1 exu_U18543(.A(bypass_sr_out_mux_n187), .Y(exu_n4730));
AND2X1 exu_U18544(.A(ffu_exu_rsr_data_m[24]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n191));
INVX1 exu_U18545(.A(bypass_sr_out_mux_n191), .Y(exu_n4731));
AND2X1 exu_U18546(.A(ffu_exu_rsr_data_m[23]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n195));
INVX1 exu_U18547(.A(bypass_sr_out_mux_n195), .Y(exu_n4732));
AND2X1 exu_U18548(.A(ffu_exu_rsr_data_m[22]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n199));
INVX1 exu_U18549(.A(bypass_sr_out_mux_n199), .Y(exu_n4733));
AND2X1 exu_U18550(.A(ffu_exu_rsr_data_m[21]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n203));
INVX1 exu_U18551(.A(bypass_sr_out_mux_n203), .Y(exu_n4734));
AND2X1 exu_U18552(.A(ffu_exu_rsr_data_m[20]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n207));
INVX1 exu_U18553(.A(bypass_sr_out_mux_n207), .Y(exu_n4735));
AND2X1 exu_U18554(.A(ffu_exu_rsr_data_m[1]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n211));
INVX1 exu_U18555(.A(bypass_sr_out_mux_n211), .Y(exu_n4736));
AND2X1 exu_U18556(.A(ffu_exu_rsr_data_m[19]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n215));
INVX1 exu_U18557(.A(bypass_sr_out_mux_n215), .Y(exu_n4737));
AND2X1 exu_U18558(.A(ffu_exu_rsr_data_m[18]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n219));
INVX1 exu_U18559(.A(bypass_sr_out_mux_n219), .Y(exu_n4738));
AND2X1 exu_U18560(.A(ffu_exu_rsr_data_m[17]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n223));
INVX1 exu_U18561(.A(bypass_sr_out_mux_n223), .Y(exu_n4739));
AND2X1 exu_U18562(.A(ffu_exu_rsr_data_m[16]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n227));
INVX1 exu_U18563(.A(bypass_sr_out_mux_n227), .Y(exu_n4740));
AND2X1 exu_U18564(.A(ffu_exu_rsr_data_m[15]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n231));
INVX1 exu_U18565(.A(bypass_sr_out_mux_n231), .Y(exu_n4741));
AND2X1 exu_U18566(.A(ffu_exu_rsr_data_m[14]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n235));
INVX1 exu_U18567(.A(bypass_sr_out_mux_n235), .Y(exu_n4742));
AND2X1 exu_U18568(.A(ffu_exu_rsr_data_m[13]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n239));
INVX1 exu_U18569(.A(bypass_sr_out_mux_n239), .Y(exu_n4743));
AND2X1 exu_U18570(.A(ffu_exu_rsr_data_m[12]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n243));
INVX1 exu_U18571(.A(bypass_sr_out_mux_n243), .Y(exu_n4744));
AND2X1 exu_U18572(.A(ffu_exu_rsr_data_m[11]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n247));
INVX1 exu_U18573(.A(bypass_sr_out_mux_n247), .Y(exu_n4745));
AND2X1 exu_U18574(.A(ffu_exu_rsr_data_m[10]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n251));
INVX1 exu_U18575(.A(bypass_sr_out_mux_n251), .Y(exu_n4746));
AND2X1 exu_U18576(.A(ffu_exu_rsr_data_m[0]), .B(ecl_byp_sel_ffusr_m), .Y(bypass_sr_out_mux_n255));
INVX1 exu_U18577(.A(bypass_sr_out_mux_n255), .Y(exu_n4747));
AND2X1 exu_U18578(.A(ecl_byp_sel_alu_e), .B(alu_byp_rd_data_e[9]), .Y(bypass_ifu_exu_sr_mux_n3));
INVX1 exu_U18579(.A(bypass_ifu_exu_sr_mux_n3), .Y(exu_n4748));
AND2X1 exu_U18580(.A(alu_byp_rd_data_e[8]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n9));
INVX1 exu_U18581(.A(bypass_ifu_exu_sr_mux_n9), .Y(exu_n4749));
AND2X1 exu_U18582(.A(alu_byp_rd_data_e[7]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n15));
INVX1 exu_U18583(.A(bypass_ifu_exu_sr_mux_n15), .Y(exu_n4750));
AND2X1 exu_U18584(.A(ecl_byp_eclpr_e[7]), .B(ecl_byp_sel_eclpr_e), .Y(bypass_ifu_exu_sr_mux_n17));
INVX1 exu_U18585(.A(bypass_ifu_exu_sr_mux_n17), .Y(exu_n4751));
AND2X1 exu_U18586(.A(alu_byp_rd_data_e[6]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n21));
INVX1 exu_U18587(.A(bypass_ifu_exu_sr_mux_n21), .Y(exu_n4752));
AND2X1 exu_U18588(.A(ecl_byp_eclpr_e[6]), .B(ecl_byp_sel_eclpr_e), .Y(bypass_ifu_exu_sr_mux_n23));
INVX1 exu_U18589(.A(bypass_ifu_exu_sr_mux_n23), .Y(exu_n4753));
AND2X1 exu_U18590(.A(exu_n11754), .B(exu_n10589), .Y(bypass_ifu_exu_sr_mux_n26));
INVX1 exu_U18591(.A(bypass_ifu_exu_sr_mux_n26), .Y(exu_n4754));
AND2X1 exu_U18592(.A(exu_n11755), .B(exu_n10590), .Y(bypass_ifu_exu_sr_mux_n32));
INVX1 exu_U18593(.A(bypass_ifu_exu_sr_mux_n32), .Y(exu_n4755));
AND2X1 exu_U18594(.A(exu_n11756), .B(exu_n10591), .Y(bypass_ifu_exu_sr_mux_n38));
INVX1 exu_U18595(.A(bypass_ifu_exu_sr_mux_n38), .Y(exu_n4756));
AND2X1 exu_U18596(.A(exu_n11757), .B(exu_n10592), .Y(bypass_ifu_exu_sr_mux_n44));
INVX1 exu_U18597(.A(bypass_ifu_exu_sr_mux_n44), .Y(exu_n4757));
AND2X1 exu_U18598(.A(alu_byp_rd_data_e[5]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n51));
INVX1 exu_U18599(.A(bypass_ifu_exu_sr_mux_n51), .Y(exu_n4758));
AND2X1 exu_U18600(.A(ecl_byp_eclpr_e[5]), .B(ecl_byp_sel_eclpr_e), .Y(bypass_ifu_exu_sr_mux_n53));
INVX1 exu_U18601(.A(bypass_ifu_exu_sr_mux_n53), .Y(exu_n4759));
AND2X1 exu_U18602(.A(exu_n11758), .B(exu_n10593), .Y(bypass_ifu_exu_sr_mux_n56));
INVX1 exu_U18603(.A(bypass_ifu_exu_sr_mux_n56), .Y(exu_n4760));
AND2X1 exu_U18604(.A(exu_n11759), .B(exu_n10594), .Y(bypass_ifu_exu_sr_mux_n62));
INVX1 exu_U18605(.A(bypass_ifu_exu_sr_mux_n62), .Y(exu_n4761));
AND2X1 exu_U18606(.A(exu_n11760), .B(exu_n10595), .Y(bypass_ifu_exu_sr_mux_n68));
INVX1 exu_U18607(.A(bypass_ifu_exu_sr_mux_n68), .Y(exu_n4762));
AND2X1 exu_U18608(.A(exu_n11761), .B(exu_n10596), .Y(bypass_ifu_exu_sr_mux_n74));
INVX1 exu_U18609(.A(bypass_ifu_exu_sr_mux_n74), .Y(exu_n4763));
AND2X1 exu_U18610(.A(exu_n11762), .B(exu_n10597), .Y(bypass_ifu_exu_sr_mux_n80));
INVX1 exu_U18611(.A(bypass_ifu_exu_sr_mux_n80), .Y(exu_n4764));
AND2X1 exu_U18612(.A(exu_n11763), .B(exu_n10598), .Y(bypass_ifu_exu_sr_mux_n86));
INVX1 exu_U18613(.A(bypass_ifu_exu_sr_mux_n86), .Y(exu_n4765));
AND2X1 exu_U18614(.A(exu_n11764), .B(exu_n10599), .Y(bypass_ifu_exu_sr_mux_n92));
INVX1 exu_U18615(.A(bypass_ifu_exu_sr_mux_n92), .Y(exu_n4766));
AND2X1 exu_U18616(.A(exu_n11765), .B(exu_n10600), .Y(bypass_ifu_exu_sr_mux_n98));
INVX1 exu_U18617(.A(bypass_ifu_exu_sr_mux_n98), .Y(exu_n4767));
AND2X1 exu_U18618(.A(exu_n11766), .B(exu_n10601), .Y(bypass_ifu_exu_sr_mux_n104));
INVX1 exu_U18619(.A(bypass_ifu_exu_sr_mux_n104), .Y(exu_n4768));
AND2X1 exu_U18620(.A(exu_n11767), .B(exu_n10602), .Y(bypass_ifu_exu_sr_mux_n110));
INVX1 exu_U18621(.A(bypass_ifu_exu_sr_mux_n110), .Y(exu_n4769));
AND2X1 exu_U18622(.A(alu_byp_rd_data_e[4]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n117));
INVX1 exu_U18623(.A(bypass_ifu_exu_sr_mux_n117), .Y(exu_n4770));
AND2X1 exu_U18624(.A(ecl_byp_eclpr_e[4]), .B(ecl_byp_sel_eclpr_e), .Y(bypass_ifu_exu_sr_mux_n119));
INVX1 exu_U18625(.A(bypass_ifu_exu_sr_mux_n119), .Y(exu_n4771));
AND2X1 exu_U18626(.A(exu_n11768), .B(exu_n10603), .Y(bypass_ifu_exu_sr_mux_n122));
INVX1 exu_U18627(.A(bypass_ifu_exu_sr_mux_n122), .Y(exu_n4772));
AND2X1 exu_U18628(.A(exu_n11769), .B(exu_n10604), .Y(bypass_ifu_exu_sr_mux_n128));
INVX1 exu_U18629(.A(bypass_ifu_exu_sr_mux_n128), .Y(exu_n4773));
AND2X1 exu_U18630(.A(exu_n11770), .B(exu_n10605), .Y(bypass_ifu_exu_sr_mux_n134));
INVX1 exu_U18631(.A(bypass_ifu_exu_sr_mux_n134), .Y(exu_n4774));
AND2X1 exu_U18632(.A(exu_n11771), .B(exu_n10606), .Y(bypass_ifu_exu_sr_mux_n140));
INVX1 exu_U18633(.A(bypass_ifu_exu_sr_mux_n140), .Y(exu_n4775));
AND2X1 exu_U18634(.A(exu_n11772), .B(exu_n10607), .Y(bypass_ifu_exu_sr_mux_n146));
INVX1 exu_U18635(.A(bypass_ifu_exu_sr_mux_n146), .Y(exu_n4776));
AND2X1 exu_U18636(.A(exu_n11773), .B(exu_n10608), .Y(bypass_ifu_exu_sr_mux_n152));
INVX1 exu_U18637(.A(bypass_ifu_exu_sr_mux_n152), .Y(exu_n4777));
AND2X1 exu_U18638(.A(exu_n11774), .B(exu_n10609), .Y(bypass_ifu_exu_sr_mux_n158));
INVX1 exu_U18639(.A(bypass_ifu_exu_sr_mux_n158), .Y(exu_n4778));
AND2X1 exu_U18640(.A(exu_n11775), .B(exu_n10610), .Y(bypass_ifu_exu_sr_mux_n164));
INVX1 exu_U18641(.A(bypass_ifu_exu_sr_mux_n164), .Y(exu_n4779));
AND2X1 exu_U18642(.A(exu_n11776), .B(exu_n10611), .Y(bypass_ifu_exu_sr_mux_n170));
INVX1 exu_U18643(.A(bypass_ifu_exu_sr_mux_n170), .Y(exu_n4780));
AND2X1 exu_U18644(.A(exu_n11777), .B(exu_n10612), .Y(bypass_ifu_exu_sr_mux_n176));
INVX1 exu_U18645(.A(bypass_ifu_exu_sr_mux_n176), .Y(exu_n4781));
AND2X1 exu_U18646(.A(alu_byp_rd_data_e[3]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n183));
INVX1 exu_U18647(.A(bypass_ifu_exu_sr_mux_n183), .Y(exu_n4782));
AND2X1 exu_U18648(.A(ecl_byp_eclpr_e[3]), .B(ecl_byp_sel_eclpr_e), .Y(bypass_ifu_exu_sr_mux_n185));
INVX1 exu_U18649(.A(bypass_ifu_exu_sr_mux_n185), .Y(exu_n4783));
AND2X1 exu_U18650(.A(exu_n11778), .B(exu_n10613), .Y(bypass_ifu_exu_sr_mux_n188));
INVX1 exu_U18651(.A(bypass_ifu_exu_sr_mux_n188), .Y(exu_n4784));
AND2X1 exu_U18652(.A(exu_n11779), .B(exu_n10614), .Y(bypass_ifu_exu_sr_mux_n194));
INVX1 exu_U18653(.A(bypass_ifu_exu_sr_mux_n194), .Y(exu_n4785));
AND2X1 exu_U18654(.A(exu_n11780), .B(exu_n10615), .Y(bypass_ifu_exu_sr_mux_n200));
INVX1 exu_U18655(.A(bypass_ifu_exu_sr_mux_n200), .Y(exu_n4786));
AND2X1 exu_U18656(.A(exu_n11781), .B(exu_n10616), .Y(bypass_ifu_exu_sr_mux_n206));
INVX1 exu_U18657(.A(bypass_ifu_exu_sr_mux_n206), .Y(exu_n4787));
AND2X1 exu_U18658(.A(exu_n11782), .B(exu_n10617), .Y(bypass_ifu_exu_sr_mux_n212));
INVX1 exu_U18659(.A(bypass_ifu_exu_sr_mux_n212), .Y(exu_n4788));
AND2X1 exu_U18660(.A(exu_n11783), .B(exu_n10618), .Y(bypass_ifu_exu_sr_mux_n218));
INVX1 exu_U18661(.A(bypass_ifu_exu_sr_mux_n218), .Y(exu_n4789));
AND2X1 exu_U18662(.A(exu_n11784), .B(exu_n10619), .Y(bypass_ifu_exu_sr_mux_n224));
INVX1 exu_U18663(.A(bypass_ifu_exu_sr_mux_n224), .Y(exu_n4790));
AND2X1 exu_U18664(.A(exu_n11785), .B(exu_n10620), .Y(bypass_ifu_exu_sr_mux_n230));
INVX1 exu_U18665(.A(bypass_ifu_exu_sr_mux_n230), .Y(exu_n4791));
AND2X1 exu_U18666(.A(alu_byp_rd_data_e[31]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n237));
INVX1 exu_U18667(.A(bypass_ifu_exu_sr_mux_n237), .Y(exu_n4792));
AND2X1 exu_U18668(.A(alu_byp_rd_data_e[30]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n243));
INVX1 exu_U18669(.A(bypass_ifu_exu_sr_mux_n243), .Y(exu_n4793));
AND2X1 exu_U18670(.A(alu_byp_rd_data_e[2]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n249));
INVX1 exu_U18671(.A(bypass_ifu_exu_sr_mux_n249), .Y(exu_n4794));
AND2X1 exu_U18672(.A(ecl_byp_eclpr_e[2]), .B(ecl_byp_sel_eclpr_e), .Y(bypass_ifu_exu_sr_mux_n251));
INVX1 exu_U18673(.A(bypass_ifu_exu_sr_mux_n251), .Y(exu_n4795));
AND2X1 exu_U18674(.A(alu_byp_rd_data_e[29]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n255));
INVX1 exu_U18675(.A(bypass_ifu_exu_sr_mux_n255), .Y(exu_n4796));
AND2X1 exu_U18676(.A(alu_byp_rd_data_e[28]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n261));
INVX1 exu_U18677(.A(bypass_ifu_exu_sr_mux_n261), .Y(exu_n4797));
AND2X1 exu_U18678(.A(alu_byp_rd_data_e[27]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n267));
INVX1 exu_U18679(.A(bypass_ifu_exu_sr_mux_n267), .Y(exu_n4798));
AND2X1 exu_U18680(.A(alu_byp_rd_data_e[26]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n273));
INVX1 exu_U18681(.A(bypass_ifu_exu_sr_mux_n273), .Y(exu_n4799));
AND2X1 exu_U18682(.A(alu_byp_rd_data_e[25]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n279));
INVX1 exu_U18683(.A(bypass_ifu_exu_sr_mux_n279), .Y(exu_n4800));
AND2X1 exu_U18684(.A(alu_byp_rd_data_e[24]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n285));
INVX1 exu_U18685(.A(bypass_ifu_exu_sr_mux_n285), .Y(exu_n4801));
AND2X1 exu_U18686(.A(alu_byp_rd_data_e[23]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n291));
INVX1 exu_U18687(.A(bypass_ifu_exu_sr_mux_n291), .Y(exu_n4802));
AND2X1 exu_U18688(.A(alu_byp_rd_data_e[22]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n297));
INVX1 exu_U18689(.A(bypass_ifu_exu_sr_mux_n297), .Y(exu_n4803));
AND2X1 exu_U18690(.A(alu_byp_rd_data_e[21]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n303));
INVX1 exu_U18691(.A(bypass_ifu_exu_sr_mux_n303), .Y(exu_n4804));
AND2X1 exu_U18692(.A(alu_byp_rd_data_e[20]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n309));
INVX1 exu_U18693(.A(bypass_ifu_exu_sr_mux_n309), .Y(exu_n4805));
AND2X1 exu_U18694(.A(alu_byp_rd_data_e[1]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n315));
INVX1 exu_U18695(.A(bypass_ifu_exu_sr_mux_n315), .Y(exu_n4806));
AND2X1 exu_U18696(.A(ecl_byp_eclpr_e[1]), .B(ecl_byp_sel_eclpr_e), .Y(bypass_ifu_exu_sr_mux_n317));
INVX1 exu_U18697(.A(bypass_ifu_exu_sr_mux_n317), .Y(exu_n4807));
AND2X1 exu_U18698(.A(alu_byp_rd_data_e[19]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n321));
INVX1 exu_U18699(.A(bypass_ifu_exu_sr_mux_n321), .Y(exu_n4808));
AND2X1 exu_U18700(.A(alu_byp_rd_data_e[18]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n327));
INVX1 exu_U18701(.A(bypass_ifu_exu_sr_mux_n327), .Y(exu_n4809));
AND2X1 exu_U18702(.A(alu_byp_rd_data_e[17]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n333));
INVX1 exu_U18703(.A(bypass_ifu_exu_sr_mux_n333), .Y(exu_n4810));
AND2X1 exu_U18704(.A(alu_byp_rd_data_e[16]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n339));
INVX1 exu_U18705(.A(bypass_ifu_exu_sr_mux_n339), .Y(exu_n4811));
AND2X1 exu_U18706(.A(alu_byp_rd_data_e[15]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n345));
INVX1 exu_U18707(.A(bypass_ifu_exu_sr_mux_n345), .Y(exu_n4812));
AND2X1 exu_U18708(.A(alu_byp_rd_data_e[14]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n351));
INVX1 exu_U18709(.A(bypass_ifu_exu_sr_mux_n351), .Y(exu_n4813));
AND2X1 exu_U18710(.A(alu_byp_rd_data_e[13]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n357));
INVX1 exu_U18711(.A(bypass_ifu_exu_sr_mux_n357), .Y(exu_n4814));
AND2X1 exu_U18712(.A(alu_byp_rd_data_e[12]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n363));
INVX1 exu_U18713(.A(bypass_ifu_exu_sr_mux_n363), .Y(exu_n4815));
AND2X1 exu_U18714(.A(alu_byp_rd_data_e[11]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n369));
INVX1 exu_U18715(.A(bypass_ifu_exu_sr_mux_n369), .Y(exu_n4816));
AND2X1 exu_U18716(.A(alu_byp_rd_data_e[10]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n375));
INVX1 exu_U18717(.A(bypass_ifu_exu_sr_mux_n375), .Y(exu_n4817));
AND2X1 exu_U18718(.A(alu_byp_rd_data_e[0]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n381));
INVX1 exu_U18719(.A(bypass_ifu_exu_sr_mux_n381), .Y(exu_n4818));
AND2X1 exu_U18720(.A(ecl_byp_eclpr_e[0]), .B(ecl_byp_sel_eclpr_e), .Y(bypass_ifu_exu_sr_mux_n383));
INVX1 exu_U18721(.A(bypass_ifu_exu_sr_mux_n383), .Y(exu_n4819));
AND2X1 exu_U18722(.A(exu_n11786), .B(exu_n10621), .Y(bypass_dfill_data_g[9]));
INVX1 exu_U18723(.A(bypass_dfill_data_g[9]), .Y(exu_n4820));
AND2X1 exu_U18724(.A(exu_n11787), .B(exu_n10622), .Y(bypass_dfill_data_g[8]));
INVX1 exu_U18725(.A(bypass_dfill_data_g[8]), .Y(exu_n4821));
AND2X1 exu_U18726(.A(exu_n11788), .B(exu_n10623), .Y(bypass_dfill_data_g[7]));
INVX1 exu_U18727(.A(bypass_dfill_data_g[7]), .Y(exu_n4822));
AND2X1 exu_U18728(.A(exu_n11789), .B(exu_n10624), .Y(bypass_dfill_data_g[6]));
INVX1 exu_U18729(.A(bypass_dfill_data_g[6]), .Y(exu_n4823));
AND2X1 exu_U18730(.A(exu_n11790), .B(exu_n10625), .Y(bypass_dfill_data_g[63]));
INVX1 exu_U18731(.A(bypass_dfill_data_g[63]), .Y(exu_n4824));
AND2X1 exu_U18732(.A(exu_n11791), .B(exu_n10626), .Y(bypass_dfill_data_g[62]));
INVX1 exu_U18733(.A(bypass_dfill_data_g[62]), .Y(exu_n4825));
AND2X1 exu_U18734(.A(exu_n11792), .B(exu_n10627), .Y(bypass_dfill_data_g[61]));
INVX1 exu_U18735(.A(bypass_dfill_data_g[61]), .Y(exu_n4826));
AND2X1 exu_U18736(.A(exu_n11793), .B(exu_n10628), .Y(bypass_dfill_data_g[60]));
INVX1 exu_U18737(.A(bypass_dfill_data_g[60]), .Y(exu_n4827));
AND2X1 exu_U18738(.A(exu_n11794), .B(exu_n10629), .Y(bypass_dfill_data_g[5]));
INVX1 exu_U18739(.A(bypass_dfill_data_g[5]), .Y(exu_n4828));
AND2X1 exu_U18740(.A(exu_n11795), .B(exu_n10630), .Y(bypass_dfill_data_g[59]));
INVX1 exu_U18741(.A(bypass_dfill_data_g[59]), .Y(exu_n4829));
AND2X1 exu_U18742(.A(exu_n11796), .B(exu_n10631), .Y(bypass_dfill_data_g[58]));
INVX1 exu_U18743(.A(bypass_dfill_data_g[58]), .Y(exu_n4830));
AND2X1 exu_U18744(.A(exu_n11797), .B(exu_n10632), .Y(bypass_dfill_data_g[57]));
INVX1 exu_U18745(.A(bypass_dfill_data_g[57]), .Y(exu_n4831));
AND2X1 exu_U18746(.A(exu_n11798), .B(exu_n10633), .Y(bypass_dfill_data_g[56]));
INVX1 exu_U18747(.A(bypass_dfill_data_g[56]), .Y(exu_n4832));
AND2X1 exu_U18748(.A(exu_n11799), .B(exu_n10634), .Y(bypass_dfill_data_g[55]));
INVX1 exu_U18749(.A(bypass_dfill_data_g[55]), .Y(exu_n4833));
AND2X1 exu_U18750(.A(exu_n11800), .B(exu_n10635), .Y(bypass_dfill_data_g[54]));
INVX1 exu_U18751(.A(bypass_dfill_data_g[54]), .Y(exu_n4834));
AND2X1 exu_U18752(.A(exu_n11801), .B(exu_n10636), .Y(bypass_dfill_data_g[53]));
INVX1 exu_U18753(.A(bypass_dfill_data_g[53]), .Y(exu_n4835));
AND2X1 exu_U18754(.A(exu_n11802), .B(exu_n10637), .Y(bypass_dfill_data_g[52]));
INVX1 exu_U18755(.A(bypass_dfill_data_g[52]), .Y(exu_n4836));
AND2X1 exu_U18756(.A(exu_n11803), .B(exu_n10638), .Y(bypass_dfill_data_g[51]));
INVX1 exu_U18757(.A(bypass_dfill_data_g[51]), .Y(exu_n4837));
AND2X1 exu_U18758(.A(exu_n11804), .B(exu_n10639), .Y(bypass_dfill_data_g[50]));
INVX1 exu_U18759(.A(bypass_dfill_data_g[50]), .Y(exu_n4838));
AND2X1 exu_U18760(.A(exu_n11805), .B(exu_n10640), .Y(bypass_dfill_data_g[4]));
INVX1 exu_U18761(.A(bypass_dfill_data_g[4]), .Y(exu_n4839));
AND2X1 exu_U18762(.A(exu_n11806), .B(exu_n10641), .Y(bypass_dfill_data_g[49]));
INVX1 exu_U18763(.A(bypass_dfill_data_g[49]), .Y(exu_n4840));
AND2X1 exu_U18764(.A(exu_n11807), .B(exu_n10642), .Y(bypass_dfill_data_g[48]));
INVX1 exu_U18765(.A(bypass_dfill_data_g[48]), .Y(exu_n4841));
AND2X1 exu_U18766(.A(exu_n11808), .B(exu_n10643), .Y(bypass_dfill_data_g[47]));
INVX1 exu_U18767(.A(bypass_dfill_data_g[47]), .Y(exu_n4842));
AND2X1 exu_U18768(.A(exu_n11809), .B(exu_n10644), .Y(bypass_dfill_data_g[46]));
INVX1 exu_U18769(.A(bypass_dfill_data_g[46]), .Y(exu_n4843));
AND2X1 exu_U18770(.A(exu_n11810), .B(exu_n10645), .Y(bypass_dfill_data_g[45]));
INVX1 exu_U18771(.A(bypass_dfill_data_g[45]), .Y(exu_n4844));
AND2X1 exu_U18772(.A(exu_n11811), .B(exu_n10646), .Y(bypass_dfill_data_g[44]));
INVX1 exu_U18773(.A(bypass_dfill_data_g[44]), .Y(exu_n4845));
AND2X1 exu_U18774(.A(exu_n11812), .B(exu_n10647), .Y(bypass_dfill_data_g[43]));
INVX1 exu_U18775(.A(bypass_dfill_data_g[43]), .Y(exu_n4846));
AND2X1 exu_U18776(.A(exu_n11813), .B(exu_n10648), .Y(bypass_dfill_data_g[42]));
INVX1 exu_U18777(.A(bypass_dfill_data_g[42]), .Y(exu_n4847));
AND2X1 exu_U18778(.A(exu_n11814), .B(exu_n10649), .Y(bypass_dfill_data_g[41]));
INVX1 exu_U18779(.A(bypass_dfill_data_g[41]), .Y(exu_n4848));
AND2X1 exu_U18780(.A(exu_n11815), .B(exu_n10650), .Y(bypass_dfill_data_g[40]));
INVX1 exu_U18781(.A(bypass_dfill_data_g[40]), .Y(exu_n4849));
AND2X1 exu_U18782(.A(exu_n11816), .B(exu_n10651), .Y(bypass_dfill_data_g[3]));
INVX1 exu_U18783(.A(bypass_dfill_data_g[3]), .Y(exu_n4850));
AND2X1 exu_U18784(.A(exu_n11817), .B(exu_n10652), .Y(bypass_dfill_data_g[39]));
INVX1 exu_U18785(.A(bypass_dfill_data_g[39]), .Y(exu_n4851));
AND2X1 exu_U18786(.A(exu_n11818), .B(exu_n10653), .Y(bypass_dfill_data_g[38]));
INVX1 exu_U18787(.A(bypass_dfill_data_g[38]), .Y(exu_n4852));
AND2X1 exu_U18788(.A(exu_n11819), .B(exu_n10654), .Y(bypass_dfill_data_g[37]));
INVX1 exu_U18789(.A(bypass_dfill_data_g[37]), .Y(exu_n4853));
AND2X1 exu_U18790(.A(exu_n11820), .B(exu_n10655), .Y(bypass_dfill_data_g[36]));
INVX1 exu_U18791(.A(bypass_dfill_data_g[36]), .Y(exu_n4854));
AND2X1 exu_U18792(.A(exu_n11821), .B(exu_n10656), .Y(bypass_dfill_data_g[35]));
INVX1 exu_U18793(.A(bypass_dfill_data_g[35]), .Y(exu_n4855));
AND2X1 exu_U18794(.A(exu_n11822), .B(exu_n10657), .Y(bypass_dfill_data_g[34]));
INVX1 exu_U18795(.A(bypass_dfill_data_g[34]), .Y(exu_n4856));
AND2X1 exu_U18796(.A(exu_n11823), .B(exu_n10658), .Y(bypass_dfill_data_g[33]));
INVX1 exu_U18797(.A(bypass_dfill_data_g[33]), .Y(exu_n4857));
AND2X1 exu_U18798(.A(exu_n11824), .B(exu_n10659), .Y(bypass_dfill_data_g[32]));
INVX1 exu_U18799(.A(bypass_dfill_data_g[32]), .Y(exu_n4858));
AND2X1 exu_U18800(.A(exu_n11825), .B(exu_n10660), .Y(bypass_dfill_data_g[31]));
INVX1 exu_U18801(.A(bypass_dfill_data_g[31]), .Y(exu_n4859));
AND2X1 exu_U18802(.A(exu_n11826), .B(exu_n10661), .Y(bypass_dfill_data_g[30]));
INVX1 exu_U18803(.A(bypass_dfill_data_g[30]), .Y(exu_n4860));
AND2X1 exu_U18804(.A(exu_n11827), .B(exu_n10662), .Y(bypass_dfill_data_g[2]));
INVX1 exu_U18805(.A(bypass_dfill_data_g[2]), .Y(exu_n4861));
AND2X1 exu_U18806(.A(exu_n11828), .B(exu_n10663), .Y(bypass_dfill_data_g[29]));
INVX1 exu_U18807(.A(bypass_dfill_data_g[29]), .Y(exu_n4862));
AND2X1 exu_U18808(.A(exu_n11829), .B(exu_n10664), .Y(bypass_dfill_data_g[28]));
INVX1 exu_U18809(.A(bypass_dfill_data_g[28]), .Y(exu_n4863));
AND2X1 exu_U18810(.A(exu_n11830), .B(exu_n10665), .Y(bypass_dfill_data_g[27]));
INVX1 exu_U18811(.A(bypass_dfill_data_g[27]), .Y(exu_n4864));
AND2X1 exu_U18812(.A(exu_n11831), .B(exu_n10666), .Y(bypass_dfill_data_g[26]));
INVX1 exu_U18813(.A(bypass_dfill_data_g[26]), .Y(exu_n4865));
AND2X1 exu_U18814(.A(exu_n11832), .B(exu_n10667), .Y(bypass_dfill_data_g[25]));
INVX1 exu_U18815(.A(bypass_dfill_data_g[25]), .Y(exu_n4866));
AND2X1 exu_U18816(.A(exu_n11833), .B(exu_n10668), .Y(bypass_dfill_data_g[24]));
INVX1 exu_U18817(.A(bypass_dfill_data_g[24]), .Y(exu_n4867));
AND2X1 exu_U18818(.A(exu_n11834), .B(exu_n10669), .Y(bypass_dfill_data_g[23]));
INVX1 exu_U18819(.A(bypass_dfill_data_g[23]), .Y(exu_n4868));
AND2X1 exu_U18820(.A(exu_n11835), .B(exu_n10670), .Y(bypass_dfill_data_g[22]));
INVX1 exu_U18821(.A(bypass_dfill_data_g[22]), .Y(exu_n4869));
AND2X1 exu_U18822(.A(exu_n11836), .B(exu_n10671), .Y(bypass_dfill_data_g[21]));
INVX1 exu_U18823(.A(bypass_dfill_data_g[21]), .Y(exu_n4870));
AND2X1 exu_U18824(.A(exu_n11837), .B(exu_n10672), .Y(bypass_dfill_data_g[20]));
INVX1 exu_U18825(.A(bypass_dfill_data_g[20]), .Y(exu_n4871));
AND2X1 exu_U18826(.A(exu_n11838), .B(exu_n10673), .Y(bypass_dfill_data_g[1]));
INVX1 exu_U18827(.A(bypass_dfill_data_g[1]), .Y(exu_n4872));
AND2X1 exu_U18828(.A(exu_n11839), .B(exu_n10674), .Y(bypass_dfill_data_g[19]));
INVX1 exu_U18829(.A(bypass_dfill_data_g[19]), .Y(exu_n4873));
AND2X1 exu_U18830(.A(exu_n11840), .B(exu_n10675), .Y(bypass_dfill_data_g[18]));
INVX1 exu_U18831(.A(bypass_dfill_data_g[18]), .Y(exu_n4874));
AND2X1 exu_U18832(.A(exu_n11841), .B(exu_n10676), .Y(bypass_dfill_data_g[17]));
INVX1 exu_U18833(.A(bypass_dfill_data_g[17]), .Y(exu_n4875));
AND2X1 exu_U18834(.A(exu_n11842), .B(exu_n10677), .Y(bypass_dfill_data_g[16]));
INVX1 exu_U18835(.A(bypass_dfill_data_g[16]), .Y(exu_n4876));
AND2X1 exu_U18836(.A(exu_n11843), .B(exu_n10678), .Y(bypass_dfill_data_g[15]));
INVX1 exu_U18837(.A(bypass_dfill_data_g[15]), .Y(exu_n4877));
AND2X1 exu_U18838(.A(exu_n11844), .B(exu_n10679), .Y(bypass_dfill_data_g[14]));
INVX1 exu_U18839(.A(bypass_dfill_data_g[14]), .Y(exu_n4878));
AND2X1 exu_U18840(.A(exu_n11845), .B(exu_n10680), .Y(bypass_dfill_data_g[13]));
INVX1 exu_U18841(.A(bypass_dfill_data_g[13]), .Y(exu_n4879));
AND2X1 exu_U18842(.A(exu_n11846), .B(exu_n10681), .Y(bypass_dfill_data_g[12]));
INVX1 exu_U18843(.A(bypass_dfill_data_g[12]), .Y(exu_n4880));
AND2X1 exu_U18844(.A(exu_n11847), .B(exu_n10682), .Y(bypass_dfill_data_g[11]));
INVX1 exu_U18845(.A(bypass_dfill_data_g[11]), .Y(exu_n4881));
AND2X1 exu_U18846(.A(exu_n11848), .B(exu_n10683), .Y(bypass_dfill_data_g[10]));
INVX1 exu_U18847(.A(bypass_dfill_data_g[10]), .Y(exu_n4882));
AND2X1 exu_U18848(.A(exu_n11849), .B(exu_n10684), .Y(bypass_dfill_data_g[0]));
INVX1 exu_U18849(.A(bypass_dfill_data_g[0]), .Y(exu_n4883));
AND2X1 exu_U18850(.A(exu_n11851), .B(exu_n15683), .Y(rml_n38));
INVX1 exu_U18851(.A(rml_n38), .Y(exu_n4884));
OR2X1 exu_U18852(.A(ifu_exu_saved_e), .B(ifu_exu_restored_e), .Y(rml_n60));
INVX1 exu_U18853(.A(rml_n60), .Y(exu_n4885));
AND2X1 exu_U18854(.A(rml_agp_thr1[1]), .B(exu_n9), .Y(rml_n64));
INVX1 exu_U18855(.A(rml_n64), .Y(exu_n4886));
AND2X1 exu_U18856(.A(rml_agp_thr3[1]), .B(rml_n70), .Y(rml_n68));
INVX1 exu_U18857(.A(rml_n68), .Y(exu_n4887));
AND2X1 exu_U18858(.A(rml_agp_thr1[0]), .B(exu_n9), .Y(rml_n73));
INVX1 exu_U18859(.A(rml_n73), .Y(exu_n4888));
AND2X1 exu_U18860(.A(rml_agp_thr3[0]), .B(rml_n70), .Y(rml_n75));
INVX1 exu_U18861(.A(rml_n75), .Y(exu_n4889));
OR2X1 exu_U18862(.A(exu_n9), .B(exu_n15470), .Y(rml_n78));
INVX1 exu_U18863(.A(rml_n78), .Y(exu_n4890));
AND2X1 exu_U18864(.A(exu_n11855), .B(exu_n10687), .Y(rml_oddwin_m[3]));
INVX1 exu_U18865(.A(rml_oddwin_m[3]), .Y(exu_n4891));
AND2X1 exu_U18866(.A(exu_n11856), .B(exu_n10689), .Y(rml_oddwin_m[2]));
INVX1 exu_U18867(.A(rml_oddwin_m[2]), .Y(exu_n4892));
AND2X1 exu_U18868(.A(exu_n11857), .B(exu_n10691), .Y(rml_oddwin_m[1]));
INVX1 exu_U18869(.A(rml_oddwin_m[1]), .Y(exu_n4893));
AND2X1 exu_U18870(.A(exu_n11858), .B(exu_n10693), .Y(rml_oddwin_m[0]));
INVX1 exu_U18871(.A(rml_oddwin_m[0]), .Y(exu_n4894));
OR2X1 exu_U18872(.A(rml_spill_m), .B(exu_n16605), .Y(rml_kill_restore_m));
INVX1 exu_U18873(.A(rml_kill_restore_m), .Y(exu_n4895));
OR2X1 exu_U18874(.A(ecl_rml_kill_e), .B(rml_n97), .Y(rml_cwp_wen_e));
INVX1 exu_U18875(.A(rml_cwp_wen_e), .Y(exu_n4896));
AND2X1 exu_U18876(.A(ifu_exu_restored_e), .B(exu_n16603), .Y(rml_n105));
INVX1 exu_U18877(.A(rml_n105), .Y(exu_n4897));
OR2X1 exu_U18878(.A(ecl_rml_kill_w), .B(exu_n14976), .Y(rml_n107));
INVX1 exu_U18879(.A(rml_n107), .Y(exu_n4898));
AND2X1 exu_U18880(.A(ifu_exu_saved_e), .B(exu_n16603), .Y(rml_n110));
INVX1 exu_U18881(.A(rml_n110), .Y(exu_n4899));
OR2X1 exu_U18882(.A(rml_n122), .B(rml_n123), .Y(rml_n115));
INVX1 exu_U18883(.A(rml_n115), .Y(exu_n4900));
AND2X1 exu_U18884(.A(rml_restore_e), .B(exu_n15344), .Y(rml_n111));
INVX1 exu_U18885(.A(rml_n111), .Y(exu_n4901));
OR2X1 exu_U18886(.A(rml_rml_ecl_canrestore_e[2]), .B(rml_rml_ecl_canrestore_e[1]), .Y(rml_n124));
INVX1 exu_U18887(.A(rml_n124), .Y(exu_n4902));
AND2X1 exu_U18888(.A(tlu_exu_agp_swap), .B(rml_agp_thr[3]), .Y(rml_n125));
INVX1 exu_U18889(.A(rml_n125), .Y(exu_n4903));
AND2X1 exu_U18890(.A(rml_agp_thr[2]), .B(tlu_exu_agp_swap), .Y(rml_n126));
INVX1 exu_U18891(.A(rml_n126), .Y(exu_n4904));
AND2X1 exu_U18892(.A(exu_n15439), .B(tlu_exu_agp_swap), .Y(rml_n127));
INVX1 exu_U18893(.A(rml_n127), .Y(exu_n4905));
AND2X1 exu_U18894(.A(exu_n15440), .B(tlu_exu_agp_swap), .Y(rml_n128));
INVX1 exu_U18895(.A(rml_n128), .Y(exu_n4906));
OR2X1 exu_U18896(.A(exu_n12034), .B(exu_n14922), .Y(div_n43));
INVX1 exu_U18897(.A(div_n43), .Y(exu_n4907));
OR2X1 exu_U18898(.A(exu_n12032), .B(exu_n14920), .Y(div_n45));
INVX1 exu_U18899(.A(div_n45), .Y(exu_n4908));
OR2X1 exu_U18900(.A(exu_n12070), .B(exu_n14979), .Y(div_n39));
INVX1 exu_U18901(.A(div_n39), .Y(exu_n4909));
OR2X1 exu_U18902(.A(exu_n12038), .B(exu_n14926), .Y(div_n49));
INVX1 exu_U18903(.A(div_n49), .Y(exu_n4910));
OR2X1 exu_U18904(.A(exu_n12036), .B(exu_n14924), .Y(div_n51));
INVX1 exu_U18905(.A(div_n51), .Y(exu_n4911));
OR2X1 exu_U18906(.A(exu_n12022), .B(exu_n14914), .Y(div_n57));
INVX1 exu_U18907(.A(div_n57), .Y(exu_n4912));
OR2X1 exu_U18908(.A(exu_n12008), .B(exu_n14896), .Y(div_n59));
INVX1 exu_U18909(.A(div_n59), .Y(exu_n4913));
OR2X1 exu_U18910(.A(exu_n12072), .B(exu_n14981), .Y(div_n53));
INVX1 exu_U18911(.A(div_n53), .Y(exu_n4914));
OR2X1 exu_U18912(.A(exu_n12030), .B(exu_n14918), .Y(div_n63));
INVX1 exu_U18913(.A(div_n63), .Y(exu_n4915));
OR2X1 exu_U18914(.A(exu_n12028), .B(exu_n14916), .Y(div_n65));
INVX1 exu_U18915(.A(div_n65), .Y(exu_n4916));
OR2X1 exu_U18916(.A(exu_n12021), .B(exu_n14909), .Y(div_n73));
INVX1 exu_U18917(.A(div_n73), .Y(exu_n4917));
OR2X1 exu_U18918(.A(exu_n12019), .B(exu_n14907), .Y(div_n75));
INVX1 exu_U18919(.A(div_n75), .Y(exu_n4918));
OR2X1 exu_U18920(.A(exu_n12074), .B(exu_n14983), .Y(div_n69));
INVX1 exu_U18921(.A(div_n69), .Y(exu_n4919));
OR2X1 exu_U18922(.A(exu_n12026), .B(exu_n14913), .Y(div_n79));
INVX1 exu_U18923(.A(div_n79), .Y(exu_n4920));
OR2X1 exu_U18924(.A(exu_n12024), .B(exu_n14911), .Y(div_n81));
INVX1 exu_U18925(.A(div_n81), .Y(exu_n4921));
OR2X1 exu_U18926(.A(exu_n12013), .B(exu_n14900), .Y(div_n87));
INVX1 exu_U18927(.A(div_n87), .Y(exu_n4922));
OR2X1 exu_U18928(.A(exu_n12010), .B(exu_n14898), .Y(div_n89));
INVX1 exu_U18929(.A(div_n89), .Y(exu_n4923));
OR2X1 exu_U18930(.A(exu_n12076), .B(exu_n14985), .Y(div_n83));
INVX1 exu_U18931(.A(div_n83), .Y(exu_n4924));
OR2X1 exu_U18932(.A(exu_n12017), .B(exu_n14905), .Y(div_n93));
INVX1 exu_U18933(.A(div_n93), .Y(exu_n4925));
OR2X1 exu_U18934(.A(exu_n12015), .B(exu_n14902), .Y(div_n95));
INVX1 exu_U18935(.A(div_n95), .Y(exu_n4926));
OR2X1 exu_U18936(.A(exu_n11986), .B(exu_n14875), .Y(alu_n75));
INVX1 exu_U18937(.A(alu_n75), .Y(exu_n4927));
OR2X1 exu_U18938(.A(exu_n11984), .B(exu_n14873), .Y(alu_n77));
INVX1 exu_U18939(.A(alu_n77), .Y(exu_n4928));
OR2X1 exu_U18940(.A(exu_n12078), .B(exu_n14987), .Y(alu_n71));
INVX1 exu_U18941(.A(alu_n71), .Y(exu_n4929));
OR2X1 exu_U18942(.A(exu_n11990), .B(exu_n14879), .Y(alu_n81));
INVX1 exu_U18943(.A(alu_n81), .Y(exu_n4930));
OR2X1 exu_U18944(.A(exu_n11988), .B(exu_n14877), .Y(alu_n83));
INVX1 exu_U18945(.A(alu_n83), .Y(exu_n4931));
OR2X1 exu_U18946(.A(exu_n11974), .B(exu_n14867), .Y(alu_n89));
INVX1 exu_U18947(.A(alu_n89), .Y(exu_n4932));
OR2X1 exu_U18948(.A(exu_n11960), .B(exu_n14849), .Y(alu_n91));
INVX1 exu_U18949(.A(alu_n91), .Y(exu_n4933));
OR2X1 exu_U18950(.A(exu_n12080), .B(exu_n14989), .Y(alu_n85));
INVX1 exu_U18951(.A(alu_n85), .Y(exu_n4934));
OR2X1 exu_U18952(.A(exu_n11982), .B(exu_n14871), .Y(alu_n95));
INVX1 exu_U18953(.A(alu_n95), .Y(exu_n4935));
OR2X1 exu_U18954(.A(exu_n11980), .B(exu_n14869), .Y(alu_n97));
INVX1 exu_U18955(.A(alu_n97), .Y(exu_n4936));
OR2X1 exu_U18956(.A(exu_n11973), .B(exu_n14862), .Y(alu_n105));
INVX1 exu_U18957(.A(alu_n105), .Y(exu_n4937));
OR2X1 exu_U18958(.A(exu_n11971), .B(exu_n14860), .Y(alu_n107));
INVX1 exu_U18959(.A(alu_n107), .Y(exu_n4938));
OR2X1 exu_U18960(.A(exu_n12082), .B(exu_n14992), .Y(alu_n101));
INVX1 exu_U18961(.A(alu_n101), .Y(exu_n4939));
OR2X1 exu_U18962(.A(exu_n11978), .B(exu_n14866), .Y(alu_n111));
INVX1 exu_U18963(.A(alu_n111), .Y(exu_n4940));
OR2X1 exu_U18964(.A(exu_n11976), .B(exu_n14864), .Y(alu_n113));
INVX1 exu_U18965(.A(alu_n113), .Y(exu_n4941));
OR2X1 exu_U18966(.A(exu_n11965), .B(exu_n14853), .Y(alu_n119));
INVX1 exu_U18967(.A(alu_n119), .Y(exu_n4942));
OR2X1 exu_U18968(.A(exu_n11962), .B(exu_n14851), .Y(alu_n121));
INVX1 exu_U18969(.A(alu_n121), .Y(exu_n4943));
OR2X1 exu_U18970(.A(exu_n12085), .B(exu_n14994), .Y(alu_n115));
INVX1 exu_U18971(.A(alu_n115), .Y(exu_n4944));
OR2X1 exu_U18972(.A(exu_n11969), .B(exu_n14858), .Y(alu_n125));
INVX1 exu_U18973(.A(alu_n125), .Y(exu_n4945));
OR2X1 exu_U18974(.A(exu_n11967), .B(exu_n14855), .Y(alu_n127));
INVX1 exu_U18975(.A(alu_n127), .Y(exu_n4946));
OR2X1 exu_U18976(.A(ecl_div_ecl_yreg_0_d), .B(exu_n16386), .Y(ecl_zero_rs2_d));
INVX1 exu_U18977(.A(ecl_zero_rs2_d), .Y(exu_n4947));
OR2X1 exu_U18978(.A(ecl_addr_mask_e), .B(exu_n16609), .Y(ecl_valid_range_check_jlret_e));
INVX1 exu_U18979(.A(ecl_valid_range_check_jlret_e), .Y(exu_n4948));
OR2X1 exu_U18980(.A(ifu_exu_rd_ffusr_e), .B(ifu_exu_rd_exusr_e), .Y(ecl_n45));
INVX1 exu_U18981(.A(ecl_n45), .Y(exu_n4949));
AND2X1 exu_U18982(.A(exu_n11922), .B(exu_n10697), .Y(ecl_perr_store_next[3]));
INVX1 exu_U18983(.A(ecl_perr_store_next[3]), .Y(exu_n4950));
AND2X1 exu_U18984(.A(exu_n11923), .B(exu_n10699), .Y(ecl_perr_store_next[2]));
INVX1 exu_U18985(.A(ecl_perr_store_next[2]), .Y(exu_n4951));
AND2X1 exu_U18986(.A(exu_n11924), .B(exu_n10701), .Y(ecl_perr_store_next[1]));
INVX1 exu_U18987(.A(ecl_perr_store_next[1]), .Y(exu_n4952));
AND2X1 exu_U18988(.A(exu_n11925), .B(exu_n10703), .Y(ecl_perr_store_next[0]));
INVX1 exu_U18989(.A(ecl_perr_store_next[0]), .Y(exu_n4953));
AND2X1 exu_U18990(.A(exu_n11926), .B(exu_n15212), .Y(ecl_part_early_flush_m));
INVX1 exu_U18991(.A(ecl_part_early_flush_m), .Y(exu_n4954));
AND2X1 exu_U18992(.A(exu_n11927), .B(exu_n10705), .Y(ecl_next_yreg_data_31));
INVX1 exu_U18993(.A(ecl_next_yreg_data_31), .Y(exu_n4955));
OR2X1 exu_U18994(.A(ecl_n65), .B(ecl_n66), .Y(ecl_ld_thr_match_sg_dff_din[0]));
INVX1 exu_U18995(.A(ecl_ld_thr_match_sg_dff_din[0]), .Y(exu_n4956));
OR2X1 exu_U18996(.A(ecl_n69), .B(exu_n16155), .Y(ecl_n67));
INVX1 exu_U18997(.A(ecl_n67), .Y(exu_n4957));
OR2X1 exu_U18998(.A(ecl_n70), .B(ecl_n71), .Y(ecl_thr_match_sd_dff_din[0]));
INVX1 exu_U18999(.A(ecl_thr_match_sd_dff_din[0]), .Y(exu_n4958));
OR2X1 exu_U19000(.A(ecl_n72), .B(ecl_n73), .Y(ecl_thr_match_se_dff_din[0]));
INVX1 exu_U19001(.A(ecl_thr_match_se_dff_din[0]), .Y(exu_n4959));
OR2X1 exu_U19002(.A(ecl_n74), .B(ecl_n75), .Y(ecl_thr_match_ew_dff_din[0]));
INVX1 exu_U19003(.A(ecl_thr_match_ew_dff_din[0]), .Y(exu_n4960));
OR2X1 exu_U19004(.A(ifu_exu_aluop_d[1]), .B(ifu_exu_aluop_d[0]), .Y(ecl_n77));
INVX1 exu_U19005(.A(ecl_n77), .Y(exu_n4961));
OR2X1 exu_U19006(.A(ecl_n79), .B(ecl_n80), .Y(ecl_ld_thr_match_sm_dff_din[0]));
INVX1 exu_U19007(.A(ecl_ld_thr_match_sm_dff_din[0]), .Y(exu_n4962));
AND2X1 exu_U19008(.A(ecl_n81), .B(exu_n15212), .Y(ecl_kill_rml_m));
INVX1 exu_U19009(.A(ecl_kill_rml_m), .Y(exu_n4963));
AND2X1 exu_U19010(.A(exu_n15922), .B(ecl_perr_store[2]), .Y(ecl_n86));
INVX1 exu_U19011(.A(ecl_n86), .Y(exu_n4964));
AND2X1 exu_U19012(.A(exu_n15924), .B(ecl_perr_store[0]), .Y(ecl_n99));
INVX1 exu_U19013(.A(ecl_n99), .Y(exu_n4965));
AND2X1 exu_U19014(.A(exu_tlu_misalign_addr_jmpl_rtn_m), .B(exu_n16403), .Y(ecl_n101));
INVX1 exu_U19015(.A(ecl_n101), .Y(exu_n4966));
OR2X1 exu_U19016(.A(ecl_ifu_exu_aluop_e[2]), .B(ecl_ifu_exu_aluop_e[1]), .Y(ecl_n123));
INVX1 exu_U19017(.A(ecl_n123), .Y(exu_n4967));
AND2X1 exu_U19018(.A(ifu_exu_dontmv_regz1_e), .B(exu_ifu_regz_e), .Y(ecl_n124));
INVX1 exu_U19019(.A(ecl_n124), .Y(exu_n4968));
AND2X1 exu_U19020(.A(exu_n11936), .B(exu_n10709), .Y(ecl_n130));
INVX1 exu_U19021(.A(ecl_n130), .Y(exu_n4969));
AND2X1 exu_U19022(.A(exu_n11939), .B(exu_n10710), .Y(ecl_n136));
INVX1 exu_U19023(.A(ecl_n136), .Y(exu_n4970));
AND2X1 exu_U19024(.A(exu_n11576), .B(exu_n10342), .Y(ecl_divcntl_inputs_neg_dff_n9));
INVX1 exu_U19025(.A(ecl_divcntl_inputs_neg_dff_n9), .Y(exu_n4971));
AND2X1 exu_U19026(.A(exu_n11585), .B(exu_n10349), .Y(ecl_writeback_restore_rd_dff_n23));
INVX1 exu_U19027(.A(ecl_writeback_restore_rd_dff_n23), .Y(exu_n4972));
AND2X1 exu_U19028(.A(exu_n11586), .B(exu_n10350), .Y(ecl_writeback_restore_rd_dff_n24));
INVX1 exu_U19029(.A(ecl_writeback_restore_rd_dff_n24), .Y(exu_n4973));
AND2X1 exu_U19030(.A(exu_n11587), .B(exu_n10351), .Y(ecl_writeback_restore_rd_dff_n25));
INVX1 exu_U19031(.A(ecl_writeback_restore_rd_dff_n25), .Y(exu_n4974));
AND2X1 exu_U19032(.A(exu_n11588), .B(exu_n10352), .Y(ecl_writeback_restore_rd_dff_n26));
INVX1 exu_U19033(.A(ecl_writeback_restore_rd_dff_n26), .Y(exu_n4975));
AND2X1 exu_U19034(.A(exu_n11589), .B(exu_n10353), .Y(ecl_writeback_restore_rd_dff_n27));
INVX1 exu_U19035(.A(ecl_writeback_restore_rd_dff_n27), .Y(exu_n4976));
AND2X1 exu_U19036(.A(exu_n11590), .B(exu_n10354), .Y(ecl_writeback_restore_tid_dff_n14));
INVX1 exu_U19037(.A(ecl_writeback_restore_tid_dff_n14), .Y(exu_n4977));
AND2X1 exu_U19038(.A(exu_n11591), .B(exu_n10355), .Y(ecl_writeback_restore_tid_dff_n15));
INVX1 exu_U19039(.A(ecl_writeback_restore_tid_dff_n15), .Y(exu_n4978));
AND2X1 exu_U19040(.A(exu_n10713), .B(exu_n9676), .Y(exu_n16633));
INVX1 exu_U19041(.A(exu_n16633), .Y(exu_n4979));
OR2X1 exu_U19042(.A(exu_n11940), .B(exu_n14822), .Y(ecl_byplog_rs1_N3));
INVX1 exu_U19043(.A(ecl_byplog_rs1_N3), .Y(exu_n4980));
AND2X1 exu_U19044(.A(exu_n10715), .B(exu_n9678), .Y(exu_n16647));
INVX1 exu_U19045(.A(exu_n16647), .Y(exu_n4981));
AND2X1 exu_U19046(.A(exu_n10717), .B(exu_n9680), .Y(exu_n16661));
INVX1 exu_U19047(.A(exu_n16661), .Y(exu_n4982));
AND2X1 exu_U19048(.A(exu_n10719), .B(exu_n9682), .Y(exu_n16675));
INVX1 exu_U19049(.A(exu_n16675), .Y(exu_n4983));
AND2X1 exu_U19050(.A(exu_n10721), .B(exu_n9684), .Y(exu_n16689));
INVX1 exu_U19051(.A(exu_n16689), .Y(exu_n4984));
OR2X1 exu_U19052(.A(exu_n11943), .B(exu_n14825), .Y(ecl_byplog_rs2_N3));
INVX1 exu_U19053(.A(ecl_byplog_rs2_N3), .Y(exu_n4985));
AND2X1 exu_U19054(.A(exu_n10723), .B(exu_n9686), .Y(exu_n16703));
INVX1 exu_U19055(.A(exu_n16703), .Y(exu_n4986));
AND2X1 exu_U19056(.A(exu_n10725), .B(exu_n9688), .Y(exu_n16717));
INVX1 exu_U19057(.A(exu_n16717), .Y(exu_n4987));
AND2X1 exu_U19058(.A(exu_n10727), .B(exu_n9690), .Y(exu_n16731));
INVX1 exu_U19059(.A(exu_n16731), .Y(exu_n4988));
AND2X1 exu_U19060(.A(exu_n15794), .B(exu_n16740), .Y(exu_n16741));
INVX1 exu_U19061(.A(exu_n16741), .Y(exu_n4989));
AND2X1 exu_U19062(.A(div_adderin2[1]), .B(exu_n16743), .Y(exu_n16744));
INVX1 exu_U19063(.A(exu_n16744), .Y(exu_n4990));
AND2X1 exu_U19064(.A(div_adderin2[2]), .B(exu_n16746), .Y(exu_n16747));
INVX1 exu_U19065(.A(exu_n16747), .Y(exu_n4991));
AND2X1 exu_U19066(.A(div_adderin2[3]), .B(exu_n16749), .Y(exu_n16750));
INVX1 exu_U19067(.A(exu_n16750), .Y(exu_n4992));
AND2X1 exu_U19068(.A(div_adderin2[4]), .B(exu_n16752), .Y(exu_n16753));
INVX1 exu_U19069(.A(exu_n16753), .Y(exu_n4993));
AND2X1 exu_U19070(.A(div_adderin2[5]), .B(exu_n16755), .Y(exu_n16756));
INVX1 exu_U19071(.A(exu_n16756), .Y(exu_n4994));
AND2X1 exu_U19072(.A(div_adderin2[6]), .B(exu_n16758), .Y(exu_n16759));
INVX1 exu_U19073(.A(exu_n16759), .Y(exu_n4995));
AND2X1 exu_U19074(.A(div_adderin2[7]), .B(exu_n16761), .Y(exu_n16762));
INVX1 exu_U19075(.A(exu_n16762), .Y(exu_n4996));
AND2X1 exu_U19076(.A(div_adderin2[8]), .B(exu_n16764), .Y(exu_n16765));
INVX1 exu_U19077(.A(exu_n16765), .Y(exu_n4997));
AND2X1 exu_U19078(.A(div_adderin2[9]), .B(exu_n16767), .Y(exu_n16768));
INVX1 exu_U19079(.A(exu_n16768), .Y(exu_n4998));
AND2X1 exu_U19080(.A(div_adderin2[10]), .B(exu_n16772), .Y(exu_n16773));
INVX1 exu_U19081(.A(exu_n16773), .Y(exu_n4999));
AND2X1 exu_U19082(.A(div_adderin2[11]), .B(exu_n16777), .Y(exu_n16778));
INVX1 exu_U19083(.A(exu_n16778), .Y(exu_n5000));
AND2X1 exu_U19084(.A(div_adderin2[12]), .B(exu_n16782), .Y(exu_n16783));
INVX1 exu_U19085(.A(exu_n16783), .Y(exu_n5001));
AND2X1 exu_U19086(.A(div_adderin2[13]), .B(exu_n16787), .Y(exu_n16788));
INVX1 exu_U19087(.A(exu_n16788), .Y(exu_n5002));
AND2X1 exu_U19088(.A(div_adderin2[14]), .B(exu_n16792), .Y(exu_n16793));
INVX1 exu_U19089(.A(exu_n16793), .Y(exu_n5003));
AND2X1 exu_U19090(.A(div_adderin2[15]), .B(exu_n16797), .Y(exu_n16798));
INVX1 exu_U19091(.A(exu_n16798), .Y(exu_n5004));
AND2X1 exu_U19092(.A(div_adderin2[16]), .B(exu_n16802), .Y(exu_n16803));
INVX1 exu_U19093(.A(exu_n16803), .Y(exu_n5005));
AND2X1 exu_U19094(.A(div_adderin2[17]), .B(exu_n16807), .Y(exu_n16808));
INVX1 exu_U19095(.A(exu_n16808), .Y(exu_n5006));
AND2X1 exu_U19096(.A(div_adderin2[18]), .B(exu_n16812), .Y(exu_n16813));
INVX1 exu_U19097(.A(exu_n16813), .Y(exu_n5007));
AND2X1 exu_U19098(.A(div_adderin2[19]), .B(exu_n16819), .Y(exu_n16820));
INVX1 exu_U19099(.A(exu_n16820), .Y(exu_n5008));
AND2X1 exu_U19100(.A(div_adderin2[20]), .B(exu_n16824), .Y(exu_n16825));
INVX1 exu_U19101(.A(exu_n16825), .Y(exu_n5009));
AND2X1 exu_U19102(.A(div_adderin2[21]), .B(exu_n16829), .Y(exu_n16830));
INVX1 exu_U19103(.A(exu_n16830), .Y(exu_n5010));
AND2X1 exu_U19104(.A(div_adderin2[22]), .B(exu_n16834), .Y(exu_n16835));
INVX1 exu_U19105(.A(exu_n16835), .Y(exu_n5011));
AND2X1 exu_U19106(.A(div_adderin2[23]), .B(exu_n16839), .Y(exu_n16840));
INVX1 exu_U19107(.A(exu_n16840), .Y(exu_n5012));
AND2X1 exu_U19108(.A(div_adderin2[24]), .B(exu_n16844), .Y(exu_n16845));
INVX1 exu_U19109(.A(exu_n16845), .Y(exu_n5013));
AND2X1 exu_U19110(.A(div_adderin2[25]), .B(exu_n16849), .Y(exu_n16850));
INVX1 exu_U19111(.A(exu_n16850), .Y(exu_n5014));
AND2X1 exu_U19112(.A(div_adderin2[26]), .B(exu_n16854), .Y(exu_n16855));
INVX1 exu_U19113(.A(exu_n16855), .Y(exu_n5015));
AND2X1 exu_U19114(.A(div_adderin2[27]), .B(exu_n16859), .Y(exu_n16860));
INVX1 exu_U19115(.A(exu_n16860), .Y(exu_n5016));
AND2X1 exu_U19116(.A(div_adderin2[28]), .B(exu_n16864), .Y(exu_n16865));
INVX1 exu_U19117(.A(exu_n16865), .Y(exu_n5017));
AND2X1 exu_U19118(.A(div_adderin2[29]), .B(exu_n16871), .Y(exu_n16872));
INVX1 exu_U19119(.A(exu_n16872), .Y(exu_n5018));
AND2X1 exu_U19120(.A(div_adderin2[30]), .B(exu_n16876), .Y(exu_n16877));
INVX1 exu_U19121(.A(exu_n16877), .Y(exu_n5019));
AND2X1 exu_U19122(.A(div_adderin2[31]), .B(exu_n16881), .Y(exu_n16882));
INVX1 exu_U19123(.A(exu_n16882), .Y(exu_n5020));
AND2X1 exu_U19124(.A(exu_n15558), .B(exu_n16899), .Y(exu_n16900));
INVX1 exu_U19125(.A(exu_n16900), .Y(exu_n5021));
AND2X1 exu_U19126(.A(div_adderin2[33]), .B(exu_n16902), .Y(exu_n16903));
INVX1 exu_U19127(.A(exu_n16903), .Y(exu_n5022));
AND2X1 exu_U19128(.A(div_adderin2[34]), .B(exu_n16905), .Y(exu_n16906));
INVX1 exu_U19129(.A(exu_n16906), .Y(exu_n5023));
AND2X1 exu_U19130(.A(div_adderin2[35]), .B(exu_n16908), .Y(exu_n16909));
INVX1 exu_U19131(.A(exu_n16909), .Y(exu_n5024));
AND2X1 exu_U19132(.A(div_adderin2[36]), .B(exu_n16911), .Y(exu_n16912));
INVX1 exu_U19133(.A(exu_n16912), .Y(exu_n5025));
AND2X1 exu_U19134(.A(div_adderin2[37]), .B(exu_n16914), .Y(exu_n16915));
INVX1 exu_U19135(.A(exu_n16915), .Y(exu_n5026));
AND2X1 exu_U19136(.A(div_adderin2[38]), .B(exu_n16917), .Y(exu_n16918));
INVX1 exu_U19137(.A(exu_n16918), .Y(exu_n5027));
AND2X1 exu_U19138(.A(div_adderin2[39]), .B(exu_n16920), .Y(exu_n16921));
INVX1 exu_U19139(.A(exu_n16921), .Y(exu_n5028));
AND2X1 exu_U19140(.A(div_adderin2[40]), .B(exu_n16923), .Y(exu_n16924));
INVX1 exu_U19141(.A(exu_n16924), .Y(exu_n5029));
AND2X1 exu_U19142(.A(div_adderin2[41]), .B(exu_n16926), .Y(exu_n16927));
INVX1 exu_U19143(.A(exu_n16927), .Y(exu_n5030));
AND2X1 exu_U19144(.A(div_adderin2[42]), .B(exu_n16931), .Y(exu_n16932));
INVX1 exu_U19145(.A(exu_n16932), .Y(exu_n5031));
AND2X1 exu_U19146(.A(div_adderin2[43]), .B(exu_n16936), .Y(exu_n16937));
INVX1 exu_U19147(.A(exu_n16937), .Y(exu_n5032));
AND2X1 exu_U19148(.A(div_adderin2[44]), .B(exu_n16941), .Y(exu_n16942));
INVX1 exu_U19149(.A(exu_n16942), .Y(exu_n5033));
AND2X1 exu_U19150(.A(div_adderin2[45]), .B(exu_n16946), .Y(exu_n16947));
INVX1 exu_U19151(.A(exu_n16947), .Y(exu_n5034));
AND2X1 exu_U19152(.A(div_adderin2[46]), .B(exu_n16951), .Y(exu_n16952));
INVX1 exu_U19153(.A(exu_n16952), .Y(exu_n5035));
AND2X1 exu_U19154(.A(div_adderin2[47]), .B(exu_n16956), .Y(exu_n16957));
INVX1 exu_U19155(.A(exu_n16957), .Y(exu_n5036));
AND2X1 exu_U19156(.A(div_adderin2[48]), .B(exu_n16961), .Y(exu_n16962));
INVX1 exu_U19157(.A(exu_n16962), .Y(exu_n5037));
AND2X1 exu_U19158(.A(div_adderin2[49]), .B(exu_n16966), .Y(exu_n16967));
INVX1 exu_U19159(.A(exu_n16967), .Y(exu_n5038));
AND2X1 exu_U19160(.A(div_adderin2[50]), .B(exu_n16971), .Y(exu_n16972));
INVX1 exu_U19161(.A(exu_n16972), .Y(exu_n5039));
AND2X1 exu_U19162(.A(div_adderin2[51]), .B(exu_n16978), .Y(exu_n16979));
INVX1 exu_U19163(.A(exu_n16979), .Y(exu_n5040));
AND2X1 exu_U19164(.A(div_adderin2[52]), .B(exu_n16983), .Y(exu_n16984));
INVX1 exu_U19165(.A(exu_n16984), .Y(exu_n5041));
AND2X1 exu_U19166(.A(div_adderin2[53]), .B(exu_n16988), .Y(exu_n16989));
INVX1 exu_U19167(.A(exu_n16989), .Y(exu_n5042));
AND2X1 exu_U19168(.A(div_adderin2[54]), .B(exu_n16993), .Y(exu_n16994));
INVX1 exu_U19169(.A(exu_n16994), .Y(exu_n5043));
AND2X1 exu_U19170(.A(div_adderin2[55]), .B(exu_n16998), .Y(exu_n16999));
INVX1 exu_U19171(.A(exu_n16999), .Y(exu_n5044));
AND2X1 exu_U19172(.A(div_adderin2[56]), .B(exu_n17003), .Y(exu_n17004));
INVX1 exu_U19173(.A(exu_n17004), .Y(exu_n5045));
AND2X1 exu_U19174(.A(div_adderin2[57]), .B(exu_n17008), .Y(exu_n17009));
INVX1 exu_U19175(.A(exu_n17009), .Y(exu_n5046));
AND2X1 exu_U19176(.A(div_adderin2[58]), .B(exu_n17013), .Y(exu_n17014));
INVX1 exu_U19177(.A(exu_n17014), .Y(exu_n5047));
AND2X1 exu_U19178(.A(div_adderin2[59]), .B(exu_n17018), .Y(exu_n17019));
INVX1 exu_U19179(.A(exu_n17019), .Y(exu_n5048));
AND2X1 exu_U19180(.A(div_adderin2[60]), .B(exu_n17023), .Y(exu_n17024));
INVX1 exu_U19181(.A(exu_n17024), .Y(exu_n5049));
AND2X1 exu_U19182(.A(div_adderin2[61]), .B(exu_n17030), .Y(exu_n17031));
INVX1 exu_U19183(.A(exu_n17031), .Y(exu_n5050));
AND2X1 exu_U19184(.A(div_adderin2[62]), .B(exu_n17035), .Y(exu_n17036));
INVX1 exu_U19185(.A(exu_n17036), .Y(exu_n5051));
AND2X1 exu_U19186(.A(div_adderin2[63]), .B(exu_n17040), .Y(exu_n17041));
INVX1 exu_U19187(.A(exu_n17041), .Y(exu_n5052));
AND2X1 exu_U19188(.A(ecl_alu_cin_e), .B(exu_n17058), .Y(exu_n17059));
INVX1 exu_U19189(.A(exu_n17059), .Y(exu_n5053));
AND2X1 exu_U19190(.A(alu_addsub_rs2_data_1), .B(exu_n17061), .Y(exu_n17062));
INVX1 exu_U19191(.A(exu_n17062), .Y(exu_n5054));
AND2X1 exu_U19192(.A(alu_addsub_rs2_data_2), .B(exu_n17064), .Y(exu_n17065));
INVX1 exu_U19193(.A(exu_n17065), .Y(exu_n5055));
AND2X1 exu_U19194(.A(alu_addsub_rs2_data_3), .B(exu_n17067), .Y(exu_n17068));
INVX1 exu_U19195(.A(exu_n17068), .Y(exu_n5056));
AND2X1 exu_U19196(.A(alu_addsub_rs2_data_4), .B(exu_n17070), .Y(exu_n17071));
INVX1 exu_U19197(.A(exu_n17071), .Y(exu_n5057));
AND2X1 exu_U19198(.A(alu_addsub_rs2_data_5), .B(exu_n17073), .Y(exu_n17074));
INVX1 exu_U19199(.A(exu_n17074), .Y(exu_n5058));
AND2X1 exu_U19200(.A(alu_addsub_rs2_data_6), .B(exu_n17076), .Y(exu_n17077));
INVX1 exu_U19201(.A(exu_n17077), .Y(exu_n5059));
AND2X1 exu_U19202(.A(alu_addsub_rs2_data_7), .B(exu_n17079), .Y(exu_n17080));
INVX1 exu_U19203(.A(exu_n17080), .Y(exu_n5060));
AND2X1 exu_U19204(.A(alu_addsub_rs2_data_8), .B(exu_n17082), .Y(exu_n17083));
INVX1 exu_U19205(.A(exu_n17083), .Y(exu_n5061));
AND2X1 exu_U19206(.A(alu_addsub_rs2_data_9), .B(exu_n17085), .Y(exu_n17086));
INVX1 exu_U19207(.A(exu_n17086), .Y(exu_n5062));
AND2X1 exu_U19208(.A(alu_addsub_rs2_data_10), .B(exu_n17090), .Y(exu_n17091));
INVX1 exu_U19209(.A(exu_n17091), .Y(exu_n5063));
AND2X1 exu_U19210(.A(alu_addsub_rs2_data_11), .B(exu_n17095), .Y(exu_n17096));
INVX1 exu_U19211(.A(exu_n17096), .Y(exu_n5064));
AND2X1 exu_U19212(.A(alu_addsub_rs2_data_12), .B(exu_n17100), .Y(exu_n17101));
INVX1 exu_U19213(.A(exu_n17101), .Y(exu_n5065));
AND2X1 exu_U19214(.A(alu_addsub_rs2_data_13), .B(exu_n17105), .Y(exu_n17106));
INVX1 exu_U19215(.A(exu_n17106), .Y(exu_n5066));
AND2X1 exu_U19216(.A(alu_addsub_rs2_data_14), .B(exu_n17110), .Y(exu_n17111));
INVX1 exu_U19217(.A(exu_n17111), .Y(exu_n5067));
AND2X1 exu_U19218(.A(alu_addsub_rs2_data_15), .B(exu_n17115), .Y(exu_n17116));
INVX1 exu_U19219(.A(exu_n17116), .Y(exu_n5068));
AND2X1 exu_U19220(.A(alu_addsub_rs2_data_16), .B(exu_n17120), .Y(exu_n17121));
INVX1 exu_U19221(.A(exu_n17121), .Y(exu_n5069));
AND2X1 exu_U19222(.A(alu_addsub_rs2_data_17), .B(exu_n17125), .Y(exu_n17126));
INVX1 exu_U19223(.A(exu_n17126), .Y(exu_n5070));
AND2X1 exu_U19224(.A(alu_addsub_rs2_data_18), .B(exu_n17130), .Y(exu_n17131));
INVX1 exu_U19225(.A(exu_n17131), .Y(exu_n5071));
AND2X1 exu_U19226(.A(alu_addsub_rs2_data_19), .B(exu_n17137), .Y(exu_n17138));
INVX1 exu_U19227(.A(exu_n17138), .Y(exu_n5072));
AND2X1 exu_U19228(.A(alu_addsub_rs2_data_20), .B(exu_n17142), .Y(exu_n17143));
INVX1 exu_U19229(.A(exu_n17143), .Y(exu_n5073));
AND2X1 exu_U19230(.A(alu_addsub_rs2_data_21), .B(exu_n17147), .Y(exu_n17148));
INVX1 exu_U19231(.A(exu_n17148), .Y(exu_n5074));
AND2X1 exu_U19232(.A(alu_addsub_rs2_data_22), .B(exu_n17152), .Y(exu_n17153));
INVX1 exu_U19233(.A(exu_n17153), .Y(exu_n5075));
AND2X1 exu_U19234(.A(alu_addsub_rs2_data_23), .B(exu_n17157), .Y(exu_n17158));
INVX1 exu_U19235(.A(exu_n17158), .Y(exu_n5076));
AND2X1 exu_U19236(.A(alu_addsub_rs2_data_24), .B(exu_n17162), .Y(exu_n17163));
INVX1 exu_U19237(.A(exu_n17163), .Y(exu_n5077));
AND2X1 exu_U19238(.A(alu_addsub_rs2_data_25), .B(exu_n17167), .Y(exu_n17168));
INVX1 exu_U19239(.A(exu_n17168), .Y(exu_n5078));
AND2X1 exu_U19240(.A(alu_addsub_rs2_data_26), .B(exu_n17172), .Y(exu_n17173));
INVX1 exu_U19241(.A(exu_n17173), .Y(exu_n5079));
AND2X1 exu_U19242(.A(alu_addsub_rs2_data_27), .B(exu_n17177), .Y(exu_n17178));
INVX1 exu_U19243(.A(exu_n17178), .Y(exu_n5080));
AND2X1 exu_U19244(.A(alu_addsub_rs2_data_28), .B(exu_n17182), .Y(exu_n17183));
INVX1 exu_U19245(.A(exu_n17183), .Y(exu_n5081));
AND2X1 exu_U19246(.A(alu_addsub_rs2_data_29), .B(exu_n17189), .Y(exu_n17190));
INVX1 exu_U19247(.A(exu_n17190), .Y(exu_n5082));
AND2X1 exu_U19248(.A(alu_addsub_rs2_data_30), .B(exu_n17194), .Y(exu_n17195));
INVX1 exu_U19249(.A(exu_n17195), .Y(exu_n5083));
AND2X1 exu_U19250(.A(alu_ecl_adderin2_31_e), .B(exu_n17199), .Y(exu_n17200));
INVX1 exu_U19251(.A(exu_n17200), .Y(exu_n5084));
AND2X1 exu_U19252(.A(exu_n15795), .B(exu_n17217), .Y(exu_n17218));
INVX1 exu_U19253(.A(exu_n17218), .Y(exu_n5085));
AND2X1 exu_U19254(.A(alu_addsub_rs2_data[33]), .B(exu_n17220), .Y(exu_n17221));
INVX1 exu_U19255(.A(exu_n17221), .Y(exu_n5086));
AND2X1 exu_U19256(.A(alu_addsub_rs2_data[34]), .B(exu_n17223), .Y(exu_n17224));
INVX1 exu_U19257(.A(exu_n17224), .Y(exu_n5087));
AND2X1 exu_U19258(.A(alu_addsub_rs2_data[35]), .B(exu_n17226), .Y(exu_n17227));
INVX1 exu_U19259(.A(exu_n17227), .Y(exu_n5088));
AND2X1 exu_U19260(.A(alu_addsub_rs2_data[36]), .B(exu_n17229), .Y(exu_n17230));
INVX1 exu_U19261(.A(exu_n17230), .Y(exu_n5089));
AND2X1 exu_U19262(.A(alu_addsub_rs2_data[37]), .B(exu_n17232), .Y(exu_n17233));
INVX1 exu_U19263(.A(exu_n17233), .Y(exu_n5090));
AND2X1 exu_U19264(.A(alu_addsub_rs2_data[38]), .B(exu_n17235), .Y(exu_n17236));
INVX1 exu_U19265(.A(exu_n17236), .Y(exu_n5091));
AND2X1 exu_U19266(.A(alu_addsub_rs2_data[39]), .B(exu_n17238), .Y(exu_n17239));
INVX1 exu_U19267(.A(exu_n17239), .Y(exu_n5092));
AND2X1 exu_U19268(.A(alu_addsub_rs2_data[40]), .B(exu_n17241), .Y(exu_n17242));
INVX1 exu_U19269(.A(exu_n17242), .Y(exu_n5093));
AND2X1 exu_U19270(.A(alu_addsub_rs2_data[41]), .B(exu_n17244), .Y(exu_n17245));
INVX1 exu_U19271(.A(exu_n17245), .Y(exu_n5094));
AND2X1 exu_U19272(.A(alu_addsub_rs2_data[42]), .B(exu_n17249), .Y(exu_n17250));
INVX1 exu_U19273(.A(exu_n17250), .Y(exu_n5095));
AND2X1 exu_U19274(.A(alu_addsub_rs2_data[43]), .B(exu_n17254), .Y(exu_n17255));
INVX1 exu_U19275(.A(exu_n17255), .Y(exu_n5096));
AND2X1 exu_U19276(.A(alu_addsub_rs2_data[44]), .B(exu_n17259), .Y(exu_n17260));
INVX1 exu_U19277(.A(exu_n17260), .Y(exu_n5097));
AND2X1 exu_U19278(.A(alu_addsub_rs2_data[45]), .B(exu_n17264), .Y(exu_n17265));
INVX1 exu_U19279(.A(exu_n17265), .Y(exu_n5098));
AND2X1 exu_U19280(.A(alu_addsub_rs2_data[46]), .B(exu_n17269), .Y(exu_n17270));
INVX1 exu_U19281(.A(exu_n17270), .Y(exu_n5099));
AND2X1 exu_U19282(.A(alu_addsub_rs2_data[47]), .B(exu_n17274), .Y(exu_n17275));
INVX1 exu_U19283(.A(exu_n17275), .Y(exu_n5100));
AND2X1 exu_U19284(.A(alu_addsub_rs2_data[48]), .B(exu_n17279), .Y(exu_n17280));
INVX1 exu_U19285(.A(exu_n17280), .Y(exu_n5101));
AND2X1 exu_U19286(.A(alu_addsub_rs2_data[49]), .B(exu_n17284), .Y(exu_n17285));
INVX1 exu_U19287(.A(exu_n17285), .Y(exu_n5102));
AND2X1 exu_U19288(.A(alu_addsub_rs2_data[50]), .B(exu_n17289), .Y(exu_n17290));
INVX1 exu_U19289(.A(exu_n17290), .Y(exu_n5103));
AND2X1 exu_U19290(.A(alu_addsub_rs2_data[51]), .B(exu_n17296), .Y(exu_n17297));
INVX1 exu_U19291(.A(exu_n17297), .Y(exu_n5104));
AND2X1 exu_U19292(.A(alu_addsub_rs2_data[52]), .B(exu_n17301), .Y(exu_n17302));
INVX1 exu_U19293(.A(exu_n17302), .Y(exu_n5105));
AND2X1 exu_U19294(.A(alu_addsub_rs2_data[53]), .B(exu_n17306), .Y(exu_n17307));
INVX1 exu_U19295(.A(exu_n17307), .Y(exu_n5106));
AND2X1 exu_U19296(.A(alu_addsub_rs2_data[54]), .B(exu_n17311), .Y(exu_n17312));
INVX1 exu_U19297(.A(exu_n17312), .Y(exu_n5107));
AND2X1 exu_U19298(.A(alu_addsub_rs2_data[55]), .B(exu_n17316), .Y(exu_n17317));
INVX1 exu_U19299(.A(exu_n17317), .Y(exu_n5108));
AND2X1 exu_U19300(.A(alu_addsub_rs2_data[56]), .B(exu_n17321), .Y(exu_n17322));
INVX1 exu_U19301(.A(exu_n17322), .Y(exu_n5109));
AND2X1 exu_U19302(.A(alu_addsub_rs2_data[57]), .B(exu_n17326), .Y(exu_n17327));
INVX1 exu_U19303(.A(exu_n17327), .Y(exu_n5110));
AND2X1 exu_U19304(.A(alu_addsub_rs2_data[58]), .B(exu_n17331), .Y(exu_n17332));
INVX1 exu_U19305(.A(exu_n17332), .Y(exu_n5111));
AND2X1 exu_U19306(.A(alu_addsub_rs2_data[59]), .B(exu_n17336), .Y(exu_n17337));
INVX1 exu_U19307(.A(exu_n17337), .Y(exu_n5112));
AND2X1 exu_U19308(.A(alu_addsub_rs2_data[60]), .B(exu_n17341), .Y(exu_n17342));
INVX1 exu_U19309(.A(exu_n17342), .Y(exu_n5113));
AND2X1 exu_U19310(.A(alu_addsub_rs2_data[61]), .B(exu_n17348), .Y(exu_n17349));
INVX1 exu_U19311(.A(exu_n17349), .Y(exu_n5114));
AND2X1 exu_U19312(.A(alu_addsub_rs2_data[62]), .B(exu_n17353), .Y(exu_n17354));
INVX1 exu_U19313(.A(exu_n17354), .Y(exu_n5115));
AND2X1 exu_U19314(.A(alu_ecl_adderin2_63_e), .B(exu_n17358), .Y(exu_n17359));
INVX1 exu_U19315(.A(exu_n17359), .Y(exu_n5116));
OR2X1 exu_U19316(.A(exu_n11946), .B(exu_n14828), .Y(ecl_byplog_rs3h_N3));
INVX1 exu_U19317(.A(ecl_byplog_rs3h_N3), .Y(exu_n5117));
AND2X1 exu_U19318(.A(exu_n10729), .B(exu_n9692), .Y(exu_n17409));
INVX1 exu_U19319(.A(exu_n17409), .Y(exu_n5118));
OR2X1 exu_U19320(.A(exu_n11949), .B(exu_n14831), .Y(ecl_byplog_rs3_N3));
INVX1 exu_U19321(.A(ecl_byplog_rs3_N3), .Y(exu_n5119));
AND2X1 exu_U19322(.A(exu_n10731), .B(exu_n9694), .Y(exu_n17423));
INVX1 exu_U19323(.A(exu_n17423), .Y(exu_n5120));
AND2X1 exu_U19324(.A(exu_n10733), .B(exu_n9696), .Y(exu_n17437));
INVX1 exu_U19325(.A(exu_n17437), .Y(exu_n5121));
AND2X1 exu_U19326(.A(exu_n10735), .B(exu_n9698), .Y(exu_n17451));
INVX1 exu_U19327(.A(exu_n17451), .Y(exu_n5122));
AND2X1 exu_U19328(.A(exu_n15851), .B(rml_cwp_n37), .Y(exu_n17516));
INVX1 exu_U19329(.A(exu_n17516), .Y(exu_n5123));
AND2X1 exu_U19330(.A(exu_n15852), .B(rml_cwp_n37), .Y(exu_n17520));
INVX1 exu_U19331(.A(exu_n17520), .Y(exu_n5124));
AND2X1 exu_U19332(.A(exu_n15853), .B(rml_cwp_n37), .Y(exu_n17524));
INVX1 exu_U19333(.A(exu_n17524), .Y(exu_n5125));
AND2X1 exu_U19334(.A(rml_rml_ecl_cwp_e[2]), .B(rml_cwp_n37), .Y(exu_n17528));
INVX1 exu_U19335(.A(exu_n17528), .Y(exu_n5126));
AND2X1 exu_U19336(.A(rml_rml_ecl_cwp_e[1]), .B(rml_cwp_n37), .Y(exu_n17532));
INVX1 exu_U19337(.A(exu_n17532), .Y(exu_n5127));
AND2X1 exu_U19338(.A(rml_rml_ecl_cwp_e[0]), .B(rml_cwp_n37), .Y(exu_n17542));
INVX1 exu_U19339(.A(exu_n17542), .Y(exu_n5128));
AND2X1 exu_U19340(.A(exu_n15851), .B(rml_cwp_n36), .Y(exu_n17553));
INVX1 exu_U19341(.A(exu_n17553), .Y(exu_n5129));
AND2X1 exu_U19342(.A(exu_n15852), .B(rml_cwp_n36), .Y(exu_n17557));
INVX1 exu_U19343(.A(exu_n17557), .Y(exu_n5130));
AND2X1 exu_U19344(.A(exu_n15853), .B(rml_cwp_n36), .Y(exu_n17561));
INVX1 exu_U19345(.A(exu_n17561), .Y(exu_n5131));
AND2X1 exu_U19346(.A(rml_rml_ecl_cwp_e[2]), .B(rml_cwp_n36), .Y(exu_n17565));
INVX1 exu_U19347(.A(exu_n17565), .Y(exu_n5132));
AND2X1 exu_U19348(.A(rml_rml_ecl_cwp_e[1]), .B(rml_cwp_n36), .Y(exu_n17569));
INVX1 exu_U19349(.A(exu_n17569), .Y(exu_n5133));
AND2X1 exu_U19350(.A(rml_rml_ecl_cwp_e[0]), .B(rml_cwp_n36), .Y(exu_n17579));
INVX1 exu_U19351(.A(exu_n17579), .Y(exu_n5134));
AND2X1 exu_U19352(.A(exu_n15851), .B(rml_cwp_n35), .Y(exu_n17590));
INVX1 exu_U19353(.A(exu_n17590), .Y(exu_n5135));
AND2X1 exu_U19354(.A(exu_n15852), .B(rml_cwp_n35), .Y(exu_n17594));
INVX1 exu_U19355(.A(exu_n17594), .Y(exu_n5136));
AND2X1 exu_U19356(.A(exu_n15853), .B(rml_cwp_n35), .Y(exu_n17598));
INVX1 exu_U19357(.A(exu_n17598), .Y(exu_n5137));
AND2X1 exu_U19358(.A(rml_rml_ecl_cwp_e[2]), .B(rml_cwp_n35), .Y(exu_n17602));
INVX1 exu_U19359(.A(exu_n17602), .Y(exu_n5138));
AND2X1 exu_U19360(.A(rml_rml_ecl_cwp_e[1]), .B(rml_cwp_n35), .Y(exu_n17606));
INVX1 exu_U19361(.A(exu_n17606), .Y(exu_n5139));
AND2X1 exu_U19362(.A(rml_rml_ecl_cwp_e[0]), .B(rml_cwp_n35), .Y(exu_n17616));
INVX1 exu_U19363(.A(exu_n17616), .Y(exu_n5140));
OR2X1 exu_U19364(.A(exu_n11952), .B(exu_n14834), .Y(exu_n17627));
INVX1 exu_U19365(.A(exu_n17627), .Y(exu_n5141));
OR2X1 exu_U19366(.A(exu_n11953), .B(exu_n14836), .Y(exu_n17639));
INVX1 exu_U19367(.A(exu_n17639), .Y(exu_n5142));
OR2X1 exu_U19368(.A(exu_n11954), .B(exu_n14838), .Y(exu_n17651));
INVX1 exu_U19369(.A(exu_n17651), .Y(exu_n5143));
OR2X1 exu_U19370(.A(exu_n11955), .B(exu_n14840), .Y(exu_n17663));
INVX1 exu_U19371(.A(exu_n17663), .Y(exu_n5144));
OR2X1 exu_U19372(.A(exu_n11956), .B(exu_n14842), .Y(exu_n17675));
INVX1 exu_U19373(.A(exu_n17675), .Y(exu_n5145));
OR2X1 exu_U19374(.A(exu_n11957), .B(exu_n14844), .Y(exu_n17687));
INVX1 exu_U19375(.A(exu_n17687), .Y(exu_n5146));
OR2X1 exu_U19376(.A(exu_n11958), .B(exu_n14846), .Y(exu_n17698));
INVX1 exu_U19377(.A(exu_n17698), .Y(exu_n5147));
AND2X1 exu_U19378(.A(ecl_ecc_log_rs3_m), .B(ecl_ifu_exu_rs3_m[4]), .Y(exu_n17709));
INVX1 exu_U19379(.A(exu_n17709), .Y(exu_n5148));
AND2X1 exu_U19380(.A(exu_n15028), .B(ecl_ifu_exu_rs1_m[4]), .Y(exu_n17711));
INVX1 exu_U19381(.A(exu_n17711), .Y(exu_n5149));
AND2X1 exu_U19382(.A(ecl_ifu_exu_rs3_m[3]), .B(ecl_ecc_log_rs3_m), .Y(exu_n17713));
INVX1 exu_U19383(.A(exu_n17713), .Y(exu_n5150));
AND2X1 exu_U19384(.A(ecl_ifu_exu_rs1_m[3]), .B(exu_n15028), .Y(exu_n17715));
INVX1 exu_U19385(.A(exu_n17715), .Y(exu_n5151));
AND2X1 exu_U19386(.A(ecl_ifu_exu_rs1_m[2]), .B(exu_n15028), .Y(exu_n17719));
INVX1 exu_U19387(.A(exu_n17719), .Y(exu_n5152));
AND2X1 exu_U19388(.A(ecl_ifu_exu_rs1_m[1]), .B(exu_n15028), .Y(exu_n17723));
INVX1 exu_U19389(.A(exu_n17723), .Y(exu_n5153));
AND2X1 exu_U19390(.A(ecl_ifu_exu_rs1_m[0]), .B(exu_n15028), .Y(exu_n17727));
INVX1 exu_U19391(.A(exu_n17727), .Y(exu_n5154));
AND2X1 exu_U19392(.A(ecl_rml_thr_w[2]), .B(exu_tlu_cwp2_w[2]), .Y(exu_n17731));
INVX1 exu_U19393(.A(exu_n17731), .Y(exu_n5155));
AND2X1 exu_U19394(.A(exu_n15959), .B(exu_tlu_cwp0_w[2]), .Y(exu_n17733));
INVX1 exu_U19395(.A(exu_n17733), .Y(exu_n5156));
AND2X1 exu_U19396(.A(exu_tlu_cwp2_w[1]), .B(ecl_rml_thr_w[2]), .Y(exu_n17737));
INVX1 exu_U19397(.A(exu_n17737), .Y(exu_n5157));
AND2X1 exu_U19398(.A(exu_tlu_cwp0_w[1]), .B(exu_n15960), .Y(exu_n17739));
INVX1 exu_U19399(.A(exu_n17739), .Y(exu_n5158));
AND2X1 exu_U19400(.A(exu_tlu_cwp2_w[0]), .B(ecl_rml_thr_w[2]), .Y(exu_n17743));
INVX1 exu_U19401(.A(exu_n17743), .Y(exu_n5159));
AND2X1 exu_U19402(.A(exu_tlu_cwp0_w[0]), .B(exu_n15960), .Y(exu_n17745));
INVX1 exu_U19403(.A(exu_n17745), .Y(exu_n5160));
AND2X1 exu_U19404(.A(exu_n15950), .B(exu_tlu_cwp2_w[2]), .Y(exu_n17749));
INVX1 exu_U19405(.A(exu_n17749), .Y(exu_n5161));
AND2X1 exu_U19406(.A(exu_n15955), .B(exu_tlu_cwp0_w[2]), .Y(exu_n17751));
INVX1 exu_U19407(.A(exu_n17751), .Y(exu_n5162));
AND2X1 exu_U19408(.A(exu_tlu_cwp2_w[1]), .B(exu_n15951), .Y(exu_n17755));
INVX1 exu_U19409(.A(exu_n17755), .Y(exu_n5163));
AND2X1 exu_U19410(.A(exu_tlu_cwp0_w[1]), .B(exu_n15956), .Y(exu_n17757));
INVX1 exu_U19411(.A(exu_n17757), .Y(exu_n5164));
AND2X1 exu_U19412(.A(exu_tlu_cwp2_w[0]), .B(exu_n3), .Y(exu_n17761));
INVX1 exu_U19413(.A(exu_n17761), .Y(exu_n5165));
AND2X1 exu_U19414(.A(exu_tlu_cwp0_w[0]), .B(exu_n4), .Y(exu_n17763));
INVX1 exu_U19415(.A(exu_n17763), .Y(exu_n5166));
AND2X1 exu_U19416(.A(rml_cwp_thr_e[2]), .B(exu_tlu_cwp2_w[2]), .Y(exu_n17767));
INVX1 exu_U19417(.A(exu_n17767), .Y(exu_n5167));
AND2X1 exu_U19418(.A(exu_n15691), .B(exu_tlu_cwp0_w[2]), .Y(exu_n17769));
INVX1 exu_U19419(.A(exu_n17769), .Y(exu_n5168));
AND2X1 exu_U19420(.A(exu_tlu_cwp2_w[1]), .B(rml_cwp_thr_e[2]), .Y(exu_n17773));
INVX1 exu_U19421(.A(exu_n17773), .Y(exu_n5169));
AND2X1 exu_U19422(.A(exu_tlu_cwp0_w[1]), .B(exu_n15691), .Y(exu_n17775));
INVX1 exu_U19423(.A(exu_n17775), .Y(exu_n5170));
AND2X1 exu_U19424(.A(exu_tlu_cwp2_w[0]), .B(rml_cwp_thr_e[2]), .Y(exu_n17779));
INVX1 exu_U19425(.A(exu_n17779), .Y(exu_n5171));
AND2X1 exu_U19426(.A(exu_tlu_cwp0_w[0]), .B(exu_n15691), .Y(exu_n17781));
INVX1 exu_U19427(.A(exu_n17781), .Y(exu_n5172));
AND2X1 exu_U19428(.A(exu_n15922), .B(exu_tlu_cwp2_w[2]), .Y(exu_n17785));
INVX1 exu_U19429(.A(exu_n17785), .Y(exu_n5173));
AND2X1 exu_U19430(.A(exu_n15924), .B(exu_tlu_cwp0_w[2]), .Y(exu_n17787));
INVX1 exu_U19431(.A(exu_n17787), .Y(exu_n5174));
AND2X1 exu_U19432(.A(exu_tlu_cwp2_w[1]), .B(exu_n15922), .Y(exu_n17791));
INVX1 exu_U19433(.A(exu_n17791), .Y(exu_n5175));
AND2X1 exu_U19434(.A(exu_tlu_cwp0_w[1]), .B(exu_n15924), .Y(exu_n17793));
INVX1 exu_U19435(.A(exu_n17793), .Y(exu_n5176));
AND2X1 exu_U19436(.A(exu_tlu_cwp2_w[0]), .B(exu_n15922), .Y(exu_n17797));
INVX1 exu_U19437(.A(exu_n17797), .Y(exu_n5177));
AND2X1 exu_U19438(.A(exu_tlu_cwp0_w[0]), .B(exu_n15924), .Y(exu_n17799));
INVX1 exu_U19439(.A(exu_n17799), .Y(exu_n5178));
AND2X1 exu_U19440(.A(exu_n15431), .B(rml_cwp_tlu_exu_cwp_w[2]), .Y(exu_n17803));
INVX1 exu_U19441(.A(exu_n17803), .Y(exu_n5179));
AND2X1 exu_U19442(.A(rml_cwp_cwp_next0_mux_sel0), .B(exu_tlu_cwp0_w[2]), .Y(exu_n17805));
INVX1 exu_U19443(.A(exu_n17805), .Y(exu_n5180));
AND2X1 exu_U19444(.A(rml_cwp_tlu_exu_cwp_w[1]), .B(exu_n15431), .Y(exu_n17809));
INVX1 exu_U19445(.A(exu_n17809), .Y(exu_n5181));
AND2X1 exu_U19446(.A(exu_tlu_cwp0_w[1]), .B(rml_cwp_cwp_next0_mux_sel0), .Y(exu_n17811));
INVX1 exu_U19447(.A(exu_n17811), .Y(exu_n5182));
AND2X1 exu_U19448(.A(rml_cwp_tlu_exu_cwp_w[0]), .B(exu_n15431), .Y(exu_n17815));
INVX1 exu_U19449(.A(exu_n17815), .Y(exu_n5183));
AND2X1 exu_U19450(.A(exu_tlu_cwp0_w[0]), .B(rml_cwp_cwp_next0_mux_sel0), .Y(exu_n17817));
INVX1 exu_U19451(.A(exu_n17817), .Y(exu_n5184));
AND2X1 exu_U19452(.A(exu_n15430), .B(rml_cwp_tlu_exu_cwp_w[2]), .Y(exu_n17821));
INVX1 exu_U19453(.A(exu_n17821), .Y(exu_n5185));
AND2X1 exu_U19454(.A(rml_cwp_cwp_next1_mux_sel0), .B(exu_tlu_cwp1_w[2]), .Y(exu_n17823));
INVX1 exu_U19455(.A(exu_n17823), .Y(exu_n5186));
AND2X1 exu_U19456(.A(rml_cwp_tlu_exu_cwp_w[1]), .B(exu_n15430), .Y(exu_n17827));
INVX1 exu_U19457(.A(exu_n17827), .Y(exu_n5187));
AND2X1 exu_U19458(.A(exu_tlu_cwp1_w[1]), .B(rml_cwp_cwp_next1_mux_sel0), .Y(exu_n17829));
INVX1 exu_U19459(.A(exu_n17829), .Y(exu_n5188));
AND2X1 exu_U19460(.A(rml_cwp_tlu_exu_cwp_w[0]), .B(exu_n15430), .Y(exu_n17833));
INVX1 exu_U19461(.A(exu_n17833), .Y(exu_n5189));
AND2X1 exu_U19462(.A(exu_tlu_cwp1_w[0]), .B(rml_cwp_cwp_next1_mux_sel0), .Y(exu_n17835));
INVX1 exu_U19463(.A(exu_n17835), .Y(exu_n5190));
AND2X1 exu_U19464(.A(exu_n15429), .B(rml_cwp_tlu_exu_cwp_w[2]), .Y(exu_n17839));
INVX1 exu_U19465(.A(exu_n17839), .Y(exu_n5191));
AND2X1 exu_U19466(.A(rml_cwp_cwp_next2_mux_sel0), .B(exu_tlu_cwp2_w[2]), .Y(exu_n17841));
INVX1 exu_U19467(.A(exu_n17841), .Y(exu_n5192));
AND2X1 exu_U19468(.A(rml_cwp_tlu_exu_cwp_w[1]), .B(exu_n15429), .Y(exu_n17845));
INVX1 exu_U19469(.A(exu_n17845), .Y(exu_n5193));
AND2X1 exu_U19470(.A(exu_tlu_cwp2_w[1]), .B(rml_cwp_cwp_next2_mux_sel0), .Y(exu_n17847));
INVX1 exu_U19471(.A(exu_n17847), .Y(exu_n5194));
AND2X1 exu_U19472(.A(rml_cwp_tlu_exu_cwp_w[0]), .B(exu_n15429), .Y(exu_n17851));
INVX1 exu_U19473(.A(exu_n17851), .Y(exu_n5195));
AND2X1 exu_U19474(.A(exu_tlu_cwp2_w[0]), .B(rml_cwp_cwp_next2_mux_sel0), .Y(exu_n17853));
INVX1 exu_U19475(.A(exu_n17853), .Y(exu_n5196));
AND2X1 exu_U19476(.A(exu_n15428), .B(rml_cwp_tlu_exu_cwp_w[2]), .Y(exu_n17857));
INVX1 exu_U19477(.A(exu_n17857), .Y(exu_n5197));
AND2X1 exu_U19478(.A(rml_cwp_cwp_next3_mux_sel0), .B(exu_tlu_cwp3_w[2]), .Y(exu_n17859));
INVX1 exu_U19479(.A(exu_n17859), .Y(exu_n5198));
AND2X1 exu_U19480(.A(rml_cwp_tlu_exu_cwp_w[1]), .B(exu_n15428), .Y(exu_n17863));
INVX1 exu_U19481(.A(exu_n17863), .Y(exu_n5199));
AND2X1 exu_U19482(.A(exu_tlu_cwp3_w[1]), .B(rml_cwp_cwp_next3_mux_sel0), .Y(exu_n17865));
INVX1 exu_U19483(.A(exu_n17865), .Y(exu_n5200));
AND2X1 exu_U19484(.A(rml_cwp_tlu_exu_cwp_w[0]), .B(exu_n15428), .Y(exu_n17869));
INVX1 exu_U19485(.A(exu_n17869), .Y(exu_n5201));
AND2X1 exu_U19486(.A(exu_tlu_cwp3_w[0]), .B(rml_cwp_cwp_next3_mux_sel0), .Y(exu_n17871));
INVX1 exu_U19487(.A(exu_n17871), .Y(exu_n5202));
AND2X1 exu_U19488(.A(exu_n15951), .B(rml_cansave_reg_data_thr2[2]), .Y(exu_n17875));
INVX1 exu_U19489(.A(exu_n17875), .Y(exu_n5203));
AND2X1 exu_U19490(.A(exu_n15956), .B(rml_cansave_reg_data_thr0[2]), .Y(exu_n17877));
INVX1 exu_U19491(.A(exu_n17877), .Y(exu_n5204));
AND2X1 exu_U19492(.A(rml_cansave_reg_data_thr2[1]), .B(exu_n15950), .Y(exu_n17881));
INVX1 exu_U19493(.A(exu_n17881), .Y(exu_n5205));
AND2X1 exu_U19494(.A(rml_cansave_reg_data_thr0[1]), .B(exu_n15955), .Y(exu_n17883));
INVX1 exu_U19495(.A(exu_n17883), .Y(exu_n5206));
AND2X1 exu_U19496(.A(rml_cansave_reg_data_thr2[0]), .B(exu_n15950), .Y(exu_n17887));
INVX1 exu_U19497(.A(exu_n17887), .Y(exu_n5207));
AND2X1 exu_U19498(.A(rml_cansave_reg_data_thr0[0]), .B(exu_n15955), .Y(exu_n17889));
INVX1 exu_U19499(.A(exu_n17889), .Y(exu_n5208));
AND2X1 exu_U19500(.A(exu_n15188), .B(rml_canrestore_reg_data_thr2[2]), .Y(exu_n17893));
INVX1 exu_U19501(.A(exu_n17893), .Y(exu_n5209));
AND2X1 exu_U19502(.A(exu_n15192), .B(rml_canrestore_reg_data_thr0[2]), .Y(exu_n17895));
INVX1 exu_U19503(.A(exu_n17895), .Y(exu_n5210));
AND2X1 exu_U19504(.A(rml_canrestore_reg_data_thr2[1]), .B(exu_n15188), .Y(exu_n17899));
INVX1 exu_U19505(.A(exu_n17899), .Y(exu_n5211));
AND2X1 exu_U19506(.A(rml_canrestore_reg_data_thr0[1]), .B(exu_n15192), .Y(exu_n17901));
INVX1 exu_U19507(.A(exu_n17901), .Y(exu_n5212));
AND2X1 exu_U19508(.A(rml_canrestore_reg_data_thr2[0]), .B(exu_n15188), .Y(exu_n17905));
INVX1 exu_U19509(.A(exu_n17905), .Y(exu_n5213));
AND2X1 exu_U19510(.A(rml_canrestore_reg_data_thr0[0]), .B(exu_n15192), .Y(exu_n17907));
INVX1 exu_U19511(.A(exu_n17907), .Y(exu_n5214));
AND2X1 exu_U19512(.A(exu_n15188), .B(rml_otherwin_reg_data_thr2[2]), .Y(exu_n17911));
INVX1 exu_U19513(.A(exu_n17911), .Y(exu_n5215));
AND2X1 exu_U19514(.A(exu_n15192), .B(rml_otherwin_reg_data_thr0[2]), .Y(exu_n17913));
INVX1 exu_U19515(.A(exu_n17913), .Y(exu_n5216));
AND2X1 exu_U19516(.A(rml_otherwin_reg_data_thr2[1]), .B(exu_n15951), .Y(exu_n17917));
INVX1 exu_U19517(.A(exu_n17917), .Y(exu_n5217));
AND2X1 exu_U19518(.A(rml_otherwin_reg_data_thr0[1]), .B(exu_n15956), .Y(exu_n17919));
INVX1 exu_U19519(.A(exu_n17919), .Y(exu_n5218));
AND2X1 exu_U19520(.A(rml_otherwin_reg_data_thr2[0]), .B(exu_n15188), .Y(exu_n17923));
INVX1 exu_U19521(.A(exu_n17923), .Y(exu_n5219));
AND2X1 exu_U19522(.A(rml_otherwin_reg_data_thr0[0]), .B(exu_n15192), .Y(exu_n17925));
INVX1 exu_U19523(.A(exu_n17925), .Y(exu_n5220));
AND2X1 exu_U19524(.A(exu_n3), .B(rml_cleanwin_reg_data_thr2[2]), .Y(exu_n17929));
INVX1 exu_U19525(.A(exu_n17929), .Y(exu_n5221));
AND2X1 exu_U19526(.A(exu_n4), .B(rml_cleanwin_reg_data_thr0[2]), .Y(exu_n17931));
INVX1 exu_U19527(.A(exu_n17931), .Y(exu_n5222));
AND2X1 exu_U19528(.A(rml_cleanwin_reg_data_thr2[1]), .B(exu_n3), .Y(exu_n17935));
INVX1 exu_U19529(.A(exu_n17935), .Y(exu_n5223));
AND2X1 exu_U19530(.A(rml_cleanwin_reg_data_thr0[1]), .B(exu_n4), .Y(exu_n17937));
INVX1 exu_U19531(.A(exu_n17937), .Y(exu_n5224));
AND2X1 exu_U19532(.A(rml_cleanwin_reg_data_thr2[0]), .B(exu_n15188), .Y(exu_n17941));
INVX1 exu_U19533(.A(exu_n17941), .Y(exu_n5225));
AND2X1 exu_U19534(.A(rml_cleanwin_reg_data_thr0[0]), .B(exu_n15192), .Y(exu_n17943));
INVX1 exu_U19535(.A(exu_n17943), .Y(exu_n5226));
AND2X1 exu_U19536(.A(exu_n15950), .B(rml_hi_wstate_reg_data_thr2[2]), .Y(exu_n17947));
INVX1 exu_U19537(.A(exu_n17947), .Y(exu_n5227));
AND2X1 exu_U19538(.A(exu_n15955), .B(rml_hi_wstate_reg_data_thr0[2]), .Y(exu_n17949));
INVX1 exu_U19539(.A(exu_n17949), .Y(exu_n5228));
AND2X1 exu_U19540(.A(rml_hi_wstate_reg_data_thr2[1]), .B(exu_n15951), .Y(exu_n17953));
INVX1 exu_U19541(.A(exu_n17953), .Y(exu_n5229));
AND2X1 exu_U19542(.A(rml_hi_wstate_reg_data_thr0[1]), .B(exu_n15956), .Y(exu_n17955));
INVX1 exu_U19543(.A(exu_n17955), .Y(exu_n5230));
AND2X1 exu_U19544(.A(rml_hi_wstate_reg_data_thr2[0]), .B(exu_n15951), .Y(exu_n17959));
INVX1 exu_U19545(.A(exu_n17959), .Y(exu_n5231));
AND2X1 exu_U19546(.A(rml_hi_wstate_reg_data_thr0[0]), .B(exu_n15956), .Y(exu_n17961));
INVX1 exu_U19547(.A(exu_n17961), .Y(exu_n5232));
AND2X1 exu_U19548(.A(exu_n3), .B(rml_lo_wstate_reg_data_thr2[2]), .Y(exu_n17965));
INVX1 exu_U19549(.A(exu_n17965), .Y(exu_n5233));
AND2X1 exu_U19550(.A(exu_n4), .B(rml_lo_wstate_reg_data_thr0[2]), .Y(exu_n17967));
INVX1 exu_U19551(.A(exu_n17967), .Y(exu_n5234));
AND2X1 exu_U19552(.A(rml_lo_wstate_reg_data_thr2[1]), .B(exu_n3), .Y(exu_n17971));
INVX1 exu_U19553(.A(exu_n17971), .Y(exu_n5235));
AND2X1 exu_U19554(.A(rml_lo_wstate_reg_data_thr0[1]), .B(exu_n4), .Y(exu_n17973));
INVX1 exu_U19555(.A(exu_n17973), .Y(exu_n5236));
AND2X1 exu_U19556(.A(rml_lo_wstate_reg_data_thr2[0]), .B(exu_n15950), .Y(exu_n17977));
INVX1 exu_U19557(.A(exu_n17977), .Y(exu_n5237));
AND2X1 exu_U19558(.A(rml_lo_wstate_reg_data_thr0[0]), .B(exu_n15955), .Y(exu_n17979));
INVX1 exu_U19559(.A(exu_n17979), .Y(exu_n5238));
AND2X1 exu_U19560(.A(ecl_byp_sel_ecc_m), .B(exu_n10347), .Y(exu_n17984));
INVX1 exu_U19561(.A(exu_n17984), .Y(exu_n5239));
AND2X1 exu_U19562(.A(exu_n16274), .B(ecl_rd_m[4]), .Y(exu_n17986));
INVX1 exu_U19563(.A(exu_n17986), .Y(exu_n5240));
AND2X1 exu_U19564(.A(exu_n11581), .B(ecl_byp_sel_ecc_m), .Y(exu_n17990));
INVX1 exu_U19565(.A(exu_n17990), .Y(exu_n5241));
AND2X1 exu_U19566(.A(ecl_rd_m[3]), .B(exu_n16274), .Y(exu_n17992));
INVX1 exu_U19567(.A(exu_n17992), .Y(exu_n5242));
AND2X1 exu_U19568(.A(exu_n11582), .B(ecl_byp_sel_ecc_m), .Y(exu_n17996));
INVX1 exu_U19569(.A(exu_n17996), .Y(exu_n5243));
AND2X1 exu_U19570(.A(ecl_rd_m[2]), .B(exu_n16274), .Y(exu_n17998));
INVX1 exu_U19571(.A(exu_n17998), .Y(exu_n5244));
AND2X1 exu_U19572(.A(exu_n11583), .B(ecl_byp_sel_ecc_m), .Y(exu_n18002));
INVX1 exu_U19573(.A(exu_n18002), .Y(exu_n5245));
AND2X1 exu_U19574(.A(ecl_rd_m[1]), .B(exu_n16274), .Y(exu_n18004));
INVX1 exu_U19575(.A(exu_n18004), .Y(exu_n5246));
AND2X1 exu_U19576(.A(exu_n11584), .B(ecl_byp_sel_ecc_m), .Y(exu_n18008));
INVX1 exu_U19577(.A(exu_n18008), .Y(exu_n5247));
AND2X1 exu_U19578(.A(ecl_rd_m[0]), .B(exu_n16274), .Y(exu_n18010));
INVX1 exu_U19579(.A(exu_n18010), .Y(exu_n5248));
AND2X1 exu_U19580(.A(rml_ecl_wstate_d[2]), .B(exu_n15824), .Y(exu_n18022));
INVX1 exu_U19581(.A(exu_n18022), .Y(exu_n5249));
AND2X1 exu_U19582(.A(exu_ifu_cc_d[2]), .B(exu_n16373), .Y(exu_n18024));
INVX1 exu_U19583(.A(exu_n18024), .Y(exu_n5250));
AND2X1 exu_U19584(.A(rml_ecl_wstate_d[1]), .B(exu_n15824), .Y(exu_n18028));
INVX1 exu_U19585(.A(exu_n18028), .Y(exu_n5251));
AND2X1 exu_U19586(.A(exu_ifu_cc_d[1]), .B(exu_n16373), .Y(exu_n18030));
INVX1 exu_U19587(.A(exu_n18030), .Y(exu_n5252));
AND2X1 exu_U19588(.A(rml_ecl_wstate_d[0]), .B(exu_n15824), .Y(exu_n18034));
INVX1 exu_U19589(.A(exu_n18034), .Y(exu_n5253));
AND2X1 exu_U19590(.A(exu_ifu_cc_d[0]), .B(exu_n16373), .Y(exu_n18036));
INVX1 exu_U19591(.A(exu_n18036), .Y(exu_n5254));
AND2X1 exu_U19592(.A(ecl_ccr_wen_thr1_w), .B(exu_n15686), .Y(exu_n18040));
INVX1 exu_U19593(.A(exu_n18040), .Y(exu_n5255));
AND2X1 exu_U19594(.A(exu_n15702), .B(ecl_ccr_wen_thr1_w), .Y(exu_n18044));
INVX1 exu_U19595(.A(exu_n18044), .Y(exu_n5256));
AND2X1 exu_U19596(.A(exu_n15699), .B(ecl_ccr_wen_thr1_w), .Y(exu_n18052));
INVX1 exu_U19597(.A(exu_n18052), .Y(exu_n5257));
AND2X1 exu_U19598(.A(exu_n15698), .B(ecl_ccr_wen_thr1_w), .Y(exu_n18056));
INVX1 exu_U19599(.A(exu_n18056), .Y(exu_n5258));
AND2X1 exu_U19600(.A(exu_n15697), .B(ecl_ccr_wen_thr1_w), .Y(exu_n18060));
INVX1 exu_U19601(.A(exu_n18060), .Y(exu_n5259));
AND2X1 exu_U19602(.A(exu_n15696), .B(ecl_ccr_wen_thr1_w), .Y(exu_n18064));
INVX1 exu_U19603(.A(exu_n18064), .Y(exu_n5260));
AND2X1 exu_U19604(.A(ecl_ccr_wen_thr2_w), .B(exu_n15686), .Y(exu_n18068));
INVX1 exu_U19605(.A(exu_n18068), .Y(exu_n5261));
AND2X1 exu_U19606(.A(exu_n15702), .B(ecl_ccr_wen_thr2_w), .Y(exu_n18072));
INVX1 exu_U19607(.A(exu_n18072), .Y(exu_n5262));
AND2X1 exu_U19608(.A(exu_n15699), .B(ecl_ccr_wen_thr2_w), .Y(exu_n18080));
INVX1 exu_U19609(.A(exu_n18080), .Y(exu_n5263));
AND2X1 exu_U19610(.A(exu_n15698), .B(ecl_ccr_wen_thr2_w), .Y(exu_n18084));
INVX1 exu_U19611(.A(exu_n18084), .Y(exu_n5264));
AND2X1 exu_U19612(.A(exu_n15697), .B(ecl_ccr_wen_thr2_w), .Y(exu_n18088));
INVX1 exu_U19613(.A(exu_n18088), .Y(exu_n5265));
AND2X1 exu_U19614(.A(exu_n15696), .B(ecl_ccr_wen_thr2_w), .Y(exu_n18092));
INVX1 exu_U19615(.A(exu_n18092), .Y(exu_n5266));
AND2X1 exu_U19616(.A(ecl_ccr_wen_thr3_w), .B(exu_n15686), .Y(exu_n18096));
INVX1 exu_U19617(.A(exu_n18096), .Y(exu_n5267));
AND2X1 exu_U19618(.A(exu_n15702), .B(ecl_ccr_wen_thr3_w), .Y(exu_n18100));
INVX1 exu_U19619(.A(exu_n18100), .Y(exu_n5268));
AND2X1 exu_U19620(.A(exu_n15699), .B(ecl_ccr_wen_thr3_w), .Y(exu_n18108));
INVX1 exu_U19621(.A(exu_n18108), .Y(exu_n5269));
AND2X1 exu_U19622(.A(exu_n15698), .B(ecl_ccr_wen_thr3_w), .Y(exu_n18112));
INVX1 exu_U19623(.A(exu_n18112), .Y(exu_n5270));
AND2X1 exu_U19624(.A(exu_n15697), .B(ecl_ccr_wen_thr3_w), .Y(exu_n18116));
INVX1 exu_U19625(.A(exu_n18116), .Y(exu_n5271));
AND2X1 exu_U19626(.A(exu_n15696), .B(ecl_ccr_wen_thr3_w), .Y(exu_n18120));
INVX1 exu_U19627(.A(exu_n18120), .Y(exu_n5272));
AND2X1 exu_U19628(.A(ecl_ccr_use_cc_w), .B(ecl_ccr_alu_cc_w[7]), .Y(exu_n18122));
INVX1 exu_U19629(.A(exu_n18122), .Y(exu_n5273));
AND2X1 exu_U19630(.A(exu_n15931), .B(ecl_ccr_ccr_d[7]), .Y(exu_n18124));
INVX1 exu_U19631(.A(exu_n18124), .Y(exu_n5274));
AND2X1 exu_U19632(.A(ecl_ccr_alu_cc_w[6]), .B(ecl_ccr_use_cc_w), .Y(exu_n18126));
INVX1 exu_U19633(.A(exu_n18126), .Y(exu_n5275));
AND2X1 exu_U19634(.A(ecl_ccr_ccr_d[6]), .B(exu_n15931), .Y(exu_n18128));
INVX1 exu_U19635(.A(exu_n18128), .Y(exu_n5276));
AND2X1 exu_U19636(.A(ecl_ccr_alu_cc_w[5]), .B(ecl_ccr_use_cc_w), .Y(exu_n18130));
INVX1 exu_U19637(.A(exu_n18130), .Y(exu_n5277));
AND2X1 exu_U19638(.A(ecl_ccr_ccr_d[5]), .B(exu_n15931), .Y(exu_n18132));
INVX1 exu_U19639(.A(exu_n18132), .Y(exu_n5278));
AND2X1 exu_U19640(.A(ecl_ccr_alu_cc_w[4]), .B(ecl_ccr_use_cc_w), .Y(exu_n18134));
INVX1 exu_U19641(.A(exu_n18134), .Y(exu_n5279));
AND2X1 exu_U19642(.A(ecl_ccr_ccr_d[4]), .B(exu_n15931), .Y(exu_n18136));
INVX1 exu_U19643(.A(exu_n18136), .Y(exu_n5280));
AND2X1 exu_U19644(.A(ecl_ccr_alu_cc_w[3]), .B(ecl_ccr_use_cc_w), .Y(exu_n18138));
INVX1 exu_U19645(.A(exu_n18138), .Y(exu_n5281));
AND2X1 exu_U19646(.A(ecl_ccr_ccr_d[3]), .B(exu_n15931), .Y(exu_n18140));
INVX1 exu_U19647(.A(exu_n18140), .Y(exu_n5282));
AND2X1 exu_U19648(.A(ecl_ccr_alu_cc_w[2]), .B(ecl_ccr_use_cc_w), .Y(exu_n18142));
INVX1 exu_U19649(.A(exu_n18142), .Y(exu_n5283));
AND2X1 exu_U19650(.A(ecl_ccr_ccr_d[2]), .B(exu_n15931), .Y(exu_n18144));
INVX1 exu_U19651(.A(exu_n18144), .Y(exu_n5284));
AND2X1 exu_U19652(.A(ecl_ccr_alu_cc_w[1]), .B(ecl_ccr_use_cc_w), .Y(exu_n18146));
INVX1 exu_U19653(.A(exu_n18146), .Y(exu_n5285));
AND2X1 exu_U19654(.A(ecl_ccr_ccr_d[1]), .B(exu_n15931), .Y(exu_n18148));
INVX1 exu_U19655(.A(exu_n18148), .Y(exu_n5286));
AND2X1 exu_U19656(.A(ecl_ccr_alu_cc_w[0]), .B(ecl_ccr_use_cc_w), .Y(exu_n18150));
INVX1 exu_U19657(.A(exu_n18150), .Y(exu_n5287));
AND2X1 exu_U19658(.A(ecl_ccr_ccr_d[0]), .B(exu_n15931), .Y(exu_n18152));
INVX1 exu_U19659(.A(exu_n18152), .Y(exu_n5288));
AND2X1 exu_U19660(.A(byp_irf_rd_data_w[0]), .B(exu_n15939), .Y(exu_n18154));
INVX1 exu_U19661(.A(exu_n18154), .Y(exu_n5289));
AND2X1 exu_U19662(.A(byp_irf_rd_data_w[1]), .B(exu_n15939), .Y(exu_n18156));
INVX1 exu_U19663(.A(exu_n18156), .Y(exu_n5290));
AND2X1 exu_U19664(.A(byp_irf_rd_data_w[2]), .B(exu_n15939), .Y(exu_n18158));
INVX1 exu_U19665(.A(exu_n18158), .Y(exu_n5291));
AND2X1 exu_U19666(.A(byp_irf_rd_data_w[3]), .B(exu_n15939), .Y(exu_n18160));
INVX1 exu_U19667(.A(exu_n18160), .Y(exu_n5292));
AND2X1 exu_U19668(.A(byp_irf_rd_data_w[4]), .B(exu_n15939), .Y(exu_n18162));
INVX1 exu_U19669(.A(exu_n18162), .Y(exu_n5293));
AND2X1 exu_U19670(.A(byp_irf_rd_data_w[5]), .B(exu_n15939), .Y(exu_n18164));
INVX1 exu_U19671(.A(exu_n18164), .Y(exu_n5294));
AND2X1 exu_U19672(.A(byp_irf_rd_data_w[6]), .B(exu_n15939), .Y(exu_n18166));
INVX1 exu_U19673(.A(exu_n18166), .Y(exu_n5295));
AND2X1 exu_U19674(.A(byp_irf_rd_data_w[7]), .B(exu_n15939), .Y(exu_n18168));
INVX1 exu_U19675(.A(exu_n18168), .Y(exu_n5296));
AND2X1 exu_U19676(.A(exu_n10777), .B(exu_n9772), .Y(ecl_divcntl_q_next_nocout[0]));
INVX1 exu_U19677(.A(ecl_divcntl_q_next_nocout[0]), .Y(exu_n5297));
AND2X1 exu_U19678(.A(exu_n16437), .B(exu_n16215), .Y(exu_n18183));
INVX1 exu_U19679(.A(exu_n18183), .Y(exu_n5298));
AND2X1 exu_U19680(.A(exu_n10780), .B(exu_n9773), .Y(ecl_divcntl_sub_next_nocout[0]));
INVX1 exu_U19681(.A(ecl_divcntl_sub_next_nocout[0]), .Y(exu_n5299));
AND2X1 exu_U19682(.A(exu_n15412), .B(exu_n18426), .Y(exu_n18425));
INVX1 exu_U19683(.A(exu_n18425), .Y(exu_n5300));
AND2X1 exu_U19684(.A(exu_n15413), .B(exu_n18431), .Y(exu_n18430));
INVX1 exu_U19685(.A(exu_n18430), .Y(exu_n5301));
AND2X1 exu_U19686(.A(ecl_div_mul_get_new_data), .B(alu_logic_rs1_data_bf1[9]), .Y(exu_n18606));
INVX1 exu_U19687(.A(exu_n18606), .Y(exu_n5302));
AND2X1 exu_U19688(.A(div_input_data_e[99]), .B(ecl_div_mul_get_new_data), .Y(exu_n18609));
INVX1 exu_U19689(.A(exu_n18609), .Y(exu_n5303));
AND2X1 exu_U19690(.A(div_input_data_e[98]), .B(exu_n16254), .Y(exu_n18612));
INVX1 exu_U19691(.A(exu_n18612), .Y(exu_n5304));
AND2X1 exu_U19692(.A(div_input_data_e[97]), .B(exu_n16254), .Y(exu_n18615));
INVX1 exu_U19693(.A(exu_n18615), .Y(exu_n5305));
AND2X1 exu_U19694(.A(div_input_data_e[96]), .B(exu_n16254), .Y(exu_n18618));
INVX1 exu_U19695(.A(exu_n18618), .Y(exu_n5306));
AND2X1 exu_U19696(.A(div_input_data_e[95]), .B(ecl_div_mul_get_new_data), .Y(exu_n18622));
INVX1 exu_U19697(.A(exu_n18622), .Y(exu_n5307));
AND2X1 exu_U19698(.A(div_input_data_e[94]), .B(exu_n16254), .Y(exu_n18626));
INVX1 exu_U19699(.A(exu_n18626), .Y(exu_n5308));
AND2X1 exu_U19700(.A(div_input_data_e[93]), .B(ecl_div_mul_get_new_data), .Y(exu_n18630));
INVX1 exu_U19701(.A(exu_n18630), .Y(exu_n5309));
AND2X1 exu_U19702(.A(div_input_data_e[92]), .B(ecl_div_mul_get_new_data), .Y(exu_n18634));
INVX1 exu_U19703(.A(exu_n18634), .Y(exu_n5310));
AND2X1 exu_U19704(.A(div_input_data_e[91]), .B(exu_n16254), .Y(exu_n18638));
INVX1 exu_U19705(.A(exu_n18638), .Y(exu_n5311));
AND2X1 exu_U19706(.A(div_input_data_e[90]), .B(exu_n16254), .Y(exu_n18642));
INVX1 exu_U19707(.A(exu_n18642), .Y(exu_n5312));
AND2X1 exu_U19708(.A(alu_logic_rs1_data_bf1[8]), .B(ecl_div_mul_get_new_data), .Y(exu_n18646));
INVX1 exu_U19709(.A(exu_n18646), .Y(exu_n5313));
AND2X1 exu_U19710(.A(div_input_data_e[89]), .B(exu_n16254), .Y(exu_n18650));
INVX1 exu_U19711(.A(exu_n18650), .Y(exu_n5314));
AND2X1 exu_U19712(.A(div_input_data_e[88]), .B(ecl_div_mul_get_new_data), .Y(exu_n18654));
INVX1 exu_U19713(.A(exu_n18654), .Y(exu_n5315));
AND2X1 exu_U19714(.A(div_input_data_e[87]), .B(exu_n16254), .Y(exu_n18658));
INVX1 exu_U19715(.A(exu_n18658), .Y(exu_n5316));
AND2X1 exu_U19716(.A(div_input_data_e[86]), .B(exu_n16254), .Y(exu_n18662));
INVX1 exu_U19717(.A(exu_n18662), .Y(exu_n5317));
AND2X1 exu_U19718(.A(div_input_data_e[85]), .B(ecl_div_mul_get_new_data), .Y(exu_n18666));
INVX1 exu_U19719(.A(exu_n18666), .Y(exu_n5318));
AND2X1 exu_U19720(.A(div_input_data_e[84]), .B(ecl_div_mul_get_new_data), .Y(exu_n18670));
INVX1 exu_U19721(.A(exu_n18670), .Y(exu_n5319));
AND2X1 exu_U19722(.A(div_input_data_e[83]), .B(exu_n16254), .Y(exu_n18674));
INVX1 exu_U19723(.A(exu_n18674), .Y(exu_n5320));
AND2X1 exu_U19724(.A(div_input_data_e[82]), .B(exu_n16254), .Y(exu_n18678));
INVX1 exu_U19725(.A(exu_n18678), .Y(exu_n5321));
AND2X1 exu_U19726(.A(div_input_data_e[81]), .B(exu_n16254), .Y(exu_n18682));
INVX1 exu_U19727(.A(exu_n18682), .Y(exu_n5322));
AND2X1 exu_U19728(.A(div_input_data_e[80]), .B(ecl_div_mul_get_new_data), .Y(exu_n18686));
INVX1 exu_U19729(.A(exu_n18686), .Y(exu_n5323));
AND2X1 exu_U19730(.A(alu_logic_rs1_data_bf1[7]), .B(ecl_div_mul_get_new_data), .Y(exu_n18690));
INVX1 exu_U19731(.A(exu_n18690), .Y(exu_n5324));
AND2X1 exu_U19732(.A(div_input_data_e[79]), .B(exu_n16254), .Y(exu_n18694));
INVX1 exu_U19733(.A(exu_n18694), .Y(exu_n5325));
AND2X1 exu_U19734(.A(div_input_data_e[78]), .B(ecl_div_mul_get_new_data), .Y(exu_n18698));
INVX1 exu_U19735(.A(exu_n18698), .Y(exu_n5326));
AND2X1 exu_U19736(.A(div_input_data_e[77]), .B(ecl_div_mul_get_new_data), .Y(exu_n18702));
INVX1 exu_U19737(.A(exu_n18702), .Y(exu_n5327));
AND2X1 exu_U19738(.A(div_input_data_e[76]), .B(ecl_div_mul_get_new_data), .Y(exu_n18706));
INVX1 exu_U19739(.A(exu_n18706), .Y(exu_n5328));
AND2X1 exu_U19740(.A(div_input_data_e[75]), .B(exu_n16254), .Y(exu_n18710));
INVX1 exu_U19741(.A(exu_n18710), .Y(exu_n5329));
AND2X1 exu_U19742(.A(div_input_data_e[74]), .B(ecl_div_mul_get_new_data), .Y(exu_n18714));
INVX1 exu_U19743(.A(exu_n18714), .Y(exu_n5330));
AND2X1 exu_U19744(.A(div_input_data_e[73]), .B(ecl_div_mul_get_new_data), .Y(exu_n18718));
INVX1 exu_U19745(.A(exu_n18718), .Y(exu_n5331));
AND2X1 exu_U19746(.A(div_input_data_e[72]), .B(ecl_div_mul_get_new_data), .Y(exu_n18722));
INVX1 exu_U19747(.A(exu_n18722), .Y(exu_n5332));
AND2X1 exu_U19748(.A(div_input_data_e[71]), .B(ecl_div_mul_get_new_data), .Y(exu_n18726));
INVX1 exu_U19749(.A(exu_n18726), .Y(exu_n5333));
AND2X1 exu_U19750(.A(div_input_data_e[70]), .B(exu_n16254), .Y(exu_n18730));
INVX1 exu_U19751(.A(exu_n18730), .Y(exu_n5334));
AND2X1 exu_U19752(.A(alu_logic_rs1_data_bf1[6]), .B(exu_n16254), .Y(exu_n18734));
INVX1 exu_U19753(.A(exu_n18734), .Y(exu_n5335));
AND2X1 exu_U19754(.A(div_input_data_e[69]), .B(ecl_div_mul_get_new_data), .Y(exu_n18738));
INVX1 exu_U19755(.A(exu_n18738), .Y(exu_n5336));
AND2X1 exu_U19756(.A(div_input_data_e[68]), .B(exu_n16254), .Y(exu_n18742));
INVX1 exu_U19757(.A(exu_n18742), .Y(exu_n5337));
AND2X1 exu_U19758(.A(div_input_data_e[67]), .B(exu_n16254), .Y(exu_n18746));
INVX1 exu_U19759(.A(exu_n18746), .Y(exu_n5338));
AND2X1 exu_U19760(.A(div_input_data_e[66]), .B(exu_n16254), .Y(exu_n18750));
INVX1 exu_U19761(.A(exu_n18750), .Y(exu_n5339));
AND2X1 exu_U19762(.A(div_input_data_e[65]), .B(exu_n16254), .Y(exu_n18754));
INVX1 exu_U19763(.A(exu_n18754), .Y(exu_n5340));
AND2X1 exu_U19764(.A(div_input_data_e[64]), .B(exu_n16254), .Y(exu_n18758));
INVX1 exu_U19765(.A(exu_n18758), .Y(exu_n5341));
AND2X1 exu_U19766(.A(alu_logic_rs1_data_bf1[63]), .B(exu_n16254), .Y(exu_n18761));
INVX1 exu_U19767(.A(exu_n18761), .Y(exu_n5342));
AND2X1 exu_U19768(.A(alu_logic_rs1_data_bf1[62]), .B(exu_n16254), .Y(exu_n18764));
INVX1 exu_U19769(.A(exu_n18764), .Y(exu_n5343));
AND2X1 exu_U19770(.A(alu_logic_rs1_data_bf1[61]), .B(exu_n16254), .Y(exu_n18767));
INVX1 exu_U19771(.A(exu_n18767), .Y(exu_n5344));
AND2X1 exu_U19772(.A(alu_logic_rs1_data_bf1[60]), .B(ecl_div_mul_get_new_data), .Y(exu_n18770));
INVX1 exu_U19773(.A(exu_n18770), .Y(exu_n5345));
AND2X1 exu_U19774(.A(alu_logic_rs1_data_bf1[5]), .B(ecl_div_mul_get_new_data), .Y(exu_n18774));
INVX1 exu_U19775(.A(exu_n18774), .Y(exu_n5346));
AND2X1 exu_U19776(.A(alu_logic_rs1_data_bf1[59]), .B(exu_n16254), .Y(exu_n18777));
INVX1 exu_U19777(.A(exu_n18777), .Y(exu_n5347));
AND2X1 exu_U19778(.A(alu_logic_rs1_data_bf1[58]), .B(exu_n16254), .Y(exu_n18780));
INVX1 exu_U19779(.A(exu_n18780), .Y(exu_n5348));
AND2X1 exu_U19780(.A(alu_logic_rs1_data_bf1[57]), .B(ecl_div_mul_get_new_data), .Y(exu_n18783));
INVX1 exu_U19781(.A(exu_n18783), .Y(exu_n5349));
AND2X1 exu_U19782(.A(alu_logic_rs1_data_bf1[56]), .B(ecl_div_mul_get_new_data), .Y(exu_n18786));
INVX1 exu_U19783(.A(exu_n18786), .Y(exu_n5350));
AND2X1 exu_U19784(.A(alu_logic_rs1_data_bf1[55]), .B(ecl_div_mul_get_new_data), .Y(exu_n18789));
INVX1 exu_U19785(.A(exu_n18789), .Y(exu_n5351));
AND2X1 exu_U19786(.A(alu_logic_rs1_data_bf1[54]), .B(exu_n16254), .Y(exu_n18792));
INVX1 exu_U19787(.A(exu_n18792), .Y(exu_n5352));
AND2X1 exu_U19788(.A(alu_logic_rs1_data_bf1[53]), .B(exu_n16254), .Y(exu_n18795));
INVX1 exu_U19789(.A(exu_n18795), .Y(exu_n5353));
AND2X1 exu_U19790(.A(alu_logic_rs1_data_bf1[52]), .B(exu_n16254), .Y(exu_n18798));
INVX1 exu_U19791(.A(exu_n18798), .Y(exu_n5354));
AND2X1 exu_U19792(.A(alu_logic_rs1_data_bf1[51]), .B(ecl_div_mul_get_new_data), .Y(exu_n18801));
INVX1 exu_U19793(.A(exu_n18801), .Y(exu_n5355));
AND2X1 exu_U19794(.A(alu_logic_rs1_data_bf1[50]), .B(exu_n16254), .Y(exu_n18804));
INVX1 exu_U19795(.A(exu_n18804), .Y(exu_n5356));
AND2X1 exu_U19796(.A(alu_logic_rs1_data_bf1[4]), .B(ecl_div_mul_get_new_data), .Y(exu_n18808));
INVX1 exu_U19797(.A(exu_n18808), .Y(exu_n5357));
AND2X1 exu_U19798(.A(alu_logic_rs1_data_bf1[49]), .B(ecl_div_mul_get_new_data), .Y(exu_n18811));
INVX1 exu_U19799(.A(exu_n18811), .Y(exu_n5358));
AND2X1 exu_U19800(.A(alu_logic_rs1_data_bf1[48]), .B(ecl_div_mul_get_new_data), .Y(exu_n18814));
INVX1 exu_U19801(.A(exu_n18814), .Y(exu_n5359));
AND2X1 exu_U19802(.A(alu_logic_rs1_data_bf1[47]), .B(ecl_div_mul_get_new_data), .Y(exu_n18817));
INVX1 exu_U19803(.A(exu_n18817), .Y(exu_n5360));
AND2X1 exu_U19804(.A(alu_logic_rs1_data_bf1[46]), .B(exu_n16254), .Y(exu_n18820));
INVX1 exu_U19805(.A(exu_n18820), .Y(exu_n5361));
AND2X1 exu_U19806(.A(alu_logic_rs1_data_bf1[45]), .B(exu_n16254), .Y(exu_n18823));
INVX1 exu_U19807(.A(exu_n18823), .Y(exu_n5362));
AND2X1 exu_U19808(.A(alu_logic_rs1_data_bf1[44]), .B(ecl_div_mul_get_new_data), .Y(exu_n18826));
INVX1 exu_U19809(.A(exu_n18826), .Y(exu_n5363));
AND2X1 exu_U19810(.A(alu_logic_rs1_data_bf1[43]), .B(exu_n16254), .Y(exu_n18829));
INVX1 exu_U19811(.A(exu_n18829), .Y(exu_n5364));
AND2X1 exu_U19812(.A(alu_logic_rs1_data_bf1[42]), .B(ecl_div_mul_get_new_data), .Y(exu_n18832));
INVX1 exu_U19813(.A(exu_n18832), .Y(exu_n5365));
AND2X1 exu_U19814(.A(alu_logic_rs1_data_bf1[41]), .B(exu_n16254), .Y(exu_n18835));
INVX1 exu_U19815(.A(exu_n18835), .Y(exu_n5366));
AND2X1 exu_U19816(.A(alu_logic_rs1_data_bf1[40]), .B(exu_n16254), .Y(exu_n18838));
INVX1 exu_U19817(.A(exu_n18838), .Y(exu_n5367));
AND2X1 exu_U19818(.A(alu_logic_rs1_data_bf1[3]), .B(ecl_div_mul_get_new_data), .Y(exu_n18842));
INVX1 exu_U19819(.A(exu_n18842), .Y(exu_n5368));
AND2X1 exu_U19820(.A(alu_logic_rs1_data_bf1[39]), .B(ecl_div_mul_get_new_data), .Y(exu_n18845));
INVX1 exu_U19821(.A(exu_n18845), .Y(exu_n5369));
AND2X1 exu_U19822(.A(alu_logic_rs1_data_bf1[38]), .B(exu_n16254), .Y(exu_n18848));
INVX1 exu_U19823(.A(exu_n18848), .Y(exu_n5370));
AND2X1 exu_U19824(.A(alu_logic_rs1_data_bf1[37]), .B(ecl_div_mul_get_new_data), .Y(exu_n18851));
INVX1 exu_U19825(.A(exu_n18851), .Y(exu_n5371));
AND2X1 exu_U19826(.A(alu_logic_rs1_data_bf1[36]), .B(ecl_div_mul_get_new_data), .Y(exu_n18854));
INVX1 exu_U19827(.A(exu_n18854), .Y(exu_n5372));
AND2X1 exu_U19828(.A(alu_logic_rs1_data_bf1[35]), .B(exu_n16254), .Y(exu_n18857));
INVX1 exu_U19829(.A(exu_n18857), .Y(exu_n5373));
AND2X1 exu_U19830(.A(alu_logic_rs1_data_bf1[34]), .B(exu_n16254), .Y(exu_n18860));
INVX1 exu_U19831(.A(exu_n18860), .Y(exu_n5374));
AND2X1 exu_U19832(.A(alu_logic_rs1_data_bf1[33]), .B(exu_n16254), .Y(exu_n18863));
INVX1 exu_U19833(.A(exu_n18863), .Y(exu_n5375));
AND2X1 exu_U19834(.A(alu_logic_rs1_data_bf1[32]), .B(exu_n16254), .Y(exu_n18867));
INVX1 exu_U19835(.A(exu_n18867), .Y(exu_n5376));
AND2X1 exu_U19836(.A(alu_logic_rs1_data_bf1[31]), .B(ecl_div_mul_get_new_data), .Y(exu_n18871));
INVX1 exu_U19837(.A(exu_n18871), .Y(exu_n5377));
AND2X1 exu_U19838(.A(alu_logic_rs1_data_bf1[30]), .B(ecl_div_mul_get_new_data), .Y(exu_n18875));
INVX1 exu_U19839(.A(exu_n18875), .Y(exu_n5378));
AND2X1 exu_U19840(.A(alu_logic_rs1_data_bf1[2]), .B(ecl_div_mul_get_new_data), .Y(exu_n18879));
INVX1 exu_U19841(.A(exu_n18879), .Y(exu_n5379));
AND2X1 exu_U19842(.A(alu_logic_rs1_data_bf1[29]), .B(ecl_div_mul_get_new_data), .Y(exu_n18883));
INVX1 exu_U19843(.A(exu_n18883), .Y(exu_n5380));
AND2X1 exu_U19844(.A(alu_logic_rs1_data_bf1[28]), .B(exu_n16254), .Y(exu_n18887));
INVX1 exu_U19845(.A(exu_n18887), .Y(exu_n5381));
AND2X1 exu_U19846(.A(alu_logic_rs1_data_bf1[27]), .B(exu_n16254), .Y(exu_n18891));
INVX1 exu_U19847(.A(exu_n18891), .Y(exu_n5382));
AND2X1 exu_U19848(.A(alu_logic_rs1_data_bf1[26]), .B(exu_n16254), .Y(exu_n18895));
INVX1 exu_U19849(.A(exu_n18895), .Y(exu_n5383));
AND2X1 exu_U19850(.A(alu_logic_rs1_data_bf1[25]), .B(exu_n16254), .Y(exu_n18899));
INVX1 exu_U19851(.A(exu_n18899), .Y(exu_n5384));
AND2X1 exu_U19852(.A(alu_logic_rs1_data_bf1[24]), .B(exu_n16254), .Y(exu_n18903));
INVX1 exu_U19853(.A(exu_n18903), .Y(exu_n5385));
AND2X1 exu_U19854(.A(alu_logic_rs1_data_bf1[23]), .B(exu_n16254), .Y(exu_n18907));
INVX1 exu_U19855(.A(exu_n18907), .Y(exu_n5386));
AND2X1 exu_U19856(.A(alu_logic_rs1_data_bf1[22]), .B(exu_n16254), .Y(exu_n18911));
INVX1 exu_U19857(.A(exu_n18911), .Y(exu_n5387));
AND2X1 exu_U19858(.A(alu_logic_rs1_data_bf1[21]), .B(exu_n16254), .Y(exu_n18915));
INVX1 exu_U19859(.A(exu_n18915), .Y(exu_n5388));
AND2X1 exu_U19860(.A(alu_logic_rs1_data_bf1[20]), .B(ecl_div_mul_get_new_data), .Y(exu_n18919));
INVX1 exu_U19861(.A(exu_n18919), .Y(exu_n5389));
AND2X1 exu_U19862(.A(alu_logic_rs1_data_bf1[1]), .B(ecl_div_mul_get_new_data), .Y(exu_n18923));
INVX1 exu_U19863(.A(exu_n18923), .Y(exu_n5390));
AND2X1 exu_U19864(.A(alu_logic_rs1_data_bf1[19]), .B(exu_n16254), .Y(exu_n18927));
INVX1 exu_U19865(.A(exu_n18927), .Y(exu_n5391));
AND2X1 exu_U19866(.A(alu_logic_rs1_data_bf1[18]), .B(ecl_div_mul_get_new_data), .Y(exu_n18931));
INVX1 exu_U19867(.A(exu_n18931), .Y(exu_n5392));
AND2X1 exu_U19868(.A(alu_logic_rs1_data_bf1[17]), .B(exu_n16254), .Y(exu_n18935));
INVX1 exu_U19869(.A(exu_n18935), .Y(exu_n5393));
AND2X1 exu_U19870(.A(alu_logic_rs1_data_bf1[16]), .B(exu_n16254), .Y(exu_n18939));
INVX1 exu_U19871(.A(exu_n18939), .Y(exu_n5394));
AND2X1 exu_U19872(.A(alu_logic_rs1_data_bf1[15]), .B(exu_n16254), .Y(exu_n18943));
INVX1 exu_U19873(.A(exu_n18943), .Y(exu_n5395));
AND2X1 exu_U19874(.A(alu_logic_rs1_data_bf1[14]), .B(exu_n16254), .Y(exu_n18947));
INVX1 exu_U19875(.A(exu_n18947), .Y(exu_n5396));
AND2X1 exu_U19876(.A(alu_logic_rs1_data_bf1[13]), .B(exu_n16254), .Y(exu_n18951));
INVX1 exu_U19877(.A(exu_n18951), .Y(exu_n5397));
AND2X1 exu_U19878(.A(alu_logic_rs1_data_bf1[12]), .B(exu_n16254), .Y(exu_n18955));
INVX1 exu_U19879(.A(exu_n18955), .Y(exu_n5398));
AND2X1 exu_U19880(.A(div_input_data_e[127]), .B(exu_n16254), .Y(exu_n18958));
INVX1 exu_U19881(.A(exu_n18958), .Y(exu_n5399));
AND2X1 exu_U19882(.A(div_input_data_e[126]), .B(exu_n16254), .Y(exu_n18961));
INVX1 exu_U19883(.A(exu_n18961), .Y(exu_n5400));
AND2X1 exu_U19884(.A(div_input_data_e[125]), .B(exu_n16254), .Y(exu_n18964));
INVX1 exu_U19885(.A(exu_n18964), .Y(exu_n5401));
AND2X1 exu_U19886(.A(div_input_data_e[124]), .B(exu_n16254), .Y(exu_n18967));
INVX1 exu_U19887(.A(exu_n18967), .Y(exu_n5402));
AND2X1 exu_U19888(.A(div_input_data_e[123]), .B(exu_n16254), .Y(exu_n18970));
INVX1 exu_U19889(.A(exu_n18970), .Y(exu_n5403));
AND2X1 exu_U19890(.A(div_input_data_e[122]), .B(exu_n16254), .Y(exu_n18973));
INVX1 exu_U19891(.A(exu_n18973), .Y(exu_n5404));
AND2X1 exu_U19892(.A(div_input_data_e[121]), .B(exu_n16254), .Y(exu_n18976));
INVX1 exu_U19893(.A(exu_n18976), .Y(exu_n5405));
AND2X1 exu_U19894(.A(div_input_data_e[120]), .B(exu_n16254), .Y(exu_n18979));
INVX1 exu_U19895(.A(exu_n18979), .Y(exu_n5406));
AND2X1 exu_U19896(.A(alu_logic_rs1_data_bf1[11]), .B(ecl_div_mul_get_new_data), .Y(exu_n18983));
INVX1 exu_U19897(.A(exu_n18983), .Y(exu_n5407));
AND2X1 exu_U19898(.A(div_input_data_e[119]), .B(ecl_div_mul_get_new_data), .Y(exu_n18986));
INVX1 exu_U19899(.A(exu_n18986), .Y(exu_n5408));
AND2X1 exu_U19900(.A(div_input_data_e[118]), .B(exu_n16254), .Y(exu_n18989));
INVX1 exu_U19901(.A(exu_n18989), .Y(exu_n5409));
AND2X1 exu_U19902(.A(div_input_data_e[117]), .B(ecl_div_mul_get_new_data), .Y(exu_n18992));
INVX1 exu_U19903(.A(exu_n18992), .Y(exu_n5410));
AND2X1 exu_U19904(.A(div_input_data_e[116]), .B(ecl_div_mul_get_new_data), .Y(exu_n18995));
INVX1 exu_U19905(.A(exu_n18995), .Y(exu_n5411));
AND2X1 exu_U19906(.A(div_input_data_e[115]), .B(ecl_div_mul_get_new_data), .Y(exu_n18998));
INVX1 exu_U19907(.A(exu_n18998), .Y(exu_n5412));
AND2X1 exu_U19908(.A(div_input_data_e[114]), .B(ecl_div_mul_get_new_data), .Y(exu_n19001));
INVX1 exu_U19909(.A(exu_n19001), .Y(exu_n5413));
AND2X1 exu_U19910(.A(div_input_data_e[113]), .B(ecl_div_mul_get_new_data), .Y(exu_n19004));
INVX1 exu_U19911(.A(exu_n19004), .Y(exu_n5414));
AND2X1 exu_U19912(.A(div_input_data_e[112]), .B(exu_n16254), .Y(exu_n19007));
INVX1 exu_U19913(.A(exu_n19007), .Y(exu_n5415));
AND2X1 exu_U19914(.A(div_input_data_e[111]), .B(ecl_div_mul_get_new_data), .Y(exu_n19010));
INVX1 exu_U19915(.A(exu_n19010), .Y(exu_n5416));
AND2X1 exu_U19916(.A(div_input_data_e[110]), .B(exu_n16254), .Y(exu_n19013));
INVX1 exu_U19917(.A(exu_n19013), .Y(exu_n5417));
AND2X1 exu_U19918(.A(alu_logic_rs1_data_bf1[10]), .B(exu_n16254), .Y(exu_n19017));
INVX1 exu_U19919(.A(exu_n19017), .Y(exu_n5418));
AND2X1 exu_U19920(.A(div_input_data_e[109]), .B(ecl_div_mul_get_new_data), .Y(exu_n19020));
INVX1 exu_U19921(.A(exu_n19020), .Y(exu_n5419));
AND2X1 exu_U19922(.A(div_input_data_e[108]), .B(ecl_div_mul_get_new_data), .Y(exu_n19023));
INVX1 exu_U19923(.A(exu_n19023), .Y(exu_n5420));
AND2X1 exu_U19924(.A(div_input_data_e[107]), .B(ecl_div_mul_get_new_data), .Y(exu_n19026));
INVX1 exu_U19925(.A(exu_n19026), .Y(exu_n5421));
AND2X1 exu_U19926(.A(div_input_data_e[106]), .B(ecl_div_mul_get_new_data), .Y(exu_n19029));
INVX1 exu_U19927(.A(exu_n19029), .Y(exu_n5422));
AND2X1 exu_U19928(.A(div_input_data_e[105]), .B(exu_n16254), .Y(exu_n19032));
INVX1 exu_U19929(.A(exu_n19032), .Y(exu_n5423));
AND2X1 exu_U19930(.A(div_input_data_e[104]), .B(ecl_div_mul_get_new_data), .Y(exu_n19035));
INVX1 exu_U19931(.A(exu_n19035), .Y(exu_n5424));
AND2X1 exu_U19932(.A(div_input_data_e[103]), .B(exu_n16254), .Y(exu_n19038));
INVX1 exu_U19933(.A(exu_n19038), .Y(exu_n5425));
AND2X1 exu_U19934(.A(div_input_data_e[102]), .B(ecl_div_mul_get_new_data), .Y(exu_n19041));
INVX1 exu_U19935(.A(exu_n19041), .Y(exu_n5426));
AND2X1 exu_U19936(.A(div_input_data_e[101]), .B(ecl_div_mul_get_new_data), .Y(exu_n19044));
INVX1 exu_U19937(.A(exu_n19044), .Y(exu_n5427));
AND2X1 exu_U19938(.A(div_input_data_e[100]), .B(ecl_div_mul_get_new_data), .Y(exu_n19048));
INVX1 exu_U19939(.A(exu_n19048), .Y(exu_n5428));
AND2X1 exu_U19940(.A(alu_logic_rs1_data_bf1[0]), .B(exu_n16254), .Y(exu_n19052));
INVX1 exu_U19941(.A(exu_n19052), .Y(exu_n5429));
AND2X1 exu_U19942(.A(div_byp_yreg_e[9]), .B(exu_n16192), .Y(exu_n19054));
INVX1 exu_U19943(.A(exu_n19054), .Y(exu_n5430));
AND2X1 exu_U19944(.A(div_byp_yreg_e[8]), .B(exu_n16192), .Y(exu_n19056));
INVX1 exu_U19945(.A(exu_n19056), .Y(exu_n5431));
AND2X1 exu_U19946(.A(div_byp_yreg_e[7]), .B(exu_n16192), .Y(exu_n19058));
INVX1 exu_U19947(.A(exu_n19058), .Y(exu_n5432));
AND2X1 exu_U19948(.A(div_byp_yreg_e[6]), .B(exu_n16192), .Y(exu_n19060));
INVX1 exu_U19949(.A(exu_n19060), .Y(exu_n5433));
AND2X1 exu_U19950(.A(div_byp_yreg_e[5]), .B(exu_n16192), .Y(exu_n19062));
INVX1 exu_U19951(.A(exu_n19062), .Y(exu_n5434));
AND2X1 exu_U19952(.A(div_byp_yreg_e[4]), .B(exu_n16192), .Y(exu_n19064));
INVX1 exu_U19953(.A(exu_n19064), .Y(exu_n5435));
AND2X1 exu_U19954(.A(div_byp_yreg_e[3]), .B(exu_n16192), .Y(exu_n19066));
INVX1 exu_U19955(.A(exu_n19066), .Y(exu_n5436));
AND2X1 exu_U19956(.A(div_byp_yreg_e[31]), .B(exu_n16192), .Y(exu_n19068));
INVX1 exu_U19957(.A(exu_n19068), .Y(exu_n5437));
AND2X1 exu_U19958(.A(div_byp_yreg_e[30]), .B(exu_n16192), .Y(exu_n19070));
INVX1 exu_U19959(.A(exu_n19070), .Y(exu_n5438));
AND2X1 exu_U19960(.A(div_byp_yreg_e[2]), .B(exu_n16192), .Y(exu_n19072));
INVX1 exu_U19961(.A(exu_n19072), .Y(exu_n5439));
AND2X1 exu_U19962(.A(div_byp_yreg_e[29]), .B(exu_n16192), .Y(exu_n19074));
INVX1 exu_U19963(.A(exu_n19074), .Y(exu_n5440));
AND2X1 exu_U19964(.A(div_byp_yreg_e[28]), .B(exu_n16192), .Y(exu_n19076));
INVX1 exu_U19965(.A(exu_n19076), .Y(exu_n5441));
AND2X1 exu_U19966(.A(div_byp_yreg_e[27]), .B(exu_n16192), .Y(exu_n19078));
INVX1 exu_U19967(.A(exu_n19078), .Y(exu_n5442));
AND2X1 exu_U19968(.A(div_byp_yreg_e[26]), .B(exu_n16192), .Y(exu_n19080));
INVX1 exu_U19969(.A(exu_n19080), .Y(exu_n5443));
AND2X1 exu_U19970(.A(div_byp_yreg_e[25]), .B(exu_n16192), .Y(exu_n19082));
INVX1 exu_U19971(.A(exu_n19082), .Y(exu_n5444));
AND2X1 exu_U19972(.A(div_byp_yreg_e[24]), .B(exu_n16192), .Y(exu_n19084));
INVX1 exu_U19973(.A(exu_n19084), .Y(exu_n5445));
AND2X1 exu_U19974(.A(div_byp_yreg_e[23]), .B(exu_n16192), .Y(exu_n19086));
INVX1 exu_U19975(.A(exu_n19086), .Y(exu_n5446));
AND2X1 exu_U19976(.A(div_byp_yreg_e[22]), .B(exu_n16192), .Y(exu_n19088));
INVX1 exu_U19977(.A(exu_n19088), .Y(exu_n5447));
AND2X1 exu_U19978(.A(div_byp_yreg_e[21]), .B(exu_n16192), .Y(exu_n19090));
INVX1 exu_U19979(.A(exu_n19090), .Y(exu_n5448));
AND2X1 exu_U19980(.A(div_byp_yreg_e[20]), .B(exu_n16192), .Y(exu_n19092));
INVX1 exu_U19981(.A(exu_n19092), .Y(exu_n5449));
AND2X1 exu_U19982(.A(div_byp_yreg_e[1]), .B(exu_n16192), .Y(exu_n19094));
INVX1 exu_U19983(.A(exu_n19094), .Y(exu_n5450));
AND2X1 exu_U19984(.A(div_byp_yreg_e[19]), .B(exu_n16192), .Y(exu_n19096));
INVX1 exu_U19985(.A(exu_n19096), .Y(exu_n5451));
AND2X1 exu_U19986(.A(div_byp_yreg_e[18]), .B(exu_n16192), .Y(exu_n19098));
INVX1 exu_U19987(.A(exu_n19098), .Y(exu_n5452));
AND2X1 exu_U19988(.A(div_byp_yreg_e[17]), .B(exu_n16192), .Y(exu_n19100));
INVX1 exu_U19989(.A(exu_n19100), .Y(exu_n5453));
AND2X1 exu_U19990(.A(div_byp_yreg_e[16]), .B(exu_n16192), .Y(exu_n19102));
INVX1 exu_U19991(.A(exu_n19102), .Y(exu_n5454));
AND2X1 exu_U19992(.A(div_byp_yreg_e[15]), .B(exu_n16192), .Y(exu_n19104));
INVX1 exu_U19993(.A(exu_n19104), .Y(exu_n5455));
AND2X1 exu_U19994(.A(div_byp_yreg_e[14]), .B(exu_n16192), .Y(exu_n19106));
INVX1 exu_U19995(.A(exu_n19106), .Y(exu_n5456));
AND2X1 exu_U19996(.A(div_byp_yreg_e[13]), .B(exu_n16192), .Y(exu_n19108));
INVX1 exu_U19997(.A(exu_n19108), .Y(exu_n5457));
AND2X1 exu_U19998(.A(div_byp_yreg_e[12]), .B(exu_n16192), .Y(exu_n19110));
INVX1 exu_U19999(.A(exu_n19110), .Y(exu_n5458));
AND2X1 exu_U20000(.A(div_byp_yreg_e[11]), .B(exu_n16192), .Y(exu_n19112));
INVX1 exu_U20001(.A(exu_n19112), .Y(exu_n5459));
AND2X1 exu_U20002(.A(div_byp_yreg_e[10]), .B(exu_n16192), .Y(exu_n19114));
INVX1 exu_U20003(.A(exu_n19114), .Y(exu_n5460));
AND2X1 exu_U20004(.A(div_byp_yreg_e[0]), .B(exu_n16192), .Y(exu_n19116));
INVX1 exu_U20005(.A(exu_n19116), .Y(exu_n5461));
INVX1 exu_U20006(.A(exu_n5465), .Y(exu_n5462));
INVX1 exu_U20007(.A(exu_n5462), .Y(exu_n5463));
INVX1 exu_U20008(.A(exu_n5467), .Y(exu_n5464));
INVX1 exu_U20009(.A(exu_n5464), .Y(exu_n5465));
INVX1 exu_U20010(.A(exu_n5469), .Y(exu_n5466));
INVX1 exu_U20011(.A(exu_n5466), .Y(exu_n5467));
INVX1 exu_U20012(.A(exu_n5471), .Y(exu_n5468));
INVX1 exu_U20013(.A(exu_n5468), .Y(exu_n5469));
INVX1 exu_U20014(.A(exu_n5473), .Y(exu_n5470));
INVX1 exu_U20015(.A(exu_n5470), .Y(exu_n5471));
INVX1 exu_U20016(.A(exu_n5475), .Y(exu_n5472));
INVX1 exu_U20017(.A(exu_n5472), .Y(exu_n5473));
INVX1 exu_U20018(.A(exu_n5477), .Y(exu_n5474));
INVX1 exu_U20019(.A(exu_n5474), .Y(exu_n5475));
INVX1 exu_U20020(.A(exu_n5479), .Y(exu_n5476));
INVX1 exu_U20021(.A(exu_n5476), .Y(exu_n5477));
INVX1 exu_U20022(.A(exu_n5481), .Y(exu_n5478));
INVX1 exu_U20023(.A(exu_n5478), .Y(exu_n5479));
INVX1 exu_U20024(.A(exu_n5483), .Y(exu_n5480));
INVX1 exu_U20025(.A(exu_n5480), .Y(exu_n5481));
INVX1 exu_U20026(.A(exu_n5485), .Y(exu_n5482));
INVX1 exu_U20027(.A(exu_n5482), .Y(exu_n5483));
INVX1 exu_U20028(.A(exu_n5487), .Y(exu_n5484));
INVX1 exu_U20029(.A(exu_n5484), .Y(exu_n5485));
INVX1 exu_U20030(.A(exu_n5489), .Y(exu_n5486));
INVX1 exu_U20031(.A(exu_n5486), .Y(exu_n5487));
INVX1 exu_U20032(.A(exu_n5491), .Y(exu_n5488));
INVX1 exu_U20033(.A(exu_n5488), .Y(exu_n5489));
INVX1 exu_U20034(.A(exu_n5493), .Y(exu_n5490));
INVX1 exu_U20035(.A(exu_n5490), .Y(exu_n5491));
INVX1 exu_U20036(.A(exu_n5494), .Y(exu_n5492));
INVX1 exu_U20037(.A(exu_n5492), .Y(exu_n5493));
AND2X1 exu_U20038(.A(exu_n16260), .B(exu_n16185), .Y(exu_n19148));
INVX1 exu_U20039(.A(exu_n19148), .Y(exu_n5494));
AND2X1 exu_U20040(.A(exu_n15814), .B(exu_n16185), .Y(exu_n19150));
INVX1 exu_U20041(.A(exu_n19150), .Y(exu_n5495));
INVX1 exu_U20042(.A(exu_n5499), .Y(exu_n5496));
INVX1 exu_U20043(.A(exu_n5496), .Y(exu_n5497));
INVX1 exu_U20044(.A(exu_n5501), .Y(exu_n5498));
INVX1 exu_U20045(.A(exu_n5498), .Y(exu_n5499));
INVX1 exu_U20046(.A(exu_n5503), .Y(exu_n5500));
INVX1 exu_U20047(.A(exu_n5500), .Y(exu_n5501));
INVX1 exu_U20048(.A(exu_n5505), .Y(exu_n5502));
INVX1 exu_U20049(.A(exu_n5502), .Y(exu_n5503));
INVX1 exu_U20050(.A(exu_n5507), .Y(exu_n5504));
INVX1 exu_U20051(.A(exu_n5504), .Y(exu_n5505));
INVX1 exu_U20052(.A(exu_n5511), .Y(exu_n5506));
INVX1 exu_U20053(.A(exu_n5506), .Y(exu_n5507));
INVX1 exu_U20054(.A(exu_n5511), .Y(exu_n5508));
INVX1 exu_U20055(.A(exu_n5508), .Y(exu_n5509));
INVX1 exu_U20056(.A(exu_n5513), .Y(exu_n5510));
INVX1 exu_U20057(.A(exu_n5510), .Y(exu_n5511));
INVX1 exu_U20058(.A(exu_n5515), .Y(exu_n5512));
INVX1 exu_U20059(.A(exu_n5512), .Y(exu_n5513));
INVX1 exu_U20060(.A(exu_n5517), .Y(exu_n5514));
INVX1 exu_U20061(.A(exu_n5514), .Y(exu_n5515));
INVX1 exu_U20062(.A(exu_n5519), .Y(exu_n5516));
INVX1 exu_U20063(.A(exu_n5516), .Y(exu_n5517));
INVX1 exu_U20064(.A(exu_n5521), .Y(exu_n5518));
INVX1 exu_U20065(.A(exu_n5518), .Y(exu_n5519));
INVX1 exu_U20066(.A(exu_n5523), .Y(exu_n5520));
INVX1 exu_U20067(.A(exu_n5520), .Y(exu_n5521));
INVX1 exu_U20068(.A(exu_n5525), .Y(exu_n5522));
INVX1 exu_U20069(.A(exu_n5522), .Y(exu_n5523));
INVX1 exu_U20070(.A(exu_n5527), .Y(exu_n5524));
INVX1 exu_U20071(.A(exu_n5524), .Y(exu_n5525));
INVX1 exu_U20072(.A(exu_n5529), .Y(exu_n5526));
INVX1 exu_U20073(.A(exu_n5526), .Y(exu_n5527));
INVX1 exu_U20074(.A(exu_n5530), .Y(exu_n5528));
INVX1 exu_U20075(.A(exu_n5528), .Y(exu_n5529));
AND2X1 exu_U20076(.A(ecl_div_xinmask), .B(exu_n16192), .Y(exu_n19183));
INVX1 exu_U20077(.A(exu_n19183), .Y(exu_n5530));
AND2X1 exu_U20078(.A(exu_n19189), .B(exu_n19190), .Y(exu_n19188));
INVX1 exu_U20079(.A(exu_n19188), .Y(exu_n5531));
AND2X1 exu_U20080(.A(exu_n15818), .B(exu_n15421), .Y(exu_n19208));
INVX1 exu_U20081(.A(exu_n19208), .Y(exu_n5532));
AND2X1 exu_U20082(.A(exu_n15462), .B(exu_n9987), .Y(exu_n19209));
INVX1 exu_U20083(.A(exu_n19209), .Y(exu_n5533));
AND2X1 exu_U20084(.A(exu_n10991), .B(exu_n9988), .Y(exu_n19216));
INVX1 exu_U20085(.A(exu_n19216), .Y(exu_n5534));
AND2X1 exu_U20086(.A(exu_n19225), .B(exu_n19226), .Y(exu_n19224));
INVX1 exu_U20087(.A(exu_n19224), .Y(exu_n5535));
AND2X1 exu_U20088(.A(exu_n15819), .B(exu_n15422), .Y(exu_n19244));
INVX1 exu_U20089(.A(exu_n19244), .Y(exu_n5536));
AND2X1 exu_U20090(.A(exu_n15463), .B(exu_n9991), .Y(exu_n19245));
INVX1 exu_U20091(.A(exu_n19245), .Y(exu_n5537));
AND2X1 exu_U20092(.A(exu_n15028), .B(ecc_rs1_err_m[6]), .Y(exu_n19925));
INVX1 exu_U20093(.A(exu_n19925), .Y(exu_n5538));
AND2X1 exu_U20094(.A(ecc_rs1_err_m[5]), .B(exu_n15028), .Y(exu_n19929));
INVX1 exu_U20095(.A(exu_n19929), .Y(exu_n5539));
AND2X1 exu_U20096(.A(ecc_rs1_err_m[4]), .B(exu_n15028), .Y(exu_n19933));
INVX1 exu_U20097(.A(exu_n19933), .Y(exu_n5540));
AND2X1 exu_U20098(.A(ecc_rs1_err_m[3]), .B(exu_n15028), .Y(exu_n19937));
INVX1 exu_U20099(.A(exu_n19937), .Y(exu_n5541));
AND2X1 exu_U20100(.A(ecc_rs1_err_m[2]), .B(exu_n15028), .Y(exu_n19941));
INVX1 exu_U20101(.A(exu_n19941), .Y(exu_n5542));
AND2X1 exu_U20102(.A(ecc_rs1_err_m[1]), .B(exu_n15028), .Y(exu_n19945));
INVX1 exu_U20103(.A(exu_n19945), .Y(exu_n5543));
AND2X1 exu_U20104(.A(ecc_rs1_err_m[0]), .B(exu_n15028), .Y(exu_n19949));
INVX1 exu_U20105(.A(exu_n19949), .Y(exu_n5544));
OR2X1 exu_U20106(.A(ecc_rs2_err_e[6]), .B(ecc_rs2_err_e[5]), .Y(exu_n20001));
INVX1 exu_U20107(.A(exu_n20001), .Y(exu_n5545));
OR2X1 exu_U20108(.A(ecc_rs3_err_e[6]), .B(ecc_rs3_err_e[5]), .Y(exu_n20137));
INVX1 exu_U20109(.A(exu_n20137), .Y(exu_n5546));
AND2X1 exu_U20110(.A(exu_n16288), .B(alu_byp_rd_data_e[9]), .Y(exu_n20479));
INVX1 exu_U20111(.A(exu_n20479), .Y(exu_n5547));
AND2X1 exu_U20112(.A(exu_n19220), .B(bypass_rs3h_data_btwn_mux[9]), .Y(exu_n20481));
INVX1 exu_U20113(.A(exu_n20481), .Y(exu_n5548));
AND2X1 exu_U20114(.A(alu_byp_rd_data_e[8]), .B(exu_n16288), .Y(exu_n20485));
INVX1 exu_U20115(.A(exu_n20485), .Y(exu_n5549));
AND2X1 exu_U20116(.A(bypass_rs3h_data_btwn_mux[8]), .B(exu_n19220), .Y(exu_n20487));
INVX1 exu_U20117(.A(exu_n20487), .Y(exu_n5550));
AND2X1 exu_U20118(.A(alu_byp_rd_data_e[7]), .B(exu_n16288), .Y(exu_n20491));
INVX1 exu_U20119(.A(exu_n20491), .Y(exu_n5551));
AND2X1 exu_U20120(.A(bypass_rs3h_data_btwn_mux[7]), .B(exu_n19220), .Y(exu_n20493));
INVX1 exu_U20121(.A(exu_n20493), .Y(exu_n5552));
AND2X1 exu_U20122(.A(alu_byp_rd_data_e[6]), .B(exu_n16288), .Y(exu_n20497));
INVX1 exu_U20123(.A(exu_n20497), .Y(exu_n5553));
AND2X1 exu_U20124(.A(bypass_rs3h_data_btwn_mux[6]), .B(exu_n19220), .Y(exu_n20499));
INVX1 exu_U20125(.A(exu_n20499), .Y(exu_n5554));
AND2X1 exu_U20126(.A(alu_byp_rd_data_e[5]), .B(exu_n16288), .Y(exu_n20503));
INVX1 exu_U20127(.A(exu_n20503), .Y(exu_n5555));
AND2X1 exu_U20128(.A(bypass_rs3h_data_btwn_mux[5]), .B(exu_n19220), .Y(exu_n20505));
INVX1 exu_U20129(.A(exu_n20505), .Y(exu_n5556));
AND2X1 exu_U20130(.A(alu_byp_rd_data_e[4]), .B(exu_n16288), .Y(exu_n20509));
INVX1 exu_U20131(.A(exu_n20509), .Y(exu_n5557));
AND2X1 exu_U20132(.A(bypass_rs3h_data_btwn_mux[4]), .B(exu_n19220), .Y(exu_n20511));
INVX1 exu_U20133(.A(exu_n20511), .Y(exu_n5558));
AND2X1 exu_U20134(.A(alu_byp_rd_data_e[3]), .B(exu_n16288), .Y(exu_n20515));
INVX1 exu_U20135(.A(exu_n20515), .Y(exu_n5559));
AND2X1 exu_U20136(.A(bypass_rs3h_data_btwn_mux[3]), .B(exu_n19220), .Y(exu_n20517));
INVX1 exu_U20137(.A(exu_n20517), .Y(exu_n5560));
AND2X1 exu_U20138(.A(alu_byp_rd_data_e[31]), .B(exu_n16288), .Y(exu_n20521));
INVX1 exu_U20139(.A(exu_n20521), .Y(exu_n5561));
AND2X1 exu_U20140(.A(bypass_rs3h_data_btwn_mux[31]), .B(exu_n19220), .Y(exu_n20523));
INVX1 exu_U20141(.A(exu_n20523), .Y(exu_n5562));
AND2X1 exu_U20142(.A(alu_byp_rd_data_e[30]), .B(exu_n16288), .Y(exu_n20527));
INVX1 exu_U20143(.A(exu_n20527), .Y(exu_n5563));
AND2X1 exu_U20144(.A(bypass_rs3h_data_btwn_mux[30]), .B(exu_n19220), .Y(exu_n20529));
INVX1 exu_U20145(.A(exu_n20529), .Y(exu_n5564));
AND2X1 exu_U20146(.A(alu_byp_rd_data_e[2]), .B(exu_n16288), .Y(exu_n20533));
INVX1 exu_U20147(.A(exu_n20533), .Y(exu_n5565));
AND2X1 exu_U20148(.A(bypass_rs3h_data_btwn_mux[2]), .B(exu_n19220), .Y(exu_n20535));
INVX1 exu_U20149(.A(exu_n20535), .Y(exu_n5566));
AND2X1 exu_U20150(.A(alu_byp_rd_data_e[29]), .B(exu_n16288), .Y(exu_n20539));
INVX1 exu_U20151(.A(exu_n20539), .Y(exu_n5567));
AND2X1 exu_U20152(.A(bypass_rs3h_data_btwn_mux[29]), .B(exu_n19220), .Y(exu_n20541));
INVX1 exu_U20153(.A(exu_n20541), .Y(exu_n5568));
AND2X1 exu_U20154(.A(alu_byp_rd_data_e[28]), .B(exu_n16288), .Y(exu_n20545));
INVX1 exu_U20155(.A(exu_n20545), .Y(exu_n5569));
AND2X1 exu_U20156(.A(bypass_rs3h_data_btwn_mux[28]), .B(exu_n19220), .Y(exu_n20547));
INVX1 exu_U20157(.A(exu_n20547), .Y(exu_n5570));
AND2X1 exu_U20158(.A(alu_byp_rd_data_e[27]), .B(exu_n16288), .Y(exu_n20551));
INVX1 exu_U20159(.A(exu_n20551), .Y(exu_n5571));
AND2X1 exu_U20160(.A(bypass_rs3h_data_btwn_mux[27]), .B(exu_n19220), .Y(exu_n20553));
INVX1 exu_U20161(.A(exu_n20553), .Y(exu_n5572));
AND2X1 exu_U20162(.A(alu_byp_rd_data_e[26]), .B(exu_n16288), .Y(exu_n20557));
INVX1 exu_U20163(.A(exu_n20557), .Y(exu_n5573));
AND2X1 exu_U20164(.A(bypass_rs3h_data_btwn_mux[26]), .B(exu_n19220), .Y(exu_n20559));
INVX1 exu_U20165(.A(exu_n20559), .Y(exu_n5574));
AND2X1 exu_U20166(.A(alu_byp_rd_data_e[25]), .B(exu_n16288), .Y(exu_n20563));
INVX1 exu_U20167(.A(exu_n20563), .Y(exu_n5575));
AND2X1 exu_U20168(.A(bypass_rs3h_data_btwn_mux[25]), .B(exu_n19220), .Y(exu_n20565));
INVX1 exu_U20169(.A(exu_n20565), .Y(exu_n5576));
AND2X1 exu_U20170(.A(alu_byp_rd_data_e[24]), .B(exu_n16288), .Y(exu_n20569));
INVX1 exu_U20171(.A(exu_n20569), .Y(exu_n5577));
AND2X1 exu_U20172(.A(bypass_rs3h_data_btwn_mux[24]), .B(exu_n19220), .Y(exu_n20571));
INVX1 exu_U20173(.A(exu_n20571), .Y(exu_n5578));
AND2X1 exu_U20174(.A(alu_byp_rd_data_e[23]), .B(exu_n16288), .Y(exu_n20575));
INVX1 exu_U20175(.A(exu_n20575), .Y(exu_n5579));
AND2X1 exu_U20176(.A(bypass_rs3h_data_btwn_mux[23]), .B(exu_n19220), .Y(exu_n20577));
INVX1 exu_U20177(.A(exu_n20577), .Y(exu_n5580));
AND2X1 exu_U20178(.A(alu_byp_rd_data_e[22]), .B(exu_n16288), .Y(exu_n20581));
INVX1 exu_U20179(.A(exu_n20581), .Y(exu_n5581));
AND2X1 exu_U20180(.A(bypass_rs3h_data_btwn_mux[22]), .B(exu_n19220), .Y(exu_n20583));
INVX1 exu_U20181(.A(exu_n20583), .Y(exu_n5582));
AND2X1 exu_U20182(.A(alu_byp_rd_data_e[21]), .B(exu_n16288), .Y(exu_n20587));
INVX1 exu_U20183(.A(exu_n20587), .Y(exu_n5583));
AND2X1 exu_U20184(.A(bypass_rs3h_data_btwn_mux[21]), .B(exu_n19220), .Y(exu_n20589));
INVX1 exu_U20185(.A(exu_n20589), .Y(exu_n5584));
AND2X1 exu_U20186(.A(alu_byp_rd_data_e[20]), .B(exu_n16288), .Y(exu_n20593));
INVX1 exu_U20187(.A(exu_n20593), .Y(exu_n5585));
AND2X1 exu_U20188(.A(bypass_rs3h_data_btwn_mux[20]), .B(exu_n19220), .Y(exu_n20595));
INVX1 exu_U20189(.A(exu_n20595), .Y(exu_n5586));
AND2X1 exu_U20190(.A(alu_byp_rd_data_e[1]), .B(exu_n16288), .Y(exu_n20599));
INVX1 exu_U20191(.A(exu_n20599), .Y(exu_n5587));
AND2X1 exu_U20192(.A(bypass_rs3h_data_btwn_mux[1]), .B(exu_n19220), .Y(exu_n20601));
INVX1 exu_U20193(.A(exu_n20601), .Y(exu_n5588));
AND2X1 exu_U20194(.A(alu_byp_rd_data_e[19]), .B(exu_n16288), .Y(exu_n20605));
INVX1 exu_U20195(.A(exu_n20605), .Y(exu_n5589));
AND2X1 exu_U20196(.A(bypass_rs3h_data_btwn_mux[19]), .B(exu_n19220), .Y(exu_n20607));
INVX1 exu_U20197(.A(exu_n20607), .Y(exu_n5590));
AND2X1 exu_U20198(.A(alu_byp_rd_data_e[18]), .B(exu_n16288), .Y(exu_n20611));
INVX1 exu_U20199(.A(exu_n20611), .Y(exu_n5591));
AND2X1 exu_U20200(.A(bypass_rs3h_data_btwn_mux[18]), .B(exu_n19220), .Y(exu_n20613));
INVX1 exu_U20201(.A(exu_n20613), .Y(exu_n5592));
AND2X1 exu_U20202(.A(alu_byp_rd_data_e[17]), .B(exu_n16288), .Y(exu_n20617));
INVX1 exu_U20203(.A(exu_n20617), .Y(exu_n5593));
AND2X1 exu_U20204(.A(bypass_rs3h_data_btwn_mux[17]), .B(exu_n19220), .Y(exu_n20619));
INVX1 exu_U20205(.A(exu_n20619), .Y(exu_n5594));
AND2X1 exu_U20206(.A(alu_byp_rd_data_e[16]), .B(exu_n16288), .Y(exu_n20623));
INVX1 exu_U20207(.A(exu_n20623), .Y(exu_n5595));
AND2X1 exu_U20208(.A(bypass_rs3h_data_btwn_mux[16]), .B(exu_n19220), .Y(exu_n20625));
INVX1 exu_U20209(.A(exu_n20625), .Y(exu_n5596));
AND2X1 exu_U20210(.A(alu_byp_rd_data_e[15]), .B(exu_n16288), .Y(exu_n20629));
INVX1 exu_U20211(.A(exu_n20629), .Y(exu_n5597));
AND2X1 exu_U20212(.A(bypass_rs3h_data_btwn_mux[15]), .B(exu_n19220), .Y(exu_n20631));
INVX1 exu_U20213(.A(exu_n20631), .Y(exu_n5598));
AND2X1 exu_U20214(.A(alu_byp_rd_data_e[14]), .B(exu_n16288), .Y(exu_n20635));
INVX1 exu_U20215(.A(exu_n20635), .Y(exu_n5599));
AND2X1 exu_U20216(.A(bypass_rs3h_data_btwn_mux[14]), .B(exu_n19220), .Y(exu_n20637));
INVX1 exu_U20217(.A(exu_n20637), .Y(exu_n5600));
AND2X1 exu_U20218(.A(alu_byp_rd_data_e[13]), .B(exu_n16288), .Y(exu_n20641));
INVX1 exu_U20219(.A(exu_n20641), .Y(exu_n5601));
AND2X1 exu_U20220(.A(bypass_rs3h_data_btwn_mux[13]), .B(exu_n19220), .Y(exu_n20643));
INVX1 exu_U20221(.A(exu_n20643), .Y(exu_n5602));
AND2X1 exu_U20222(.A(alu_byp_rd_data_e[12]), .B(exu_n16288), .Y(exu_n20647));
INVX1 exu_U20223(.A(exu_n20647), .Y(exu_n5603));
AND2X1 exu_U20224(.A(bypass_rs3h_data_btwn_mux[12]), .B(exu_n19220), .Y(exu_n20649));
INVX1 exu_U20225(.A(exu_n20649), .Y(exu_n5604));
AND2X1 exu_U20226(.A(alu_byp_rd_data_e[11]), .B(exu_n16288), .Y(exu_n20653));
INVX1 exu_U20227(.A(exu_n20653), .Y(exu_n5605));
AND2X1 exu_U20228(.A(bypass_rs3h_data_btwn_mux[11]), .B(exu_n19220), .Y(exu_n20655));
INVX1 exu_U20229(.A(exu_n20655), .Y(exu_n5606));
AND2X1 exu_U20230(.A(alu_byp_rd_data_e[10]), .B(exu_n16288), .Y(exu_n20659));
INVX1 exu_U20231(.A(exu_n20659), .Y(exu_n5607));
AND2X1 exu_U20232(.A(bypass_rs3h_data_btwn_mux[10]), .B(exu_n19220), .Y(exu_n20661));
INVX1 exu_U20233(.A(exu_n20661), .Y(exu_n5608));
AND2X1 exu_U20234(.A(alu_byp_rd_data_e[0]), .B(exu_n16288), .Y(exu_n20665));
INVX1 exu_U20235(.A(exu_n20665), .Y(exu_n5609));
AND2X1 exu_U20236(.A(bypass_rs3h_data_btwn_mux[0]), .B(exu_n19220), .Y(exu_n20667));
INVX1 exu_U20237(.A(exu_n20667), .Y(exu_n5610));
AND2X1 exu_U20238(.A(exu_n16222), .B(div_yreg_yreg_thr2[9]), .Y(exu_n20671));
INVX1 exu_U20239(.A(exu_n20671), .Y(exu_n5611));
AND2X1 exu_U20240(.A(exu_n16220), .B(div_yreg_yreg_thr0[9]), .Y(exu_n20673));
INVX1 exu_U20241(.A(exu_n20673), .Y(exu_n5612));
AND2X1 exu_U20242(.A(div_yreg_yreg_thr2[8]), .B(exu_n16222), .Y(exu_n20677));
INVX1 exu_U20243(.A(exu_n20677), .Y(exu_n5613));
AND2X1 exu_U20244(.A(div_yreg_yreg_thr0[8]), .B(exu_n16220), .Y(exu_n20679));
INVX1 exu_U20245(.A(exu_n20679), .Y(exu_n5614));
AND2X1 exu_U20246(.A(div_yreg_yreg_thr2[7]), .B(exu_n16222), .Y(exu_n20683));
INVX1 exu_U20247(.A(exu_n20683), .Y(exu_n5615));
AND2X1 exu_U20248(.A(div_yreg_yreg_thr0[7]), .B(exu_n16220), .Y(exu_n20685));
INVX1 exu_U20249(.A(exu_n20685), .Y(exu_n5616));
AND2X1 exu_U20250(.A(div_yreg_yreg_thr2[6]), .B(exu_n16222), .Y(exu_n20689));
INVX1 exu_U20251(.A(exu_n20689), .Y(exu_n5617));
AND2X1 exu_U20252(.A(div_yreg_yreg_thr0[6]), .B(exu_n16220), .Y(exu_n20691));
INVX1 exu_U20253(.A(exu_n20691), .Y(exu_n5618));
AND2X1 exu_U20254(.A(div_yreg_yreg_thr2[5]), .B(exu_n16222), .Y(exu_n20695));
INVX1 exu_U20255(.A(exu_n20695), .Y(exu_n5619));
AND2X1 exu_U20256(.A(div_yreg_yreg_thr0[5]), .B(exu_n16220), .Y(exu_n20697));
INVX1 exu_U20257(.A(exu_n20697), .Y(exu_n5620));
AND2X1 exu_U20258(.A(div_yreg_yreg_thr2[4]), .B(exu_n16222), .Y(exu_n20701));
INVX1 exu_U20259(.A(exu_n20701), .Y(exu_n5621));
AND2X1 exu_U20260(.A(div_yreg_yreg_thr0[4]), .B(exu_n16220), .Y(exu_n20703));
INVX1 exu_U20261(.A(exu_n20703), .Y(exu_n5622));
AND2X1 exu_U20262(.A(div_yreg_yreg_thr2[3]), .B(exu_n16222), .Y(exu_n20707));
INVX1 exu_U20263(.A(exu_n20707), .Y(exu_n5623));
AND2X1 exu_U20264(.A(div_yreg_yreg_thr0[3]), .B(exu_n16220), .Y(exu_n20709));
INVX1 exu_U20265(.A(exu_n20709), .Y(exu_n5624));
AND2X1 exu_U20266(.A(div_yreg_yreg_thr2[31]), .B(exu_n16222), .Y(exu_n20713));
INVX1 exu_U20267(.A(exu_n20713), .Y(exu_n5625));
AND2X1 exu_U20268(.A(div_yreg_yreg_thr0[31]), .B(exu_n16220), .Y(exu_n20715));
INVX1 exu_U20269(.A(exu_n20715), .Y(exu_n5626));
AND2X1 exu_U20270(.A(div_yreg_yreg_thr2[30]), .B(exu_n16222), .Y(exu_n20719));
INVX1 exu_U20271(.A(exu_n20719), .Y(exu_n5627));
AND2X1 exu_U20272(.A(div_yreg_yreg_thr0[30]), .B(exu_n16220), .Y(exu_n20721));
INVX1 exu_U20273(.A(exu_n20721), .Y(exu_n5628));
AND2X1 exu_U20274(.A(div_yreg_yreg_thr2[2]), .B(exu_n16222), .Y(exu_n20725));
INVX1 exu_U20275(.A(exu_n20725), .Y(exu_n5629));
AND2X1 exu_U20276(.A(div_yreg_yreg_thr0[2]), .B(exu_n16220), .Y(exu_n20727));
INVX1 exu_U20277(.A(exu_n20727), .Y(exu_n5630));
AND2X1 exu_U20278(.A(div_yreg_yreg_thr2[29]), .B(exu_n16222), .Y(exu_n20731));
INVX1 exu_U20279(.A(exu_n20731), .Y(exu_n5631));
AND2X1 exu_U20280(.A(div_yreg_yreg_thr0[29]), .B(exu_n16220), .Y(exu_n20733));
INVX1 exu_U20281(.A(exu_n20733), .Y(exu_n5632));
AND2X1 exu_U20282(.A(div_yreg_yreg_thr2[28]), .B(exu_n16222), .Y(exu_n20737));
INVX1 exu_U20283(.A(exu_n20737), .Y(exu_n5633));
AND2X1 exu_U20284(.A(div_yreg_yreg_thr0[28]), .B(exu_n16220), .Y(exu_n20739));
INVX1 exu_U20285(.A(exu_n20739), .Y(exu_n5634));
AND2X1 exu_U20286(.A(div_yreg_yreg_thr2[27]), .B(exu_n16222), .Y(exu_n20743));
INVX1 exu_U20287(.A(exu_n20743), .Y(exu_n5635));
AND2X1 exu_U20288(.A(div_yreg_yreg_thr0[27]), .B(exu_n16220), .Y(exu_n20745));
INVX1 exu_U20289(.A(exu_n20745), .Y(exu_n5636));
AND2X1 exu_U20290(.A(div_yreg_yreg_thr2[26]), .B(exu_n16222), .Y(exu_n20749));
INVX1 exu_U20291(.A(exu_n20749), .Y(exu_n5637));
AND2X1 exu_U20292(.A(div_yreg_yreg_thr0[26]), .B(exu_n16220), .Y(exu_n20751));
INVX1 exu_U20293(.A(exu_n20751), .Y(exu_n5638));
AND2X1 exu_U20294(.A(div_yreg_yreg_thr2[25]), .B(exu_n16222), .Y(exu_n20755));
INVX1 exu_U20295(.A(exu_n20755), .Y(exu_n5639));
AND2X1 exu_U20296(.A(div_yreg_yreg_thr0[25]), .B(exu_n16220), .Y(exu_n20757));
INVX1 exu_U20297(.A(exu_n20757), .Y(exu_n5640));
AND2X1 exu_U20298(.A(div_yreg_yreg_thr2[24]), .B(exu_n16222), .Y(exu_n20761));
INVX1 exu_U20299(.A(exu_n20761), .Y(exu_n5641));
AND2X1 exu_U20300(.A(div_yreg_yreg_thr0[24]), .B(exu_n16220), .Y(exu_n20763));
INVX1 exu_U20301(.A(exu_n20763), .Y(exu_n5642));
AND2X1 exu_U20302(.A(div_yreg_yreg_thr2[23]), .B(exu_n16222), .Y(exu_n20767));
INVX1 exu_U20303(.A(exu_n20767), .Y(exu_n5643));
AND2X1 exu_U20304(.A(div_yreg_yreg_thr0[23]), .B(exu_n16220), .Y(exu_n20769));
INVX1 exu_U20305(.A(exu_n20769), .Y(exu_n5644));
AND2X1 exu_U20306(.A(div_yreg_yreg_thr2[22]), .B(exu_n16222), .Y(exu_n20773));
INVX1 exu_U20307(.A(exu_n20773), .Y(exu_n5645));
AND2X1 exu_U20308(.A(div_yreg_yreg_thr0[22]), .B(exu_n16220), .Y(exu_n20775));
INVX1 exu_U20309(.A(exu_n20775), .Y(exu_n5646));
AND2X1 exu_U20310(.A(div_yreg_yreg_thr2[21]), .B(exu_n16222), .Y(exu_n20779));
INVX1 exu_U20311(.A(exu_n20779), .Y(exu_n5647));
AND2X1 exu_U20312(.A(div_yreg_yreg_thr0[21]), .B(exu_n16220), .Y(exu_n20781));
INVX1 exu_U20313(.A(exu_n20781), .Y(exu_n5648));
AND2X1 exu_U20314(.A(div_yreg_yreg_thr2[20]), .B(exu_n16222), .Y(exu_n20785));
INVX1 exu_U20315(.A(exu_n20785), .Y(exu_n5649));
AND2X1 exu_U20316(.A(div_yreg_yreg_thr0[20]), .B(exu_n16220), .Y(exu_n20787));
INVX1 exu_U20317(.A(exu_n20787), .Y(exu_n5650));
AND2X1 exu_U20318(.A(div_yreg_yreg_thr2[1]), .B(exu_n16222), .Y(exu_n20791));
INVX1 exu_U20319(.A(exu_n20791), .Y(exu_n5651));
AND2X1 exu_U20320(.A(div_yreg_yreg_thr0[1]), .B(exu_n16220), .Y(exu_n20793));
INVX1 exu_U20321(.A(exu_n20793), .Y(exu_n5652));
AND2X1 exu_U20322(.A(div_yreg_yreg_thr2[19]), .B(exu_n16222), .Y(exu_n20797));
INVX1 exu_U20323(.A(exu_n20797), .Y(exu_n5653));
AND2X1 exu_U20324(.A(div_yreg_yreg_thr0[19]), .B(exu_n16220), .Y(exu_n20799));
INVX1 exu_U20325(.A(exu_n20799), .Y(exu_n5654));
AND2X1 exu_U20326(.A(div_yreg_yreg_thr2[18]), .B(exu_n16222), .Y(exu_n20803));
INVX1 exu_U20327(.A(exu_n20803), .Y(exu_n5655));
AND2X1 exu_U20328(.A(div_yreg_yreg_thr0[18]), .B(exu_n16220), .Y(exu_n20805));
INVX1 exu_U20329(.A(exu_n20805), .Y(exu_n5656));
AND2X1 exu_U20330(.A(div_yreg_yreg_thr2[17]), .B(exu_n16222), .Y(exu_n20809));
INVX1 exu_U20331(.A(exu_n20809), .Y(exu_n5657));
AND2X1 exu_U20332(.A(div_yreg_yreg_thr0[17]), .B(exu_n16220), .Y(exu_n20811));
INVX1 exu_U20333(.A(exu_n20811), .Y(exu_n5658));
AND2X1 exu_U20334(.A(div_yreg_yreg_thr2[16]), .B(exu_n16222), .Y(exu_n20815));
INVX1 exu_U20335(.A(exu_n20815), .Y(exu_n5659));
AND2X1 exu_U20336(.A(div_yreg_yreg_thr0[16]), .B(exu_n16220), .Y(exu_n20817));
INVX1 exu_U20337(.A(exu_n20817), .Y(exu_n5660));
AND2X1 exu_U20338(.A(div_yreg_yreg_thr2[15]), .B(exu_n16222), .Y(exu_n20821));
INVX1 exu_U20339(.A(exu_n20821), .Y(exu_n5661));
AND2X1 exu_U20340(.A(div_yreg_yreg_thr0[15]), .B(exu_n16220), .Y(exu_n20823));
INVX1 exu_U20341(.A(exu_n20823), .Y(exu_n5662));
AND2X1 exu_U20342(.A(div_yreg_yreg_thr2[14]), .B(exu_n16222), .Y(exu_n20827));
INVX1 exu_U20343(.A(exu_n20827), .Y(exu_n5663));
AND2X1 exu_U20344(.A(div_yreg_yreg_thr0[14]), .B(exu_n16220), .Y(exu_n20829));
INVX1 exu_U20345(.A(exu_n20829), .Y(exu_n5664));
AND2X1 exu_U20346(.A(div_yreg_yreg_thr2[13]), .B(exu_n16222), .Y(exu_n20833));
INVX1 exu_U20347(.A(exu_n20833), .Y(exu_n5665));
AND2X1 exu_U20348(.A(div_yreg_yreg_thr0[13]), .B(exu_n16220), .Y(exu_n20835));
INVX1 exu_U20349(.A(exu_n20835), .Y(exu_n5666));
AND2X1 exu_U20350(.A(div_yreg_yreg_thr2[12]), .B(exu_n16222), .Y(exu_n20839));
INVX1 exu_U20351(.A(exu_n20839), .Y(exu_n5667));
AND2X1 exu_U20352(.A(div_yreg_yreg_thr0[12]), .B(exu_n16220), .Y(exu_n20841));
INVX1 exu_U20353(.A(exu_n20841), .Y(exu_n5668));
AND2X1 exu_U20354(.A(div_yreg_yreg_thr2[11]), .B(exu_n16222), .Y(exu_n20845));
INVX1 exu_U20355(.A(exu_n20845), .Y(exu_n5669));
AND2X1 exu_U20356(.A(div_yreg_yreg_thr0[11]), .B(exu_n16220), .Y(exu_n20847));
INVX1 exu_U20357(.A(exu_n20847), .Y(exu_n5670));
AND2X1 exu_U20358(.A(div_yreg_yreg_thr2[10]), .B(exu_n16222), .Y(exu_n20851));
INVX1 exu_U20359(.A(exu_n20851), .Y(exu_n5671));
AND2X1 exu_U20360(.A(div_yreg_yreg_thr0[10]), .B(exu_n16220), .Y(exu_n20853));
INVX1 exu_U20361(.A(exu_n20853), .Y(exu_n5672));
AND2X1 exu_U20362(.A(div_yreg_div_ecl_yreg_0[2]), .B(exu_n16222), .Y(exu_n20857));
INVX1 exu_U20363(.A(exu_n20857), .Y(exu_n5673));
AND2X1 exu_U20364(.A(div_yreg_div_ecl_yreg_0[0]), .B(exu_n16220), .Y(exu_n20859));
INVX1 exu_U20365(.A(exu_n20859), .Y(exu_n5674));
AND2X1 exu_U20366(.A(ecl_div_yreg_wen_l[0]), .B(div_yreg_yreg_thr0[9]), .Y(exu_n20863));
INVX1 exu_U20367(.A(exu_n20863), .Y(exu_n5675));
AND2X1 exu_U20368(.A(exu_n16241), .B(div_yreg_yreg_data_w1[9]), .Y(exu_n20865));
INVX1 exu_U20369(.A(exu_n20865), .Y(exu_n5676));
AND2X1 exu_U20370(.A(div_yreg_yreg_thr0[8]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20869));
INVX1 exu_U20371(.A(exu_n20869), .Y(exu_n5677));
AND2X1 exu_U20372(.A(div_yreg_yreg_data_w1[8]), .B(exu_n16241), .Y(exu_n20871));
INVX1 exu_U20373(.A(exu_n20871), .Y(exu_n5678));
AND2X1 exu_U20374(.A(div_yreg_yreg_thr0[7]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20875));
INVX1 exu_U20375(.A(exu_n20875), .Y(exu_n5679));
AND2X1 exu_U20376(.A(div_yreg_yreg_data_w1[7]), .B(exu_n16241), .Y(exu_n20877));
INVX1 exu_U20377(.A(exu_n20877), .Y(exu_n5680));
AND2X1 exu_U20378(.A(div_yreg_yreg_thr0[6]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20881));
INVX1 exu_U20379(.A(exu_n20881), .Y(exu_n5681));
AND2X1 exu_U20380(.A(div_yreg_yreg_data_w1[6]), .B(exu_n16241), .Y(exu_n20883));
INVX1 exu_U20381(.A(exu_n20883), .Y(exu_n5682));
AND2X1 exu_U20382(.A(div_yreg_yreg_thr0[5]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20887));
INVX1 exu_U20383(.A(exu_n20887), .Y(exu_n5683));
AND2X1 exu_U20384(.A(div_yreg_yreg_data_w1[5]), .B(exu_n16241), .Y(exu_n20889));
INVX1 exu_U20385(.A(exu_n20889), .Y(exu_n5684));
AND2X1 exu_U20386(.A(div_yreg_yreg_thr0[4]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20893));
INVX1 exu_U20387(.A(exu_n20893), .Y(exu_n5685));
AND2X1 exu_U20388(.A(div_yreg_yreg_data_w1[4]), .B(exu_n16241), .Y(exu_n20895));
INVX1 exu_U20389(.A(exu_n20895), .Y(exu_n5686));
AND2X1 exu_U20390(.A(div_yreg_yreg_thr0[3]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20899));
INVX1 exu_U20391(.A(exu_n20899), .Y(exu_n5687));
AND2X1 exu_U20392(.A(div_yreg_yreg_data_w1[3]), .B(exu_n16241), .Y(exu_n20901));
INVX1 exu_U20393(.A(exu_n20901), .Y(exu_n5688));
AND2X1 exu_U20394(.A(div_yreg_yreg_thr0[31]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20905));
INVX1 exu_U20395(.A(exu_n20905), .Y(exu_n5689));
AND2X1 exu_U20396(.A(div_yreg_yreg_data_w1[31]), .B(exu_n16241), .Y(exu_n20907));
INVX1 exu_U20397(.A(exu_n20907), .Y(exu_n5690));
AND2X1 exu_U20398(.A(div_yreg_yreg_thr0[30]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20911));
INVX1 exu_U20399(.A(exu_n20911), .Y(exu_n5691));
AND2X1 exu_U20400(.A(div_yreg_yreg_data_w1[30]), .B(exu_n16241), .Y(exu_n20913));
INVX1 exu_U20401(.A(exu_n20913), .Y(exu_n5692));
AND2X1 exu_U20402(.A(div_yreg_yreg_thr0[2]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20917));
INVX1 exu_U20403(.A(exu_n20917), .Y(exu_n5693));
AND2X1 exu_U20404(.A(div_yreg_yreg_data_w1[2]), .B(exu_n16241), .Y(exu_n20919));
INVX1 exu_U20405(.A(exu_n20919), .Y(exu_n5694));
AND2X1 exu_U20406(.A(div_yreg_yreg_thr0[29]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20923));
INVX1 exu_U20407(.A(exu_n20923), .Y(exu_n5695));
AND2X1 exu_U20408(.A(div_yreg_yreg_data_w1[29]), .B(exu_n16241), .Y(exu_n20925));
INVX1 exu_U20409(.A(exu_n20925), .Y(exu_n5696));
AND2X1 exu_U20410(.A(div_yreg_yreg_thr0[28]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20929));
INVX1 exu_U20411(.A(exu_n20929), .Y(exu_n5697));
AND2X1 exu_U20412(.A(div_yreg_yreg_data_w1[28]), .B(exu_n16241), .Y(exu_n20931));
INVX1 exu_U20413(.A(exu_n20931), .Y(exu_n5698));
AND2X1 exu_U20414(.A(div_yreg_yreg_thr0[27]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20935));
INVX1 exu_U20415(.A(exu_n20935), .Y(exu_n5699));
AND2X1 exu_U20416(.A(div_yreg_yreg_data_w1[27]), .B(exu_n16241), .Y(exu_n20937));
INVX1 exu_U20417(.A(exu_n20937), .Y(exu_n5700));
AND2X1 exu_U20418(.A(div_yreg_yreg_thr0[26]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20941));
INVX1 exu_U20419(.A(exu_n20941), .Y(exu_n5701));
AND2X1 exu_U20420(.A(div_yreg_yreg_data_w1[26]), .B(exu_n16241), .Y(exu_n20943));
INVX1 exu_U20421(.A(exu_n20943), .Y(exu_n5702));
AND2X1 exu_U20422(.A(div_yreg_yreg_thr0[25]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20947));
INVX1 exu_U20423(.A(exu_n20947), .Y(exu_n5703));
AND2X1 exu_U20424(.A(div_yreg_yreg_data_w1[25]), .B(exu_n16241), .Y(exu_n20949));
INVX1 exu_U20425(.A(exu_n20949), .Y(exu_n5704));
AND2X1 exu_U20426(.A(div_yreg_yreg_thr0[24]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20953));
INVX1 exu_U20427(.A(exu_n20953), .Y(exu_n5705));
AND2X1 exu_U20428(.A(div_yreg_yreg_data_w1[24]), .B(exu_n16241), .Y(exu_n20955));
INVX1 exu_U20429(.A(exu_n20955), .Y(exu_n5706));
AND2X1 exu_U20430(.A(div_yreg_yreg_thr0[23]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20959));
INVX1 exu_U20431(.A(exu_n20959), .Y(exu_n5707));
AND2X1 exu_U20432(.A(div_yreg_yreg_data_w1[23]), .B(exu_n16241), .Y(exu_n20961));
INVX1 exu_U20433(.A(exu_n20961), .Y(exu_n5708));
AND2X1 exu_U20434(.A(div_yreg_yreg_thr0[22]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20965));
INVX1 exu_U20435(.A(exu_n20965), .Y(exu_n5709));
AND2X1 exu_U20436(.A(div_yreg_yreg_data_w1[22]), .B(exu_n16241), .Y(exu_n20967));
INVX1 exu_U20437(.A(exu_n20967), .Y(exu_n5710));
AND2X1 exu_U20438(.A(div_yreg_yreg_thr0[21]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20971));
INVX1 exu_U20439(.A(exu_n20971), .Y(exu_n5711));
AND2X1 exu_U20440(.A(div_yreg_yreg_data_w1[21]), .B(exu_n16241), .Y(exu_n20973));
INVX1 exu_U20441(.A(exu_n20973), .Y(exu_n5712));
AND2X1 exu_U20442(.A(div_yreg_yreg_thr0[20]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20977));
INVX1 exu_U20443(.A(exu_n20977), .Y(exu_n5713));
AND2X1 exu_U20444(.A(div_yreg_yreg_data_w1[20]), .B(exu_n16241), .Y(exu_n20979));
INVX1 exu_U20445(.A(exu_n20979), .Y(exu_n5714));
AND2X1 exu_U20446(.A(div_yreg_yreg_thr0[1]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20983));
INVX1 exu_U20447(.A(exu_n20983), .Y(exu_n5715));
AND2X1 exu_U20448(.A(div_yreg_yreg_data_w1[1]), .B(exu_n16241), .Y(exu_n20985));
INVX1 exu_U20449(.A(exu_n20985), .Y(exu_n5716));
AND2X1 exu_U20450(.A(div_yreg_yreg_thr0[19]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20989));
INVX1 exu_U20451(.A(exu_n20989), .Y(exu_n5717));
AND2X1 exu_U20452(.A(div_yreg_yreg_data_w1[19]), .B(exu_n16241), .Y(exu_n20991));
INVX1 exu_U20453(.A(exu_n20991), .Y(exu_n5718));
AND2X1 exu_U20454(.A(div_yreg_yreg_thr0[18]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n20995));
INVX1 exu_U20455(.A(exu_n20995), .Y(exu_n5719));
AND2X1 exu_U20456(.A(div_yreg_yreg_data_w1[18]), .B(exu_n16241), .Y(exu_n20997));
INVX1 exu_U20457(.A(exu_n20997), .Y(exu_n5720));
AND2X1 exu_U20458(.A(div_yreg_yreg_thr0[17]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n21001));
INVX1 exu_U20459(.A(exu_n21001), .Y(exu_n5721));
AND2X1 exu_U20460(.A(div_yreg_yreg_data_w1[17]), .B(exu_n16241), .Y(exu_n21003));
INVX1 exu_U20461(.A(exu_n21003), .Y(exu_n5722));
AND2X1 exu_U20462(.A(div_yreg_yreg_thr0[16]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n21007));
INVX1 exu_U20463(.A(exu_n21007), .Y(exu_n5723));
AND2X1 exu_U20464(.A(div_yreg_yreg_data_w1[16]), .B(exu_n16241), .Y(exu_n21009));
INVX1 exu_U20465(.A(exu_n21009), .Y(exu_n5724));
AND2X1 exu_U20466(.A(div_yreg_yreg_thr0[15]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n21013));
INVX1 exu_U20467(.A(exu_n21013), .Y(exu_n5725));
AND2X1 exu_U20468(.A(div_yreg_yreg_data_w1[15]), .B(exu_n16241), .Y(exu_n21015));
INVX1 exu_U20469(.A(exu_n21015), .Y(exu_n5726));
AND2X1 exu_U20470(.A(div_yreg_yreg_thr0[14]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n21019));
INVX1 exu_U20471(.A(exu_n21019), .Y(exu_n5727));
AND2X1 exu_U20472(.A(div_yreg_yreg_data_w1[14]), .B(exu_n16241), .Y(exu_n21021));
INVX1 exu_U20473(.A(exu_n21021), .Y(exu_n5728));
AND2X1 exu_U20474(.A(div_yreg_yreg_thr0[13]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n21025));
INVX1 exu_U20475(.A(exu_n21025), .Y(exu_n5729));
AND2X1 exu_U20476(.A(div_yreg_yreg_data_w1[13]), .B(exu_n16241), .Y(exu_n21027));
INVX1 exu_U20477(.A(exu_n21027), .Y(exu_n5730));
AND2X1 exu_U20478(.A(div_yreg_yreg_thr0[12]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n21031));
INVX1 exu_U20479(.A(exu_n21031), .Y(exu_n5731));
AND2X1 exu_U20480(.A(div_yreg_yreg_data_w1[12]), .B(exu_n16241), .Y(exu_n21033));
INVX1 exu_U20481(.A(exu_n21033), .Y(exu_n5732));
AND2X1 exu_U20482(.A(div_yreg_yreg_thr0[11]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n21037));
INVX1 exu_U20483(.A(exu_n21037), .Y(exu_n5733));
AND2X1 exu_U20484(.A(div_yreg_yreg_data_w1[11]), .B(exu_n16241), .Y(exu_n21039));
INVX1 exu_U20485(.A(exu_n21039), .Y(exu_n5734));
AND2X1 exu_U20486(.A(div_yreg_yreg_thr0[10]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n21043));
INVX1 exu_U20487(.A(exu_n21043), .Y(exu_n5735));
AND2X1 exu_U20488(.A(div_yreg_yreg_data_w1[10]), .B(exu_n16241), .Y(exu_n21045));
INVX1 exu_U20489(.A(exu_n21045), .Y(exu_n5736));
AND2X1 exu_U20490(.A(div_yreg_div_ecl_yreg_0[0]), .B(ecl_div_yreg_wen_l[0]), .Y(exu_n21049));
INVX1 exu_U20491(.A(exu_n21049), .Y(exu_n5737));
AND2X1 exu_U20492(.A(div_yreg_yreg_data_w1[0]), .B(exu_n16241), .Y(exu_n21051));
INVX1 exu_U20493(.A(exu_n21051), .Y(exu_n5738));
AND2X1 exu_U20494(.A(exu_n16242), .B(div_yreg_yreg_thr1[9]), .Y(exu_n21055));
INVX1 exu_U20495(.A(exu_n21055), .Y(exu_n5739));
AND2X1 exu_U20496(.A(ecl_div_yreg_wen_w[1]), .B(div_yreg_yreg_data_w1[9]), .Y(exu_n21057));
INVX1 exu_U20497(.A(exu_n21057), .Y(exu_n5740));
AND2X1 exu_U20498(.A(div_yreg_yreg_thr1[8]), .B(exu_n16242), .Y(exu_n21061));
INVX1 exu_U20499(.A(exu_n21061), .Y(exu_n5741));
AND2X1 exu_U20500(.A(div_yreg_yreg_data_w1[8]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21063));
INVX1 exu_U20501(.A(exu_n21063), .Y(exu_n5742));
AND2X1 exu_U20502(.A(div_yreg_yreg_thr1[7]), .B(exu_n16242), .Y(exu_n21067));
INVX1 exu_U20503(.A(exu_n21067), .Y(exu_n5743));
AND2X1 exu_U20504(.A(div_yreg_yreg_data_w1[7]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21069));
INVX1 exu_U20505(.A(exu_n21069), .Y(exu_n5744));
AND2X1 exu_U20506(.A(div_yreg_yreg_thr1[6]), .B(exu_n16242), .Y(exu_n21073));
INVX1 exu_U20507(.A(exu_n21073), .Y(exu_n5745));
AND2X1 exu_U20508(.A(div_yreg_yreg_data_w1[6]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21075));
INVX1 exu_U20509(.A(exu_n21075), .Y(exu_n5746));
AND2X1 exu_U20510(.A(div_yreg_yreg_thr1[5]), .B(exu_n16242), .Y(exu_n21079));
INVX1 exu_U20511(.A(exu_n21079), .Y(exu_n5747));
AND2X1 exu_U20512(.A(div_yreg_yreg_data_w1[5]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21081));
INVX1 exu_U20513(.A(exu_n21081), .Y(exu_n5748));
AND2X1 exu_U20514(.A(div_yreg_yreg_thr1[4]), .B(exu_n16242), .Y(exu_n21085));
INVX1 exu_U20515(.A(exu_n21085), .Y(exu_n5749));
AND2X1 exu_U20516(.A(div_yreg_yreg_data_w1[4]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21087));
INVX1 exu_U20517(.A(exu_n21087), .Y(exu_n5750));
AND2X1 exu_U20518(.A(div_yreg_yreg_thr1[3]), .B(exu_n16242), .Y(exu_n21091));
INVX1 exu_U20519(.A(exu_n21091), .Y(exu_n5751));
AND2X1 exu_U20520(.A(div_yreg_yreg_data_w1[3]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21093));
INVX1 exu_U20521(.A(exu_n21093), .Y(exu_n5752));
AND2X1 exu_U20522(.A(div_yreg_yreg_thr1[31]), .B(exu_n16242), .Y(exu_n21097));
INVX1 exu_U20523(.A(exu_n21097), .Y(exu_n5753));
AND2X1 exu_U20524(.A(div_yreg_yreg_data_w1[31]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21099));
INVX1 exu_U20525(.A(exu_n21099), .Y(exu_n5754));
AND2X1 exu_U20526(.A(div_yreg_yreg_thr1[30]), .B(exu_n16242), .Y(exu_n21103));
INVX1 exu_U20527(.A(exu_n21103), .Y(exu_n5755));
AND2X1 exu_U20528(.A(div_yreg_yreg_data_w1[30]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21105));
INVX1 exu_U20529(.A(exu_n21105), .Y(exu_n5756));
AND2X1 exu_U20530(.A(div_yreg_yreg_thr1[2]), .B(exu_n16242), .Y(exu_n21109));
INVX1 exu_U20531(.A(exu_n21109), .Y(exu_n5757));
AND2X1 exu_U20532(.A(div_yreg_yreg_data_w1[2]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21111));
INVX1 exu_U20533(.A(exu_n21111), .Y(exu_n5758));
AND2X1 exu_U20534(.A(div_yreg_yreg_thr1[29]), .B(exu_n16242), .Y(exu_n21115));
INVX1 exu_U20535(.A(exu_n21115), .Y(exu_n5759));
AND2X1 exu_U20536(.A(div_yreg_yreg_data_w1[29]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21117));
INVX1 exu_U20537(.A(exu_n21117), .Y(exu_n5760));
AND2X1 exu_U20538(.A(div_yreg_yreg_thr1[28]), .B(exu_n16242), .Y(exu_n21121));
INVX1 exu_U20539(.A(exu_n21121), .Y(exu_n5761));
AND2X1 exu_U20540(.A(div_yreg_yreg_data_w1[28]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21123));
INVX1 exu_U20541(.A(exu_n21123), .Y(exu_n5762));
AND2X1 exu_U20542(.A(div_yreg_yreg_thr1[27]), .B(exu_n16242), .Y(exu_n21127));
INVX1 exu_U20543(.A(exu_n21127), .Y(exu_n5763));
AND2X1 exu_U20544(.A(div_yreg_yreg_data_w1[27]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21129));
INVX1 exu_U20545(.A(exu_n21129), .Y(exu_n5764));
AND2X1 exu_U20546(.A(div_yreg_yreg_thr1[26]), .B(exu_n16242), .Y(exu_n21133));
INVX1 exu_U20547(.A(exu_n21133), .Y(exu_n5765));
AND2X1 exu_U20548(.A(div_yreg_yreg_data_w1[26]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21135));
INVX1 exu_U20549(.A(exu_n21135), .Y(exu_n5766));
AND2X1 exu_U20550(.A(div_yreg_yreg_thr1[25]), .B(exu_n16242), .Y(exu_n21139));
INVX1 exu_U20551(.A(exu_n21139), .Y(exu_n5767));
AND2X1 exu_U20552(.A(div_yreg_yreg_data_w1[25]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21141));
INVX1 exu_U20553(.A(exu_n21141), .Y(exu_n5768));
AND2X1 exu_U20554(.A(div_yreg_yreg_thr1[24]), .B(exu_n16242), .Y(exu_n21145));
INVX1 exu_U20555(.A(exu_n21145), .Y(exu_n5769));
AND2X1 exu_U20556(.A(div_yreg_yreg_data_w1[24]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21147));
INVX1 exu_U20557(.A(exu_n21147), .Y(exu_n5770));
AND2X1 exu_U20558(.A(div_yreg_yreg_thr1[23]), .B(exu_n16242), .Y(exu_n21151));
INVX1 exu_U20559(.A(exu_n21151), .Y(exu_n5771));
AND2X1 exu_U20560(.A(div_yreg_yreg_data_w1[23]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21153));
INVX1 exu_U20561(.A(exu_n21153), .Y(exu_n5772));
AND2X1 exu_U20562(.A(div_yreg_yreg_thr1[22]), .B(exu_n16242), .Y(exu_n21157));
INVX1 exu_U20563(.A(exu_n21157), .Y(exu_n5773));
AND2X1 exu_U20564(.A(div_yreg_yreg_data_w1[22]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21159));
INVX1 exu_U20565(.A(exu_n21159), .Y(exu_n5774));
AND2X1 exu_U20566(.A(div_yreg_yreg_thr1[21]), .B(exu_n16242), .Y(exu_n21163));
INVX1 exu_U20567(.A(exu_n21163), .Y(exu_n5775));
AND2X1 exu_U20568(.A(div_yreg_yreg_data_w1[21]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21165));
INVX1 exu_U20569(.A(exu_n21165), .Y(exu_n5776));
AND2X1 exu_U20570(.A(div_yreg_yreg_thr1[20]), .B(exu_n16242), .Y(exu_n21169));
INVX1 exu_U20571(.A(exu_n21169), .Y(exu_n5777));
AND2X1 exu_U20572(.A(div_yreg_yreg_data_w1[20]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21171));
INVX1 exu_U20573(.A(exu_n21171), .Y(exu_n5778));
AND2X1 exu_U20574(.A(div_yreg_yreg_thr1[1]), .B(exu_n16242), .Y(exu_n21175));
INVX1 exu_U20575(.A(exu_n21175), .Y(exu_n5779));
AND2X1 exu_U20576(.A(div_yreg_yreg_data_w1[1]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21177));
INVX1 exu_U20577(.A(exu_n21177), .Y(exu_n5780));
AND2X1 exu_U20578(.A(div_yreg_yreg_thr1[19]), .B(exu_n16242), .Y(exu_n21181));
INVX1 exu_U20579(.A(exu_n21181), .Y(exu_n5781));
AND2X1 exu_U20580(.A(div_yreg_yreg_data_w1[19]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21183));
INVX1 exu_U20581(.A(exu_n21183), .Y(exu_n5782));
AND2X1 exu_U20582(.A(div_yreg_yreg_thr1[18]), .B(exu_n16242), .Y(exu_n21187));
INVX1 exu_U20583(.A(exu_n21187), .Y(exu_n5783));
AND2X1 exu_U20584(.A(div_yreg_yreg_data_w1[18]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21189));
INVX1 exu_U20585(.A(exu_n21189), .Y(exu_n5784));
AND2X1 exu_U20586(.A(div_yreg_yreg_thr1[17]), .B(exu_n16242), .Y(exu_n21193));
INVX1 exu_U20587(.A(exu_n21193), .Y(exu_n5785));
AND2X1 exu_U20588(.A(div_yreg_yreg_data_w1[17]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21195));
INVX1 exu_U20589(.A(exu_n21195), .Y(exu_n5786));
AND2X1 exu_U20590(.A(div_yreg_yreg_thr1[16]), .B(exu_n16242), .Y(exu_n21199));
INVX1 exu_U20591(.A(exu_n21199), .Y(exu_n5787));
AND2X1 exu_U20592(.A(div_yreg_yreg_data_w1[16]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21201));
INVX1 exu_U20593(.A(exu_n21201), .Y(exu_n5788));
AND2X1 exu_U20594(.A(div_yreg_yreg_thr1[15]), .B(exu_n16242), .Y(exu_n21205));
INVX1 exu_U20595(.A(exu_n21205), .Y(exu_n5789));
AND2X1 exu_U20596(.A(div_yreg_yreg_data_w1[15]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21207));
INVX1 exu_U20597(.A(exu_n21207), .Y(exu_n5790));
AND2X1 exu_U20598(.A(div_yreg_yreg_thr1[14]), .B(exu_n16242), .Y(exu_n21211));
INVX1 exu_U20599(.A(exu_n21211), .Y(exu_n5791));
AND2X1 exu_U20600(.A(div_yreg_yreg_data_w1[14]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21213));
INVX1 exu_U20601(.A(exu_n21213), .Y(exu_n5792));
AND2X1 exu_U20602(.A(div_yreg_yreg_thr1[13]), .B(exu_n16242), .Y(exu_n21217));
INVX1 exu_U20603(.A(exu_n21217), .Y(exu_n5793));
AND2X1 exu_U20604(.A(div_yreg_yreg_data_w1[13]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21219));
INVX1 exu_U20605(.A(exu_n21219), .Y(exu_n5794));
AND2X1 exu_U20606(.A(div_yreg_yreg_thr1[12]), .B(exu_n16242), .Y(exu_n21223));
INVX1 exu_U20607(.A(exu_n21223), .Y(exu_n5795));
AND2X1 exu_U20608(.A(div_yreg_yreg_data_w1[12]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21225));
INVX1 exu_U20609(.A(exu_n21225), .Y(exu_n5796));
AND2X1 exu_U20610(.A(div_yreg_yreg_thr1[11]), .B(exu_n16242), .Y(exu_n21229));
INVX1 exu_U20611(.A(exu_n21229), .Y(exu_n5797));
AND2X1 exu_U20612(.A(div_yreg_yreg_data_w1[11]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21231));
INVX1 exu_U20613(.A(exu_n21231), .Y(exu_n5798));
AND2X1 exu_U20614(.A(div_yreg_yreg_thr1[10]), .B(exu_n16242), .Y(exu_n21235));
INVX1 exu_U20615(.A(exu_n21235), .Y(exu_n5799));
AND2X1 exu_U20616(.A(div_yreg_yreg_data_w1[10]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21237));
INVX1 exu_U20617(.A(exu_n21237), .Y(exu_n5800));
AND2X1 exu_U20618(.A(div_yreg_div_ecl_yreg_0[1]), .B(exu_n16242), .Y(exu_n21241));
INVX1 exu_U20619(.A(exu_n21241), .Y(exu_n5801));
AND2X1 exu_U20620(.A(div_yreg_yreg_data_w1[0]), .B(ecl_div_yreg_wen_w[1]), .Y(exu_n21243));
INVX1 exu_U20621(.A(exu_n21243), .Y(exu_n5802));
AND2X1 exu_U20622(.A(exu_n16243), .B(div_yreg_yreg_thr2[9]), .Y(exu_n21247));
INVX1 exu_U20623(.A(exu_n21247), .Y(exu_n5803));
AND2X1 exu_U20624(.A(ecl_div_yreg_wen_w[2]), .B(div_yreg_yreg_data_w1[9]), .Y(exu_n21249));
INVX1 exu_U20625(.A(exu_n21249), .Y(exu_n5804));
AND2X1 exu_U20626(.A(div_yreg_yreg_thr2[8]), .B(exu_n16243), .Y(exu_n21253));
INVX1 exu_U20627(.A(exu_n21253), .Y(exu_n5805));
AND2X1 exu_U20628(.A(div_yreg_yreg_data_w1[8]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21255));
INVX1 exu_U20629(.A(exu_n21255), .Y(exu_n5806));
AND2X1 exu_U20630(.A(div_yreg_yreg_thr2[7]), .B(exu_n16243), .Y(exu_n21259));
INVX1 exu_U20631(.A(exu_n21259), .Y(exu_n5807));
AND2X1 exu_U20632(.A(div_yreg_yreg_data_w1[7]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21261));
INVX1 exu_U20633(.A(exu_n21261), .Y(exu_n5808));
AND2X1 exu_U20634(.A(div_yreg_yreg_thr2[6]), .B(exu_n16243), .Y(exu_n21265));
INVX1 exu_U20635(.A(exu_n21265), .Y(exu_n5809));
AND2X1 exu_U20636(.A(div_yreg_yreg_data_w1[6]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21267));
INVX1 exu_U20637(.A(exu_n21267), .Y(exu_n5810));
AND2X1 exu_U20638(.A(div_yreg_yreg_thr2[5]), .B(exu_n16243), .Y(exu_n21271));
INVX1 exu_U20639(.A(exu_n21271), .Y(exu_n5811));
AND2X1 exu_U20640(.A(div_yreg_yreg_data_w1[5]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21273));
INVX1 exu_U20641(.A(exu_n21273), .Y(exu_n5812));
AND2X1 exu_U20642(.A(div_yreg_yreg_thr2[4]), .B(exu_n16243), .Y(exu_n21277));
INVX1 exu_U20643(.A(exu_n21277), .Y(exu_n5813));
AND2X1 exu_U20644(.A(div_yreg_yreg_data_w1[4]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21279));
INVX1 exu_U20645(.A(exu_n21279), .Y(exu_n5814));
AND2X1 exu_U20646(.A(div_yreg_yreg_thr2[3]), .B(exu_n16243), .Y(exu_n21283));
INVX1 exu_U20647(.A(exu_n21283), .Y(exu_n5815));
AND2X1 exu_U20648(.A(div_yreg_yreg_data_w1[3]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21285));
INVX1 exu_U20649(.A(exu_n21285), .Y(exu_n5816));
AND2X1 exu_U20650(.A(div_yreg_yreg_thr2[31]), .B(exu_n16243), .Y(exu_n21289));
INVX1 exu_U20651(.A(exu_n21289), .Y(exu_n5817));
AND2X1 exu_U20652(.A(div_yreg_yreg_data_w1[31]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21291));
INVX1 exu_U20653(.A(exu_n21291), .Y(exu_n5818));
AND2X1 exu_U20654(.A(div_yreg_yreg_thr2[30]), .B(exu_n16243), .Y(exu_n21295));
INVX1 exu_U20655(.A(exu_n21295), .Y(exu_n5819));
AND2X1 exu_U20656(.A(div_yreg_yreg_data_w1[30]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21297));
INVX1 exu_U20657(.A(exu_n21297), .Y(exu_n5820));
AND2X1 exu_U20658(.A(div_yreg_yreg_thr2[2]), .B(exu_n16243), .Y(exu_n21301));
INVX1 exu_U20659(.A(exu_n21301), .Y(exu_n5821));
AND2X1 exu_U20660(.A(div_yreg_yreg_data_w1[2]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21303));
INVX1 exu_U20661(.A(exu_n21303), .Y(exu_n5822));
AND2X1 exu_U20662(.A(div_yreg_yreg_thr2[29]), .B(exu_n16243), .Y(exu_n21307));
INVX1 exu_U20663(.A(exu_n21307), .Y(exu_n5823));
AND2X1 exu_U20664(.A(div_yreg_yreg_data_w1[29]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21309));
INVX1 exu_U20665(.A(exu_n21309), .Y(exu_n5824));
AND2X1 exu_U20666(.A(div_yreg_yreg_thr2[28]), .B(exu_n16243), .Y(exu_n21313));
INVX1 exu_U20667(.A(exu_n21313), .Y(exu_n5825));
AND2X1 exu_U20668(.A(div_yreg_yreg_data_w1[28]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21315));
INVX1 exu_U20669(.A(exu_n21315), .Y(exu_n5826));
AND2X1 exu_U20670(.A(div_yreg_yreg_thr2[27]), .B(exu_n16243), .Y(exu_n21319));
INVX1 exu_U20671(.A(exu_n21319), .Y(exu_n5827));
AND2X1 exu_U20672(.A(div_yreg_yreg_data_w1[27]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21321));
INVX1 exu_U20673(.A(exu_n21321), .Y(exu_n5828));
AND2X1 exu_U20674(.A(div_yreg_yreg_thr2[26]), .B(exu_n16243), .Y(exu_n21325));
INVX1 exu_U20675(.A(exu_n21325), .Y(exu_n5829));
AND2X1 exu_U20676(.A(div_yreg_yreg_data_w1[26]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21327));
INVX1 exu_U20677(.A(exu_n21327), .Y(exu_n5830));
AND2X1 exu_U20678(.A(div_yreg_yreg_thr2[25]), .B(exu_n16243), .Y(exu_n21331));
INVX1 exu_U20679(.A(exu_n21331), .Y(exu_n5831));
AND2X1 exu_U20680(.A(div_yreg_yreg_data_w1[25]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21333));
INVX1 exu_U20681(.A(exu_n21333), .Y(exu_n5832));
AND2X1 exu_U20682(.A(div_yreg_yreg_thr2[24]), .B(exu_n16243), .Y(exu_n21337));
INVX1 exu_U20683(.A(exu_n21337), .Y(exu_n5833));
AND2X1 exu_U20684(.A(div_yreg_yreg_data_w1[24]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21339));
INVX1 exu_U20685(.A(exu_n21339), .Y(exu_n5834));
AND2X1 exu_U20686(.A(div_yreg_yreg_thr2[23]), .B(exu_n16243), .Y(exu_n21343));
INVX1 exu_U20687(.A(exu_n21343), .Y(exu_n5835));
AND2X1 exu_U20688(.A(div_yreg_yreg_data_w1[23]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21345));
INVX1 exu_U20689(.A(exu_n21345), .Y(exu_n5836));
AND2X1 exu_U20690(.A(div_yreg_yreg_thr2[22]), .B(exu_n16243), .Y(exu_n21349));
INVX1 exu_U20691(.A(exu_n21349), .Y(exu_n5837));
AND2X1 exu_U20692(.A(div_yreg_yreg_data_w1[22]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21351));
INVX1 exu_U20693(.A(exu_n21351), .Y(exu_n5838));
AND2X1 exu_U20694(.A(div_yreg_yreg_thr2[21]), .B(exu_n16243), .Y(exu_n21355));
INVX1 exu_U20695(.A(exu_n21355), .Y(exu_n5839));
AND2X1 exu_U20696(.A(div_yreg_yreg_data_w1[21]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21357));
INVX1 exu_U20697(.A(exu_n21357), .Y(exu_n5840));
AND2X1 exu_U20698(.A(div_yreg_yreg_thr2[20]), .B(exu_n16243), .Y(exu_n21361));
INVX1 exu_U20699(.A(exu_n21361), .Y(exu_n5841));
AND2X1 exu_U20700(.A(div_yreg_yreg_data_w1[20]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21363));
INVX1 exu_U20701(.A(exu_n21363), .Y(exu_n5842));
AND2X1 exu_U20702(.A(div_yreg_yreg_thr2[1]), .B(exu_n16243), .Y(exu_n21367));
INVX1 exu_U20703(.A(exu_n21367), .Y(exu_n5843));
AND2X1 exu_U20704(.A(div_yreg_yreg_data_w1[1]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21369));
INVX1 exu_U20705(.A(exu_n21369), .Y(exu_n5844));
AND2X1 exu_U20706(.A(div_yreg_yreg_thr2[19]), .B(exu_n16243), .Y(exu_n21373));
INVX1 exu_U20707(.A(exu_n21373), .Y(exu_n5845));
AND2X1 exu_U20708(.A(div_yreg_yreg_data_w1[19]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21375));
INVX1 exu_U20709(.A(exu_n21375), .Y(exu_n5846));
AND2X1 exu_U20710(.A(div_yreg_yreg_thr2[18]), .B(exu_n16243), .Y(exu_n21379));
INVX1 exu_U20711(.A(exu_n21379), .Y(exu_n5847));
AND2X1 exu_U20712(.A(div_yreg_yreg_data_w1[18]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21381));
INVX1 exu_U20713(.A(exu_n21381), .Y(exu_n5848));
AND2X1 exu_U20714(.A(div_yreg_yreg_thr2[17]), .B(exu_n16243), .Y(exu_n21385));
INVX1 exu_U20715(.A(exu_n21385), .Y(exu_n5849));
AND2X1 exu_U20716(.A(div_yreg_yreg_data_w1[17]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21387));
INVX1 exu_U20717(.A(exu_n21387), .Y(exu_n5850));
AND2X1 exu_U20718(.A(div_yreg_yreg_thr2[16]), .B(exu_n16243), .Y(exu_n21391));
INVX1 exu_U20719(.A(exu_n21391), .Y(exu_n5851));
AND2X1 exu_U20720(.A(div_yreg_yreg_data_w1[16]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21393));
INVX1 exu_U20721(.A(exu_n21393), .Y(exu_n5852));
AND2X1 exu_U20722(.A(div_yreg_yreg_thr2[15]), .B(exu_n16243), .Y(exu_n21397));
INVX1 exu_U20723(.A(exu_n21397), .Y(exu_n5853));
AND2X1 exu_U20724(.A(div_yreg_yreg_data_w1[15]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21399));
INVX1 exu_U20725(.A(exu_n21399), .Y(exu_n5854));
AND2X1 exu_U20726(.A(div_yreg_yreg_thr2[14]), .B(exu_n16243), .Y(exu_n21403));
INVX1 exu_U20727(.A(exu_n21403), .Y(exu_n5855));
AND2X1 exu_U20728(.A(div_yreg_yreg_data_w1[14]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21405));
INVX1 exu_U20729(.A(exu_n21405), .Y(exu_n5856));
AND2X1 exu_U20730(.A(div_yreg_yreg_thr2[13]), .B(exu_n16243), .Y(exu_n21409));
INVX1 exu_U20731(.A(exu_n21409), .Y(exu_n5857));
AND2X1 exu_U20732(.A(div_yreg_yreg_data_w1[13]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21411));
INVX1 exu_U20733(.A(exu_n21411), .Y(exu_n5858));
AND2X1 exu_U20734(.A(div_yreg_yreg_thr2[12]), .B(exu_n16243), .Y(exu_n21415));
INVX1 exu_U20735(.A(exu_n21415), .Y(exu_n5859));
AND2X1 exu_U20736(.A(div_yreg_yreg_data_w1[12]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21417));
INVX1 exu_U20737(.A(exu_n21417), .Y(exu_n5860));
AND2X1 exu_U20738(.A(div_yreg_yreg_thr2[11]), .B(exu_n16243), .Y(exu_n21421));
INVX1 exu_U20739(.A(exu_n21421), .Y(exu_n5861));
AND2X1 exu_U20740(.A(div_yreg_yreg_data_w1[11]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21423));
INVX1 exu_U20741(.A(exu_n21423), .Y(exu_n5862));
AND2X1 exu_U20742(.A(div_yreg_yreg_thr2[10]), .B(exu_n16243), .Y(exu_n21427));
INVX1 exu_U20743(.A(exu_n21427), .Y(exu_n5863));
AND2X1 exu_U20744(.A(div_yreg_yreg_data_w1[10]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21429));
INVX1 exu_U20745(.A(exu_n21429), .Y(exu_n5864));
AND2X1 exu_U20746(.A(div_yreg_div_ecl_yreg_0[2]), .B(exu_n16243), .Y(exu_n21433));
INVX1 exu_U20747(.A(exu_n21433), .Y(exu_n5865));
AND2X1 exu_U20748(.A(div_yreg_yreg_data_w1[0]), .B(ecl_div_yreg_wen_w[2]), .Y(exu_n21435));
INVX1 exu_U20749(.A(exu_n21435), .Y(exu_n5866));
AND2X1 exu_U20750(.A(exu_n16244), .B(div_yreg_yreg_thr3[9]), .Y(exu_n21439));
INVX1 exu_U20751(.A(exu_n21439), .Y(exu_n5867));
AND2X1 exu_U20752(.A(ecl_div_yreg_wen_w[3]), .B(div_yreg_yreg_data_w1[9]), .Y(exu_n21441));
INVX1 exu_U20753(.A(exu_n21441), .Y(exu_n5868));
AND2X1 exu_U20754(.A(div_yreg_yreg_thr3[8]), .B(exu_n16244), .Y(exu_n21445));
INVX1 exu_U20755(.A(exu_n21445), .Y(exu_n5869));
AND2X1 exu_U20756(.A(div_yreg_yreg_data_w1[8]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21447));
INVX1 exu_U20757(.A(exu_n21447), .Y(exu_n5870));
AND2X1 exu_U20758(.A(div_yreg_yreg_thr3[7]), .B(exu_n16244), .Y(exu_n21451));
INVX1 exu_U20759(.A(exu_n21451), .Y(exu_n5871));
AND2X1 exu_U20760(.A(div_yreg_yreg_data_w1[7]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21453));
INVX1 exu_U20761(.A(exu_n21453), .Y(exu_n5872));
AND2X1 exu_U20762(.A(div_yreg_yreg_thr3[6]), .B(exu_n16244), .Y(exu_n21457));
INVX1 exu_U20763(.A(exu_n21457), .Y(exu_n5873));
AND2X1 exu_U20764(.A(div_yreg_yreg_data_w1[6]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21459));
INVX1 exu_U20765(.A(exu_n21459), .Y(exu_n5874));
AND2X1 exu_U20766(.A(div_yreg_yreg_thr3[5]), .B(exu_n16244), .Y(exu_n21463));
INVX1 exu_U20767(.A(exu_n21463), .Y(exu_n5875));
AND2X1 exu_U20768(.A(div_yreg_yreg_data_w1[5]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21465));
INVX1 exu_U20769(.A(exu_n21465), .Y(exu_n5876));
AND2X1 exu_U20770(.A(div_yreg_yreg_thr3[4]), .B(exu_n16244), .Y(exu_n21469));
INVX1 exu_U20771(.A(exu_n21469), .Y(exu_n5877));
AND2X1 exu_U20772(.A(div_yreg_yreg_data_w1[4]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21471));
INVX1 exu_U20773(.A(exu_n21471), .Y(exu_n5878));
AND2X1 exu_U20774(.A(div_yreg_yreg_thr3[3]), .B(exu_n16244), .Y(exu_n21475));
INVX1 exu_U20775(.A(exu_n21475), .Y(exu_n5879));
AND2X1 exu_U20776(.A(div_yreg_yreg_data_w1[3]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21477));
INVX1 exu_U20777(.A(exu_n21477), .Y(exu_n5880));
AND2X1 exu_U20778(.A(div_yreg_yreg_thr3[31]), .B(exu_n16244), .Y(exu_n21481));
INVX1 exu_U20779(.A(exu_n21481), .Y(exu_n5881));
AND2X1 exu_U20780(.A(div_yreg_yreg_data_w1[31]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21483));
INVX1 exu_U20781(.A(exu_n21483), .Y(exu_n5882));
AND2X1 exu_U20782(.A(div_yreg_yreg_thr3[30]), .B(exu_n16244), .Y(exu_n21487));
INVX1 exu_U20783(.A(exu_n21487), .Y(exu_n5883));
AND2X1 exu_U20784(.A(div_yreg_yreg_data_w1[30]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21489));
INVX1 exu_U20785(.A(exu_n21489), .Y(exu_n5884));
AND2X1 exu_U20786(.A(div_yreg_yreg_thr3[2]), .B(exu_n16244), .Y(exu_n21493));
INVX1 exu_U20787(.A(exu_n21493), .Y(exu_n5885));
AND2X1 exu_U20788(.A(div_yreg_yreg_data_w1[2]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21495));
INVX1 exu_U20789(.A(exu_n21495), .Y(exu_n5886));
AND2X1 exu_U20790(.A(div_yreg_yreg_thr3[29]), .B(exu_n16244), .Y(exu_n21499));
INVX1 exu_U20791(.A(exu_n21499), .Y(exu_n5887));
AND2X1 exu_U20792(.A(div_yreg_yreg_data_w1[29]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21501));
INVX1 exu_U20793(.A(exu_n21501), .Y(exu_n5888));
AND2X1 exu_U20794(.A(div_yreg_yreg_thr3[28]), .B(exu_n16244), .Y(exu_n21505));
INVX1 exu_U20795(.A(exu_n21505), .Y(exu_n5889));
AND2X1 exu_U20796(.A(div_yreg_yreg_data_w1[28]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21507));
INVX1 exu_U20797(.A(exu_n21507), .Y(exu_n5890));
AND2X1 exu_U20798(.A(div_yreg_yreg_thr3[27]), .B(exu_n16244), .Y(exu_n21511));
INVX1 exu_U20799(.A(exu_n21511), .Y(exu_n5891));
AND2X1 exu_U20800(.A(div_yreg_yreg_data_w1[27]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21513));
INVX1 exu_U20801(.A(exu_n21513), .Y(exu_n5892));
AND2X1 exu_U20802(.A(div_yreg_yreg_thr3[26]), .B(exu_n16244), .Y(exu_n21517));
INVX1 exu_U20803(.A(exu_n21517), .Y(exu_n5893));
AND2X1 exu_U20804(.A(div_yreg_yreg_data_w1[26]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21519));
INVX1 exu_U20805(.A(exu_n21519), .Y(exu_n5894));
AND2X1 exu_U20806(.A(div_yreg_yreg_thr3[25]), .B(exu_n16244), .Y(exu_n21523));
INVX1 exu_U20807(.A(exu_n21523), .Y(exu_n5895));
AND2X1 exu_U20808(.A(div_yreg_yreg_data_w1[25]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21525));
INVX1 exu_U20809(.A(exu_n21525), .Y(exu_n5896));
AND2X1 exu_U20810(.A(div_yreg_yreg_thr3[24]), .B(exu_n16244), .Y(exu_n21529));
INVX1 exu_U20811(.A(exu_n21529), .Y(exu_n5897));
AND2X1 exu_U20812(.A(div_yreg_yreg_data_w1[24]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21531));
INVX1 exu_U20813(.A(exu_n21531), .Y(exu_n5898));
AND2X1 exu_U20814(.A(div_yreg_yreg_thr3[23]), .B(exu_n16244), .Y(exu_n21535));
INVX1 exu_U20815(.A(exu_n21535), .Y(exu_n5899));
AND2X1 exu_U20816(.A(div_yreg_yreg_data_w1[23]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21537));
INVX1 exu_U20817(.A(exu_n21537), .Y(exu_n5900));
AND2X1 exu_U20818(.A(div_yreg_yreg_thr3[22]), .B(exu_n16244), .Y(exu_n21541));
INVX1 exu_U20819(.A(exu_n21541), .Y(exu_n5901));
AND2X1 exu_U20820(.A(div_yreg_yreg_data_w1[22]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21543));
INVX1 exu_U20821(.A(exu_n21543), .Y(exu_n5902));
AND2X1 exu_U20822(.A(div_yreg_yreg_thr3[21]), .B(exu_n16244), .Y(exu_n21547));
INVX1 exu_U20823(.A(exu_n21547), .Y(exu_n5903));
AND2X1 exu_U20824(.A(div_yreg_yreg_data_w1[21]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21549));
INVX1 exu_U20825(.A(exu_n21549), .Y(exu_n5904));
AND2X1 exu_U20826(.A(div_yreg_yreg_thr3[20]), .B(exu_n16244), .Y(exu_n21553));
INVX1 exu_U20827(.A(exu_n21553), .Y(exu_n5905));
AND2X1 exu_U20828(.A(div_yreg_yreg_data_w1[20]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21555));
INVX1 exu_U20829(.A(exu_n21555), .Y(exu_n5906));
AND2X1 exu_U20830(.A(div_yreg_yreg_thr3[1]), .B(exu_n16244), .Y(exu_n21559));
INVX1 exu_U20831(.A(exu_n21559), .Y(exu_n5907));
AND2X1 exu_U20832(.A(div_yreg_yreg_data_w1[1]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21561));
INVX1 exu_U20833(.A(exu_n21561), .Y(exu_n5908));
AND2X1 exu_U20834(.A(div_yreg_yreg_thr3[19]), .B(exu_n16244), .Y(exu_n21565));
INVX1 exu_U20835(.A(exu_n21565), .Y(exu_n5909));
AND2X1 exu_U20836(.A(div_yreg_yreg_data_w1[19]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21567));
INVX1 exu_U20837(.A(exu_n21567), .Y(exu_n5910));
AND2X1 exu_U20838(.A(div_yreg_yreg_thr3[18]), .B(exu_n16244), .Y(exu_n21571));
INVX1 exu_U20839(.A(exu_n21571), .Y(exu_n5911));
AND2X1 exu_U20840(.A(div_yreg_yreg_data_w1[18]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21573));
INVX1 exu_U20841(.A(exu_n21573), .Y(exu_n5912));
AND2X1 exu_U20842(.A(div_yreg_yreg_thr3[17]), .B(exu_n16244), .Y(exu_n21577));
INVX1 exu_U20843(.A(exu_n21577), .Y(exu_n5913));
AND2X1 exu_U20844(.A(div_yreg_yreg_data_w1[17]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21579));
INVX1 exu_U20845(.A(exu_n21579), .Y(exu_n5914));
AND2X1 exu_U20846(.A(div_yreg_yreg_thr3[16]), .B(exu_n16244), .Y(exu_n21583));
INVX1 exu_U20847(.A(exu_n21583), .Y(exu_n5915));
AND2X1 exu_U20848(.A(div_yreg_yreg_data_w1[16]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21585));
INVX1 exu_U20849(.A(exu_n21585), .Y(exu_n5916));
AND2X1 exu_U20850(.A(div_yreg_yreg_thr3[15]), .B(exu_n16244), .Y(exu_n21589));
INVX1 exu_U20851(.A(exu_n21589), .Y(exu_n5917));
AND2X1 exu_U20852(.A(div_yreg_yreg_data_w1[15]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21591));
INVX1 exu_U20853(.A(exu_n21591), .Y(exu_n5918));
AND2X1 exu_U20854(.A(div_yreg_yreg_thr3[14]), .B(exu_n16244), .Y(exu_n21595));
INVX1 exu_U20855(.A(exu_n21595), .Y(exu_n5919));
AND2X1 exu_U20856(.A(div_yreg_yreg_data_w1[14]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21597));
INVX1 exu_U20857(.A(exu_n21597), .Y(exu_n5920));
AND2X1 exu_U20858(.A(div_yreg_yreg_thr3[13]), .B(exu_n16244), .Y(exu_n21601));
INVX1 exu_U20859(.A(exu_n21601), .Y(exu_n5921));
AND2X1 exu_U20860(.A(div_yreg_yreg_data_w1[13]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21603));
INVX1 exu_U20861(.A(exu_n21603), .Y(exu_n5922));
AND2X1 exu_U20862(.A(div_yreg_yreg_thr3[12]), .B(exu_n16244), .Y(exu_n21607));
INVX1 exu_U20863(.A(exu_n21607), .Y(exu_n5923));
AND2X1 exu_U20864(.A(div_yreg_yreg_data_w1[12]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21609));
INVX1 exu_U20865(.A(exu_n21609), .Y(exu_n5924));
AND2X1 exu_U20866(.A(div_yreg_yreg_thr3[11]), .B(exu_n16244), .Y(exu_n21613));
INVX1 exu_U20867(.A(exu_n21613), .Y(exu_n5925));
AND2X1 exu_U20868(.A(div_yreg_yreg_data_w1[11]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21615));
INVX1 exu_U20869(.A(exu_n21615), .Y(exu_n5926));
AND2X1 exu_U20870(.A(div_yreg_yreg_thr3[10]), .B(exu_n16244), .Y(exu_n21619));
INVX1 exu_U20871(.A(exu_n21619), .Y(exu_n5927));
AND2X1 exu_U20872(.A(div_yreg_yreg_data_w1[10]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21621));
INVX1 exu_U20873(.A(exu_n21621), .Y(exu_n5928));
AND2X1 exu_U20874(.A(div_yreg_div_ecl_yreg_0[3]), .B(exu_n16244), .Y(exu_n21625));
INVX1 exu_U20875(.A(exu_n21625), .Y(exu_n5929));
AND2X1 exu_U20876(.A(div_yreg_yreg_data_w1[0]), .B(ecl_div_yreg_wen_w[3]), .Y(exu_n21627));
INVX1 exu_U20877(.A(exu_n21627), .Y(exu_n5930));
AND2X1 exu_U20878(.A(exu_n15967), .B(lsu_exu_ldxa_data_g[9]), .Y(exu_n21794));
INVX1 exu_U20879(.A(exu_n21794), .Y(exu_n5931));
AND2X1 exu_U20880(.A(exu_n16282), .B(byp_irf_rd_data_w2[9]), .Y(exu_n21796));
INVX1 exu_U20881(.A(exu_n21796), .Y(exu_n5932));
AND2X1 exu_U20882(.A(lsu_exu_ldxa_data_g[8]), .B(exu_n15967), .Y(exu_n21798));
INVX1 exu_U20883(.A(exu_n21798), .Y(exu_n5933));
AND2X1 exu_U20884(.A(byp_irf_rd_data_w2[8]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21800));
INVX1 exu_U20885(.A(exu_n21800), .Y(exu_n5934));
AND2X1 exu_U20886(.A(lsu_exu_ldxa_data_g[7]), .B(exu_n15967), .Y(exu_n21802));
INVX1 exu_U20887(.A(exu_n21802), .Y(exu_n5935));
AND2X1 exu_U20888(.A(byp_irf_rd_data_w2[7]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21804));
INVX1 exu_U20889(.A(exu_n21804), .Y(exu_n5936));
AND2X1 exu_U20890(.A(lsu_exu_ldxa_data_g[6]), .B(exu_n15967), .Y(exu_n21806));
INVX1 exu_U20891(.A(exu_n21806), .Y(exu_n5937));
AND2X1 exu_U20892(.A(byp_irf_rd_data_w2[6]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21808));
INVX1 exu_U20893(.A(exu_n21808), .Y(exu_n5938));
AND2X1 exu_U20894(.A(lsu_exu_ldxa_data_g[63]), .B(exu_n15967), .Y(exu_n21810));
INVX1 exu_U20895(.A(exu_n21810), .Y(exu_n5939));
AND2X1 exu_U20896(.A(byp_irf_rd_data_w2[63]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21812));
INVX1 exu_U20897(.A(exu_n21812), .Y(exu_n5940));
AND2X1 exu_U20898(.A(lsu_exu_ldxa_data_g[62]), .B(exu_n15967), .Y(exu_n21814));
INVX1 exu_U20899(.A(exu_n21814), .Y(exu_n5941));
AND2X1 exu_U20900(.A(byp_irf_rd_data_w2[62]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21816));
INVX1 exu_U20901(.A(exu_n21816), .Y(exu_n5942));
AND2X1 exu_U20902(.A(lsu_exu_ldxa_data_g[61]), .B(exu_n15967), .Y(exu_n21818));
INVX1 exu_U20903(.A(exu_n21818), .Y(exu_n5943));
AND2X1 exu_U20904(.A(byp_irf_rd_data_w2[61]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21820));
INVX1 exu_U20905(.A(exu_n21820), .Y(exu_n5944));
AND2X1 exu_U20906(.A(lsu_exu_ldxa_data_g[60]), .B(exu_n15967), .Y(exu_n21822));
INVX1 exu_U20907(.A(exu_n21822), .Y(exu_n5945));
AND2X1 exu_U20908(.A(byp_irf_rd_data_w2[60]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21824));
INVX1 exu_U20909(.A(exu_n21824), .Y(exu_n5946));
AND2X1 exu_U20910(.A(lsu_exu_ldxa_data_g[5]), .B(exu_n15967), .Y(exu_n21826));
INVX1 exu_U20911(.A(exu_n21826), .Y(exu_n5947));
AND2X1 exu_U20912(.A(byp_irf_rd_data_w2[5]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21828));
INVX1 exu_U20913(.A(exu_n21828), .Y(exu_n5948));
AND2X1 exu_U20914(.A(lsu_exu_ldxa_data_g[59]), .B(exu_n15967), .Y(exu_n21830));
INVX1 exu_U20915(.A(exu_n21830), .Y(exu_n5949));
AND2X1 exu_U20916(.A(byp_irf_rd_data_w2[59]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21832));
INVX1 exu_U20917(.A(exu_n21832), .Y(exu_n5950));
AND2X1 exu_U20918(.A(lsu_exu_ldxa_data_g[58]), .B(exu_n15967), .Y(exu_n21834));
INVX1 exu_U20919(.A(exu_n21834), .Y(exu_n5951));
AND2X1 exu_U20920(.A(byp_irf_rd_data_w2[58]), .B(exu_n16282), .Y(exu_n21836));
INVX1 exu_U20921(.A(exu_n21836), .Y(exu_n5952));
AND2X1 exu_U20922(.A(lsu_exu_ldxa_data_g[57]), .B(exu_n15967), .Y(exu_n21838));
INVX1 exu_U20923(.A(exu_n21838), .Y(exu_n5953));
AND2X1 exu_U20924(.A(byp_irf_rd_data_w2[57]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21840));
INVX1 exu_U20925(.A(exu_n21840), .Y(exu_n5954));
AND2X1 exu_U20926(.A(lsu_exu_ldxa_data_g[56]), .B(exu_n15967), .Y(exu_n21842));
INVX1 exu_U20927(.A(exu_n21842), .Y(exu_n5955));
AND2X1 exu_U20928(.A(byp_irf_rd_data_w2[56]), .B(exu_n16282), .Y(exu_n21844));
INVX1 exu_U20929(.A(exu_n21844), .Y(exu_n5956));
AND2X1 exu_U20930(.A(lsu_exu_ldxa_data_g[55]), .B(ecl_byplog_rs1_n22), .Y(exu_n21846));
INVX1 exu_U20931(.A(exu_n21846), .Y(exu_n5957));
AND2X1 exu_U20932(.A(byp_irf_rd_data_w2[55]), .B(exu_n16282), .Y(exu_n21848));
INVX1 exu_U20933(.A(exu_n21848), .Y(exu_n5958));
AND2X1 exu_U20934(.A(lsu_exu_ldxa_data_g[54]), .B(ecl_byplog_rs1_n22), .Y(exu_n21850));
INVX1 exu_U20935(.A(exu_n21850), .Y(exu_n5959));
AND2X1 exu_U20936(.A(byp_irf_rd_data_w2[54]), .B(exu_n16282), .Y(exu_n21852));
INVX1 exu_U20937(.A(exu_n21852), .Y(exu_n5960));
AND2X1 exu_U20938(.A(lsu_exu_ldxa_data_g[53]), .B(ecl_byplog_rs1_n22), .Y(exu_n21854));
INVX1 exu_U20939(.A(exu_n21854), .Y(exu_n5961));
AND2X1 exu_U20940(.A(byp_irf_rd_data_w2[53]), .B(exu_n16282), .Y(exu_n21856));
INVX1 exu_U20941(.A(exu_n21856), .Y(exu_n5962));
AND2X1 exu_U20942(.A(lsu_exu_ldxa_data_g[52]), .B(exu_n15967), .Y(exu_n21858));
INVX1 exu_U20943(.A(exu_n21858), .Y(exu_n5963));
AND2X1 exu_U20944(.A(byp_irf_rd_data_w2[52]), .B(exu_n16282), .Y(exu_n21860));
INVX1 exu_U20945(.A(exu_n21860), .Y(exu_n5964));
AND2X1 exu_U20946(.A(lsu_exu_ldxa_data_g[51]), .B(ecl_byplog_rs1_n22), .Y(exu_n21862));
INVX1 exu_U20947(.A(exu_n21862), .Y(exu_n5965));
AND2X1 exu_U20948(.A(byp_irf_rd_data_w2[51]), .B(exu_n16282), .Y(exu_n21864));
INVX1 exu_U20949(.A(exu_n21864), .Y(exu_n5966));
AND2X1 exu_U20950(.A(lsu_exu_ldxa_data_g[50]), .B(ecl_byplog_rs1_n22), .Y(exu_n21866));
INVX1 exu_U20951(.A(exu_n21866), .Y(exu_n5967));
AND2X1 exu_U20952(.A(byp_irf_rd_data_w2[50]), .B(exu_n16282), .Y(exu_n21868));
INVX1 exu_U20953(.A(exu_n21868), .Y(exu_n5968));
AND2X1 exu_U20954(.A(lsu_exu_ldxa_data_g[4]), .B(ecl_byplog_rs1_n22), .Y(exu_n21870));
INVX1 exu_U20955(.A(exu_n21870), .Y(exu_n5969));
AND2X1 exu_U20956(.A(byp_irf_rd_data_w2[4]), .B(exu_n16282), .Y(exu_n21872));
INVX1 exu_U20957(.A(exu_n21872), .Y(exu_n5970));
AND2X1 exu_U20958(.A(lsu_exu_ldxa_data_g[49]), .B(exu_n15967), .Y(exu_n21874));
INVX1 exu_U20959(.A(exu_n21874), .Y(exu_n5971));
AND2X1 exu_U20960(.A(byp_irf_rd_data_w2[49]), .B(exu_n16282), .Y(exu_n21876));
INVX1 exu_U20961(.A(exu_n21876), .Y(exu_n5972));
AND2X1 exu_U20962(.A(lsu_exu_ldxa_data_g[48]), .B(ecl_byplog_rs1_n22), .Y(exu_n21878));
INVX1 exu_U20963(.A(exu_n21878), .Y(exu_n5973));
AND2X1 exu_U20964(.A(byp_irf_rd_data_w2[48]), .B(exu_n16282), .Y(exu_n21880));
INVX1 exu_U20965(.A(exu_n21880), .Y(exu_n5974));
AND2X1 exu_U20966(.A(lsu_exu_ldxa_data_g[47]), .B(ecl_byplog_rs1_n22), .Y(exu_n21882));
INVX1 exu_U20967(.A(exu_n21882), .Y(exu_n5975));
AND2X1 exu_U20968(.A(byp_irf_rd_data_w2[47]), .B(exu_n16282), .Y(exu_n21884));
INVX1 exu_U20969(.A(exu_n21884), .Y(exu_n5976));
AND2X1 exu_U20970(.A(lsu_exu_ldxa_data_g[46]), .B(ecl_byplog_rs1_n22), .Y(exu_n21886));
INVX1 exu_U20971(.A(exu_n21886), .Y(exu_n5977));
AND2X1 exu_U20972(.A(byp_irf_rd_data_w2[46]), .B(exu_n16282), .Y(exu_n21888));
INVX1 exu_U20973(.A(exu_n21888), .Y(exu_n5978));
AND2X1 exu_U20974(.A(lsu_exu_ldxa_data_g[45]), .B(exu_n15967), .Y(exu_n21890));
INVX1 exu_U20975(.A(exu_n21890), .Y(exu_n5979));
AND2X1 exu_U20976(.A(byp_irf_rd_data_w2[45]), .B(exu_n16282), .Y(exu_n21892));
INVX1 exu_U20977(.A(exu_n21892), .Y(exu_n5980));
AND2X1 exu_U20978(.A(lsu_exu_ldxa_data_g[44]), .B(ecl_byplog_rs1_n22), .Y(exu_n21894));
INVX1 exu_U20979(.A(exu_n21894), .Y(exu_n5981));
AND2X1 exu_U20980(.A(byp_irf_rd_data_w2[44]), .B(exu_n16282), .Y(exu_n21896));
INVX1 exu_U20981(.A(exu_n21896), .Y(exu_n5982));
AND2X1 exu_U20982(.A(lsu_exu_ldxa_data_g[43]), .B(ecl_byplog_rs1_n22), .Y(exu_n21898));
INVX1 exu_U20983(.A(exu_n21898), .Y(exu_n5983));
AND2X1 exu_U20984(.A(byp_irf_rd_data_w2[43]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21900));
INVX1 exu_U20985(.A(exu_n21900), .Y(exu_n5984));
AND2X1 exu_U20986(.A(lsu_exu_ldxa_data_g[42]), .B(ecl_byplog_rs1_n22), .Y(exu_n21902));
INVX1 exu_U20987(.A(exu_n21902), .Y(exu_n5985));
AND2X1 exu_U20988(.A(byp_irf_rd_data_w2[42]), .B(exu_n16282), .Y(exu_n21904));
INVX1 exu_U20989(.A(exu_n21904), .Y(exu_n5986));
AND2X1 exu_U20990(.A(lsu_exu_ldxa_data_g[41]), .B(exu_n15967), .Y(exu_n21906));
INVX1 exu_U20991(.A(exu_n21906), .Y(exu_n5987));
AND2X1 exu_U20992(.A(byp_irf_rd_data_w2[41]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21908));
INVX1 exu_U20993(.A(exu_n21908), .Y(exu_n5988));
AND2X1 exu_U20994(.A(lsu_exu_ldxa_data_g[40]), .B(ecl_byplog_rs1_n22), .Y(exu_n21910));
INVX1 exu_U20995(.A(exu_n21910), .Y(exu_n5989));
AND2X1 exu_U20996(.A(byp_irf_rd_data_w2[40]), .B(exu_n16282), .Y(exu_n21912));
INVX1 exu_U20997(.A(exu_n21912), .Y(exu_n5990));
AND2X1 exu_U20998(.A(lsu_exu_ldxa_data_g[3]), .B(exu_n15967), .Y(exu_n21914));
INVX1 exu_U20999(.A(exu_n21914), .Y(exu_n5991));
AND2X1 exu_U21000(.A(byp_irf_rd_data_w2[3]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21916));
INVX1 exu_U21001(.A(exu_n21916), .Y(exu_n5992));
AND2X1 exu_U21002(.A(lsu_exu_ldxa_data_g[39]), .B(exu_n15967), .Y(exu_n21918));
INVX1 exu_U21003(.A(exu_n21918), .Y(exu_n5993));
AND2X1 exu_U21004(.A(byp_irf_rd_data_w2[39]), .B(exu_n16282), .Y(exu_n21920));
INVX1 exu_U21005(.A(exu_n21920), .Y(exu_n5994));
AND2X1 exu_U21006(.A(lsu_exu_ldxa_data_g[38]), .B(ecl_byplog_rs1_n22), .Y(exu_n21922));
INVX1 exu_U21007(.A(exu_n21922), .Y(exu_n5995));
AND2X1 exu_U21008(.A(byp_irf_rd_data_w2[38]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21924));
INVX1 exu_U21009(.A(exu_n21924), .Y(exu_n5996));
AND2X1 exu_U21010(.A(lsu_exu_ldxa_data_g[37]), .B(ecl_byplog_rs1_n22), .Y(exu_n21926));
INVX1 exu_U21011(.A(exu_n21926), .Y(exu_n5997));
AND2X1 exu_U21012(.A(byp_irf_rd_data_w2[37]), .B(exu_n16282), .Y(exu_n21928));
INVX1 exu_U21013(.A(exu_n21928), .Y(exu_n5998));
AND2X1 exu_U21014(.A(lsu_exu_ldxa_data_g[36]), .B(exu_n15967), .Y(exu_n21930));
INVX1 exu_U21015(.A(exu_n21930), .Y(exu_n5999));
AND2X1 exu_U21016(.A(byp_irf_rd_data_w2[36]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21932));
INVX1 exu_U21017(.A(exu_n21932), .Y(exu_n6000));
AND2X1 exu_U21018(.A(lsu_exu_ldxa_data_g[35]), .B(ecl_byplog_rs1_n22), .Y(exu_n21934));
INVX1 exu_U21019(.A(exu_n21934), .Y(exu_n6001));
AND2X1 exu_U21020(.A(byp_irf_rd_data_w2[35]), .B(exu_n16282), .Y(exu_n21936));
INVX1 exu_U21021(.A(exu_n21936), .Y(exu_n6002));
AND2X1 exu_U21022(.A(lsu_exu_ldxa_data_g[34]), .B(exu_n15967), .Y(exu_n21938));
INVX1 exu_U21023(.A(exu_n21938), .Y(exu_n6003));
AND2X1 exu_U21024(.A(byp_irf_rd_data_w2[34]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21940));
INVX1 exu_U21025(.A(exu_n21940), .Y(exu_n6004));
AND2X1 exu_U21026(.A(lsu_exu_ldxa_data_g[33]), .B(exu_n15967), .Y(exu_n21942));
INVX1 exu_U21027(.A(exu_n21942), .Y(exu_n6005));
AND2X1 exu_U21028(.A(byp_irf_rd_data_w2[33]), .B(exu_n16282), .Y(exu_n21944));
INVX1 exu_U21029(.A(exu_n21944), .Y(exu_n6006));
AND2X1 exu_U21030(.A(lsu_exu_ldxa_data_g[32]), .B(ecl_byplog_rs1_n22), .Y(exu_n21946));
INVX1 exu_U21031(.A(exu_n21946), .Y(exu_n6007));
AND2X1 exu_U21032(.A(byp_irf_rd_data_w2[32]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21948));
INVX1 exu_U21033(.A(exu_n21948), .Y(exu_n6008));
AND2X1 exu_U21034(.A(lsu_exu_ldxa_data_g[31]), .B(ecl_byplog_rs1_n22), .Y(exu_n21950));
INVX1 exu_U21035(.A(exu_n21950), .Y(exu_n6009));
AND2X1 exu_U21036(.A(byp_irf_rd_data_w2[31]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21952));
INVX1 exu_U21037(.A(exu_n21952), .Y(exu_n6010));
AND2X1 exu_U21038(.A(lsu_exu_ldxa_data_g[30]), .B(exu_n15967), .Y(exu_n21954));
INVX1 exu_U21039(.A(exu_n21954), .Y(exu_n6011));
AND2X1 exu_U21040(.A(byp_irf_rd_data_w2[30]), .B(exu_n16282), .Y(exu_n21956));
INVX1 exu_U21041(.A(exu_n21956), .Y(exu_n6012));
AND2X1 exu_U21042(.A(lsu_exu_ldxa_data_g[2]), .B(exu_n15967), .Y(exu_n21958));
INVX1 exu_U21043(.A(exu_n21958), .Y(exu_n6013));
AND2X1 exu_U21044(.A(byp_irf_rd_data_w2[2]), .B(exu_n16282), .Y(exu_n21960));
INVX1 exu_U21045(.A(exu_n21960), .Y(exu_n6014));
AND2X1 exu_U21046(.A(lsu_exu_ldxa_data_g[29]), .B(ecl_byplog_rs1_n22), .Y(exu_n21962));
INVX1 exu_U21047(.A(exu_n21962), .Y(exu_n6015));
AND2X1 exu_U21048(.A(byp_irf_rd_data_w2[29]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21964));
INVX1 exu_U21049(.A(exu_n21964), .Y(exu_n6016));
AND2X1 exu_U21050(.A(lsu_exu_ldxa_data_g[28]), .B(ecl_byplog_rs1_n22), .Y(exu_n21966));
INVX1 exu_U21051(.A(exu_n21966), .Y(exu_n6017));
AND2X1 exu_U21052(.A(byp_irf_rd_data_w2[28]), .B(exu_n16282), .Y(exu_n21968));
INVX1 exu_U21053(.A(exu_n21968), .Y(exu_n6018));
AND2X1 exu_U21054(.A(lsu_exu_ldxa_data_g[27]), .B(ecl_byplog_rs1_n22), .Y(exu_n21970));
INVX1 exu_U21055(.A(exu_n21970), .Y(exu_n6019));
AND2X1 exu_U21056(.A(byp_irf_rd_data_w2[27]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21972));
INVX1 exu_U21057(.A(exu_n21972), .Y(exu_n6020));
AND2X1 exu_U21058(.A(lsu_exu_ldxa_data_g[26]), .B(exu_n15967), .Y(exu_n21974));
INVX1 exu_U21059(.A(exu_n21974), .Y(exu_n6021));
AND2X1 exu_U21060(.A(byp_irf_rd_data_w2[26]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21976));
INVX1 exu_U21061(.A(exu_n21976), .Y(exu_n6022));
AND2X1 exu_U21062(.A(lsu_exu_ldxa_data_g[25]), .B(ecl_byplog_rs1_n22), .Y(exu_n21978));
INVX1 exu_U21063(.A(exu_n21978), .Y(exu_n6023));
AND2X1 exu_U21064(.A(byp_irf_rd_data_w2[25]), .B(exu_n16282), .Y(exu_n21980));
INVX1 exu_U21065(.A(exu_n21980), .Y(exu_n6024));
AND2X1 exu_U21066(.A(lsu_exu_ldxa_data_g[24]), .B(exu_n15967), .Y(exu_n21982));
INVX1 exu_U21067(.A(exu_n21982), .Y(exu_n6025));
AND2X1 exu_U21068(.A(byp_irf_rd_data_w2[24]), .B(exu_n16282), .Y(exu_n21984));
INVX1 exu_U21069(.A(exu_n21984), .Y(exu_n6026));
AND2X1 exu_U21070(.A(lsu_exu_ldxa_data_g[23]), .B(ecl_byplog_rs1_n22), .Y(exu_n21986));
INVX1 exu_U21071(.A(exu_n21986), .Y(exu_n6027));
AND2X1 exu_U21072(.A(byp_irf_rd_data_w2[23]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21988));
INVX1 exu_U21073(.A(exu_n21988), .Y(exu_n6028));
AND2X1 exu_U21074(.A(lsu_exu_ldxa_data_g[22]), .B(ecl_byplog_rs1_n22), .Y(exu_n21990));
INVX1 exu_U21075(.A(exu_n21990), .Y(exu_n6029));
AND2X1 exu_U21076(.A(byp_irf_rd_data_w2[22]), .B(exu_n16282), .Y(exu_n21992));
INVX1 exu_U21077(.A(exu_n21992), .Y(exu_n6030));
AND2X1 exu_U21078(.A(lsu_exu_ldxa_data_g[21]), .B(exu_n15967), .Y(exu_n21994));
INVX1 exu_U21079(.A(exu_n21994), .Y(exu_n6031));
AND2X1 exu_U21080(.A(byp_irf_rd_data_w2[21]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n21996));
INVX1 exu_U21081(.A(exu_n21996), .Y(exu_n6032));
AND2X1 exu_U21082(.A(lsu_exu_ldxa_data_g[20]), .B(exu_n15967), .Y(exu_n21998));
INVX1 exu_U21083(.A(exu_n21998), .Y(exu_n6033));
AND2X1 exu_U21084(.A(byp_irf_rd_data_w2[20]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n22000));
INVX1 exu_U21085(.A(exu_n22000), .Y(exu_n6034));
AND2X1 exu_U21086(.A(lsu_exu_ldxa_data_g[1]), .B(ecl_byplog_rs1_n22), .Y(exu_n22002));
INVX1 exu_U21087(.A(exu_n22002), .Y(exu_n6035));
AND2X1 exu_U21088(.A(byp_irf_rd_data_w2[1]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n22004));
INVX1 exu_U21089(.A(exu_n22004), .Y(exu_n6036));
AND2X1 exu_U21090(.A(lsu_exu_ldxa_data_g[19]), .B(exu_n15967), .Y(exu_n22006));
INVX1 exu_U21091(.A(exu_n22006), .Y(exu_n6037));
AND2X1 exu_U21092(.A(byp_irf_rd_data_w2[19]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n22008));
INVX1 exu_U21093(.A(exu_n22008), .Y(exu_n6038));
AND2X1 exu_U21094(.A(lsu_exu_ldxa_data_g[18]), .B(ecl_byplog_rs1_n22), .Y(exu_n22010));
INVX1 exu_U21095(.A(exu_n22010), .Y(exu_n6039));
AND2X1 exu_U21096(.A(byp_irf_rd_data_w2[18]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n22012));
INVX1 exu_U21097(.A(exu_n22012), .Y(exu_n6040));
AND2X1 exu_U21098(.A(lsu_exu_ldxa_data_g[17]), .B(exu_n15967), .Y(exu_n22014));
INVX1 exu_U21099(.A(exu_n22014), .Y(exu_n6041));
AND2X1 exu_U21100(.A(byp_irf_rd_data_w2[17]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n22016));
INVX1 exu_U21101(.A(exu_n22016), .Y(exu_n6042));
AND2X1 exu_U21102(.A(lsu_exu_ldxa_data_g[16]), .B(ecl_byplog_rs1_n22), .Y(exu_n22018));
INVX1 exu_U21103(.A(exu_n22018), .Y(exu_n6043));
AND2X1 exu_U21104(.A(byp_irf_rd_data_w2[16]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n22020));
INVX1 exu_U21105(.A(exu_n22020), .Y(exu_n6044));
AND2X1 exu_U21106(.A(lsu_exu_ldxa_data_g[15]), .B(ecl_byplog_rs1_n22), .Y(exu_n22022));
INVX1 exu_U21107(.A(exu_n22022), .Y(exu_n6045));
AND2X1 exu_U21108(.A(byp_irf_rd_data_w2[15]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n22024));
INVX1 exu_U21109(.A(exu_n22024), .Y(exu_n6046));
AND2X1 exu_U21110(.A(lsu_exu_ldxa_data_g[14]), .B(ecl_byplog_rs1_n22), .Y(exu_n22026));
INVX1 exu_U21111(.A(exu_n22026), .Y(exu_n6047));
AND2X1 exu_U21112(.A(byp_irf_rd_data_w2[14]), .B(exu_n16282), .Y(exu_n22028));
INVX1 exu_U21113(.A(exu_n22028), .Y(exu_n6048));
AND2X1 exu_U21114(.A(lsu_exu_ldxa_data_g[13]), .B(exu_n15967), .Y(exu_n22030));
INVX1 exu_U21115(.A(exu_n22030), .Y(exu_n6049));
AND2X1 exu_U21116(.A(byp_irf_rd_data_w2[13]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n22032));
INVX1 exu_U21117(.A(exu_n22032), .Y(exu_n6050));
AND2X1 exu_U21118(.A(lsu_exu_ldxa_data_g[12]), .B(ecl_byplog_rs1_n22), .Y(exu_n22034));
INVX1 exu_U21119(.A(exu_n22034), .Y(exu_n6051));
AND2X1 exu_U21120(.A(byp_irf_rd_data_w2[12]), .B(exu_n16282), .Y(exu_n22036));
INVX1 exu_U21121(.A(exu_n22036), .Y(exu_n6052));
AND2X1 exu_U21122(.A(lsu_exu_ldxa_data_g[11]), .B(ecl_byplog_rs1_n22), .Y(exu_n22038));
INVX1 exu_U21123(.A(exu_n22038), .Y(exu_n6053));
AND2X1 exu_U21124(.A(byp_irf_rd_data_w2[11]), .B(exu_n16282), .Y(exu_n22040));
INVX1 exu_U21125(.A(exu_n22040), .Y(exu_n6054));
AND2X1 exu_U21126(.A(lsu_exu_ldxa_data_g[10]), .B(ecl_byplog_rs1_n22), .Y(exu_n22042));
INVX1 exu_U21127(.A(exu_n22042), .Y(exu_n6055));
AND2X1 exu_U21128(.A(byp_irf_rd_data_w2[10]), .B(exu_n16282), .Y(exu_n22044));
INVX1 exu_U21129(.A(exu_n22044), .Y(exu_n6056));
AND2X1 exu_U21130(.A(lsu_exu_ldxa_data_g[0]), .B(exu_n15967), .Y(exu_n22046));
INVX1 exu_U21131(.A(exu_n22046), .Y(exu_n6057));
AND2X1 exu_U21132(.A(byp_irf_rd_data_w2[0]), .B(ecl_byp_rs1_longmux_sel_w2), .Y(exu_n22048));
INVX1 exu_U21133(.A(exu_n22048), .Y(exu_n6058));
AND2X1 exu_U21134(.A(exu_n16279), .B(byp_irf_rd_data_w2[9]), .Y(exu_n22052));
INVX1 exu_U21135(.A(exu_n22052), .Y(exu_n6059));
AND2X1 exu_U21136(.A(lsu_exu_ldxa_data_g[8]), .B(exu_n15966), .Y(exu_n22054));
INVX1 exu_U21137(.A(exu_n22054), .Y(exu_n6060));
AND2X1 exu_U21138(.A(byp_irf_rd_data_w2[8]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22056));
INVX1 exu_U21139(.A(exu_n22056), .Y(exu_n6061));
AND2X1 exu_U21140(.A(lsu_exu_ldxa_data_g[7]), .B(exu_n15966), .Y(exu_n22058));
INVX1 exu_U21141(.A(exu_n22058), .Y(exu_n6062));
AND2X1 exu_U21142(.A(byp_irf_rd_data_w2[7]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22060));
INVX1 exu_U21143(.A(exu_n22060), .Y(exu_n6063));
AND2X1 exu_U21144(.A(lsu_exu_ldxa_data_g[6]), .B(exu_n15966), .Y(exu_n22062));
INVX1 exu_U21145(.A(exu_n22062), .Y(exu_n6064));
AND2X1 exu_U21146(.A(byp_irf_rd_data_w2[6]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22064));
INVX1 exu_U21147(.A(exu_n22064), .Y(exu_n6065));
AND2X1 exu_U21148(.A(lsu_exu_ldxa_data_g[63]), .B(exu_n15966), .Y(exu_n22066));
INVX1 exu_U21149(.A(exu_n22066), .Y(exu_n6066));
AND2X1 exu_U21150(.A(byp_irf_rd_data_w2[63]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22068));
INVX1 exu_U21151(.A(exu_n22068), .Y(exu_n6067));
AND2X1 exu_U21152(.A(lsu_exu_ldxa_data_g[62]), .B(exu_n15966), .Y(exu_n22070));
INVX1 exu_U21153(.A(exu_n22070), .Y(exu_n6068));
AND2X1 exu_U21154(.A(byp_irf_rd_data_w2[62]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22072));
INVX1 exu_U21155(.A(exu_n22072), .Y(exu_n6069));
AND2X1 exu_U21156(.A(lsu_exu_ldxa_data_g[61]), .B(exu_n15966), .Y(exu_n22074));
INVX1 exu_U21157(.A(exu_n22074), .Y(exu_n6070));
AND2X1 exu_U21158(.A(byp_irf_rd_data_w2[61]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22076));
INVX1 exu_U21159(.A(exu_n22076), .Y(exu_n6071));
AND2X1 exu_U21160(.A(lsu_exu_ldxa_data_g[60]), .B(exu_n15966), .Y(exu_n22078));
INVX1 exu_U21161(.A(exu_n22078), .Y(exu_n6072));
AND2X1 exu_U21162(.A(byp_irf_rd_data_w2[60]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22080));
INVX1 exu_U21163(.A(exu_n22080), .Y(exu_n6073));
AND2X1 exu_U21164(.A(lsu_exu_ldxa_data_g[5]), .B(exu_n15966), .Y(exu_n22082));
INVX1 exu_U21165(.A(exu_n22082), .Y(exu_n6074));
AND2X1 exu_U21166(.A(byp_irf_rd_data_w2[5]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22084));
INVX1 exu_U21167(.A(exu_n22084), .Y(exu_n6075));
AND2X1 exu_U21168(.A(lsu_exu_ldxa_data_g[59]), .B(exu_n15966), .Y(exu_n22086));
INVX1 exu_U21169(.A(exu_n22086), .Y(exu_n6076));
AND2X1 exu_U21170(.A(byp_irf_rd_data_w2[59]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22088));
INVX1 exu_U21171(.A(exu_n22088), .Y(exu_n6077));
AND2X1 exu_U21172(.A(lsu_exu_ldxa_data_g[58]), .B(exu_n15966), .Y(exu_n22090));
INVX1 exu_U21173(.A(exu_n22090), .Y(exu_n6078));
AND2X1 exu_U21174(.A(byp_irf_rd_data_w2[58]), .B(exu_n16279), .Y(exu_n22092));
INVX1 exu_U21175(.A(exu_n22092), .Y(exu_n6079));
AND2X1 exu_U21176(.A(lsu_exu_ldxa_data_g[57]), .B(exu_n15966), .Y(exu_n22094));
INVX1 exu_U21177(.A(exu_n22094), .Y(exu_n6080));
AND2X1 exu_U21178(.A(byp_irf_rd_data_w2[57]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22096));
INVX1 exu_U21179(.A(exu_n22096), .Y(exu_n6081));
AND2X1 exu_U21180(.A(lsu_exu_ldxa_data_g[56]), .B(exu_n15966), .Y(exu_n22098));
INVX1 exu_U21181(.A(exu_n22098), .Y(exu_n6082));
AND2X1 exu_U21182(.A(byp_irf_rd_data_w2[56]), .B(exu_n16279), .Y(exu_n22100));
INVX1 exu_U21183(.A(exu_n22100), .Y(exu_n6083));
AND2X1 exu_U21184(.A(lsu_exu_ldxa_data_g[55]), .B(ecl_byplog_rs2_n20), .Y(exu_n22102));
INVX1 exu_U21185(.A(exu_n22102), .Y(exu_n6084));
AND2X1 exu_U21186(.A(byp_irf_rd_data_w2[55]), .B(exu_n16279), .Y(exu_n22104));
INVX1 exu_U21187(.A(exu_n22104), .Y(exu_n6085));
AND2X1 exu_U21188(.A(lsu_exu_ldxa_data_g[54]), .B(exu_n15966), .Y(exu_n22106));
INVX1 exu_U21189(.A(exu_n22106), .Y(exu_n6086));
AND2X1 exu_U21190(.A(byp_irf_rd_data_w2[54]), .B(exu_n16279), .Y(exu_n22108));
INVX1 exu_U21191(.A(exu_n22108), .Y(exu_n6087));
AND2X1 exu_U21192(.A(lsu_exu_ldxa_data_g[53]), .B(ecl_byplog_rs2_n20), .Y(exu_n22110));
INVX1 exu_U21193(.A(exu_n22110), .Y(exu_n6088));
AND2X1 exu_U21194(.A(byp_irf_rd_data_w2[53]), .B(exu_n16279), .Y(exu_n22112));
INVX1 exu_U21195(.A(exu_n22112), .Y(exu_n6089));
AND2X1 exu_U21196(.A(lsu_exu_ldxa_data_g[52]), .B(ecl_byplog_rs2_n20), .Y(exu_n22114));
INVX1 exu_U21197(.A(exu_n22114), .Y(exu_n6090));
AND2X1 exu_U21198(.A(byp_irf_rd_data_w2[52]), .B(exu_n16279), .Y(exu_n22116));
INVX1 exu_U21199(.A(exu_n22116), .Y(exu_n6091));
AND2X1 exu_U21200(.A(lsu_exu_ldxa_data_g[51]), .B(ecl_byplog_rs2_n20), .Y(exu_n22118));
INVX1 exu_U21201(.A(exu_n22118), .Y(exu_n6092));
AND2X1 exu_U21202(.A(byp_irf_rd_data_w2[51]), .B(exu_n16279), .Y(exu_n22120));
INVX1 exu_U21203(.A(exu_n22120), .Y(exu_n6093));
AND2X1 exu_U21204(.A(lsu_exu_ldxa_data_g[50]), .B(ecl_byplog_rs2_n20), .Y(exu_n22122));
INVX1 exu_U21205(.A(exu_n22122), .Y(exu_n6094));
AND2X1 exu_U21206(.A(byp_irf_rd_data_w2[50]), .B(exu_n16279), .Y(exu_n22124));
INVX1 exu_U21207(.A(exu_n22124), .Y(exu_n6095));
AND2X1 exu_U21208(.A(lsu_exu_ldxa_data_g[4]), .B(ecl_byplog_rs2_n20), .Y(exu_n22126));
INVX1 exu_U21209(.A(exu_n22126), .Y(exu_n6096));
AND2X1 exu_U21210(.A(byp_irf_rd_data_w2[4]), .B(exu_n16279), .Y(exu_n22128));
INVX1 exu_U21211(.A(exu_n22128), .Y(exu_n6097));
AND2X1 exu_U21212(.A(lsu_exu_ldxa_data_g[49]), .B(exu_n15966), .Y(exu_n22130));
INVX1 exu_U21213(.A(exu_n22130), .Y(exu_n6098));
AND2X1 exu_U21214(.A(byp_irf_rd_data_w2[49]), .B(exu_n16279), .Y(exu_n22132));
INVX1 exu_U21215(.A(exu_n22132), .Y(exu_n6099));
AND2X1 exu_U21216(.A(lsu_exu_ldxa_data_g[48]), .B(exu_n15966), .Y(exu_n22134));
INVX1 exu_U21217(.A(exu_n22134), .Y(exu_n6100));
AND2X1 exu_U21218(.A(byp_irf_rd_data_w2[48]), .B(exu_n16279), .Y(exu_n22136));
INVX1 exu_U21219(.A(exu_n22136), .Y(exu_n6101));
AND2X1 exu_U21220(.A(lsu_exu_ldxa_data_g[47]), .B(ecl_byplog_rs2_n20), .Y(exu_n22138));
INVX1 exu_U21221(.A(exu_n22138), .Y(exu_n6102));
AND2X1 exu_U21222(.A(byp_irf_rd_data_w2[47]), .B(exu_n16279), .Y(exu_n22140));
INVX1 exu_U21223(.A(exu_n22140), .Y(exu_n6103));
AND2X1 exu_U21224(.A(lsu_exu_ldxa_data_g[46]), .B(ecl_byplog_rs2_n20), .Y(exu_n22142));
INVX1 exu_U21225(.A(exu_n22142), .Y(exu_n6104));
AND2X1 exu_U21226(.A(byp_irf_rd_data_w2[46]), .B(exu_n16279), .Y(exu_n22144));
INVX1 exu_U21227(.A(exu_n22144), .Y(exu_n6105));
AND2X1 exu_U21228(.A(lsu_exu_ldxa_data_g[45]), .B(ecl_byplog_rs2_n20), .Y(exu_n22146));
INVX1 exu_U21229(.A(exu_n22146), .Y(exu_n6106));
AND2X1 exu_U21230(.A(byp_irf_rd_data_w2[45]), .B(exu_n16279), .Y(exu_n22148));
INVX1 exu_U21231(.A(exu_n22148), .Y(exu_n6107));
AND2X1 exu_U21232(.A(lsu_exu_ldxa_data_g[44]), .B(ecl_byplog_rs2_n20), .Y(exu_n22150));
INVX1 exu_U21233(.A(exu_n22150), .Y(exu_n6108));
AND2X1 exu_U21234(.A(byp_irf_rd_data_w2[44]), .B(exu_n16279), .Y(exu_n22152));
INVX1 exu_U21235(.A(exu_n22152), .Y(exu_n6109));
AND2X1 exu_U21236(.A(lsu_exu_ldxa_data_g[43]), .B(exu_n15966), .Y(exu_n22154));
INVX1 exu_U21237(.A(exu_n22154), .Y(exu_n6110));
AND2X1 exu_U21238(.A(byp_irf_rd_data_w2[43]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22156));
INVX1 exu_U21239(.A(exu_n22156), .Y(exu_n6111));
AND2X1 exu_U21240(.A(lsu_exu_ldxa_data_g[42]), .B(exu_n15966), .Y(exu_n22158));
INVX1 exu_U21241(.A(exu_n22158), .Y(exu_n6112));
AND2X1 exu_U21242(.A(byp_irf_rd_data_w2[42]), .B(exu_n16279), .Y(exu_n22160));
INVX1 exu_U21243(.A(exu_n22160), .Y(exu_n6113));
AND2X1 exu_U21244(.A(lsu_exu_ldxa_data_g[41]), .B(ecl_byplog_rs2_n20), .Y(exu_n22162));
INVX1 exu_U21245(.A(exu_n22162), .Y(exu_n6114));
AND2X1 exu_U21246(.A(byp_irf_rd_data_w2[41]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22164));
INVX1 exu_U21247(.A(exu_n22164), .Y(exu_n6115));
AND2X1 exu_U21248(.A(lsu_exu_ldxa_data_g[40]), .B(ecl_byplog_rs2_n20), .Y(exu_n22166));
INVX1 exu_U21249(.A(exu_n22166), .Y(exu_n6116));
AND2X1 exu_U21250(.A(byp_irf_rd_data_w2[40]), .B(exu_n16279), .Y(exu_n22168));
INVX1 exu_U21251(.A(exu_n22168), .Y(exu_n6117));
AND2X1 exu_U21252(.A(lsu_exu_ldxa_data_g[3]), .B(exu_n15966), .Y(exu_n22170));
INVX1 exu_U21253(.A(exu_n22170), .Y(exu_n6118));
AND2X1 exu_U21254(.A(byp_irf_rd_data_w2[3]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22172));
INVX1 exu_U21255(.A(exu_n22172), .Y(exu_n6119));
AND2X1 exu_U21256(.A(lsu_exu_ldxa_data_g[39]), .B(ecl_byplog_rs2_n20), .Y(exu_n22174));
INVX1 exu_U21257(.A(exu_n22174), .Y(exu_n6120));
AND2X1 exu_U21258(.A(byp_irf_rd_data_w2[39]), .B(exu_n16279), .Y(exu_n22176));
INVX1 exu_U21259(.A(exu_n22176), .Y(exu_n6121));
AND2X1 exu_U21260(.A(lsu_exu_ldxa_data_g[38]), .B(exu_n15966), .Y(exu_n22178));
INVX1 exu_U21261(.A(exu_n22178), .Y(exu_n6122));
AND2X1 exu_U21262(.A(byp_irf_rd_data_w2[38]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22180));
INVX1 exu_U21263(.A(exu_n22180), .Y(exu_n6123));
AND2X1 exu_U21264(.A(lsu_exu_ldxa_data_g[37]), .B(ecl_byplog_rs2_n20), .Y(exu_n22182));
INVX1 exu_U21265(.A(exu_n22182), .Y(exu_n6124));
AND2X1 exu_U21266(.A(byp_irf_rd_data_w2[37]), .B(exu_n16279), .Y(exu_n22184));
INVX1 exu_U21267(.A(exu_n22184), .Y(exu_n6125));
AND2X1 exu_U21268(.A(lsu_exu_ldxa_data_g[36]), .B(exu_n15966), .Y(exu_n22186));
INVX1 exu_U21269(.A(exu_n22186), .Y(exu_n6126));
AND2X1 exu_U21270(.A(byp_irf_rd_data_w2[36]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22188));
INVX1 exu_U21271(.A(exu_n22188), .Y(exu_n6127));
AND2X1 exu_U21272(.A(lsu_exu_ldxa_data_g[35]), .B(ecl_byplog_rs2_n20), .Y(exu_n22190));
INVX1 exu_U21273(.A(exu_n22190), .Y(exu_n6128));
AND2X1 exu_U21274(.A(byp_irf_rd_data_w2[35]), .B(exu_n16279), .Y(exu_n22192));
INVX1 exu_U21275(.A(exu_n22192), .Y(exu_n6129));
AND2X1 exu_U21276(.A(lsu_exu_ldxa_data_g[34]), .B(ecl_byplog_rs2_n20), .Y(exu_n22194));
INVX1 exu_U21277(.A(exu_n22194), .Y(exu_n6130));
AND2X1 exu_U21278(.A(byp_irf_rd_data_w2[34]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22196));
INVX1 exu_U21279(.A(exu_n22196), .Y(exu_n6131));
AND2X1 exu_U21280(.A(lsu_exu_ldxa_data_g[33]), .B(ecl_byplog_rs2_n20), .Y(exu_n22198));
INVX1 exu_U21281(.A(exu_n22198), .Y(exu_n6132));
AND2X1 exu_U21282(.A(byp_irf_rd_data_w2[33]), .B(exu_n16279), .Y(exu_n22200));
INVX1 exu_U21283(.A(exu_n22200), .Y(exu_n6133));
AND2X1 exu_U21284(.A(lsu_exu_ldxa_data_g[32]), .B(exu_n15966), .Y(exu_n22202));
INVX1 exu_U21285(.A(exu_n22202), .Y(exu_n6134));
AND2X1 exu_U21286(.A(byp_irf_rd_data_w2[32]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22204));
INVX1 exu_U21287(.A(exu_n22204), .Y(exu_n6135));
AND2X1 exu_U21288(.A(lsu_exu_ldxa_data_g[31]), .B(ecl_byplog_rs2_n20), .Y(exu_n22206));
INVX1 exu_U21289(.A(exu_n22206), .Y(exu_n6136));
AND2X1 exu_U21290(.A(byp_irf_rd_data_w2[31]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22208));
INVX1 exu_U21291(.A(exu_n22208), .Y(exu_n6137));
AND2X1 exu_U21292(.A(lsu_exu_ldxa_data_g[30]), .B(exu_n15966), .Y(exu_n22210));
INVX1 exu_U21293(.A(exu_n22210), .Y(exu_n6138));
AND2X1 exu_U21294(.A(byp_irf_rd_data_w2[30]), .B(exu_n16279), .Y(exu_n22212));
INVX1 exu_U21295(.A(exu_n22212), .Y(exu_n6139));
AND2X1 exu_U21296(.A(lsu_exu_ldxa_data_g[2]), .B(ecl_byplog_rs2_n20), .Y(exu_n22214));
INVX1 exu_U21297(.A(exu_n22214), .Y(exu_n6140));
AND2X1 exu_U21298(.A(byp_irf_rd_data_w2[2]), .B(exu_n16279), .Y(exu_n22216));
INVX1 exu_U21299(.A(exu_n22216), .Y(exu_n6141));
AND2X1 exu_U21300(.A(lsu_exu_ldxa_data_g[29]), .B(exu_n15966), .Y(exu_n22218));
INVX1 exu_U21301(.A(exu_n22218), .Y(exu_n6142));
AND2X1 exu_U21302(.A(byp_irf_rd_data_w2[29]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22220));
INVX1 exu_U21303(.A(exu_n22220), .Y(exu_n6143));
AND2X1 exu_U21304(.A(lsu_exu_ldxa_data_g[28]), .B(ecl_byplog_rs2_n20), .Y(exu_n22222));
INVX1 exu_U21305(.A(exu_n22222), .Y(exu_n6144));
AND2X1 exu_U21306(.A(byp_irf_rd_data_w2[28]), .B(exu_n16279), .Y(exu_n22224));
INVX1 exu_U21307(.A(exu_n22224), .Y(exu_n6145));
AND2X1 exu_U21308(.A(lsu_exu_ldxa_data_g[27]), .B(exu_n15966), .Y(exu_n22226));
INVX1 exu_U21309(.A(exu_n22226), .Y(exu_n6146));
AND2X1 exu_U21310(.A(byp_irf_rd_data_w2[27]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22228));
INVX1 exu_U21311(.A(exu_n22228), .Y(exu_n6147));
AND2X1 exu_U21312(.A(lsu_exu_ldxa_data_g[26]), .B(exu_n15966), .Y(exu_n22230));
INVX1 exu_U21313(.A(exu_n22230), .Y(exu_n6148));
AND2X1 exu_U21314(.A(byp_irf_rd_data_w2[26]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22232));
INVX1 exu_U21315(.A(exu_n22232), .Y(exu_n6149));
AND2X1 exu_U21316(.A(lsu_exu_ldxa_data_g[25]), .B(ecl_byplog_rs2_n20), .Y(exu_n22234));
INVX1 exu_U21317(.A(exu_n22234), .Y(exu_n6150));
AND2X1 exu_U21318(.A(byp_irf_rd_data_w2[25]), .B(exu_n16279), .Y(exu_n22236));
INVX1 exu_U21319(.A(exu_n22236), .Y(exu_n6151));
AND2X1 exu_U21320(.A(lsu_exu_ldxa_data_g[24]), .B(ecl_byplog_rs2_n20), .Y(exu_n22238));
INVX1 exu_U21321(.A(exu_n22238), .Y(exu_n6152));
AND2X1 exu_U21322(.A(byp_irf_rd_data_w2[24]), .B(exu_n16279), .Y(exu_n22240));
INVX1 exu_U21323(.A(exu_n22240), .Y(exu_n6153));
AND2X1 exu_U21324(.A(lsu_exu_ldxa_data_g[23]), .B(ecl_byplog_rs2_n20), .Y(exu_n22242));
INVX1 exu_U21325(.A(exu_n22242), .Y(exu_n6154));
AND2X1 exu_U21326(.A(byp_irf_rd_data_w2[23]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22244));
INVX1 exu_U21327(.A(exu_n22244), .Y(exu_n6155));
AND2X1 exu_U21328(.A(lsu_exu_ldxa_data_g[22]), .B(exu_n15966), .Y(exu_n22246));
INVX1 exu_U21329(.A(exu_n22246), .Y(exu_n6156));
AND2X1 exu_U21330(.A(byp_irf_rd_data_w2[22]), .B(exu_n16279), .Y(exu_n22248));
INVX1 exu_U21331(.A(exu_n22248), .Y(exu_n6157));
AND2X1 exu_U21332(.A(lsu_exu_ldxa_data_g[21]), .B(ecl_byplog_rs2_n20), .Y(exu_n22250));
INVX1 exu_U21333(.A(exu_n22250), .Y(exu_n6158));
AND2X1 exu_U21334(.A(byp_irf_rd_data_w2[21]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22252));
INVX1 exu_U21335(.A(exu_n22252), .Y(exu_n6159));
AND2X1 exu_U21336(.A(lsu_exu_ldxa_data_g[20]), .B(exu_n15966), .Y(exu_n22254));
INVX1 exu_U21337(.A(exu_n22254), .Y(exu_n6160));
AND2X1 exu_U21338(.A(byp_irf_rd_data_w2[20]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22256));
INVX1 exu_U21339(.A(exu_n22256), .Y(exu_n6161));
AND2X1 exu_U21340(.A(lsu_exu_ldxa_data_g[1]), .B(ecl_byplog_rs2_n20), .Y(exu_n22258));
INVX1 exu_U21341(.A(exu_n22258), .Y(exu_n6162));
AND2X1 exu_U21342(.A(byp_irf_rd_data_w2[1]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22260));
INVX1 exu_U21343(.A(exu_n22260), .Y(exu_n6163));
AND2X1 exu_U21344(.A(lsu_exu_ldxa_data_g[19]), .B(ecl_byplog_rs2_n20), .Y(exu_n22262));
INVX1 exu_U21345(.A(exu_n22262), .Y(exu_n6164));
AND2X1 exu_U21346(.A(byp_irf_rd_data_w2[19]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22264));
INVX1 exu_U21347(.A(exu_n22264), .Y(exu_n6165));
AND2X1 exu_U21348(.A(lsu_exu_ldxa_data_g[18]), .B(exu_n15966), .Y(exu_n22266));
INVX1 exu_U21349(.A(exu_n22266), .Y(exu_n6166));
AND2X1 exu_U21350(.A(byp_irf_rd_data_w2[18]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22268));
INVX1 exu_U21351(.A(exu_n22268), .Y(exu_n6167));
AND2X1 exu_U21352(.A(lsu_exu_ldxa_data_g[17]), .B(exu_n15966), .Y(exu_n22270));
INVX1 exu_U21353(.A(exu_n22270), .Y(exu_n6168));
AND2X1 exu_U21354(.A(byp_irf_rd_data_w2[17]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22272));
INVX1 exu_U21355(.A(exu_n22272), .Y(exu_n6169));
AND2X1 exu_U21356(.A(lsu_exu_ldxa_data_g[16]), .B(ecl_byplog_rs2_n20), .Y(exu_n22274));
INVX1 exu_U21357(.A(exu_n22274), .Y(exu_n6170));
AND2X1 exu_U21358(.A(byp_irf_rd_data_w2[16]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22276));
INVX1 exu_U21359(.A(exu_n22276), .Y(exu_n6171));
AND2X1 exu_U21360(.A(lsu_exu_ldxa_data_g[15]), .B(exu_n15966), .Y(exu_n22278));
INVX1 exu_U21361(.A(exu_n22278), .Y(exu_n6172));
AND2X1 exu_U21362(.A(byp_irf_rd_data_w2[15]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22280));
INVX1 exu_U21363(.A(exu_n22280), .Y(exu_n6173));
AND2X1 exu_U21364(.A(lsu_exu_ldxa_data_g[14]), .B(ecl_byplog_rs2_n20), .Y(exu_n22282));
INVX1 exu_U21365(.A(exu_n22282), .Y(exu_n6174));
AND2X1 exu_U21366(.A(byp_irf_rd_data_w2[14]), .B(exu_n16279), .Y(exu_n22284));
INVX1 exu_U21367(.A(exu_n22284), .Y(exu_n6175));
AND2X1 exu_U21368(.A(lsu_exu_ldxa_data_g[13]), .B(ecl_byplog_rs2_n20), .Y(exu_n22286));
INVX1 exu_U21369(.A(exu_n22286), .Y(exu_n6176));
AND2X1 exu_U21370(.A(byp_irf_rd_data_w2[13]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22288));
INVX1 exu_U21371(.A(exu_n22288), .Y(exu_n6177));
AND2X1 exu_U21372(.A(lsu_exu_ldxa_data_g[12]), .B(ecl_byplog_rs2_n20), .Y(exu_n22290));
INVX1 exu_U21373(.A(exu_n22290), .Y(exu_n6178));
AND2X1 exu_U21374(.A(byp_irf_rd_data_w2[12]), .B(exu_n16279), .Y(exu_n22292));
INVX1 exu_U21375(.A(exu_n22292), .Y(exu_n6179));
AND2X1 exu_U21376(.A(lsu_exu_ldxa_data_g[11]), .B(ecl_byplog_rs2_n20), .Y(exu_n22294));
INVX1 exu_U21377(.A(exu_n22294), .Y(exu_n6180));
AND2X1 exu_U21378(.A(byp_irf_rd_data_w2[11]), .B(exu_n16279), .Y(exu_n22296));
INVX1 exu_U21379(.A(exu_n22296), .Y(exu_n6181));
AND2X1 exu_U21380(.A(lsu_exu_ldxa_data_g[10]), .B(ecl_byplog_rs2_n20), .Y(exu_n22298));
INVX1 exu_U21381(.A(exu_n22298), .Y(exu_n6182));
AND2X1 exu_U21382(.A(byp_irf_rd_data_w2[10]), .B(exu_n16279), .Y(exu_n22300));
INVX1 exu_U21383(.A(exu_n22300), .Y(exu_n6183));
AND2X1 exu_U21384(.A(lsu_exu_ldxa_data_g[0]), .B(exu_n15966), .Y(exu_n22302));
INVX1 exu_U21385(.A(exu_n22302), .Y(exu_n6184));
AND2X1 exu_U21386(.A(byp_irf_rd_data_w2[0]), .B(ecl_byp_rs2_longmux_sel_w2), .Y(exu_n22304));
INVX1 exu_U21387(.A(exu_n22304), .Y(exu_n6185));
AND2X1 exu_U21388(.A(exu_n22305), .B(exu_n10001), .Y(bypass_rs3_data_w2[9]));
INVX1 exu_U21389(.A(bypass_rs3_data_w2[9]), .Y(exu_n6186));
AND2X1 exu_U21390(.A(exu_n16276), .B(byp_irf_rd_data_w2[9]), .Y(exu_n22308));
INVX1 exu_U21391(.A(exu_n22308), .Y(exu_n6187));
AND2X1 exu_U21392(.A(byp_irf_rd_data_w2[8]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22312));
INVX1 exu_U21393(.A(exu_n22312), .Y(exu_n6188));
AND2X1 exu_U21394(.A(byp_irf_rd_data_w2[7]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22316));
INVX1 exu_U21395(.A(exu_n22316), .Y(exu_n6189));
AND2X1 exu_U21396(.A(byp_irf_rd_data_w2[6]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22320));
INVX1 exu_U21397(.A(exu_n22320), .Y(exu_n6190));
AND2X1 exu_U21398(.A(byp_irf_rd_data_w2[63]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22324));
INVX1 exu_U21399(.A(exu_n22324), .Y(exu_n6191));
AND2X1 exu_U21400(.A(byp_irf_rd_data_w2[62]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22328));
INVX1 exu_U21401(.A(exu_n22328), .Y(exu_n6192));
AND2X1 exu_U21402(.A(byp_irf_rd_data_w2[61]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22332));
INVX1 exu_U21403(.A(exu_n22332), .Y(exu_n6193));
AND2X1 exu_U21404(.A(byp_irf_rd_data_w2[60]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22336));
INVX1 exu_U21405(.A(exu_n22336), .Y(exu_n6194));
AND2X1 exu_U21406(.A(byp_irf_rd_data_w2[5]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22340));
INVX1 exu_U21407(.A(exu_n22340), .Y(exu_n6195));
AND2X1 exu_U21408(.A(byp_irf_rd_data_w2[59]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22344));
INVX1 exu_U21409(.A(exu_n22344), .Y(exu_n6196));
AND2X1 exu_U21410(.A(byp_irf_rd_data_w2[58]), .B(exu_n16276), .Y(exu_n22348));
INVX1 exu_U21411(.A(exu_n22348), .Y(exu_n6197));
AND2X1 exu_U21412(.A(byp_irf_rd_data_w2[57]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22352));
INVX1 exu_U21413(.A(exu_n22352), .Y(exu_n6198));
AND2X1 exu_U21414(.A(byp_irf_rd_data_w2[56]), .B(exu_n16276), .Y(exu_n22356));
INVX1 exu_U21415(.A(exu_n22356), .Y(exu_n6199));
AND2X1 exu_U21416(.A(byp_irf_rd_data_w2[55]), .B(exu_n16276), .Y(exu_n22360));
INVX1 exu_U21417(.A(exu_n22360), .Y(exu_n6200));
AND2X1 exu_U21418(.A(byp_irf_rd_data_w2[54]), .B(exu_n16276), .Y(exu_n22364));
INVX1 exu_U21419(.A(exu_n22364), .Y(exu_n6201));
AND2X1 exu_U21420(.A(byp_irf_rd_data_w2[53]), .B(exu_n16276), .Y(exu_n22368));
INVX1 exu_U21421(.A(exu_n22368), .Y(exu_n6202));
AND2X1 exu_U21422(.A(byp_irf_rd_data_w2[52]), .B(exu_n16276), .Y(exu_n22372));
INVX1 exu_U21423(.A(exu_n22372), .Y(exu_n6203));
AND2X1 exu_U21424(.A(byp_irf_rd_data_w2[51]), .B(exu_n16276), .Y(exu_n22376));
INVX1 exu_U21425(.A(exu_n22376), .Y(exu_n6204));
AND2X1 exu_U21426(.A(byp_irf_rd_data_w2[50]), .B(exu_n16276), .Y(exu_n22380));
INVX1 exu_U21427(.A(exu_n22380), .Y(exu_n6205));
AND2X1 exu_U21428(.A(byp_irf_rd_data_w2[4]), .B(exu_n16276), .Y(exu_n22384));
INVX1 exu_U21429(.A(exu_n22384), .Y(exu_n6206));
AND2X1 exu_U21430(.A(byp_irf_rd_data_w2[49]), .B(exu_n16276), .Y(exu_n22388));
INVX1 exu_U21431(.A(exu_n22388), .Y(exu_n6207));
AND2X1 exu_U21432(.A(byp_irf_rd_data_w2[48]), .B(exu_n16276), .Y(exu_n22392));
INVX1 exu_U21433(.A(exu_n22392), .Y(exu_n6208));
AND2X1 exu_U21434(.A(byp_irf_rd_data_w2[47]), .B(exu_n16276), .Y(exu_n22396));
INVX1 exu_U21435(.A(exu_n22396), .Y(exu_n6209));
AND2X1 exu_U21436(.A(byp_irf_rd_data_w2[46]), .B(exu_n16276), .Y(exu_n22400));
INVX1 exu_U21437(.A(exu_n22400), .Y(exu_n6210));
AND2X1 exu_U21438(.A(byp_irf_rd_data_w2[45]), .B(exu_n16276), .Y(exu_n22404));
INVX1 exu_U21439(.A(exu_n22404), .Y(exu_n6211));
AND2X1 exu_U21440(.A(byp_irf_rd_data_w2[44]), .B(exu_n16276), .Y(exu_n22408));
INVX1 exu_U21441(.A(exu_n22408), .Y(exu_n6212));
AND2X1 exu_U21442(.A(byp_irf_rd_data_w2[43]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22412));
INVX1 exu_U21443(.A(exu_n22412), .Y(exu_n6213));
AND2X1 exu_U21444(.A(byp_irf_rd_data_w2[42]), .B(exu_n16276), .Y(exu_n22416));
INVX1 exu_U21445(.A(exu_n22416), .Y(exu_n6214));
AND2X1 exu_U21446(.A(byp_irf_rd_data_w2[41]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22420));
INVX1 exu_U21447(.A(exu_n22420), .Y(exu_n6215));
AND2X1 exu_U21448(.A(byp_irf_rd_data_w2[40]), .B(exu_n16276), .Y(exu_n22424));
INVX1 exu_U21449(.A(exu_n22424), .Y(exu_n6216));
AND2X1 exu_U21450(.A(byp_irf_rd_data_w2[3]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22428));
INVX1 exu_U21451(.A(exu_n22428), .Y(exu_n6217));
AND2X1 exu_U21452(.A(byp_irf_rd_data_w2[39]), .B(exu_n16276), .Y(exu_n22432));
INVX1 exu_U21453(.A(exu_n22432), .Y(exu_n6218));
AND2X1 exu_U21454(.A(byp_irf_rd_data_w2[38]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22436));
INVX1 exu_U21455(.A(exu_n22436), .Y(exu_n6219));
AND2X1 exu_U21456(.A(byp_irf_rd_data_w2[37]), .B(exu_n16276), .Y(exu_n22440));
INVX1 exu_U21457(.A(exu_n22440), .Y(exu_n6220));
AND2X1 exu_U21458(.A(byp_irf_rd_data_w2[36]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22444));
INVX1 exu_U21459(.A(exu_n22444), .Y(exu_n6221));
AND2X1 exu_U21460(.A(byp_irf_rd_data_w2[35]), .B(exu_n16276), .Y(exu_n22448));
INVX1 exu_U21461(.A(exu_n22448), .Y(exu_n6222));
AND2X1 exu_U21462(.A(byp_irf_rd_data_w2[34]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22452));
INVX1 exu_U21463(.A(exu_n22452), .Y(exu_n6223));
AND2X1 exu_U21464(.A(byp_irf_rd_data_w2[33]), .B(exu_n16276), .Y(exu_n22456));
INVX1 exu_U21465(.A(exu_n22456), .Y(exu_n6224));
AND2X1 exu_U21466(.A(byp_irf_rd_data_w2[32]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22460));
INVX1 exu_U21467(.A(exu_n22460), .Y(exu_n6225));
AND2X1 exu_U21468(.A(byp_irf_rd_data_w2[31]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22464));
INVX1 exu_U21469(.A(exu_n22464), .Y(exu_n6226));
AND2X1 exu_U21470(.A(byp_irf_rd_data_w2[30]), .B(exu_n16276), .Y(exu_n22468));
INVX1 exu_U21471(.A(exu_n22468), .Y(exu_n6227));
AND2X1 exu_U21472(.A(byp_irf_rd_data_w2[2]), .B(exu_n16276), .Y(exu_n22472));
INVX1 exu_U21473(.A(exu_n22472), .Y(exu_n6228));
AND2X1 exu_U21474(.A(byp_irf_rd_data_w2[29]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22476));
INVX1 exu_U21475(.A(exu_n22476), .Y(exu_n6229));
AND2X1 exu_U21476(.A(byp_irf_rd_data_w2[28]), .B(exu_n16276), .Y(exu_n22480));
INVX1 exu_U21477(.A(exu_n22480), .Y(exu_n6230));
AND2X1 exu_U21478(.A(byp_irf_rd_data_w2[27]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22484));
INVX1 exu_U21479(.A(exu_n22484), .Y(exu_n6231));
AND2X1 exu_U21480(.A(byp_irf_rd_data_w2[26]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22488));
INVX1 exu_U21481(.A(exu_n22488), .Y(exu_n6232));
AND2X1 exu_U21482(.A(byp_irf_rd_data_w2[25]), .B(exu_n16276), .Y(exu_n22492));
INVX1 exu_U21483(.A(exu_n22492), .Y(exu_n6233));
AND2X1 exu_U21484(.A(byp_irf_rd_data_w2[24]), .B(exu_n16276), .Y(exu_n22496));
INVX1 exu_U21485(.A(exu_n22496), .Y(exu_n6234));
AND2X1 exu_U21486(.A(byp_irf_rd_data_w2[23]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22500));
INVX1 exu_U21487(.A(exu_n22500), .Y(exu_n6235));
AND2X1 exu_U21488(.A(byp_irf_rd_data_w2[22]), .B(exu_n16276), .Y(exu_n22504));
INVX1 exu_U21489(.A(exu_n22504), .Y(exu_n6236));
AND2X1 exu_U21490(.A(byp_irf_rd_data_w2[21]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22508));
INVX1 exu_U21491(.A(exu_n22508), .Y(exu_n6237));
AND2X1 exu_U21492(.A(byp_irf_rd_data_w2[20]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22512));
INVX1 exu_U21493(.A(exu_n22512), .Y(exu_n6238));
AND2X1 exu_U21494(.A(byp_irf_rd_data_w2[1]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22516));
INVX1 exu_U21495(.A(exu_n22516), .Y(exu_n6239));
AND2X1 exu_U21496(.A(byp_irf_rd_data_w2[19]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22520));
INVX1 exu_U21497(.A(exu_n22520), .Y(exu_n6240));
AND2X1 exu_U21498(.A(byp_irf_rd_data_w2[18]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22524));
INVX1 exu_U21499(.A(exu_n22524), .Y(exu_n6241));
AND2X1 exu_U21500(.A(byp_irf_rd_data_w2[17]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22528));
INVX1 exu_U21501(.A(exu_n22528), .Y(exu_n6242));
AND2X1 exu_U21502(.A(byp_irf_rd_data_w2[16]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22532));
INVX1 exu_U21503(.A(exu_n22532), .Y(exu_n6243));
AND2X1 exu_U21504(.A(byp_irf_rd_data_w2[15]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22536));
INVX1 exu_U21505(.A(exu_n22536), .Y(exu_n6244));
AND2X1 exu_U21506(.A(byp_irf_rd_data_w2[14]), .B(exu_n16276), .Y(exu_n22540));
INVX1 exu_U21507(.A(exu_n22540), .Y(exu_n6245));
AND2X1 exu_U21508(.A(byp_irf_rd_data_w2[13]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22544));
INVX1 exu_U21509(.A(exu_n22544), .Y(exu_n6246));
AND2X1 exu_U21510(.A(byp_irf_rd_data_w2[12]), .B(exu_n16276), .Y(exu_n22548));
INVX1 exu_U21511(.A(exu_n22548), .Y(exu_n6247));
AND2X1 exu_U21512(.A(byp_irf_rd_data_w2[11]), .B(exu_n16276), .Y(exu_n22552));
INVX1 exu_U21513(.A(exu_n22552), .Y(exu_n6248));
AND2X1 exu_U21514(.A(byp_irf_rd_data_w2[10]), .B(exu_n16276), .Y(exu_n22556));
INVX1 exu_U21515(.A(exu_n22556), .Y(exu_n6249));
AND2X1 exu_U21516(.A(byp_irf_rd_data_w2[0]), .B(ecl_byp_rs3_longmux_sel_w2), .Y(exu_n22560));
INVX1 exu_U21517(.A(exu_n22560), .Y(exu_n6250));
AND2X1 exu_U21518(.A(ecl_writeback_n129), .B(bypass_restore_rd_data[9]), .Y(exu_n22562));
INVX1 exu_U21519(.A(exu_n22562), .Y(exu_n6251));
AND2X1 exu_U21520(.A(exu_n15398), .B(exu_n10242), .Y(exu_n22564));
INVX1 exu_U21521(.A(exu_n22564), .Y(exu_n6252));
AND2X1 exu_U21522(.A(bypass_restore_rd_data[8]), .B(exu_n15988), .Y(exu_n22566));
INVX1 exu_U21523(.A(exu_n22566), .Y(exu_n6253));
AND2X1 exu_U21524(.A(exu_n11362), .B(exu_n15398), .Y(exu_n22568));
INVX1 exu_U21525(.A(exu_n22568), .Y(exu_n6254));
AND2X1 exu_U21526(.A(bypass_restore_rd_data[7]), .B(exu_n15988), .Y(exu_n22570));
INVX1 exu_U21527(.A(exu_n22570), .Y(exu_n6255));
AND2X1 exu_U21528(.A(exu_n11364), .B(exu_n15398), .Y(exu_n22572));
INVX1 exu_U21529(.A(exu_n22572), .Y(exu_n6256));
AND2X1 exu_U21530(.A(bypass_restore_rd_data[6]), .B(exu_n15988), .Y(exu_n22574));
INVX1 exu_U21531(.A(exu_n22574), .Y(exu_n6257));
AND2X1 exu_U21532(.A(exu_n11366), .B(exu_n15398), .Y(exu_n22576));
INVX1 exu_U21533(.A(exu_n22576), .Y(exu_n6258));
AND2X1 exu_U21534(.A(bypass_restore_rd_data[63]), .B(exu_n15988), .Y(exu_n22578));
INVX1 exu_U21535(.A(exu_n22578), .Y(exu_n6259));
AND2X1 exu_U21536(.A(exu_n11368), .B(exu_n15398), .Y(exu_n22580));
INVX1 exu_U21537(.A(exu_n22580), .Y(exu_n6260));
AND2X1 exu_U21538(.A(bypass_restore_rd_data[62]), .B(exu_n15988), .Y(exu_n22582));
INVX1 exu_U21539(.A(exu_n22582), .Y(exu_n6261));
AND2X1 exu_U21540(.A(exu_n11370), .B(exu_n15398), .Y(exu_n22584));
INVX1 exu_U21541(.A(exu_n22584), .Y(exu_n6262));
AND2X1 exu_U21542(.A(bypass_restore_rd_data[61]), .B(exu_n15988), .Y(exu_n22586));
INVX1 exu_U21543(.A(exu_n22586), .Y(exu_n6263));
AND2X1 exu_U21544(.A(exu_n11372), .B(exu_n15398), .Y(exu_n22588));
INVX1 exu_U21545(.A(exu_n22588), .Y(exu_n6264));
AND2X1 exu_U21546(.A(bypass_restore_rd_data[60]), .B(exu_n15988), .Y(exu_n22590));
INVX1 exu_U21547(.A(exu_n22590), .Y(exu_n6265));
AND2X1 exu_U21548(.A(exu_n11374), .B(exu_n15398), .Y(exu_n22592));
INVX1 exu_U21549(.A(exu_n22592), .Y(exu_n6266));
AND2X1 exu_U21550(.A(bypass_restore_rd_data[5]), .B(exu_n15988), .Y(exu_n22594));
INVX1 exu_U21551(.A(exu_n22594), .Y(exu_n6267));
AND2X1 exu_U21552(.A(exu_n11376), .B(exu_n15398), .Y(exu_n22596));
INVX1 exu_U21553(.A(exu_n22596), .Y(exu_n6268));
AND2X1 exu_U21554(.A(bypass_restore_rd_data[59]), .B(exu_n15988), .Y(exu_n22598));
INVX1 exu_U21555(.A(exu_n22598), .Y(exu_n6269));
AND2X1 exu_U21556(.A(exu_n11378), .B(exu_n15398), .Y(exu_n22600));
INVX1 exu_U21557(.A(exu_n22600), .Y(exu_n6270));
AND2X1 exu_U21558(.A(bypass_restore_rd_data[58]), .B(exu_n15988), .Y(exu_n22602));
INVX1 exu_U21559(.A(exu_n22602), .Y(exu_n6271));
AND2X1 exu_U21560(.A(exu_n11380), .B(exu_n15398), .Y(exu_n22604));
INVX1 exu_U21561(.A(exu_n22604), .Y(exu_n6272));
AND2X1 exu_U21562(.A(bypass_restore_rd_data[57]), .B(exu_n15988), .Y(exu_n22606));
INVX1 exu_U21563(.A(exu_n22606), .Y(exu_n6273));
AND2X1 exu_U21564(.A(exu_n11382), .B(exu_n15398), .Y(exu_n22608));
INVX1 exu_U21565(.A(exu_n22608), .Y(exu_n6274));
AND2X1 exu_U21566(.A(bypass_restore_rd_data[56]), .B(exu_n15988), .Y(exu_n22610));
INVX1 exu_U21567(.A(exu_n22610), .Y(exu_n6275));
AND2X1 exu_U21568(.A(exu_n11384), .B(exu_n15398), .Y(exu_n22612));
INVX1 exu_U21569(.A(exu_n22612), .Y(exu_n6276));
AND2X1 exu_U21570(.A(bypass_restore_rd_data[55]), .B(exu_n15988), .Y(exu_n22614));
INVX1 exu_U21571(.A(exu_n22614), .Y(exu_n6277));
AND2X1 exu_U21572(.A(exu_n11386), .B(exu_n15398), .Y(exu_n22616));
INVX1 exu_U21573(.A(exu_n22616), .Y(exu_n6278));
AND2X1 exu_U21574(.A(bypass_restore_rd_data[54]), .B(ecl_writeback_n129), .Y(exu_n22618));
INVX1 exu_U21575(.A(exu_n22618), .Y(exu_n6279));
AND2X1 exu_U21576(.A(exu_n11388), .B(exu_n15398), .Y(exu_n22620));
INVX1 exu_U21577(.A(exu_n22620), .Y(exu_n6280));
AND2X1 exu_U21578(.A(bypass_restore_rd_data[53]), .B(exu_n15988), .Y(exu_n22622));
INVX1 exu_U21579(.A(exu_n22622), .Y(exu_n6281));
AND2X1 exu_U21580(.A(exu_n11390), .B(exu_n15398), .Y(exu_n22624));
INVX1 exu_U21581(.A(exu_n22624), .Y(exu_n6282));
AND2X1 exu_U21582(.A(bypass_restore_rd_data[52]), .B(ecl_writeback_n129), .Y(exu_n22626));
INVX1 exu_U21583(.A(exu_n22626), .Y(exu_n6283));
AND2X1 exu_U21584(.A(exu_n11392), .B(exu_n15398), .Y(exu_n22628));
INVX1 exu_U21585(.A(exu_n22628), .Y(exu_n6284));
AND2X1 exu_U21586(.A(bypass_restore_rd_data[51]), .B(exu_n15988), .Y(exu_n22630));
INVX1 exu_U21587(.A(exu_n22630), .Y(exu_n6285));
AND2X1 exu_U21588(.A(exu_n11394), .B(exu_n15398), .Y(exu_n22632));
INVX1 exu_U21589(.A(exu_n22632), .Y(exu_n6286));
AND2X1 exu_U21590(.A(bypass_restore_rd_data[50]), .B(ecl_writeback_n129), .Y(exu_n22634));
INVX1 exu_U21591(.A(exu_n22634), .Y(exu_n6287));
AND2X1 exu_U21592(.A(exu_n11396), .B(exu_n15398), .Y(exu_n22636));
INVX1 exu_U21593(.A(exu_n22636), .Y(exu_n6288));
AND2X1 exu_U21594(.A(bypass_restore_rd_data[4]), .B(exu_n15988), .Y(exu_n22638));
INVX1 exu_U21595(.A(exu_n22638), .Y(exu_n6289));
AND2X1 exu_U21596(.A(exu_n11398), .B(exu_n15398), .Y(exu_n22640));
INVX1 exu_U21597(.A(exu_n22640), .Y(exu_n6290));
AND2X1 exu_U21598(.A(bypass_restore_rd_data[49]), .B(ecl_writeback_n129), .Y(exu_n22642));
INVX1 exu_U21599(.A(exu_n22642), .Y(exu_n6291));
AND2X1 exu_U21600(.A(exu_n11400), .B(exu_n15398), .Y(exu_n22644));
INVX1 exu_U21601(.A(exu_n22644), .Y(exu_n6292));
AND2X1 exu_U21602(.A(bypass_restore_rd_data[48]), .B(exu_n15988), .Y(exu_n22646));
INVX1 exu_U21603(.A(exu_n22646), .Y(exu_n6293));
AND2X1 exu_U21604(.A(exu_n11402), .B(exu_n15398), .Y(exu_n22648));
INVX1 exu_U21605(.A(exu_n22648), .Y(exu_n6294));
AND2X1 exu_U21606(.A(bypass_restore_rd_data[47]), .B(ecl_writeback_n129), .Y(exu_n22650));
INVX1 exu_U21607(.A(exu_n22650), .Y(exu_n6295));
AND2X1 exu_U21608(.A(exu_n11404), .B(exu_n15398), .Y(exu_n22652));
INVX1 exu_U21609(.A(exu_n22652), .Y(exu_n6296));
AND2X1 exu_U21610(.A(bypass_restore_rd_data[46]), .B(exu_n15988), .Y(exu_n22654));
INVX1 exu_U21611(.A(exu_n22654), .Y(exu_n6297));
AND2X1 exu_U21612(.A(exu_n11406), .B(exu_n15398), .Y(exu_n22656));
INVX1 exu_U21613(.A(exu_n22656), .Y(exu_n6298));
AND2X1 exu_U21614(.A(bypass_restore_rd_data[45]), .B(ecl_writeback_n129), .Y(exu_n22658));
INVX1 exu_U21615(.A(exu_n22658), .Y(exu_n6299));
AND2X1 exu_U21616(.A(exu_n11408), .B(exu_n15398), .Y(exu_n22660));
INVX1 exu_U21617(.A(exu_n22660), .Y(exu_n6300));
AND2X1 exu_U21618(.A(bypass_restore_rd_data[44]), .B(exu_n15988), .Y(exu_n22662));
INVX1 exu_U21619(.A(exu_n22662), .Y(exu_n6301));
AND2X1 exu_U21620(.A(exu_n11410), .B(exu_n15398), .Y(exu_n22664));
INVX1 exu_U21621(.A(exu_n22664), .Y(exu_n6302));
AND2X1 exu_U21622(.A(bypass_restore_rd_data[43]), .B(ecl_writeback_n129), .Y(exu_n22666));
INVX1 exu_U21623(.A(exu_n22666), .Y(exu_n6303));
AND2X1 exu_U21624(.A(exu_n11412), .B(exu_n15398), .Y(exu_n22668));
INVX1 exu_U21625(.A(exu_n22668), .Y(exu_n6304));
AND2X1 exu_U21626(.A(bypass_restore_rd_data[42]), .B(exu_n15988), .Y(exu_n22670));
INVX1 exu_U21627(.A(exu_n22670), .Y(exu_n6305));
AND2X1 exu_U21628(.A(exu_n11414), .B(exu_n15398), .Y(exu_n22672));
INVX1 exu_U21629(.A(exu_n22672), .Y(exu_n6306));
AND2X1 exu_U21630(.A(bypass_restore_rd_data[41]), .B(ecl_writeback_n129), .Y(exu_n22674));
INVX1 exu_U21631(.A(exu_n22674), .Y(exu_n6307));
AND2X1 exu_U21632(.A(exu_n11416), .B(exu_n15398), .Y(exu_n22676));
INVX1 exu_U21633(.A(exu_n22676), .Y(exu_n6308));
AND2X1 exu_U21634(.A(bypass_restore_rd_data[40]), .B(ecl_writeback_n129), .Y(exu_n22678));
INVX1 exu_U21635(.A(exu_n22678), .Y(exu_n6309));
AND2X1 exu_U21636(.A(exu_n11418), .B(exu_n15398), .Y(exu_n22680));
INVX1 exu_U21637(.A(exu_n22680), .Y(exu_n6310));
AND2X1 exu_U21638(.A(bypass_restore_rd_data[3]), .B(ecl_writeback_n129), .Y(exu_n22682));
INVX1 exu_U21639(.A(exu_n22682), .Y(exu_n6311));
AND2X1 exu_U21640(.A(exu_n11420), .B(exu_n15398), .Y(exu_n22684));
INVX1 exu_U21641(.A(exu_n22684), .Y(exu_n6312));
AND2X1 exu_U21642(.A(bypass_restore_rd_data[39]), .B(exu_n15988), .Y(exu_n22686));
INVX1 exu_U21643(.A(exu_n22686), .Y(exu_n6313));
AND2X1 exu_U21644(.A(exu_n11422), .B(exu_n15398), .Y(exu_n22688));
INVX1 exu_U21645(.A(exu_n22688), .Y(exu_n6314));
AND2X1 exu_U21646(.A(bypass_restore_rd_data[38]), .B(ecl_writeback_n129), .Y(exu_n22690));
INVX1 exu_U21647(.A(exu_n22690), .Y(exu_n6315));
AND2X1 exu_U21648(.A(exu_n11424), .B(exu_n15398), .Y(exu_n22692));
INVX1 exu_U21649(.A(exu_n22692), .Y(exu_n6316));
AND2X1 exu_U21650(.A(bypass_restore_rd_data[37]), .B(exu_n15988), .Y(exu_n22694));
INVX1 exu_U21651(.A(exu_n22694), .Y(exu_n6317));
AND2X1 exu_U21652(.A(exu_n11426), .B(exu_n15398), .Y(exu_n22696));
INVX1 exu_U21653(.A(exu_n22696), .Y(exu_n6318));
AND2X1 exu_U21654(.A(bypass_restore_rd_data[36]), .B(ecl_writeback_n129), .Y(exu_n22698));
INVX1 exu_U21655(.A(exu_n22698), .Y(exu_n6319));
AND2X1 exu_U21656(.A(exu_n11428), .B(exu_n15398), .Y(exu_n22700));
INVX1 exu_U21657(.A(exu_n22700), .Y(exu_n6320));
AND2X1 exu_U21658(.A(bypass_restore_rd_data[35]), .B(ecl_writeback_n129), .Y(exu_n22702));
INVX1 exu_U21659(.A(exu_n22702), .Y(exu_n6321));
AND2X1 exu_U21660(.A(exu_n11430), .B(exu_n15398), .Y(exu_n22704));
INVX1 exu_U21661(.A(exu_n22704), .Y(exu_n6322));
AND2X1 exu_U21662(.A(bypass_restore_rd_data[34]), .B(ecl_writeback_n129), .Y(exu_n22706));
INVX1 exu_U21663(.A(exu_n22706), .Y(exu_n6323));
AND2X1 exu_U21664(.A(exu_n11432), .B(exu_n15398), .Y(exu_n22708));
INVX1 exu_U21665(.A(exu_n22708), .Y(exu_n6324));
AND2X1 exu_U21666(.A(bypass_restore_rd_data[33]), .B(exu_n15988), .Y(exu_n22710));
INVX1 exu_U21667(.A(exu_n22710), .Y(exu_n6325));
AND2X1 exu_U21668(.A(exu_n11434), .B(exu_n15398), .Y(exu_n22712));
INVX1 exu_U21669(.A(exu_n22712), .Y(exu_n6326));
AND2X1 exu_U21670(.A(bypass_restore_rd_data[32]), .B(exu_n15988), .Y(exu_n22714));
INVX1 exu_U21671(.A(exu_n22714), .Y(exu_n6327));
AND2X1 exu_U21672(.A(exu_n11436), .B(exu_n15398), .Y(exu_n22716));
INVX1 exu_U21673(.A(exu_n22716), .Y(exu_n6328));
AND2X1 exu_U21674(.A(bypass_restore_rd_data[31]), .B(exu_n15988), .Y(exu_n22718));
INVX1 exu_U21675(.A(exu_n22718), .Y(exu_n6329));
AND2X1 exu_U21676(.A(exu_n11438), .B(exu_n15398), .Y(exu_n22720));
INVX1 exu_U21677(.A(exu_n22720), .Y(exu_n6330));
AND2X1 exu_U21678(.A(bypass_restore_rd_data[30]), .B(exu_n15988), .Y(exu_n22722));
INVX1 exu_U21679(.A(exu_n22722), .Y(exu_n6331));
AND2X1 exu_U21680(.A(exu_n11440), .B(exu_n15398), .Y(exu_n22724));
INVX1 exu_U21681(.A(exu_n22724), .Y(exu_n6332));
AND2X1 exu_U21682(.A(bypass_restore_rd_data[2]), .B(ecl_writeback_n129), .Y(exu_n22726));
INVX1 exu_U21683(.A(exu_n22726), .Y(exu_n6333));
AND2X1 exu_U21684(.A(exu_n11442), .B(exu_n15398), .Y(exu_n22728));
INVX1 exu_U21685(.A(exu_n22728), .Y(exu_n6334));
AND2X1 exu_U21686(.A(bypass_restore_rd_data[29]), .B(exu_n15988), .Y(exu_n22730));
INVX1 exu_U21687(.A(exu_n22730), .Y(exu_n6335));
AND2X1 exu_U21688(.A(exu_n11444), .B(exu_n15398), .Y(exu_n22732));
INVX1 exu_U21689(.A(exu_n22732), .Y(exu_n6336));
AND2X1 exu_U21690(.A(bypass_restore_rd_data[28]), .B(exu_n15988), .Y(exu_n22734));
INVX1 exu_U21691(.A(exu_n22734), .Y(exu_n6337));
AND2X1 exu_U21692(.A(exu_n11446), .B(exu_n15398), .Y(exu_n22736));
INVX1 exu_U21693(.A(exu_n22736), .Y(exu_n6338));
AND2X1 exu_U21694(.A(bypass_restore_rd_data[27]), .B(ecl_writeback_n129), .Y(exu_n22738));
INVX1 exu_U21695(.A(exu_n22738), .Y(exu_n6339));
AND2X1 exu_U21696(.A(exu_n11448), .B(exu_n15398), .Y(exu_n22740));
INVX1 exu_U21697(.A(exu_n22740), .Y(exu_n6340));
AND2X1 exu_U21698(.A(bypass_restore_rd_data[26]), .B(ecl_writeback_n129), .Y(exu_n22742));
INVX1 exu_U21699(.A(exu_n22742), .Y(exu_n6341));
AND2X1 exu_U21700(.A(exu_n11450), .B(exu_n15398), .Y(exu_n22744));
INVX1 exu_U21701(.A(exu_n22744), .Y(exu_n6342));
AND2X1 exu_U21702(.A(bypass_restore_rd_data[25]), .B(ecl_writeback_n129), .Y(exu_n22746));
INVX1 exu_U21703(.A(exu_n22746), .Y(exu_n6343));
AND2X1 exu_U21704(.A(exu_n11452), .B(exu_n15398), .Y(exu_n22748));
INVX1 exu_U21705(.A(exu_n22748), .Y(exu_n6344));
AND2X1 exu_U21706(.A(bypass_restore_rd_data[24]), .B(exu_n15988), .Y(exu_n22750));
INVX1 exu_U21707(.A(exu_n22750), .Y(exu_n6345));
AND2X1 exu_U21708(.A(exu_n11454), .B(exu_n15398), .Y(exu_n22752));
INVX1 exu_U21709(.A(exu_n22752), .Y(exu_n6346));
AND2X1 exu_U21710(.A(bypass_restore_rd_data[23]), .B(exu_n15988), .Y(exu_n22754));
INVX1 exu_U21711(.A(exu_n22754), .Y(exu_n6347));
AND2X1 exu_U21712(.A(exu_n11456), .B(exu_n15398), .Y(exu_n22756));
INVX1 exu_U21713(.A(exu_n22756), .Y(exu_n6348));
AND2X1 exu_U21714(.A(bypass_restore_rd_data[22]), .B(ecl_writeback_n129), .Y(exu_n22758));
INVX1 exu_U21715(.A(exu_n22758), .Y(exu_n6349));
AND2X1 exu_U21716(.A(exu_n11458), .B(exu_n15398), .Y(exu_n22760));
INVX1 exu_U21717(.A(exu_n22760), .Y(exu_n6350));
AND2X1 exu_U21718(.A(bypass_restore_rd_data[21]), .B(exu_n15988), .Y(exu_n22762));
INVX1 exu_U21719(.A(exu_n22762), .Y(exu_n6351));
AND2X1 exu_U21720(.A(exu_n11460), .B(exu_n15398), .Y(exu_n22764));
INVX1 exu_U21721(.A(exu_n22764), .Y(exu_n6352));
AND2X1 exu_U21722(.A(bypass_restore_rd_data[20]), .B(exu_n15988), .Y(exu_n22766));
INVX1 exu_U21723(.A(exu_n22766), .Y(exu_n6353));
AND2X1 exu_U21724(.A(exu_n11462), .B(exu_n15398), .Y(exu_n22768));
INVX1 exu_U21725(.A(exu_n22768), .Y(exu_n6354));
AND2X1 exu_U21726(.A(bypass_restore_rd_data[1]), .B(ecl_writeback_n129), .Y(exu_n22770));
INVX1 exu_U21727(.A(exu_n22770), .Y(exu_n6355));
AND2X1 exu_U21728(.A(exu_n11464), .B(exu_n15398), .Y(exu_n22772));
INVX1 exu_U21729(.A(exu_n22772), .Y(exu_n6356));
AND2X1 exu_U21730(.A(bypass_restore_rd_data[19]), .B(ecl_writeback_n129), .Y(exu_n22774));
INVX1 exu_U21731(.A(exu_n22774), .Y(exu_n6357));
AND2X1 exu_U21732(.A(exu_n11466), .B(exu_n15398), .Y(exu_n22776));
INVX1 exu_U21733(.A(exu_n22776), .Y(exu_n6358));
AND2X1 exu_U21734(.A(bypass_restore_rd_data[18]), .B(ecl_writeback_n129), .Y(exu_n22778));
INVX1 exu_U21735(.A(exu_n22778), .Y(exu_n6359));
AND2X1 exu_U21736(.A(exu_n11468), .B(exu_n15398), .Y(exu_n22780));
INVX1 exu_U21737(.A(exu_n22780), .Y(exu_n6360));
AND2X1 exu_U21738(.A(bypass_restore_rd_data[17]), .B(ecl_writeback_n129), .Y(exu_n22782));
INVX1 exu_U21739(.A(exu_n22782), .Y(exu_n6361));
AND2X1 exu_U21740(.A(exu_n11470), .B(exu_n15398), .Y(exu_n22784));
INVX1 exu_U21741(.A(exu_n22784), .Y(exu_n6362));
AND2X1 exu_U21742(.A(bypass_restore_rd_data[16]), .B(exu_n15988), .Y(exu_n22786));
INVX1 exu_U21743(.A(exu_n22786), .Y(exu_n6363));
AND2X1 exu_U21744(.A(exu_n11472), .B(exu_n15398), .Y(exu_n22788));
INVX1 exu_U21745(.A(exu_n22788), .Y(exu_n6364));
AND2X1 exu_U21746(.A(bypass_restore_rd_data[15]), .B(ecl_writeback_n129), .Y(exu_n22790));
INVX1 exu_U21747(.A(exu_n22790), .Y(exu_n6365));
AND2X1 exu_U21748(.A(exu_n11474), .B(exu_n15398), .Y(exu_n22792));
INVX1 exu_U21749(.A(exu_n22792), .Y(exu_n6366));
AND2X1 exu_U21750(.A(bypass_restore_rd_data[14]), .B(exu_n15988), .Y(exu_n22794));
INVX1 exu_U21751(.A(exu_n22794), .Y(exu_n6367));
AND2X1 exu_U21752(.A(exu_n11476), .B(exu_n15398), .Y(exu_n22796));
INVX1 exu_U21753(.A(exu_n22796), .Y(exu_n6368));
AND2X1 exu_U21754(.A(bypass_restore_rd_data[13]), .B(ecl_writeback_n129), .Y(exu_n22798));
INVX1 exu_U21755(.A(exu_n22798), .Y(exu_n6369));
AND2X1 exu_U21756(.A(exu_n11478), .B(exu_n15398), .Y(exu_n22800));
INVX1 exu_U21757(.A(exu_n22800), .Y(exu_n6370));
AND2X1 exu_U21758(.A(bypass_restore_rd_data[12]), .B(ecl_writeback_n129), .Y(exu_n22802));
INVX1 exu_U21759(.A(exu_n22802), .Y(exu_n6371));
AND2X1 exu_U21760(.A(exu_n11480), .B(exu_n15398), .Y(exu_n22804));
INVX1 exu_U21761(.A(exu_n22804), .Y(exu_n6372));
AND2X1 exu_U21762(.A(bypass_restore_rd_data[11]), .B(ecl_writeback_n129), .Y(exu_n22806));
INVX1 exu_U21763(.A(exu_n22806), .Y(exu_n6373));
AND2X1 exu_U21764(.A(exu_n11482), .B(exu_n15398), .Y(exu_n22808));
INVX1 exu_U21765(.A(exu_n22808), .Y(exu_n6374));
AND2X1 exu_U21766(.A(bypass_restore_rd_data[10]), .B(ecl_writeback_n129), .Y(exu_n22810));
INVX1 exu_U21767(.A(exu_n22810), .Y(exu_n6375));
AND2X1 exu_U21768(.A(exu_n11484), .B(exu_n15398), .Y(exu_n22812));
INVX1 exu_U21769(.A(exu_n22812), .Y(exu_n6376));
AND2X1 exu_U21770(.A(bypass_restore_rd_data[0]), .B(ecl_writeback_n129), .Y(exu_n22814));
INVX1 exu_U21771(.A(exu_n22814), .Y(exu_n6377));
AND2X1 exu_U21772(.A(exu_n11486), .B(exu_n15398), .Y(exu_n22816));
INVX1 exu_U21773(.A(exu_n22816), .Y(exu_n6378));
AND2X1 exu_U21774(.A(exu_n15973), .B(ecc_exu_lsu_rs3_data_m[9]), .Y(exu_n22818));
INVX1 exu_U21775(.A(exu_n22818), .Y(exu_n6379));
AND2X1 exu_U21776(.A(exu_n15975), .B(ecc_byp_ecc_rcc_data_m[9]), .Y(exu_n22820));
INVX1 exu_U21777(.A(exu_n22820), .Y(exu_n6380));
AND2X1 exu_U21778(.A(ecc_exu_lsu_rs3_data_m[8]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22822));
INVX1 exu_U21779(.A(exu_n22822), .Y(exu_n6381));
AND2X1 exu_U21780(.A(ecc_byp_ecc_rcc_data_m[8]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22824));
INVX1 exu_U21781(.A(exu_n22824), .Y(exu_n6382));
AND2X1 exu_U21782(.A(ecc_exu_lsu_rs3_data_m[7]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22826));
INVX1 exu_U21783(.A(exu_n22826), .Y(exu_n6383));
AND2X1 exu_U21784(.A(ecc_byp_ecc_rcc_data_m[7]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22828));
INVX1 exu_U21785(.A(exu_n22828), .Y(exu_n6384));
AND2X1 exu_U21786(.A(ecc_exu_lsu_rs3_data_m[6]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22830));
INVX1 exu_U21787(.A(exu_n22830), .Y(exu_n6385));
AND2X1 exu_U21788(.A(ecc_byp_ecc_rcc_data_m[6]), .B(exu_n15975), .Y(exu_n22832));
INVX1 exu_U21789(.A(exu_n22832), .Y(exu_n6386));
AND2X1 exu_U21790(.A(ecc_exu_lsu_rs3_data_m[63]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22834));
INVX1 exu_U21791(.A(exu_n22834), .Y(exu_n6387));
AND2X1 exu_U21792(.A(ecc_byp_ecc_rcc_data_m[63]), .B(exu_n15975), .Y(exu_n22836));
INVX1 exu_U21793(.A(exu_n22836), .Y(exu_n6388));
AND2X1 exu_U21794(.A(ecc_exu_lsu_rs3_data_m[62]), .B(exu_n15973), .Y(exu_n22838));
INVX1 exu_U21795(.A(exu_n22838), .Y(exu_n6389));
AND2X1 exu_U21796(.A(ecc_byp_ecc_rcc_data_m[62]), .B(exu_n15975), .Y(exu_n22840));
INVX1 exu_U21797(.A(exu_n22840), .Y(exu_n6390));
AND2X1 exu_U21798(.A(ecc_exu_lsu_rs3_data_m[61]), .B(exu_n15973), .Y(exu_n22842));
INVX1 exu_U21799(.A(exu_n22842), .Y(exu_n6391));
AND2X1 exu_U21800(.A(ecc_byp_ecc_rcc_data_m[61]), .B(exu_n15975), .Y(exu_n22844));
INVX1 exu_U21801(.A(exu_n22844), .Y(exu_n6392));
AND2X1 exu_U21802(.A(ecc_exu_lsu_rs3_data_m[60]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22846));
INVX1 exu_U21803(.A(exu_n22846), .Y(exu_n6393));
AND2X1 exu_U21804(.A(ecc_byp_ecc_rcc_data_m[60]), .B(exu_n15975), .Y(exu_n22848));
INVX1 exu_U21805(.A(exu_n22848), .Y(exu_n6394));
AND2X1 exu_U21806(.A(ecc_exu_lsu_rs3_data_m[5]), .B(exu_n15973), .Y(exu_n22850));
INVX1 exu_U21807(.A(exu_n22850), .Y(exu_n6395));
AND2X1 exu_U21808(.A(ecc_byp_ecc_rcc_data_m[5]), .B(exu_n15975), .Y(exu_n22852));
INVX1 exu_U21809(.A(exu_n22852), .Y(exu_n6396));
AND2X1 exu_U21810(.A(ecc_exu_lsu_rs3_data_m[59]), .B(exu_n15973), .Y(exu_n22854));
INVX1 exu_U21811(.A(exu_n22854), .Y(exu_n6397));
AND2X1 exu_U21812(.A(ecc_byp_ecc_rcc_data_m[59]), .B(exu_n15975), .Y(exu_n22856));
INVX1 exu_U21813(.A(exu_n22856), .Y(exu_n6398));
AND2X1 exu_U21814(.A(ecc_exu_lsu_rs3_data_m[58]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22858));
INVX1 exu_U21815(.A(exu_n22858), .Y(exu_n6399));
AND2X1 exu_U21816(.A(ecc_byp_ecc_rcc_data_m[58]), .B(exu_n15975), .Y(exu_n22860));
INVX1 exu_U21817(.A(exu_n22860), .Y(exu_n6400));
AND2X1 exu_U21818(.A(ecc_exu_lsu_rs3_data_m[57]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22862));
INVX1 exu_U21819(.A(exu_n22862), .Y(exu_n6401));
AND2X1 exu_U21820(.A(ecc_byp_ecc_rcc_data_m[57]), .B(exu_n15975), .Y(exu_n22864));
INVX1 exu_U21821(.A(exu_n22864), .Y(exu_n6402));
AND2X1 exu_U21822(.A(ecc_exu_lsu_rs3_data_m[56]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22866));
INVX1 exu_U21823(.A(exu_n22866), .Y(exu_n6403));
AND2X1 exu_U21824(.A(ecc_byp_ecc_rcc_data_m[56]), .B(exu_n15975), .Y(exu_n22868));
INVX1 exu_U21825(.A(exu_n22868), .Y(exu_n6404));
AND2X1 exu_U21826(.A(ecc_exu_lsu_rs3_data_m[55]), .B(exu_n15973), .Y(exu_n22870));
INVX1 exu_U21827(.A(exu_n22870), .Y(exu_n6405));
AND2X1 exu_U21828(.A(ecc_byp_ecc_rcc_data_m[55]), .B(exu_n15975), .Y(exu_n22872));
INVX1 exu_U21829(.A(exu_n22872), .Y(exu_n6406));
AND2X1 exu_U21830(.A(ecc_exu_lsu_rs3_data_m[54]), .B(exu_n15973), .Y(exu_n22874));
INVX1 exu_U21831(.A(exu_n22874), .Y(exu_n6407));
AND2X1 exu_U21832(.A(ecc_byp_ecc_rcc_data_m[54]), .B(exu_n15975), .Y(exu_n22876));
INVX1 exu_U21833(.A(exu_n22876), .Y(exu_n6408));
AND2X1 exu_U21834(.A(ecc_exu_lsu_rs3_data_m[53]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22878));
INVX1 exu_U21835(.A(exu_n22878), .Y(exu_n6409));
AND2X1 exu_U21836(.A(ecc_byp_ecc_rcc_data_m[53]), .B(exu_n15975), .Y(exu_n22880));
INVX1 exu_U21837(.A(exu_n22880), .Y(exu_n6410));
AND2X1 exu_U21838(.A(ecc_exu_lsu_rs3_data_m[52]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22882));
INVX1 exu_U21839(.A(exu_n22882), .Y(exu_n6411));
AND2X1 exu_U21840(.A(ecc_byp_ecc_rcc_data_m[52]), .B(exu_n15975), .Y(exu_n22884));
INVX1 exu_U21841(.A(exu_n22884), .Y(exu_n6412));
AND2X1 exu_U21842(.A(ecc_exu_lsu_rs3_data_m[51]), .B(exu_n15973), .Y(exu_n22886));
INVX1 exu_U21843(.A(exu_n22886), .Y(exu_n6413));
AND2X1 exu_U21844(.A(ecc_byp_ecc_rcc_data_m[51]), .B(exu_n15975), .Y(exu_n22888));
INVX1 exu_U21845(.A(exu_n22888), .Y(exu_n6414));
AND2X1 exu_U21846(.A(ecc_exu_lsu_rs3_data_m[50]), .B(exu_n15973), .Y(exu_n22890));
INVX1 exu_U21847(.A(exu_n22890), .Y(exu_n6415));
AND2X1 exu_U21848(.A(ecc_byp_ecc_rcc_data_m[50]), .B(exu_n15975), .Y(exu_n22892));
INVX1 exu_U21849(.A(exu_n22892), .Y(exu_n6416));
AND2X1 exu_U21850(.A(ecc_exu_lsu_rs3_data_m[4]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22894));
INVX1 exu_U21851(.A(exu_n22894), .Y(exu_n6417));
AND2X1 exu_U21852(.A(ecc_byp_ecc_rcc_data_m[4]), .B(exu_n15975), .Y(exu_n22896));
INVX1 exu_U21853(.A(exu_n22896), .Y(exu_n6418));
AND2X1 exu_U21854(.A(ecc_exu_lsu_rs3_data_m[49]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22898));
INVX1 exu_U21855(.A(exu_n22898), .Y(exu_n6419));
AND2X1 exu_U21856(.A(ecc_byp_ecc_rcc_data_m[49]), .B(exu_n15975), .Y(exu_n22900));
INVX1 exu_U21857(.A(exu_n22900), .Y(exu_n6420));
AND2X1 exu_U21858(.A(ecc_exu_lsu_rs3_data_m[48]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22902));
INVX1 exu_U21859(.A(exu_n22902), .Y(exu_n6421));
AND2X1 exu_U21860(.A(ecc_byp_ecc_rcc_data_m[48]), .B(exu_n15975), .Y(exu_n22904));
INVX1 exu_U21861(.A(exu_n22904), .Y(exu_n6422));
AND2X1 exu_U21862(.A(ecc_exu_lsu_rs3_data_m[47]), .B(exu_n15973), .Y(exu_n22906));
INVX1 exu_U21863(.A(exu_n22906), .Y(exu_n6423));
AND2X1 exu_U21864(.A(ecc_byp_ecc_rcc_data_m[47]), .B(exu_n15975), .Y(exu_n22908));
INVX1 exu_U21865(.A(exu_n22908), .Y(exu_n6424));
AND2X1 exu_U21866(.A(ecc_exu_lsu_rs3_data_m[46]), .B(exu_n15973), .Y(exu_n22910));
INVX1 exu_U21867(.A(exu_n22910), .Y(exu_n6425));
AND2X1 exu_U21868(.A(ecc_byp_ecc_rcc_data_m[46]), .B(exu_n15975), .Y(exu_n22912));
INVX1 exu_U21869(.A(exu_n22912), .Y(exu_n6426));
AND2X1 exu_U21870(.A(ecc_exu_lsu_rs3_data_m[45]), .B(exu_n15973), .Y(exu_n22914));
INVX1 exu_U21871(.A(exu_n22914), .Y(exu_n6427));
AND2X1 exu_U21872(.A(ecc_byp_ecc_rcc_data_m[45]), .B(exu_n15975), .Y(exu_n22916));
INVX1 exu_U21873(.A(exu_n22916), .Y(exu_n6428));
AND2X1 exu_U21874(.A(ecc_exu_lsu_rs3_data_m[44]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22918));
INVX1 exu_U21875(.A(exu_n22918), .Y(exu_n6429));
AND2X1 exu_U21876(.A(ecc_byp_ecc_rcc_data_m[44]), .B(exu_n15975), .Y(exu_n22920));
INVX1 exu_U21877(.A(exu_n22920), .Y(exu_n6430));
AND2X1 exu_U21878(.A(ecc_exu_lsu_rs3_data_m[43]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22922));
INVX1 exu_U21879(.A(exu_n22922), .Y(exu_n6431));
AND2X1 exu_U21880(.A(ecc_byp_ecc_rcc_data_m[43]), .B(exu_n15975), .Y(exu_n22924));
INVX1 exu_U21881(.A(exu_n22924), .Y(exu_n6432));
AND2X1 exu_U21882(.A(ecc_exu_lsu_rs3_data_m[42]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22926));
INVX1 exu_U21883(.A(exu_n22926), .Y(exu_n6433));
AND2X1 exu_U21884(.A(ecc_byp_ecc_rcc_data_m[42]), .B(exu_n15975), .Y(exu_n22928));
INVX1 exu_U21885(.A(exu_n22928), .Y(exu_n6434));
AND2X1 exu_U21886(.A(ecc_exu_lsu_rs3_data_m[41]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22930));
INVX1 exu_U21887(.A(exu_n22930), .Y(exu_n6435));
AND2X1 exu_U21888(.A(ecc_byp_ecc_rcc_data_m[41]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22932));
INVX1 exu_U21889(.A(exu_n22932), .Y(exu_n6436));
AND2X1 exu_U21890(.A(ecc_exu_lsu_rs3_data_m[40]), .B(exu_n15973), .Y(exu_n22934));
INVX1 exu_U21891(.A(exu_n22934), .Y(exu_n6437));
AND2X1 exu_U21892(.A(ecc_byp_ecc_rcc_data_m[40]), .B(exu_n15975), .Y(exu_n22936));
INVX1 exu_U21893(.A(exu_n22936), .Y(exu_n6438));
AND2X1 exu_U21894(.A(ecc_exu_lsu_rs3_data_m[3]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22938));
INVX1 exu_U21895(.A(exu_n22938), .Y(exu_n6439));
AND2X1 exu_U21896(.A(ecc_byp_ecc_rcc_data_m[3]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22940));
INVX1 exu_U21897(.A(exu_n22940), .Y(exu_n6440));
AND2X1 exu_U21898(.A(ecc_exu_lsu_rs3_data_m[39]), .B(exu_n15973), .Y(exu_n22942));
INVX1 exu_U21899(.A(exu_n22942), .Y(exu_n6441));
AND2X1 exu_U21900(.A(ecc_byp_ecc_rcc_data_m[39]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22944));
INVX1 exu_U21901(.A(exu_n22944), .Y(exu_n6442));
AND2X1 exu_U21902(.A(ecc_exu_lsu_rs3_data_m[38]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22946));
INVX1 exu_U21903(.A(exu_n22946), .Y(exu_n6443));
AND2X1 exu_U21904(.A(ecc_byp_ecc_rcc_data_m[38]), .B(exu_n15975), .Y(exu_n22948));
INVX1 exu_U21905(.A(exu_n22948), .Y(exu_n6444));
AND2X1 exu_U21906(.A(ecc_exu_lsu_rs3_data_m[37]), .B(exu_n15973), .Y(exu_n22950));
INVX1 exu_U21907(.A(exu_n22950), .Y(exu_n6445));
AND2X1 exu_U21908(.A(ecc_byp_ecc_rcc_data_m[37]), .B(exu_n15975), .Y(exu_n22952));
INVX1 exu_U21909(.A(exu_n22952), .Y(exu_n6446));
AND2X1 exu_U21910(.A(ecc_exu_lsu_rs3_data_m[36]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22954));
INVX1 exu_U21911(.A(exu_n22954), .Y(exu_n6447));
AND2X1 exu_U21912(.A(ecc_byp_ecc_rcc_data_m[36]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22956));
INVX1 exu_U21913(.A(exu_n22956), .Y(exu_n6448));
AND2X1 exu_U21914(.A(ecc_exu_lsu_rs3_data_m[35]), .B(exu_n15973), .Y(exu_n22958));
INVX1 exu_U21915(.A(exu_n22958), .Y(exu_n6449));
AND2X1 exu_U21916(.A(ecc_byp_ecc_rcc_data_m[35]), .B(exu_n15975), .Y(exu_n22960));
INVX1 exu_U21917(.A(exu_n22960), .Y(exu_n6450));
AND2X1 exu_U21918(.A(ecc_exu_lsu_rs3_data_m[34]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22962));
INVX1 exu_U21919(.A(exu_n22962), .Y(exu_n6451));
AND2X1 exu_U21920(.A(ecc_byp_ecc_rcc_data_m[34]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22964));
INVX1 exu_U21921(.A(exu_n22964), .Y(exu_n6452));
AND2X1 exu_U21922(.A(ecc_exu_lsu_rs3_data_m[33]), .B(exu_n15973), .Y(exu_n22966));
INVX1 exu_U21923(.A(exu_n22966), .Y(exu_n6453));
AND2X1 exu_U21924(.A(ecc_byp_ecc_rcc_data_m[33]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22968));
INVX1 exu_U21925(.A(exu_n22968), .Y(exu_n6454));
AND2X1 exu_U21926(.A(ecc_exu_lsu_rs3_data_m[32]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22970));
INVX1 exu_U21927(.A(exu_n22970), .Y(exu_n6455));
AND2X1 exu_U21928(.A(ecc_byp_ecc_rcc_data_m[32]), .B(exu_n15975), .Y(exu_n22972));
INVX1 exu_U21929(.A(exu_n22972), .Y(exu_n6456));
AND2X1 exu_U21930(.A(ecc_exu_lsu_rs3_data_m[31]), .B(exu_n15973), .Y(exu_n22974));
INVX1 exu_U21931(.A(exu_n22974), .Y(exu_n6457));
AND2X1 exu_U21932(.A(ecc_byp_ecc_rcc_data_m[31]), .B(exu_n15975), .Y(exu_n22976));
INVX1 exu_U21933(.A(exu_n22976), .Y(exu_n6458));
AND2X1 exu_U21934(.A(ecc_exu_lsu_rs3_data_m[30]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n22978));
INVX1 exu_U21935(.A(exu_n22978), .Y(exu_n6459));
AND2X1 exu_U21936(.A(ecc_byp_ecc_rcc_data_m[30]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22980));
INVX1 exu_U21937(.A(exu_n22980), .Y(exu_n6460));
AND2X1 exu_U21938(.A(ecc_exu_lsu_rs3_data_m[2]), .B(exu_n15973), .Y(exu_n22982));
INVX1 exu_U21939(.A(exu_n22982), .Y(exu_n6461));
AND2X1 exu_U21940(.A(ecc_byp_ecc_rcc_data_m[2]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22984));
INVX1 exu_U21941(.A(exu_n22984), .Y(exu_n6462));
AND2X1 exu_U21942(.A(ecc_exu_lsu_rs3_data_m[29]), .B(exu_n15973), .Y(exu_n22986));
INVX1 exu_U21943(.A(exu_n22986), .Y(exu_n6463));
AND2X1 exu_U21944(.A(ecc_byp_ecc_rcc_data_m[29]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22988));
INVX1 exu_U21945(.A(exu_n22988), .Y(exu_n6464));
AND2X1 exu_U21946(.A(ecc_exu_lsu_rs3_data_m[28]), .B(exu_n15973), .Y(exu_n22990));
INVX1 exu_U21947(.A(exu_n22990), .Y(exu_n6465));
AND2X1 exu_U21948(.A(ecc_byp_ecc_rcc_data_m[28]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n22992));
INVX1 exu_U21949(.A(exu_n22992), .Y(exu_n6466));
AND2X1 exu_U21950(.A(ecc_exu_lsu_rs3_data_m[27]), .B(exu_n15973), .Y(exu_n22994));
INVX1 exu_U21951(.A(exu_n22994), .Y(exu_n6467));
AND2X1 exu_U21952(.A(ecc_byp_ecc_rcc_data_m[27]), .B(exu_n15975), .Y(exu_n22996));
INVX1 exu_U21953(.A(exu_n22996), .Y(exu_n6468));
AND2X1 exu_U21954(.A(ecc_exu_lsu_rs3_data_m[26]), .B(exu_n15973), .Y(exu_n22998));
INVX1 exu_U21955(.A(exu_n22998), .Y(exu_n6469));
AND2X1 exu_U21956(.A(ecc_byp_ecc_rcc_data_m[26]), .B(exu_n15975), .Y(exu_n23000));
INVX1 exu_U21957(.A(exu_n23000), .Y(exu_n6470));
AND2X1 exu_U21958(.A(ecc_exu_lsu_rs3_data_m[25]), .B(exu_n15973), .Y(exu_n23002));
INVX1 exu_U21959(.A(exu_n23002), .Y(exu_n6471));
AND2X1 exu_U21960(.A(ecc_byp_ecc_rcc_data_m[25]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n23004));
INVX1 exu_U21961(.A(exu_n23004), .Y(exu_n6472));
AND2X1 exu_U21962(.A(ecc_exu_lsu_rs3_data_m[24]), .B(exu_n15973), .Y(exu_n23006));
INVX1 exu_U21963(.A(exu_n23006), .Y(exu_n6473));
AND2X1 exu_U21964(.A(ecc_byp_ecc_rcc_data_m[24]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n23008));
INVX1 exu_U21965(.A(exu_n23008), .Y(exu_n6474));
AND2X1 exu_U21966(.A(ecc_exu_lsu_rs3_data_m[23]), .B(exu_n15973), .Y(exu_n23010));
INVX1 exu_U21967(.A(exu_n23010), .Y(exu_n6475));
AND2X1 exu_U21968(.A(ecc_byp_ecc_rcc_data_m[23]), .B(exu_n15975), .Y(exu_n23012));
INVX1 exu_U21969(.A(exu_n23012), .Y(exu_n6476));
AND2X1 exu_U21970(.A(ecc_exu_lsu_rs3_data_m[22]), .B(exu_n15973), .Y(exu_n23014));
INVX1 exu_U21971(.A(exu_n23014), .Y(exu_n6477));
AND2X1 exu_U21972(.A(ecc_byp_ecc_rcc_data_m[22]), .B(exu_n15975), .Y(exu_n23016));
INVX1 exu_U21973(.A(exu_n23016), .Y(exu_n6478));
AND2X1 exu_U21974(.A(ecc_exu_lsu_rs3_data_m[21]), .B(exu_n15973), .Y(exu_n23018));
INVX1 exu_U21975(.A(exu_n23018), .Y(exu_n6479));
AND2X1 exu_U21976(.A(ecc_byp_ecc_rcc_data_m[21]), .B(exu_n15975), .Y(exu_n23020));
INVX1 exu_U21977(.A(exu_n23020), .Y(exu_n6480));
AND2X1 exu_U21978(.A(ecc_exu_lsu_rs3_data_m[20]), .B(exu_n15973), .Y(exu_n23022));
INVX1 exu_U21979(.A(exu_n23022), .Y(exu_n6481));
AND2X1 exu_U21980(.A(ecc_byp_ecc_rcc_data_m[20]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n23024));
INVX1 exu_U21981(.A(exu_n23024), .Y(exu_n6482));
AND2X1 exu_U21982(.A(ecc_exu_lsu_rs3_data_m[1]), .B(exu_n15973), .Y(exu_n23026));
INVX1 exu_U21983(.A(exu_n23026), .Y(exu_n6483));
AND2X1 exu_U21984(.A(ecc_byp_ecc_rcc_data_m[1]), .B(exu_n15975), .Y(exu_n23028));
INVX1 exu_U21985(.A(exu_n23028), .Y(exu_n6484));
AND2X1 exu_U21986(.A(ecc_exu_lsu_rs3_data_m[19]), .B(exu_n15973), .Y(exu_n23030));
INVX1 exu_U21987(.A(exu_n23030), .Y(exu_n6485));
AND2X1 exu_U21988(.A(ecc_byp_ecc_rcc_data_m[19]), .B(exu_n15975), .Y(exu_n23032));
INVX1 exu_U21989(.A(exu_n23032), .Y(exu_n6486));
AND2X1 exu_U21990(.A(ecc_exu_lsu_rs3_data_m[18]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n23034));
INVX1 exu_U21991(.A(exu_n23034), .Y(exu_n6487));
AND2X1 exu_U21992(.A(ecc_byp_ecc_rcc_data_m[18]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n23036));
INVX1 exu_U21993(.A(exu_n23036), .Y(exu_n6488));
AND2X1 exu_U21994(.A(ecc_exu_lsu_rs3_data_m[17]), .B(exu_n15973), .Y(exu_n23038));
INVX1 exu_U21995(.A(exu_n23038), .Y(exu_n6489));
AND2X1 exu_U21996(.A(ecc_byp_ecc_rcc_data_m[17]), .B(exu_n15975), .Y(exu_n23040));
INVX1 exu_U21997(.A(exu_n23040), .Y(exu_n6490));
AND2X1 exu_U21998(.A(ecc_exu_lsu_rs3_data_m[16]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n23042));
INVX1 exu_U21999(.A(exu_n23042), .Y(exu_n6491));
AND2X1 exu_U22000(.A(ecc_byp_ecc_rcc_data_m[16]), .B(exu_n15975), .Y(exu_n23044));
INVX1 exu_U22001(.A(exu_n23044), .Y(exu_n6492));
AND2X1 exu_U22002(.A(ecc_exu_lsu_rs3_data_m[15]), .B(exu_n15973), .Y(exu_n23046));
INVX1 exu_U22003(.A(exu_n23046), .Y(exu_n6493));
AND2X1 exu_U22004(.A(ecc_byp_ecc_rcc_data_m[15]), .B(exu_n15975), .Y(exu_n23048));
INVX1 exu_U22005(.A(exu_n23048), .Y(exu_n6494));
AND2X1 exu_U22006(.A(ecc_exu_lsu_rs3_data_m[14]), .B(exu_n15973), .Y(exu_n23050));
INVX1 exu_U22007(.A(exu_n23050), .Y(exu_n6495));
AND2X1 exu_U22008(.A(ecc_byp_ecc_rcc_data_m[14]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n23052));
INVX1 exu_U22009(.A(exu_n23052), .Y(exu_n6496));
AND2X1 exu_U22010(.A(ecc_exu_lsu_rs3_data_m[13]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n23054));
INVX1 exu_U22011(.A(exu_n23054), .Y(exu_n6497));
AND2X1 exu_U22012(.A(ecc_byp_ecc_rcc_data_m[13]), .B(exu_n15975), .Y(exu_n23056));
INVX1 exu_U22013(.A(exu_n23056), .Y(exu_n6498));
AND2X1 exu_U22014(.A(ecc_exu_lsu_rs3_data_m[12]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n23058));
INVX1 exu_U22015(.A(exu_n23058), .Y(exu_n6499));
AND2X1 exu_U22016(.A(ecc_byp_ecc_rcc_data_m[12]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n23060));
INVX1 exu_U22017(.A(exu_n23060), .Y(exu_n6500));
AND2X1 exu_U22018(.A(ecc_exu_lsu_rs3_data_m[11]), .B(exu_n15973), .Y(exu_n23062));
INVX1 exu_U22019(.A(exu_n23062), .Y(exu_n6501));
AND2X1 exu_U22020(.A(ecc_byp_ecc_rcc_data_m[11]), .B(exu_n15975), .Y(exu_n23064));
INVX1 exu_U22021(.A(exu_n23064), .Y(exu_n6502));
AND2X1 exu_U22022(.A(ecc_exu_lsu_rs3_data_m[10]), .B(ecl_ecc_sel_rs3_m_l), .Y(exu_n23066));
INVX1 exu_U22023(.A(exu_n23066), .Y(exu_n6503));
AND2X1 exu_U22024(.A(ecc_byp_ecc_rcc_data_m[10]), .B(ecl_ecc_sel_rs1_m_l), .Y(exu_n23068));
INVX1 exu_U22025(.A(exu_n23068), .Y(exu_n6504));
AND2X1 exu_U22026(.A(ecc_exu_lsu_rs3_data_m[0]), .B(exu_n15973), .Y(exu_n23070));
INVX1 exu_U22027(.A(exu_n23070), .Y(exu_n6505));
AND2X1 exu_U22028(.A(ecc_byp_ecc_rcc_data_m[0]), .B(exu_n15975), .Y(exu_n23072));
INVX1 exu_U22029(.A(exu_n23072), .Y(exu_n6506));
AND2X1 exu_U22030(.A(ecl_divcntl_N56), .B(div_x[9]), .Y(exu_n23074));
INVX1 exu_U22031(.A(exu_n23074), .Y(exu_n6507));
AND2X1 exu_U22032(.A(div_x[8]), .B(ecl_divcntl_N56), .Y(exu_n23076));
INVX1 exu_U22033(.A(exu_n23076), .Y(exu_n6508));
AND2X1 exu_U22034(.A(div_x[7]), .B(ecl_divcntl_N56), .Y(exu_n23078));
INVX1 exu_U22035(.A(exu_n23078), .Y(exu_n6509));
AND2X1 exu_U22036(.A(div_x[6]), .B(exu_n15978), .Y(exu_n23080));
INVX1 exu_U22037(.A(exu_n23080), .Y(exu_n6510));
AND2X1 exu_U22038(.A(div_ecl_x_msb), .B(ecl_divcntl_N56), .Y(exu_n23082));
INVX1 exu_U22039(.A(exu_n23082), .Y(exu_n6511));
AND2X1 exu_U22040(.A(div_x[62]), .B(exu_n15978), .Y(exu_n23084));
INVX1 exu_U22041(.A(exu_n23084), .Y(exu_n6512));
AND2X1 exu_U22042(.A(div_x[61]), .B(exu_n15978), .Y(exu_n23086));
INVX1 exu_U22043(.A(exu_n23086), .Y(exu_n6513));
AND2X1 exu_U22044(.A(div_x[60]), .B(ecl_divcntl_N56), .Y(exu_n23088));
INVX1 exu_U22045(.A(exu_n23088), .Y(exu_n6514));
AND2X1 exu_U22046(.A(div_x[5]), .B(ecl_divcntl_N56), .Y(exu_n23090));
INVX1 exu_U22047(.A(exu_n23090), .Y(exu_n6515));
AND2X1 exu_U22048(.A(div_x[59]), .B(exu_n15978), .Y(exu_n23092));
INVX1 exu_U22049(.A(exu_n23092), .Y(exu_n6516));
AND2X1 exu_U22050(.A(div_x[58]), .B(ecl_divcntl_N56), .Y(exu_n23094));
INVX1 exu_U22051(.A(exu_n23094), .Y(exu_n6517));
AND2X1 exu_U22052(.A(div_x[57]), .B(exu_n15978), .Y(exu_n23096));
INVX1 exu_U22053(.A(exu_n23096), .Y(exu_n6518));
AND2X1 exu_U22054(.A(div_x[56]), .B(exu_n15978), .Y(exu_n23098));
INVX1 exu_U22055(.A(exu_n23098), .Y(exu_n6519));
AND2X1 exu_U22056(.A(div_x[55]), .B(ecl_divcntl_N56), .Y(exu_n23100));
INVX1 exu_U22057(.A(exu_n23100), .Y(exu_n6520));
AND2X1 exu_U22058(.A(div_x[54]), .B(ecl_divcntl_N56), .Y(exu_n23102));
INVX1 exu_U22059(.A(exu_n23102), .Y(exu_n6521));
AND2X1 exu_U22060(.A(div_x[53]), .B(ecl_divcntl_N56), .Y(exu_n23104));
INVX1 exu_U22061(.A(exu_n23104), .Y(exu_n6522));
AND2X1 exu_U22062(.A(div_x[52]), .B(ecl_divcntl_N56), .Y(exu_n23106));
INVX1 exu_U22063(.A(exu_n23106), .Y(exu_n6523));
AND2X1 exu_U22064(.A(div_x[51]), .B(ecl_divcntl_N56), .Y(exu_n23108));
INVX1 exu_U22065(.A(exu_n23108), .Y(exu_n6524));
AND2X1 exu_U22066(.A(div_x[50]), .B(ecl_divcntl_N56), .Y(exu_n23110));
INVX1 exu_U22067(.A(exu_n23110), .Y(exu_n6525));
AND2X1 exu_U22068(.A(div_x[4]), .B(ecl_divcntl_N56), .Y(exu_n23112));
INVX1 exu_U22069(.A(exu_n23112), .Y(exu_n6526));
AND2X1 exu_U22070(.A(div_x[49]), .B(ecl_divcntl_N56), .Y(exu_n23114));
INVX1 exu_U22071(.A(exu_n23114), .Y(exu_n6527));
AND2X1 exu_U22072(.A(div_x[48]), .B(ecl_divcntl_N56), .Y(exu_n23116));
INVX1 exu_U22073(.A(exu_n23116), .Y(exu_n6528));
AND2X1 exu_U22074(.A(div_x[47]), .B(ecl_divcntl_N56), .Y(exu_n23118));
INVX1 exu_U22075(.A(exu_n23118), .Y(exu_n6529));
AND2X1 exu_U22076(.A(div_x[46]), .B(exu_n15978), .Y(exu_n23120));
INVX1 exu_U22077(.A(exu_n23120), .Y(exu_n6530));
AND2X1 exu_U22078(.A(div_x[45]), .B(ecl_divcntl_N56), .Y(exu_n23122));
INVX1 exu_U22079(.A(exu_n23122), .Y(exu_n6531));
AND2X1 exu_U22080(.A(div_x[44]), .B(exu_n15978), .Y(exu_n23124));
INVX1 exu_U22081(.A(exu_n23124), .Y(exu_n6532));
AND2X1 exu_U22082(.A(div_x[43]), .B(ecl_divcntl_N56), .Y(exu_n23126));
INVX1 exu_U22083(.A(exu_n23126), .Y(exu_n6533));
AND2X1 exu_U22084(.A(div_x[42]), .B(ecl_divcntl_N56), .Y(exu_n23128));
INVX1 exu_U22085(.A(exu_n23128), .Y(exu_n6534));
AND2X1 exu_U22086(.A(div_x[41]), .B(ecl_divcntl_N56), .Y(exu_n23130));
INVX1 exu_U22087(.A(exu_n23130), .Y(exu_n6535));
AND2X1 exu_U22088(.A(div_x[40]), .B(exu_n15978), .Y(exu_n23132));
INVX1 exu_U22089(.A(exu_n23132), .Y(exu_n6536));
AND2X1 exu_U22090(.A(div_x[3]), .B(exu_n15978), .Y(exu_n23134));
INVX1 exu_U22091(.A(exu_n23134), .Y(exu_n6537));
AND2X1 exu_U22092(.A(div_x[39]), .B(ecl_divcntl_N56), .Y(exu_n23136));
INVX1 exu_U22093(.A(exu_n23136), .Y(exu_n6538));
AND2X1 exu_U22094(.A(div_x[38]), .B(ecl_divcntl_N56), .Y(exu_n23138));
INVX1 exu_U22095(.A(exu_n23138), .Y(exu_n6539));
AND2X1 exu_U22096(.A(div_x[37]), .B(exu_n15978), .Y(exu_n23140));
INVX1 exu_U22097(.A(exu_n23140), .Y(exu_n6540));
AND2X1 exu_U22098(.A(div_x[36]), .B(ecl_divcntl_N56), .Y(exu_n23142));
INVX1 exu_U22099(.A(exu_n23142), .Y(exu_n6541));
AND2X1 exu_U22100(.A(div_x[35]), .B(ecl_divcntl_N56), .Y(exu_n23144));
INVX1 exu_U22101(.A(exu_n23144), .Y(exu_n6542));
AND2X1 exu_U22102(.A(div_x[34]), .B(exu_n15978), .Y(exu_n23146));
INVX1 exu_U22103(.A(exu_n23146), .Y(exu_n6543));
AND2X1 exu_U22104(.A(div_x[33]), .B(exu_n15978), .Y(exu_n23148));
INVX1 exu_U22105(.A(exu_n23148), .Y(exu_n6544));
AND2X1 exu_U22106(.A(div_x[32]), .B(exu_n15978), .Y(exu_n23150));
INVX1 exu_U22107(.A(exu_n23150), .Y(exu_n6545));
AND2X1 exu_U22108(.A(div_x[31]), .B(exu_n15978), .Y(exu_n23152));
INVX1 exu_U22109(.A(exu_n23152), .Y(exu_n6546));
AND2X1 exu_U22110(.A(div_x[30]), .B(exu_n15978), .Y(exu_n23154));
INVX1 exu_U22111(.A(exu_n23154), .Y(exu_n6547));
AND2X1 exu_U22112(.A(div_x[2]), .B(exu_n15978), .Y(exu_n23156));
INVX1 exu_U22113(.A(exu_n23156), .Y(exu_n6548));
AND2X1 exu_U22114(.A(div_x[29]), .B(exu_n15978), .Y(exu_n23158));
INVX1 exu_U22115(.A(exu_n23158), .Y(exu_n6549));
AND2X1 exu_U22116(.A(div_x[28]), .B(exu_n15978), .Y(exu_n23160));
INVX1 exu_U22117(.A(exu_n23160), .Y(exu_n6550));
AND2X1 exu_U22118(.A(div_x[27]), .B(exu_n15978), .Y(exu_n23162));
INVX1 exu_U22119(.A(exu_n23162), .Y(exu_n6551));
AND2X1 exu_U22120(.A(div_x[26]), .B(exu_n15978), .Y(exu_n23164));
INVX1 exu_U22121(.A(exu_n23164), .Y(exu_n6552));
AND2X1 exu_U22122(.A(div_x[25]), .B(exu_n15978), .Y(exu_n23166));
INVX1 exu_U22123(.A(exu_n23166), .Y(exu_n6553));
AND2X1 exu_U22124(.A(div_x[24]), .B(exu_n15978), .Y(exu_n23168));
INVX1 exu_U22125(.A(exu_n23168), .Y(exu_n6554));
AND2X1 exu_U22126(.A(div_x[23]), .B(exu_n15978), .Y(exu_n23170));
INVX1 exu_U22127(.A(exu_n23170), .Y(exu_n6555));
AND2X1 exu_U22128(.A(div_x[22]), .B(exu_n15978), .Y(exu_n23172));
INVX1 exu_U22129(.A(exu_n23172), .Y(exu_n6556));
AND2X1 exu_U22130(.A(div_x[21]), .B(exu_n15978), .Y(exu_n23174));
INVX1 exu_U22131(.A(exu_n23174), .Y(exu_n6557));
AND2X1 exu_U22132(.A(div_x[20]), .B(exu_n15978), .Y(exu_n23176));
INVX1 exu_U22133(.A(exu_n23176), .Y(exu_n6558));
AND2X1 exu_U22134(.A(div_x[1]), .B(ecl_divcntl_N56), .Y(exu_n23178));
INVX1 exu_U22135(.A(exu_n23178), .Y(exu_n6559));
AND2X1 exu_U22136(.A(div_x[19]), .B(exu_n15978), .Y(exu_n23180));
INVX1 exu_U22137(.A(exu_n23180), .Y(exu_n6560));
AND2X1 exu_U22138(.A(div_x[18]), .B(ecl_divcntl_N56), .Y(exu_n23182));
INVX1 exu_U22139(.A(exu_n23182), .Y(exu_n6561));
AND2X1 exu_U22140(.A(div_x[17]), .B(exu_n15978), .Y(exu_n23184));
INVX1 exu_U22141(.A(exu_n23184), .Y(exu_n6562));
AND2X1 exu_U22142(.A(div_x[16]), .B(ecl_divcntl_N56), .Y(exu_n23186));
INVX1 exu_U22143(.A(exu_n23186), .Y(exu_n6563));
AND2X1 exu_U22144(.A(div_x[15]), .B(exu_n15978), .Y(exu_n23188));
INVX1 exu_U22145(.A(exu_n23188), .Y(exu_n6564));
AND2X1 exu_U22146(.A(div_x[14]), .B(ecl_divcntl_N56), .Y(exu_n23190));
INVX1 exu_U22147(.A(exu_n23190), .Y(exu_n6565));
AND2X1 exu_U22148(.A(div_x[13]), .B(exu_n15978), .Y(exu_n23192));
INVX1 exu_U22149(.A(exu_n23192), .Y(exu_n6566));
AND2X1 exu_U22150(.A(div_x[12]), .B(ecl_divcntl_N56), .Y(exu_n23194));
INVX1 exu_U22151(.A(exu_n23194), .Y(exu_n6567));
AND2X1 exu_U22152(.A(div_x[11]), .B(exu_n15978), .Y(exu_n23196));
INVX1 exu_U22153(.A(exu_n23196), .Y(exu_n6568));
AND2X1 exu_U22154(.A(div_x[10]), .B(ecl_divcntl_N56), .Y(exu_n23198));
INVX1 exu_U22155(.A(exu_n23198), .Y(exu_n6569));
AND2X1 exu_U22156(.A(div_x[0]), .B(exu_n15978), .Y(exu_n23200));
INVX1 exu_U22157(.A(exu_n23200), .Y(exu_n6570));
AND2X1 exu_U22158(.A(ecl_byp_sel_ecc_m), .B(ecc_byp_ecc_result_m[9]), .Y(exu_n23204));
INVX1 exu_U22159(.A(exu_n23204), .Y(exu_n6571));
AND2X1 exu_U22160(.A(exu_n16274), .B(exu_n10587), .Y(exu_n23206));
INVX1 exu_U22161(.A(exu_n23206), .Y(exu_n6572));
AND2X1 exu_U22162(.A(ecc_byp_ecc_result_m[8]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23210));
INVX1 exu_U22163(.A(exu_n23210), .Y(exu_n6573));
AND2X1 exu_U22164(.A(exu_n11691), .B(exu_n16274), .Y(exu_n23212));
INVX1 exu_U22165(.A(exu_n23212), .Y(exu_n6574));
AND2X1 exu_U22166(.A(ecc_byp_ecc_result_m[7]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23216));
INVX1 exu_U22167(.A(exu_n23216), .Y(exu_n6575));
AND2X1 exu_U22168(.A(exu_n11692), .B(exu_n16274), .Y(exu_n23218));
INVX1 exu_U22169(.A(exu_n23218), .Y(exu_n6576));
AND2X1 exu_U22170(.A(ecc_byp_ecc_result_m[6]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23222));
INVX1 exu_U22171(.A(exu_n23222), .Y(exu_n6577));
AND2X1 exu_U22172(.A(exu_n11693), .B(exu_n16274), .Y(exu_n23224));
INVX1 exu_U22173(.A(exu_n23224), .Y(exu_n6578));
AND2X1 exu_U22174(.A(ecc_byp_ecc_result_m[63]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23228));
INVX1 exu_U22175(.A(exu_n23228), .Y(exu_n6579));
AND2X1 exu_U22176(.A(exu_n11694), .B(exu_n16274), .Y(exu_n23230));
INVX1 exu_U22177(.A(exu_n23230), .Y(exu_n6580));
AND2X1 exu_U22178(.A(ecc_byp_ecc_result_m[62]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23234));
INVX1 exu_U22179(.A(exu_n23234), .Y(exu_n6581));
AND2X1 exu_U22180(.A(exu_n11695), .B(exu_n16274), .Y(exu_n23236));
INVX1 exu_U22181(.A(exu_n23236), .Y(exu_n6582));
AND2X1 exu_U22182(.A(ecc_byp_ecc_result_m[61]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23240));
INVX1 exu_U22183(.A(exu_n23240), .Y(exu_n6583));
AND2X1 exu_U22184(.A(exu_n11696), .B(exu_n16274), .Y(exu_n23242));
INVX1 exu_U22185(.A(exu_n23242), .Y(exu_n6584));
AND2X1 exu_U22186(.A(ecc_byp_ecc_result_m[60]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23246));
INVX1 exu_U22187(.A(exu_n23246), .Y(exu_n6585));
AND2X1 exu_U22188(.A(exu_n11697), .B(exu_n16274), .Y(exu_n23248));
INVX1 exu_U22189(.A(exu_n23248), .Y(exu_n6586));
AND2X1 exu_U22190(.A(ecc_byp_ecc_result_m[5]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23252));
INVX1 exu_U22191(.A(exu_n23252), .Y(exu_n6587));
AND2X1 exu_U22192(.A(exu_n11698), .B(exu_n16274), .Y(exu_n23254));
INVX1 exu_U22193(.A(exu_n23254), .Y(exu_n6588));
AND2X1 exu_U22194(.A(ecc_byp_ecc_result_m[59]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23258));
INVX1 exu_U22195(.A(exu_n23258), .Y(exu_n6589));
AND2X1 exu_U22196(.A(exu_n11699), .B(exu_n16274), .Y(exu_n23260));
INVX1 exu_U22197(.A(exu_n23260), .Y(exu_n6590));
AND2X1 exu_U22198(.A(ecc_byp_ecc_result_m[58]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23264));
INVX1 exu_U22199(.A(exu_n23264), .Y(exu_n6591));
AND2X1 exu_U22200(.A(exu_n11700), .B(exu_n16274), .Y(exu_n23266));
INVX1 exu_U22201(.A(exu_n23266), .Y(exu_n6592));
AND2X1 exu_U22202(.A(ecc_byp_ecc_result_m[57]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23270));
INVX1 exu_U22203(.A(exu_n23270), .Y(exu_n6593));
AND2X1 exu_U22204(.A(exu_n11701), .B(exu_n16274), .Y(exu_n23272));
INVX1 exu_U22205(.A(exu_n23272), .Y(exu_n6594));
AND2X1 exu_U22206(.A(ecc_byp_ecc_result_m[56]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23276));
INVX1 exu_U22207(.A(exu_n23276), .Y(exu_n6595));
AND2X1 exu_U22208(.A(exu_n11702), .B(exu_n16274), .Y(exu_n23278));
INVX1 exu_U22209(.A(exu_n23278), .Y(exu_n6596));
AND2X1 exu_U22210(.A(ecc_byp_ecc_result_m[55]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23282));
INVX1 exu_U22211(.A(exu_n23282), .Y(exu_n6597));
AND2X1 exu_U22212(.A(exu_n11703), .B(exu_n16274), .Y(exu_n23284));
INVX1 exu_U22213(.A(exu_n23284), .Y(exu_n6598));
AND2X1 exu_U22214(.A(ecc_byp_ecc_result_m[54]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23288));
INVX1 exu_U22215(.A(exu_n23288), .Y(exu_n6599));
AND2X1 exu_U22216(.A(exu_n11704), .B(exu_n16274), .Y(exu_n23290));
INVX1 exu_U22217(.A(exu_n23290), .Y(exu_n6600));
AND2X1 exu_U22218(.A(ecc_byp_ecc_result_m[53]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23294));
INVX1 exu_U22219(.A(exu_n23294), .Y(exu_n6601));
AND2X1 exu_U22220(.A(exu_n11705), .B(exu_n16274), .Y(exu_n23296));
INVX1 exu_U22221(.A(exu_n23296), .Y(exu_n6602));
AND2X1 exu_U22222(.A(ecc_byp_ecc_result_m[52]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23300));
INVX1 exu_U22223(.A(exu_n23300), .Y(exu_n6603));
AND2X1 exu_U22224(.A(exu_n11706), .B(exu_n16274), .Y(exu_n23302));
INVX1 exu_U22225(.A(exu_n23302), .Y(exu_n6604));
AND2X1 exu_U22226(.A(ecc_byp_ecc_result_m[51]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23306));
INVX1 exu_U22227(.A(exu_n23306), .Y(exu_n6605));
AND2X1 exu_U22228(.A(exu_n11707), .B(exu_n16274), .Y(exu_n23308));
INVX1 exu_U22229(.A(exu_n23308), .Y(exu_n6606));
AND2X1 exu_U22230(.A(ecc_byp_ecc_result_m[50]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23312));
INVX1 exu_U22231(.A(exu_n23312), .Y(exu_n6607));
AND2X1 exu_U22232(.A(exu_n11708), .B(exu_n16274), .Y(exu_n23314));
INVX1 exu_U22233(.A(exu_n23314), .Y(exu_n6608));
AND2X1 exu_U22234(.A(ecc_byp_ecc_result_m[4]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23318));
INVX1 exu_U22235(.A(exu_n23318), .Y(exu_n6609));
AND2X1 exu_U22236(.A(exu_n11709), .B(exu_n16274), .Y(exu_n23320));
INVX1 exu_U22237(.A(exu_n23320), .Y(exu_n6610));
AND2X1 exu_U22238(.A(ecc_byp_ecc_result_m[49]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23324));
INVX1 exu_U22239(.A(exu_n23324), .Y(exu_n6611));
AND2X1 exu_U22240(.A(exu_n11710), .B(exu_n16274), .Y(exu_n23326));
INVX1 exu_U22241(.A(exu_n23326), .Y(exu_n6612));
AND2X1 exu_U22242(.A(ecc_byp_ecc_result_m[48]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23330));
INVX1 exu_U22243(.A(exu_n23330), .Y(exu_n6613));
AND2X1 exu_U22244(.A(exu_n11711), .B(exu_n16274), .Y(exu_n23332));
INVX1 exu_U22245(.A(exu_n23332), .Y(exu_n6614));
AND2X1 exu_U22246(.A(ecc_byp_ecc_result_m[47]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23336));
INVX1 exu_U22247(.A(exu_n23336), .Y(exu_n6615));
AND2X1 exu_U22248(.A(exu_n11712), .B(exu_n16274), .Y(exu_n23338));
INVX1 exu_U22249(.A(exu_n23338), .Y(exu_n6616));
AND2X1 exu_U22250(.A(ecc_byp_ecc_result_m[46]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23342));
INVX1 exu_U22251(.A(exu_n23342), .Y(exu_n6617));
AND2X1 exu_U22252(.A(exu_n11713), .B(exu_n16274), .Y(exu_n23344));
INVX1 exu_U22253(.A(exu_n23344), .Y(exu_n6618));
AND2X1 exu_U22254(.A(ecc_byp_ecc_result_m[45]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23348));
INVX1 exu_U22255(.A(exu_n23348), .Y(exu_n6619));
AND2X1 exu_U22256(.A(exu_n11714), .B(exu_n16274), .Y(exu_n23350));
INVX1 exu_U22257(.A(exu_n23350), .Y(exu_n6620));
AND2X1 exu_U22258(.A(ecc_byp_ecc_result_m[44]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23354));
INVX1 exu_U22259(.A(exu_n23354), .Y(exu_n6621));
AND2X1 exu_U22260(.A(exu_n11715), .B(exu_n16274), .Y(exu_n23356));
INVX1 exu_U22261(.A(exu_n23356), .Y(exu_n6622));
AND2X1 exu_U22262(.A(ecc_byp_ecc_result_m[43]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23360));
INVX1 exu_U22263(.A(exu_n23360), .Y(exu_n6623));
AND2X1 exu_U22264(.A(exu_n11716), .B(exu_n16274), .Y(exu_n23362));
INVX1 exu_U22265(.A(exu_n23362), .Y(exu_n6624));
AND2X1 exu_U22266(.A(ecc_byp_ecc_result_m[42]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23366));
INVX1 exu_U22267(.A(exu_n23366), .Y(exu_n6625));
AND2X1 exu_U22268(.A(exu_n11717), .B(exu_n16274), .Y(exu_n23368));
INVX1 exu_U22269(.A(exu_n23368), .Y(exu_n6626));
AND2X1 exu_U22270(.A(ecc_byp_ecc_result_m[41]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23372));
INVX1 exu_U22271(.A(exu_n23372), .Y(exu_n6627));
AND2X1 exu_U22272(.A(exu_n11718), .B(exu_n16274), .Y(exu_n23374));
INVX1 exu_U22273(.A(exu_n23374), .Y(exu_n6628));
AND2X1 exu_U22274(.A(ecc_byp_ecc_result_m[40]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23378));
INVX1 exu_U22275(.A(exu_n23378), .Y(exu_n6629));
AND2X1 exu_U22276(.A(exu_n11719), .B(exu_n16274), .Y(exu_n23380));
INVX1 exu_U22277(.A(exu_n23380), .Y(exu_n6630));
AND2X1 exu_U22278(.A(ecc_byp_ecc_result_m[3]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23384));
INVX1 exu_U22279(.A(exu_n23384), .Y(exu_n6631));
AND2X1 exu_U22280(.A(exu_n11720), .B(exu_n16274), .Y(exu_n23386));
INVX1 exu_U22281(.A(exu_n23386), .Y(exu_n6632));
AND2X1 exu_U22282(.A(ecc_byp_ecc_result_m[39]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23390));
INVX1 exu_U22283(.A(exu_n23390), .Y(exu_n6633));
AND2X1 exu_U22284(.A(exu_n11721), .B(exu_n16274), .Y(exu_n23392));
INVX1 exu_U22285(.A(exu_n23392), .Y(exu_n6634));
AND2X1 exu_U22286(.A(ecc_byp_ecc_result_m[38]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23396));
INVX1 exu_U22287(.A(exu_n23396), .Y(exu_n6635));
AND2X1 exu_U22288(.A(exu_n11722), .B(exu_n16274), .Y(exu_n23398));
INVX1 exu_U22289(.A(exu_n23398), .Y(exu_n6636));
AND2X1 exu_U22290(.A(ecc_byp_ecc_result_m[37]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23402));
INVX1 exu_U22291(.A(exu_n23402), .Y(exu_n6637));
AND2X1 exu_U22292(.A(exu_n11723), .B(exu_n16274), .Y(exu_n23404));
INVX1 exu_U22293(.A(exu_n23404), .Y(exu_n6638));
AND2X1 exu_U22294(.A(ecc_byp_ecc_result_m[36]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23408));
INVX1 exu_U22295(.A(exu_n23408), .Y(exu_n6639));
AND2X1 exu_U22296(.A(exu_n11724), .B(exu_n16274), .Y(exu_n23410));
INVX1 exu_U22297(.A(exu_n23410), .Y(exu_n6640));
AND2X1 exu_U22298(.A(ecc_byp_ecc_result_m[35]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23414));
INVX1 exu_U22299(.A(exu_n23414), .Y(exu_n6641));
AND2X1 exu_U22300(.A(exu_n11725), .B(exu_n16274), .Y(exu_n23416));
INVX1 exu_U22301(.A(exu_n23416), .Y(exu_n6642));
AND2X1 exu_U22302(.A(ecc_byp_ecc_result_m[34]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23420));
INVX1 exu_U22303(.A(exu_n23420), .Y(exu_n6643));
AND2X1 exu_U22304(.A(exu_n11726), .B(exu_n16274), .Y(exu_n23422));
INVX1 exu_U22305(.A(exu_n23422), .Y(exu_n6644));
AND2X1 exu_U22306(.A(ecc_byp_ecc_result_m[33]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23426));
INVX1 exu_U22307(.A(exu_n23426), .Y(exu_n6645));
AND2X1 exu_U22308(.A(exu_n11727), .B(exu_n16274), .Y(exu_n23428));
INVX1 exu_U22309(.A(exu_n23428), .Y(exu_n6646));
AND2X1 exu_U22310(.A(ecc_byp_ecc_result_m[32]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23432));
INVX1 exu_U22311(.A(exu_n23432), .Y(exu_n6647));
AND2X1 exu_U22312(.A(exu_n11728), .B(exu_n16274), .Y(exu_n23434));
INVX1 exu_U22313(.A(exu_n23434), .Y(exu_n6648));
AND2X1 exu_U22314(.A(ecc_byp_ecc_result_m[31]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23438));
INVX1 exu_U22315(.A(exu_n23438), .Y(exu_n6649));
AND2X1 exu_U22316(.A(exu_n11729), .B(exu_n16274), .Y(exu_n23440));
INVX1 exu_U22317(.A(exu_n23440), .Y(exu_n6650));
AND2X1 exu_U22318(.A(ecc_byp_ecc_result_m[30]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23444));
INVX1 exu_U22319(.A(exu_n23444), .Y(exu_n6651));
AND2X1 exu_U22320(.A(exu_n11730), .B(exu_n16274), .Y(exu_n23446));
INVX1 exu_U22321(.A(exu_n23446), .Y(exu_n6652));
AND2X1 exu_U22322(.A(ecc_byp_ecc_result_m[2]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23450));
INVX1 exu_U22323(.A(exu_n23450), .Y(exu_n6653));
AND2X1 exu_U22324(.A(exu_n11731), .B(exu_n16274), .Y(exu_n23452));
INVX1 exu_U22325(.A(exu_n23452), .Y(exu_n6654));
AND2X1 exu_U22326(.A(ecc_byp_ecc_result_m[29]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23456));
INVX1 exu_U22327(.A(exu_n23456), .Y(exu_n6655));
AND2X1 exu_U22328(.A(exu_n11732), .B(exu_n16274), .Y(exu_n23458));
INVX1 exu_U22329(.A(exu_n23458), .Y(exu_n6656));
AND2X1 exu_U22330(.A(ecc_byp_ecc_result_m[28]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23462));
INVX1 exu_U22331(.A(exu_n23462), .Y(exu_n6657));
AND2X1 exu_U22332(.A(exu_n11733), .B(exu_n16274), .Y(exu_n23464));
INVX1 exu_U22333(.A(exu_n23464), .Y(exu_n6658));
AND2X1 exu_U22334(.A(ecc_byp_ecc_result_m[27]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23468));
INVX1 exu_U22335(.A(exu_n23468), .Y(exu_n6659));
AND2X1 exu_U22336(.A(exu_n11734), .B(exu_n16274), .Y(exu_n23470));
INVX1 exu_U22337(.A(exu_n23470), .Y(exu_n6660));
AND2X1 exu_U22338(.A(ecc_byp_ecc_result_m[26]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23474));
INVX1 exu_U22339(.A(exu_n23474), .Y(exu_n6661));
AND2X1 exu_U22340(.A(exu_n11735), .B(exu_n16274), .Y(exu_n23476));
INVX1 exu_U22341(.A(exu_n23476), .Y(exu_n6662));
AND2X1 exu_U22342(.A(ecc_byp_ecc_result_m[25]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23480));
INVX1 exu_U22343(.A(exu_n23480), .Y(exu_n6663));
AND2X1 exu_U22344(.A(exu_n11736), .B(exu_n16274), .Y(exu_n23482));
INVX1 exu_U22345(.A(exu_n23482), .Y(exu_n6664));
AND2X1 exu_U22346(.A(ecc_byp_ecc_result_m[24]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23486));
INVX1 exu_U22347(.A(exu_n23486), .Y(exu_n6665));
AND2X1 exu_U22348(.A(exu_n11737), .B(exu_n16274), .Y(exu_n23488));
INVX1 exu_U22349(.A(exu_n23488), .Y(exu_n6666));
AND2X1 exu_U22350(.A(ecc_byp_ecc_result_m[23]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23492));
INVX1 exu_U22351(.A(exu_n23492), .Y(exu_n6667));
AND2X1 exu_U22352(.A(exu_n11738), .B(exu_n16274), .Y(exu_n23494));
INVX1 exu_U22353(.A(exu_n23494), .Y(exu_n6668));
AND2X1 exu_U22354(.A(ecc_byp_ecc_result_m[22]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23498));
INVX1 exu_U22355(.A(exu_n23498), .Y(exu_n6669));
AND2X1 exu_U22356(.A(exu_n11739), .B(exu_n16274), .Y(exu_n23500));
INVX1 exu_U22357(.A(exu_n23500), .Y(exu_n6670));
AND2X1 exu_U22358(.A(ecc_byp_ecc_result_m[21]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23504));
INVX1 exu_U22359(.A(exu_n23504), .Y(exu_n6671));
AND2X1 exu_U22360(.A(exu_n11740), .B(exu_n16274), .Y(exu_n23506));
INVX1 exu_U22361(.A(exu_n23506), .Y(exu_n6672));
AND2X1 exu_U22362(.A(ecc_byp_ecc_result_m[20]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23510));
INVX1 exu_U22363(.A(exu_n23510), .Y(exu_n6673));
AND2X1 exu_U22364(.A(exu_n11741), .B(exu_n16274), .Y(exu_n23512));
INVX1 exu_U22365(.A(exu_n23512), .Y(exu_n6674));
AND2X1 exu_U22366(.A(ecc_byp_ecc_result_m[1]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23516));
INVX1 exu_U22367(.A(exu_n23516), .Y(exu_n6675));
AND2X1 exu_U22368(.A(exu_n11742), .B(exu_n16274), .Y(exu_n23518));
INVX1 exu_U22369(.A(exu_n23518), .Y(exu_n6676));
AND2X1 exu_U22370(.A(ecc_byp_ecc_result_m[19]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23522));
INVX1 exu_U22371(.A(exu_n23522), .Y(exu_n6677));
AND2X1 exu_U22372(.A(exu_n11743), .B(exu_n16274), .Y(exu_n23524));
INVX1 exu_U22373(.A(exu_n23524), .Y(exu_n6678));
AND2X1 exu_U22374(.A(ecc_byp_ecc_result_m[18]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23528));
INVX1 exu_U22375(.A(exu_n23528), .Y(exu_n6679));
AND2X1 exu_U22376(.A(exu_n11744), .B(exu_n16274), .Y(exu_n23530));
INVX1 exu_U22377(.A(exu_n23530), .Y(exu_n6680));
AND2X1 exu_U22378(.A(ecc_byp_ecc_result_m[17]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23534));
INVX1 exu_U22379(.A(exu_n23534), .Y(exu_n6681));
AND2X1 exu_U22380(.A(exu_n11745), .B(exu_n16274), .Y(exu_n23536));
INVX1 exu_U22381(.A(exu_n23536), .Y(exu_n6682));
AND2X1 exu_U22382(.A(ecc_byp_ecc_result_m[16]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23540));
INVX1 exu_U22383(.A(exu_n23540), .Y(exu_n6683));
AND2X1 exu_U22384(.A(exu_n11746), .B(exu_n16274), .Y(exu_n23542));
INVX1 exu_U22385(.A(exu_n23542), .Y(exu_n6684));
AND2X1 exu_U22386(.A(ecc_byp_ecc_result_m[15]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23546));
INVX1 exu_U22387(.A(exu_n23546), .Y(exu_n6685));
AND2X1 exu_U22388(.A(exu_n11747), .B(exu_n16274), .Y(exu_n23548));
INVX1 exu_U22389(.A(exu_n23548), .Y(exu_n6686));
AND2X1 exu_U22390(.A(ecc_byp_ecc_result_m[14]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23552));
INVX1 exu_U22391(.A(exu_n23552), .Y(exu_n6687));
AND2X1 exu_U22392(.A(exu_n11748), .B(exu_n16274), .Y(exu_n23554));
INVX1 exu_U22393(.A(exu_n23554), .Y(exu_n6688));
AND2X1 exu_U22394(.A(ecc_byp_ecc_result_m[13]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23558));
INVX1 exu_U22395(.A(exu_n23558), .Y(exu_n6689));
AND2X1 exu_U22396(.A(exu_n11749), .B(exu_n16274), .Y(exu_n23560));
INVX1 exu_U22397(.A(exu_n23560), .Y(exu_n6690));
AND2X1 exu_U22398(.A(ecc_byp_ecc_result_m[12]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23564));
INVX1 exu_U22399(.A(exu_n23564), .Y(exu_n6691));
AND2X1 exu_U22400(.A(exu_n11750), .B(exu_n16274), .Y(exu_n23566));
INVX1 exu_U22401(.A(exu_n23566), .Y(exu_n6692));
AND2X1 exu_U22402(.A(ecc_byp_ecc_result_m[11]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23570));
INVX1 exu_U22403(.A(exu_n23570), .Y(exu_n6693));
AND2X1 exu_U22404(.A(exu_n11751), .B(exu_n16274), .Y(exu_n23572));
INVX1 exu_U22405(.A(exu_n23572), .Y(exu_n6694));
AND2X1 exu_U22406(.A(ecc_byp_ecc_result_m[10]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23576));
INVX1 exu_U22407(.A(exu_n23576), .Y(exu_n6695));
AND2X1 exu_U22408(.A(exu_n11752), .B(exu_n16274), .Y(exu_n23578));
INVX1 exu_U22409(.A(exu_n23578), .Y(exu_n6696));
AND2X1 exu_U22410(.A(ecc_byp_ecc_result_m[0]), .B(ecl_byp_sel_ecc_m), .Y(exu_n23582));
INVX1 exu_U22411(.A(exu_n23582), .Y(exu_n6697));
AND2X1 exu_U22412(.A(exu_n11753), .B(exu_n16274), .Y(exu_n23584));
INVX1 exu_U22413(.A(exu_n23584), .Y(exu_n6698));
AND2X1 exu_U22414(.A(exu_n16307), .B(exu_n15211), .Y(exu_n23588));
INVX1 exu_U22415(.A(exu_n23588), .Y(exu_n6699));
AND2X1 exu_U22416(.A(exu_n16310), .B(exu_tlu_wsr_data_m[9]), .Y(exu_n23590));
INVX1 exu_U22417(.A(exu_n23590), .Y(exu_n6700));
AND2X1 exu_U22418(.A(exu_n15271), .B(exu_n16307), .Y(exu_n23594));
INVX1 exu_U22419(.A(exu_n23594), .Y(exu_n6701));
AND2X1 exu_U22420(.A(exu_tlu_wsr_data_m[8]), .B(exu_n16310), .Y(exu_n23596));
INVX1 exu_U22421(.A(exu_n23596), .Y(exu_n6702));
AND2X1 exu_U22422(.A(exu_n15272), .B(exu_n16307), .Y(exu_n23600));
INVX1 exu_U22423(.A(exu_n23600), .Y(exu_n6703));
AND2X1 exu_U22424(.A(exu_tlu_wsr_data_m[7]), .B(exu_n16310), .Y(exu_n23602));
INVX1 exu_U22425(.A(exu_n23602), .Y(exu_n6704));
AND2X1 exu_U22426(.A(exu_n15273), .B(exu_n16307), .Y(exu_n23606));
INVX1 exu_U22427(.A(exu_n23606), .Y(exu_n6705));
AND2X1 exu_U22428(.A(exu_tlu_wsr_data_m[6]), .B(exu_n16310), .Y(exu_n23608));
INVX1 exu_U22429(.A(exu_n23608), .Y(exu_n6706));
AND2X1 exu_U22430(.A(exu_n15274), .B(exu_n16307), .Y(exu_n23611));
INVX1 exu_U22431(.A(exu_n23611), .Y(exu_n6707));
AND2X1 exu_U22432(.A(exu_tlu_wsr_data_m[63]), .B(exu_n16310), .Y(exu_n23613));
INVX1 exu_U22433(.A(exu_n23613), .Y(exu_n6708));
AND2X1 exu_U22434(.A(exu_n15275), .B(exu_n16307), .Y(exu_n23616));
INVX1 exu_U22435(.A(exu_n23616), .Y(exu_n6709));
AND2X1 exu_U22436(.A(exu_tlu_wsr_data_m[62]), .B(exu_n16310), .Y(exu_n23618));
INVX1 exu_U22437(.A(exu_n23618), .Y(exu_n6710));
AND2X1 exu_U22438(.A(exu_n15276), .B(exu_n16307), .Y(exu_n23621));
INVX1 exu_U22439(.A(exu_n23621), .Y(exu_n6711));
AND2X1 exu_U22440(.A(exu_tlu_wsr_data_m[61]), .B(exu_n16310), .Y(exu_n23623));
INVX1 exu_U22441(.A(exu_n23623), .Y(exu_n6712));
AND2X1 exu_U22442(.A(exu_n15277), .B(exu_n16307), .Y(exu_n23626));
INVX1 exu_U22443(.A(exu_n23626), .Y(exu_n6713));
AND2X1 exu_U22444(.A(exu_tlu_wsr_data_m[60]), .B(exu_n16310), .Y(exu_n23628));
INVX1 exu_U22445(.A(exu_n23628), .Y(exu_n6714));
AND2X1 exu_U22446(.A(exu_n15278), .B(exu_n16307), .Y(exu_n23632));
INVX1 exu_U22447(.A(exu_n23632), .Y(exu_n6715));
AND2X1 exu_U22448(.A(exu_tlu_wsr_data_m[5]), .B(exu_n16310), .Y(exu_n23634));
INVX1 exu_U22449(.A(exu_n23634), .Y(exu_n6716));
AND2X1 exu_U22450(.A(exu_n15279), .B(exu_n16307), .Y(exu_n23637));
INVX1 exu_U22451(.A(exu_n23637), .Y(exu_n6717));
AND2X1 exu_U22452(.A(exu_tlu_wsr_data_m[59]), .B(exu_n16310), .Y(exu_n23639));
INVX1 exu_U22453(.A(exu_n23639), .Y(exu_n6718));
AND2X1 exu_U22454(.A(exu_n15280), .B(exu_n16307), .Y(exu_n23642));
INVX1 exu_U22455(.A(exu_n23642), .Y(exu_n6719));
AND2X1 exu_U22456(.A(exu_tlu_wsr_data_m[58]), .B(exu_n16310), .Y(exu_n23644));
INVX1 exu_U22457(.A(exu_n23644), .Y(exu_n6720));
AND2X1 exu_U22458(.A(exu_n15281), .B(exu_n16307), .Y(exu_n23647));
INVX1 exu_U22459(.A(exu_n23647), .Y(exu_n6721));
AND2X1 exu_U22460(.A(exu_tlu_wsr_data_m[57]), .B(exu_n16310), .Y(exu_n23649));
INVX1 exu_U22461(.A(exu_n23649), .Y(exu_n6722));
AND2X1 exu_U22462(.A(exu_n15282), .B(exu_n16307), .Y(exu_n23652));
INVX1 exu_U22463(.A(exu_n23652), .Y(exu_n6723));
AND2X1 exu_U22464(.A(exu_tlu_wsr_data_m[56]), .B(exu_n16310), .Y(exu_n23654));
INVX1 exu_U22465(.A(exu_n23654), .Y(exu_n6724));
AND2X1 exu_U22466(.A(exu_n15283), .B(exu_n16307), .Y(exu_n23657));
INVX1 exu_U22467(.A(exu_n23657), .Y(exu_n6725));
AND2X1 exu_U22468(.A(exu_tlu_wsr_data_m[55]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23659));
INVX1 exu_U22469(.A(exu_n23659), .Y(exu_n6726));
AND2X1 exu_U22470(.A(exu_n15284), .B(exu_n16307), .Y(exu_n23662));
INVX1 exu_U22471(.A(exu_n23662), .Y(exu_n6727));
AND2X1 exu_U22472(.A(exu_tlu_wsr_data_m[54]), .B(exu_n16310), .Y(exu_n23664));
INVX1 exu_U22473(.A(exu_n23664), .Y(exu_n6728));
AND2X1 exu_U22474(.A(exu_n15285), .B(exu_n16307), .Y(exu_n23667));
INVX1 exu_U22475(.A(exu_n23667), .Y(exu_n6729));
AND2X1 exu_U22476(.A(exu_tlu_wsr_data_m[53]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23669));
INVX1 exu_U22477(.A(exu_n23669), .Y(exu_n6730));
AND2X1 exu_U22478(.A(exu_n15286), .B(exu_n16307), .Y(exu_n23672));
INVX1 exu_U22479(.A(exu_n23672), .Y(exu_n6731));
AND2X1 exu_U22480(.A(exu_tlu_wsr_data_m[52]), .B(exu_n16310), .Y(exu_n23674));
INVX1 exu_U22481(.A(exu_n23674), .Y(exu_n6732));
AND2X1 exu_U22482(.A(exu_n15287), .B(exu_n16307), .Y(exu_n23677));
INVX1 exu_U22483(.A(exu_n23677), .Y(exu_n6733));
AND2X1 exu_U22484(.A(exu_tlu_wsr_data_m[51]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23679));
INVX1 exu_U22485(.A(exu_n23679), .Y(exu_n6734));
AND2X1 exu_U22486(.A(exu_n15288), .B(exu_n16307), .Y(exu_n23682));
INVX1 exu_U22487(.A(exu_n23682), .Y(exu_n6735));
AND2X1 exu_U22488(.A(exu_tlu_wsr_data_m[50]), .B(exu_n16310), .Y(exu_n23684));
INVX1 exu_U22489(.A(exu_n23684), .Y(exu_n6736));
AND2X1 exu_U22490(.A(exu_n15289), .B(exu_n16307), .Y(exu_n23688));
INVX1 exu_U22491(.A(exu_n23688), .Y(exu_n6737));
AND2X1 exu_U22492(.A(exu_tlu_wsr_data_m[4]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23690));
INVX1 exu_U22493(.A(exu_n23690), .Y(exu_n6738));
AND2X1 exu_U22494(.A(exu_n15290), .B(exu_n16307), .Y(exu_n23693));
INVX1 exu_U22495(.A(exu_n23693), .Y(exu_n6739));
AND2X1 exu_U22496(.A(exu_tlu_wsr_data_m[49]), .B(exu_n16310), .Y(exu_n23695));
INVX1 exu_U22497(.A(exu_n23695), .Y(exu_n6740));
AND2X1 exu_U22498(.A(exu_n15291), .B(exu_n16307), .Y(exu_n23698));
INVX1 exu_U22499(.A(exu_n23698), .Y(exu_n6741));
AND2X1 exu_U22500(.A(exu_tlu_wsr_data_m[48]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23700));
INVX1 exu_U22501(.A(exu_n23700), .Y(exu_n6742));
AND2X1 exu_U22502(.A(exu_n15292), .B(exu_n16307), .Y(exu_n23704));
INVX1 exu_U22503(.A(exu_n23704), .Y(exu_n6743));
AND2X1 exu_U22504(.A(exu_tlu_wsr_data_m[47]), .B(exu_n16310), .Y(exu_n23706));
INVX1 exu_U22505(.A(exu_n23706), .Y(exu_n6744));
AND2X1 exu_U22506(.A(exu_n15293), .B(exu_n16307), .Y(exu_n23710));
INVX1 exu_U22507(.A(exu_n23710), .Y(exu_n6745));
AND2X1 exu_U22508(.A(exu_tlu_wsr_data_m[46]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23712));
INVX1 exu_U22509(.A(exu_n23712), .Y(exu_n6746));
AND2X1 exu_U22510(.A(exu_n15294), .B(exu_n16307), .Y(exu_n23716));
INVX1 exu_U22511(.A(exu_n23716), .Y(exu_n6747));
AND2X1 exu_U22512(.A(exu_tlu_wsr_data_m[45]), .B(exu_n16310), .Y(exu_n23718));
INVX1 exu_U22513(.A(exu_n23718), .Y(exu_n6748));
AND2X1 exu_U22514(.A(exu_n15295), .B(exu_n16307), .Y(exu_n23722));
INVX1 exu_U22515(.A(exu_n23722), .Y(exu_n6749));
AND2X1 exu_U22516(.A(exu_tlu_wsr_data_m[44]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23724));
INVX1 exu_U22517(.A(exu_n23724), .Y(exu_n6750));
AND2X1 exu_U22518(.A(exu_n15296), .B(exu_n16307), .Y(exu_n23728));
INVX1 exu_U22519(.A(exu_n23728), .Y(exu_n6751));
AND2X1 exu_U22520(.A(exu_tlu_wsr_data_m[43]), .B(exu_n16310), .Y(exu_n23730));
INVX1 exu_U22521(.A(exu_n23730), .Y(exu_n6752));
AND2X1 exu_U22522(.A(exu_n15297), .B(exu_n16307), .Y(exu_n23734));
INVX1 exu_U22523(.A(exu_n23734), .Y(exu_n6753));
AND2X1 exu_U22524(.A(exu_tlu_wsr_data_m[42]), .B(exu_n16310), .Y(exu_n23736));
INVX1 exu_U22525(.A(exu_n23736), .Y(exu_n6754));
AND2X1 exu_U22526(.A(exu_n15298), .B(exu_n16307), .Y(exu_n23740));
INVX1 exu_U22527(.A(exu_n23740), .Y(exu_n6755));
AND2X1 exu_U22528(.A(exu_tlu_wsr_data_m[41]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23742));
INVX1 exu_U22529(.A(exu_n23742), .Y(exu_n6756));
AND2X1 exu_U22530(.A(exu_n15299), .B(exu_n16307), .Y(exu_n23746));
INVX1 exu_U22531(.A(exu_n23746), .Y(exu_n6757));
AND2X1 exu_U22532(.A(exu_tlu_wsr_data_m[40]), .B(exu_n16310), .Y(exu_n23748));
INVX1 exu_U22533(.A(exu_n23748), .Y(exu_n6758));
AND2X1 exu_U22534(.A(exu_n15300), .B(exu_n16307), .Y(exu_n23752));
INVX1 exu_U22535(.A(exu_n23752), .Y(exu_n6759));
AND2X1 exu_U22536(.A(exu_tlu_wsr_data_m[3]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23754));
INVX1 exu_U22537(.A(exu_n23754), .Y(exu_n6760));
AND2X1 exu_U22538(.A(exu_n15301), .B(exu_n16307), .Y(exu_n23758));
INVX1 exu_U22539(.A(exu_n23758), .Y(exu_n6761));
AND2X1 exu_U22540(.A(exu_tlu_wsr_data_m[39]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23760));
INVX1 exu_U22541(.A(exu_n23760), .Y(exu_n6762));
AND2X1 exu_U22542(.A(exu_n15302), .B(exu_n16307), .Y(exu_n23764));
INVX1 exu_U22543(.A(exu_n23764), .Y(exu_n6763));
AND2X1 exu_U22544(.A(exu_tlu_wsr_data_m[38]), .B(exu_n16310), .Y(exu_n23766));
INVX1 exu_U22545(.A(exu_n23766), .Y(exu_n6764));
AND2X1 exu_U22546(.A(exu_n15303), .B(exu_n16307), .Y(exu_n23770));
INVX1 exu_U22547(.A(exu_n23770), .Y(exu_n6765));
AND2X1 exu_U22548(.A(exu_tlu_wsr_data_m[37]), .B(exu_n16310), .Y(exu_n23772));
INVX1 exu_U22549(.A(exu_n23772), .Y(exu_n6766));
AND2X1 exu_U22550(.A(exu_n15304), .B(exu_n16307), .Y(exu_n23776));
INVX1 exu_U22551(.A(exu_n23776), .Y(exu_n6767));
AND2X1 exu_U22552(.A(exu_tlu_wsr_data_m[36]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23778));
INVX1 exu_U22553(.A(exu_n23778), .Y(exu_n6768));
AND2X1 exu_U22554(.A(exu_n15305), .B(exu_n16307), .Y(exu_n23782));
INVX1 exu_U22555(.A(exu_n23782), .Y(exu_n6769));
AND2X1 exu_U22556(.A(exu_tlu_wsr_data_m[35]), .B(exu_n16310), .Y(exu_n23784));
INVX1 exu_U22557(.A(exu_n23784), .Y(exu_n6770));
AND2X1 exu_U22558(.A(exu_n15306), .B(exu_n16307), .Y(exu_n23788));
INVX1 exu_U22559(.A(exu_n23788), .Y(exu_n6771));
AND2X1 exu_U22560(.A(exu_tlu_wsr_data_m[34]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23790));
INVX1 exu_U22561(.A(exu_n23790), .Y(exu_n6772));
AND2X1 exu_U22562(.A(exu_n15307), .B(exu_n16307), .Y(exu_n23794));
INVX1 exu_U22563(.A(exu_n23794), .Y(exu_n6773));
AND2X1 exu_U22564(.A(exu_tlu_wsr_data_m[33]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23796));
INVX1 exu_U22565(.A(exu_n23796), .Y(exu_n6774));
AND2X1 exu_U22566(.A(exu_n15308), .B(exu_n16307), .Y(exu_n23800));
INVX1 exu_U22567(.A(exu_n23800), .Y(exu_n6775));
AND2X1 exu_U22568(.A(exu_tlu_wsr_data_m[32]), .B(exu_n16310), .Y(exu_n23802));
INVX1 exu_U22569(.A(exu_n23802), .Y(exu_n6776));
AND2X1 exu_U22570(.A(exu_n15309), .B(exu_n16307), .Y(exu_n23806));
INVX1 exu_U22571(.A(exu_n23806), .Y(exu_n6777));
AND2X1 exu_U22572(.A(exu_tlu_wsr_data_m[31]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23808));
INVX1 exu_U22573(.A(exu_n23808), .Y(exu_n6778));
AND2X1 exu_U22574(.A(exu_n15310), .B(exu_n16307), .Y(exu_n23812));
INVX1 exu_U22575(.A(exu_n23812), .Y(exu_n6779));
AND2X1 exu_U22576(.A(exu_tlu_wsr_data_m[30]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23814));
INVX1 exu_U22577(.A(exu_n23814), .Y(exu_n6780));
AND2X1 exu_U22578(.A(exu_n15311), .B(exu_n16307), .Y(exu_n23818));
INVX1 exu_U22579(.A(exu_n23818), .Y(exu_n6781));
AND2X1 exu_U22580(.A(exu_tlu_wsr_data_m[2]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23820));
INVX1 exu_U22581(.A(exu_n23820), .Y(exu_n6782));
AND2X1 exu_U22582(.A(exu_n15312), .B(exu_n16307), .Y(exu_n23824));
INVX1 exu_U22583(.A(exu_n23824), .Y(exu_n6783));
AND2X1 exu_U22584(.A(exu_tlu_wsr_data_m[29]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23826));
INVX1 exu_U22585(.A(exu_n23826), .Y(exu_n6784));
AND2X1 exu_U22586(.A(exu_n15313), .B(exu_n16307), .Y(exu_n23830));
INVX1 exu_U22587(.A(exu_n23830), .Y(exu_n6785));
AND2X1 exu_U22588(.A(exu_tlu_wsr_data_m[28]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23832));
INVX1 exu_U22589(.A(exu_n23832), .Y(exu_n6786));
AND2X1 exu_U22590(.A(exu_n15314), .B(exu_n16307), .Y(exu_n23836));
INVX1 exu_U22591(.A(exu_n23836), .Y(exu_n6787));
AND2X1 exu_U22592(.A(exu_tlu_wsr_data_m[27]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23838));
INVX1 exu_U22593(.A(exu_n23838), .Y(exu_n6788));
AND2X1 exu_U22594(.A(exu_n15315), .B(exu_n16307), .Y(exu_n23842));
INVX1 exu_U22595(.A(exu_n23842), .Y(exu_n6789));
AND2X1 exu_U22596(.A(exu_tlu_wsr_data_m[26]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23844));
INVX1 exu_U22597(.A(exu_n23844), .Y(exu_n6790));
AND2X1 exu_U22598(.A(exu_n15316), .B(exu_n16307), .Y(exu_n23848));
INVX1 exu_U22599(.A(exu_n23848), .Y(exu_n6791));
AND2X1 exu_U22600(.A(exu_tlu_wsr_data_m[25]), .B(exu_n16310), .Y(exu_n23850));
INVX1 exu_U22601(.A(exu_n23850), .Y(exu_n6792));
AND2X1 exu_U22602(.A(exu_n15317), .B(exu_n16307), .Y(exu_n23854));
INVX1 exu_U22603(.A(exu_n23854), .Y(exu_n6793));
AND2X1 exu_U22604(.A(exu_tlu_wsr_data_m[24]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23856));
INVX1 exu_U22605(.A(exu_n23856), .Y(exu_n6794));
AND2X1 exu_U22606(.A(exu_n15318), .B(exu_n16307), .Y(exu_n23860));
INVX1 exu_U22607(.A(exu_n23860), .Y(exu_n6795));
AND2X1 exu_U22608(.A(exu_tlu_wsr_data_m[23]), .B(exu_n16310), .Y(exu_n23862));
INVX1 exu_U22609(.A(exu_n23862), .Y(exu_n6796));
AND2X1 exu_U22610(.A(exu_n15319), .B(exu_n16307), .Y(exu_n23866));
INVX1 exu_U22611(.A(exu_n23866), .Y(exu_n6797));
AND2X1 exu_U22612(.A(exu_tlu_wsr_data_m[22]), .B(exu_n16310), .Y(exu_n23868));
INVX1 exu_U22613(.A(exu_n23868), .Y(exu_n6798));
AND2X1 exu_U22614(.A(exu_n15320), .B(exu_n16307), .Y(exu_n23872));
INVX1 exu_U22615(.A(exu_n23872), .Y(exu_n6799));
AND2X1 exu_U22616(.A(exu_tlu_wsr_data_m[21]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23874));
INVX1 exu_U22617(.A(exu_n23874), .Y(exu_n6800));
AND2X1 exu_U22618(.A(exu_n15321), .B(exu_n16307), .Y(exu_n23878));
INVX1 exu_U22619(.A(exu_n23878), .Y(exu_n6801));
AND2X1 exu_U22620(.A(exu_tlu_wsr_data_m[20]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23880));
INVX1 exu_U22621(.A(exu_n23880), .Y(exu_n6802));
AND2X1 exu_U22622(.A(exu_n15322), .B(exu_n16307), .Y(exu_n23884));
INVX1 exu_U22623(.A(exu_n23884), .Y(exu_n6803));
AND2X1 exu_U22624(.A(exu_tlu_wsr_data_m[1]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23886));
INVX1 exu_U22625(.A(exu_n23886), .Y(exu_n6804));
AND2X1 exu_U22626(.A(exu_n15323), .B(exu_n16307), .Y(exu_n23890));
INVX1 exu_U22627(.A(exu_n23890), .Y(exu_n6805));
AND2X1 exu_U22628(.A(exu_tlu_wsr_data_m[19]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23892));
INVX1 exu_U22629(.A(exu_n23892), .Y(exu_n6806));
AND2X1 exu_U22630(.A(exu_n15324), .B(exu_n16307), .Y(exu_n23896));
INVX1 exu_U22631(.A(exu_n23896), .Y(exu_n6807));
AND2X1 exu_U22632(.A(exu_tlu_wsr_data_m[18]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23898));
INVX1 exu_U22633(.A(exu_n23898), .Y(exu_n6808));
AND2X1 exu_U22634(.A(exu_n15325), .B(exu_n16307), .Y(exu_n23902));
INVX1 exu_U22635(.A(exu_n23902), .Y(exu_n6809));
AND2X1 exu_U22636(.A(exu_tlu_wsr_data_m[17]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23904));
INVX1 exu_U22637(.A(exu_n23904), .Y(exu_n6810));
AND2X1 exu_U22638(.A(exu_n15326), .B(exu_n16307), .Y(exu_n23908));
INVX1 exu_U22639(.A(exu_n23908), .Y(exu_n6811));
AND2X1 exu_U22640(.A(exu_tlu_wsr_data_m[16]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23910));
INVX1 exu_U22641(.A(exu_n23910), .Y(exu_n6812));
AND2X1 exu_U22642(.A(exu_n15327), .B(exu_n16307), .Y(exu_n23914));
INVX1 exu_U22643(.A(exu_n23914), .Y(exu_n6813));
AND2X1 exu_U22644(.A(exu_tlu_wsr_data_m[15]), .B(exu_n16310), .Y(exu_n23916));
INVX1 exu_U22645(.A(exu_n23916), .Y(exu_n6814));
AND2X1 exu_U22646(.A(exu_n15328), .B(exu_n16307), .Y(exu_n23920));
INVX1 exu_U22647(.A(exu_n23920), .Y(exu_n6815));
AND2X1 exu_U22648(.A(exu_tlu_wsr_data_m[14]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23922));
INVX1 exu_U22649(.A(exu_n23922), .Y(exu_n6816));
AND2X1 exu_U22650(.A(exu_n15329), .B(exu_n16307), .Y(exu_n23926));
INVX1 exu_U22651(.A(exu_n23926), .Y(exu_n6817));
AND2X1 exu_U22652(.A(exu_tlu_wsr_data_m[13]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23928));
INVX1 exu_U22653(.A(exu_n23928), .Y(exu_n6818));
AND2X1 exu_U22654(.A(exu_n15330), .B(exu_n16307), .Y(exu_n23932));
INVX1 exu_U22655(.A(exu_n23932), .Y(exu_n6819));
AND2X1 exu_U22656(.A(exu_tlu_wsr_data_m[12]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23934));
INVX1 exu_U22657(.A(exu_n23934), .Y(exu_n6820));
AND2X1 exu_U22658(.A(exu_n15331), .B(exu_n16307), .Y(exu_n23938));
INVX1 exu_U22659(.A(exu_n23938), .Y(exu_n6821));
AND2X1 exu_U22660(.A(exu_tlu_wsr_data_m[11]), .B(ecl_byp_rs1_mux1_sel_m), .Y(exu_n23940));
INVX1 exu_U22661(.A(exu_n23940), .Y(exu_n6822));
AND2X1 exu_U22662(.A(exu_n15332), .B(exu_n16307), .Y(exu_n23944));
INVX1 exu_U22663(.A(exu_n23944), .Y(exu_n6823));
AND2X1 exu_U22664(.A(exu_tlu_wsr_data_m[10]), .B(exu_n16310), .Y(exu_n23946));
INVX1 exu_U22665(.A(exu_n23946), .Y(exu_n6824));
AND2X1 exu_U22666(.A(exu_n15333), .B(exu_n16307), .Y(exu_n23950));
INVX1 exu_U22667(.A(exu_n23950), .Y(exu_n6825));
AND2X1 exu_U22668(.A(exu_tlu_wsr_data_m[0]), .B(exu_n16310), .Y(exu_n23952));
INVX1 exu_U22669(.A(exu_n23952), .Y(exu_n6826));
AND2X1 exu_U22670(.A(exu_n16316), .B(alu_byp_rd_data_e[9]), .Y(exu_n23956));
INVX1 exu_U22671(.A(exu_n23956), .Y(exu_n6827));
AND2X1 exu_U22672(.A(exu_n16312), .B(bypass_rs1_data_btwn_mux[9]), .Y(exu_n23958));
INVX1 exu_U22673(.A(exu_n23958), .Y(exu_n6828));
AND2X1 exu_U22674(.A(alu_byp_rd_data_e[8]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n23962));
INVX1 exu_U22675(.A(exu_n23962), .Y(exu_n6829));
AND2X1 exu_U22676(.A(bypass_rs1_data_btwn_mux[8]), .B(exu_n16312), .Y(exu_n23964));
INVX1 exu_U22677(.A(exu_n23964), .Y(exu_n6830));
AND2X1 exu_U22678(.A(alu_byp_rd_data_e[7]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n23968));
INVX1 exu_U22679(.A(exu_n23968), .Y(exu_n6831));
AND2X1 exu_U22680(.A(bypass_rs1_data_btwn_mux[7]), .B(exu_n16312), .Y(exu_n23970));
INVX1 exu_U22681(.A(exu_n23970), .Y(exu_n6832));
AND2X1 exu_U22682(.A(alu_byp_rd_data_e[6]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n23974));
INVX1 exu_U22683(.A(exu_n23974), .Y(exu_n6833));
AND2X1 exu_U22684(.A(bypass_rs1_data_btwn_mux[6]), .B(exu_n16312), .Y(exu_n23976));
INVX1 exu_U22685(.A(exu_n23976), .Y(exu_n6834));
AND2X1 exu_U22686(.A(alu_byp_rd_data_e[63]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n23980));
INVX1 exu_U22687(.A(exu_n23980), .Y(exu_n6835));
AND2X1 exu_U22688(.A(bypass_rs1_data_btwn_mux[63]), .B(exu_n16312), .Y(exu_n23982));
INVX1 exu_U22689(.A(exu_n23982), .Y(exu_n6836));
AND2X1 exu_U22690(.A(alu_byp_rd_data_e[62]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n23986));
INVX1 exu_U22691(.A(exu_n23986), .Y(exu_n6837));
AND2X1 exu_U22692(.A(bypass_rs1_data_btwn_mux[62]), .B(exu_n16312), .Y(exu_n23988));
INVX1 exu_U22693(.A(exu_n23988), .Y(exu_n6838));
AND2X1 exu_U22694(.A(alu_byp_rd_data_e[61]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n23992));
INVX1 exu_U22695(.A(exu_n23992), .Y(exu_n6839));
AND2X1 exu_U22696(.A(bypass_rs1_data_btwn_mux[61]), .B(exu_n16312), .Y(exu_n23994));
INVX1 exu_U22697(.A(exu_n23994), .Y(exu_n6840));
AND2X1 exu_U22698(.A(alu_byp_rd_data_e[60]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n23998));
INVX1 exu_U22699(.A(exu_n23998), .Y(exu_n6841));
AND2X1 exu_U22700(.A(bypass_rs1_data_btwn_mux[60]), .B(exu_n16312), .Y(exu_n24000));
INVX1 exu_U22701(.A(exu_n24000), .Y(exu_n6842));
AND2X1 exu_U22702(.A(alu_byp_rd_data_e[5]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24004));
INVX1 exu_U22703(.A(exu_n24004), .Y(exu_n6843));
AND2X1 exu_U22704(.A(bypass_rs1_data_btwn_mux[5]), .B(exu_n16312), .Y(exu_n24006));
INVX1 exu_U22705(.A(exu_n24006), .Y(exu_n6844));
AND2X1 exu_U22706(.A(alu_byp_rd_data_e[59]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24010));
INVX1 exu_U22707(.A(exu_n24010), .Y(exu_n6845));
AND2X1 exu_U22708(.A(bypass_rs1_data_btwn_mux[59]), .B(exu_n16312), .Y(exu_n24012));
INVX1 exu_U22709(.A(exu_n24012), .Y(exu_n6846));
AND2X1 exu_U22710(.A(alu_byp_rd_data_e[58]), .B(exu_n16316), .Y(exu_n24016));
INVX1 exu_U22711(.A(exu_n24016), .Y(exu_n6847));
AND2X1 exu_U22712(.A(bypass_rs1_data_btwn_mux[58]), .B(exu_n16312), .Y(exu_n24018));
INVX1 exu_U22713(.A(exu_n24018), .Y(exu_n6848));
AND2X1 exu_U22714(.A(alu_byp_rd_data_e[57]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24022));
INVX1 exu_U22715(.A(exu_n24022), .Y(exu_n6849));
AND2X1 exu_U22716(.A(bypass_rs1_data_btwn_mux[57]), .B(exu_n16312), .Y(exu_n24024));
INVX1 exu_U22717(.A(exu_n24024), .Y(exu_n6850));
AND2X1 exu_U22718(.A(alu_byp_rd_data_e[56]), .B(exu_n16316), .Y(exu_n24028));
INVX1 exu_U22719(.A(exu_n24028), .Y(exu_n6851));
AND2X1 exu_U22720(.A(bypass_rs1_data_btwn_mux[56]), .B(exu_n16312), .Y(exu_n24030));
INVX1 exu_U22721(.A(exu_n24030), .Y(exu_n6852));
AND2X1 exu_U22722(.A(alu_byp_rd_data_e[55]), .B(exu_n16316), .Y(exu_n24034));
INVX1 exu_U22723(.A(exu_n24034), .Y(exu_n6853));
AND2X1 exu_U22724(.A(bypass_rs1_data_btwn_mux[55]), .B(exu_n16312), .Y(exu_n24036));
INVX1 exu_U22725(.A(exu_n24036), .Y(exu_n6854));
AND2X1 exu_U22726(.A(alu_byp_rd_data_e[54]), .B(exu_n16316), .Y(exu_n24040));
INVX1 exu_U22727(.A(exu_n24040), .Y(exu_n6855));
AND2X1 exu_U22728(.A(bypass_rs1_data_btwn_mux[54]), .B(exu_n16312), .Y(exu_n24042));
INVX1 exu_U22729(.A(exu_n24042), .Y(exu_n6856));
AND2X1 exu_U22730(.A(alu_byp_rd_data_e[53]), .B(exu_n16316), .Y(exu_n24046));
INVX1 exu_U22731(.A(exu_n24046), .Y(exu_n6857));
AND2X1 exu_U22732(.A(bypass_rs1_data_btwn_mux[53]), .B(exu_n16312), .Y(exu_n24048));
INVX1 exu_U22733(.A(exu_n24048), .Y(exu_n6858));
AND2X1 exu_U22734(.A(alu_byp_rd_data_e[52]), .B(exu_n16316), .Y(exu_n24052));
INVX1 exu_U22735(.A(exu_n24052), .Y(exu_n6859));
AND2X1 exu_U22736(.A(bypass_rs1_data_btwn_mux[52]), .B(exu_n16312), .Y(exu_n24054));
INVX1 exu_U22737(.A(exu_n24054), .Y(exu_n6860));
AND2X1 exu_U22738(.A(alu_byp_rd_data_e[51]), .B(exu_n16316), .Y(exu_n24058));
INVX1 exu_U22739(.A(exu_n24058), .Y(exu_n6861));
AND2X1 exu_U22740(.A(bypass_rs1_data_btwn_mux[51]), .B(exu_n16312), .Y(exu_n24060));
INVX1 exu_U22741(.A(exu_n24060), .Y(exu_n6862));
AND2X1 exu_U22742(.A(alu_byp_rd_data_e[50]), .B(exu_n16316), .Y(exu_n24064));
INVX1 exu_U22743(.A(exu_n24064), .Y(exu_n6863));
AND2X1 exu_U22744(.A(bypass_rs1_data_btwn_mux[50]), .B(exu_n16312), .Y(exu_n24066));
INVX1 exu_U22745(.A(exu_n24066), .Y(exu_n6864));
AND2X1 exu_U22746(.A(alu_byp_rd_data_e[4]), .B(exu_n16316), .Y(exu_n24070));
INVX1 exu_U22747(.A(exu_n24070), .Y(exu_n6865));
AND2X1 exu_U22748(.A(bypass_rs1_data_btwn_mux[4]), .B(exu_n16312), .Y(exu_n24072));
INVX1 exu_U22749(.A(exu_n24072), .Y(exu_n6866));
AND2X1 exu_U22750(.A(alu_byp_rd_data_e[49]), .B(exu_n16316), .Y(exu_n24076));
INVX1 exu_U22751(.A(exu_n24076), .Y(exu_n6867));
AND2X1 exu_U22752(.A(bypass_rs1_data_btwn_mux[49]), .B(exu_n16312), .Y(exu_n24078));
INVX1 exu_U22753(.A(exu_n24078), .Y(exu_n6868));
AND2X1 exu_U22754(.A(alu_byp_rd_data_e[48]), .B(exu_n16316), .Y(exu_n24082));
INVX1 exu_U22755(.A(exu_n24082), .Y(exu_n6869));
AND2X1 exu_U22756(.A(bypass_rs1_data_btwn_mux[48]), .B(exu_n16312), .Y(exu_n24084));
INVX1 exu_U22757(.A(exu_n24084), .Y(exu_n6870));
AND2X1 exu_U22758(.A(alu_byp_rd_data_e[47]), .B(exu_n16316), .Y(exu_n24088));
INVX1 exu_U22759(.A(exu_n24088), .Y(exu_n6871));
AND2X1 exu_U22760(.A(bypass_rs1_data_btwn_mux[47]), .B(exu_n16312), .Y(exu_n24090));
INVX1 exu_U22761(.A(exu_n24090), .Y(exu_n6872));
AND2X1 exu_U22762(.A(alu_byp_rd_data_e[46]), .B(exu_n16316), .Y(exu_n24094));
INVX1 exu_U22763(.A(exu_n24094), .Y(exu_n6873));
AND2X1 exu_U22764(.A(bypass_rs1_data_btwn_mux[46]), .B(exu_n16312), .Y(exu_n24096));
INVX1 exu_U22765(.A(exu_n24096), .Y(exu_n6874));
AND2X1 exu_U22766(.A(alu_byp_rd_data_e[45]), .B(exu_n16316), .Y(exu_n24100));
INVX1 exu_U22767(.A(exu_n24100), .Y(exu_n6875));
AND2X1 exu_U22768(.A(bypass_rs1_data_btwn_mux[45]), .B(exu_n16312), .Y(exu_n24102));
INVX1 exu_U22769(.A(exu_n24102), .Y(exu_n6876));
AND2X1 exu_U22770(.A(alu_byp_rd_data_e[44]), .B(exu_n16316), .Y(exu_n24106));
INVX1 exu_U22771(.A(exu_n24106), .Y(exu_n6877));
AND2X1 exu_U22772(.A(bypass_rs1_data_btwn_mux[44]), .B(exu_n16312), .Y(exu_n24108));
INVX1 exu_U22773(.A(exu_n24108), .Y(exu_n6878));
AND2X1 exu_U22774(.A(alu_byp_rd_data_e[43]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24112));
INVX1 exu_U22775(.A(exu_n24112), .Y(exu_n6879));
AND2X1 exu_U22776(.A(bypass_rs1_data_btwn_mux[43]), .B(exu_n16312), .Y(exu_n24114));
INVX1 exu_U22777(.A(exu_n24114), .Y(exu_n6880));
AND2X1 exu_U22778(.A(alu_byp_rd_data_e[42]), .B(exu_n16316), .Y(exu_n24118));
INVX1 exu_U22779(.A(exu_n24118), .Y(exu_n6881));
AND2X1 exu_U22780(.A(bypass_rs1_data_btwn_mux[42]), .B(exu_n16312), .Y(exu_n24120));
INVX1 exu_U22781(.A(exu_n24120), .Y(exu_n6882));
AND2X1 exu_U22782(.A(alu_byp_rd_data_e[41]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24124));
INVX1 exu_U22783(.A(exu_n24124), .Y(exu_n6883));
AND2X1 exu_U22784(.A(bypass_rs1_data_btwn_mux[41]), .B(exu_n16312), .Y(exu_n24126));
INVX1 exu_U22785(.A(exu_n24126), .Y(exu_n6884));
AND2X1 exu_U22786(.A(alu_byp_rd_data_e[40]), .B(exu_n16316), .Y(exu_n24130));
INVX1 exu_U22787(.A(exu_n24130), .Y(exu_n6885));
AND2X1 exu_U22788(.A(bypass_rs1_data_btwn_mux[40]), .B(exu_n16312), .Y(exu_n24132));
INVX1 exu_U22789(.A(exu_n24132), .Y(exu_n6886));
AND2X1 exu_U22790(.A(alu_byp_rd_data_e[3]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24136));
INVX1 exu_U22791(.A(exu_n24136), .Y(exu_n6887));
AND2X1 exu_U22792(.A(bypass_rs1_data_btwn_mux[3]), .B(exu_n16312), .Y(exu_n24138));
INVX1 exu_U22793(.A(exu_n24138), .Y(exu_n6888));
AND2X1 exu_U22794(.A(alu_byp_rd_data_e[39]), .B(exu_n16316), .Y(exu_n24142));
INVX1 exu_U22795(.A(exu_n24142), .Y(exu_n6889));
AND2X1 exu_U22796(.A(bypass_rs1_data_btwn_mux[39]), .B(exu_n16312), .Y(exu_n24144));
INVX1 exu_U22797(.A(exu_n24144), .Y(exu_n6890));
AND2X1 exu_U22798(.A(alu_byp_rd_data_e[38]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24148));
INVX1 exu_U22799(.A(exu_n24148), .Y(exu_n6891));
AND2X1 exu_U22800(.A(bypass_rs1_data_btwn_mux[38]), .B(exu_n16312), .Y(exu_n24150));
INVX1 exu_U22801(.A(exu_n24150), .Y(exu_n6892));
AND2X1 exu_U22802(.A(alu_byp_rd_data_e[37]), .B(exu_n16316), .Y(exu_n24154));
INVX1 exu_U22803(.A(exu_n24154), .Y(exu_n6893));
AND2X1 exu_U22804(.A(bypass_rs1_data_btwn_mux[37]), .B(exu_n16312), .Y(exu_n24156));
INVX1 exu_U22805(.A(exu_n24156), .Y(exu_n6894));
AND2X1 exu_U22806(.A(alu_byp_rd_data_e[36]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24160));
INVX1 exu_U22807(.A(exu_n24160), .Y(exu_n6895));
AND2X1 exu_U22808(.A(bypass_rs1_data_btwn_mux[36]), .B(exu_n16312), .Y(exu_n24162));
INVX1 exu_U22809(.A(exu_n24162), .Y(exu_n6896));
AND2X1 exu_U22810(.A(alu_byp_rd_data_e[35]), .B(exu_n16316), .Y(exu_n24166));
INVX1 exu_U22811(.A(exu_n24166), .Y(exu_n6897));
AND2X1 exu_U22812(.A(bypass_rs1_data_btwn_mux[35]), .B(exu_n16312), .Y(exu_n24168));
INVX1 exu_U22813(.A(exu_n24168), .Y(exu_n6898));
AND2X1 exu_U22814(.A(alu_byp_rd_data_e[34]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24172));
INVX1 exu_U22815(.A(exu_n24172), .Y(exu_n6899));
AND2X1 exu_U22816(.A(bypass_rs1_data_btwn_mux[34]), .B(exu_n16312), .Y(exu_n24174));
INVX1 exu_U22817(.A(exu_n24174), .Y(exu_n6900));
AND2X1 exu_U22818(.A(alu_byp_rd_data_e[33]), .B(exu_n16316), .Y(exu_n24178));
INVX1 exu_U22819(.A(exu_n24178), .Y(exu_n6901));
AND2X1 exu_U22820(.A(bypass_rs1_data_btwn_mux[33]), .B(exu_n16312), .Y(exu_n24180));
INVX1 exu_U22821(.A(exu_n24180), .Y(exu_n6902));
AND2X1 exu_U22822(.A(alu_byp_rd_data_e[32]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24184));
INVX1 exu_U22823(.A(exu_n24184), .Y(exu_n6903));
AND2X1 exu_U22824(.A(bypass_rs1_data_btwn_mux[32]), .B(exu_n16312), .Y(exu_n24186));
INVX1 exu_U22825(.A(exu_n24186), .Y(exu_n6904));
AND2X1 exu_U22826(.A(alu_byp_rd_data_e[31]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24190));
INVX1 exu_U22827(.A(exu_n24190), .Y(exu_n6905));
AND2X1 exu_U22828(.A(bypass_rs1_data_btwn_mux[31]), .B(exu_n16312), .Y(exu_n24192));
INVX1 exu_U22829(.A(exu_n24192), .Y(exu_n6906));
AND2X1 exu_U22830(.A(alu_byp_rd_data_e[30]), .B(exu_n16316), .Y(exu_n24196));
INVX1 exu_U22831(.A(exu_n24196), .Y(exu_n6907));
AND2X1 exu_U22832(.A(bypass_rs1_data_btwn_mux[30]), .B(exu_n16312), .Y(exu_n24198));
INVX1 exu_U22833(.A(exu_n24198), .Y(exu_n6908));
AND2X1 exu_U22834(.A(alu_byp_rd_data_e[2]), .B(exu_n16316), .Y(exu_n24202));
INVX1 exu_U22835(.A(exu_n24202), .Y(exu_n6909));
AND2X1 exu_U22836(.A(bypass_rs1_data_btwn_mux[2]), .B(exu_n16312), .Y(exu_n24204));
INVX1 exu_U22837(.A(exu_n24204), .Y(exu_n6910));
AND2X1 exu_U22838(.A(alu_byp_rd_data_e[29]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24208));
INVX1 exu_U22839(.A(exu_n24208), .Y(exu_n6911));
AND2X1 exu_U22840(.A(bypass_rs1_data_btwn_mux[29]), .B(exu_n16312), .Y(exu_n24210));
INVX1 exu_U22841(.A(exu_n24210), .Y(exu_n6912));
AND2X1 exu_U22842(.A(alu_byp_rd_data_e[28]), .B(exu_n16316), .Y(exu_n24214));
INVX1 exu_U22843(.A(exu_n24214), .Y(exu_n6913));
AND2X1 exu_U22844(.A(bypass_rs1_data_btwn_mux[28]), .B(exu_n16312), .Y(exu_n24216));
INVX1 exu_U22845(.A(exu_n24216), .Y(exu_n6914));
AND2X1 exu_U22846(.A(alu_byp_rd_data_e[27]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24220));
INVX1 exu_U22847(.A(exu_n24220), .Y(exu_n6915));
AND2X1 exu_U22848(.A(bypass_rs1_data_btwn_mux[27]), .B(exu_n16312), .Y(exu_n24222));
INVX1 exu_U22849(.A(exu_n24222), .Y(exu_n6916));
AND2X1 exu_U22850(.A(alu_byp_rd_data_e[26]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24226));
INVX1 exu_U22851(.A(exu_n24226), .Y(exu_n6917));
AND2X1 exu_U22852(.A(bypass_rs1_data_btwn_mux[26]), .B(exu_n16312), .Y(exu_n24228));
INVX1 exu_U22853(.A(exu_n24228), .Y(exu_n6918));
AND2X1 exu_U22854(.A(alu_byp_rd_data_e[25]), .B(exu_n16316), .Y(exu_n24232));
INVX1 exu_U22855(.A(exu_n24232), .Y(exu_n6919));
AND2X1 exu_U22856(.A(bypass_rs1_data_btwn_mux[25]), .B(exu_n16312), .Y(exu_n24234));
INVX1 exu_U22857(.A(exu_n24234), .Y(exu_n6920));
AND2X1 exu_U22858(.A(alu_byp_rd_data_e[24]), .B(exu_n16316), .Y(exu_n24238));
INVX1 exu_U22859(.A(exu_n24238), .Y(exu_n6921));
AND2X1 exu_U22860(.A(bypass_rs1_data_btwn_mux[24]), .B(exu_n16312), .Y(exu_n24240));
INVX1 exu_U22861(.A(exu_n24240), .Y(exu_n6922));
AND2X1 exu_U22862(.A(alu_byp_rd_data_e[23]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24244));
INVX1 exu_U22863(.A(exu_n24244), .Y(exu_n6923));
AND2X1 exu_U22864(.A(bypass_rs1_data_btwn_mux[23]), .B(exu_n16312), .Y(exu_n24246));
INVX1 exu_U22865(.A(exu_n24246), .Y(exu_n6924));
AND2X1 exu_U22866(.A(alu_byp_rd_data_e[22]), .B(exu_n16316), .Y(exu_n24250));
INVX1 exu_U22867(.A(exu_n24250), .Y(exu_n6925));
AND2X1 exu_U22868(.A(bypass_rs1_data_btwn_mux[22]), .B(exu_n16312), .Y(exu_n24252));
INVX1 exu_U22869(.A(exu_n24252), .Y(exu_n6926));
AND2X1 exu_U22870(.A(alu_byp_rd_data_e[21]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24256));
INVX1 exu_U22871(.A(exu_n24256), .Y(exu_n6927));
AND2X1 exu_U22872(.A(bypass_rs1_data_btwn_mux[21]), .B(exu_n16312), .Y(exu_n24258));
INVX1 exu_U22873(.A(exu_n24258), .Y(exu_n6928));
AND2X1 exu_U22874(.A(alu_byp_rd_data_e[20]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24262));
INVX1 exu_U22875(.A(exu_n24262), .Y(exu_n6929));
AND2X1 exu_U22876(.A(bypass_rs1_data_btwn_mux[20]), .B(exu_n16312), .Y(exu_n24264));
INVX1 exu_U22877(.A(exu_n24264), .Y(exu_n6930));
AND2X1 exu_U22878(.A(alu_byp_rd_data_e[1]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24268));
INVX1 exu_U22879(.A(exu_n24268), .Y(exu_n6931));
AND2X1 exu_U22880(.A(bypass_rs1_data_btwn_mux[1]), .B(exu_n16312), .Y(exu_n24270));
INVX1 exu_U22881(.A(exu_n24270), .Y(exu_n6932));
AND2X1 exu_U22882(.A(alu_byp_rd_data_e[19]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24274));
INVX1 exu_U22883(.A(exu_n24274), .Y(exu_n6933));
AND2X1 exu_U22884(.A(bypass_rs1_data_btwn_mux[19]), .B(exu_n16312), .Y(exu_n24276));
INVX1 exu_U22885(.A(exu_n24276), .Y(exu_n6934));
AND2X1 exu_U22886(.A(alu_byp_rd_data_e[18]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24280));
INVX1 exu_U22887(.A(exu_n24280), .Y(exu_n6935));
AND2X1 exu_U22888(.A(bypass_rs1_data_btwn_mux[18]), .B(exu_n16312), .Y(exu_n24282));
INVX1 exu_U22889(.A(exu_n24282), .Y(exu_n6936));
AND2X1 exu_U22890(.A(alu_byp_rd_data_e[17]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24286));
INVX1 exu_U22891(.A(exu_n24286), .Y(exu_n6937));
AND2X1 exu_U22892(.A(bypass_rs1_data_btwn_mux[17]), .B(exu_n16312), .Y(exu_n24288));
INVX1 exu_U22893(.A(exu_n24288), .Y(exu_n6938));
AND2X1 exu_U22894(.A(alu_byp_rd_data_e[16]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24292));
INVX1 exu_U22895(.A(exu_n24292), .Y(exu_n6939));
AND2X1 exu_U22896(.A(bypass_rs1_data_btwn_mux[16]), .B(exu_n16312), .Y(exu_n24294));
INVX1 exu_U22897(.A(exu_n24294), .Y(exu_n6940));
AND2X1 exu_U22898(.A(alu_byp_rd_data_e[15]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24298));
INVX1 exu_U22899(.A(exu_n24298), .Y(exu_n6941));
AND2X1 exu_U22900(.A(bypass_rs1_data_btwn_mux[15]), .B(exu_n16312), .Y(exu_n24300));
INVX1 exu_U22901(.A(exu_n24300), .Y(exu_n6942));
AND2X1 exu_U22902(.A(alu_byp_rd_data_e[14]), .B(exu_n16316), .Y(exu_n24304));
INVX1 exu_U22903(.A(exu_n24304), .Y(exu_n6943));
AND2X1 exu_U22904(.A(bypass_rs1_data_btwn_mux[14]), .B(exu_n16312), .Y(exu_n24306));
INVX1 exu_U22905(.A(exu_n24306), .Y(exu_n6944));
AND2X1 exu_U22906(.A(alu_byp_rd_data_e[13]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24310));
INVX1 exu_U22907(.A(exu_n24310), .Y(exu_n6945));
AND2X1 exu_U22908(.A(bypass_rs1_data_btwn_mux[13]), .B(exu_n16312), .Y(exu_n24312));
INVX1 exu_U22909(.A(exu_n24312), .Y(exu_n6946));
AND2X1 exu_U22910(.A(alu_byp_rd_data_e[12]), .B(exu_n16316), .Y(exu_n24316));
INVX1 exu_U22911(.A(exu_n24316), .Y(exu_n6947));
AND2X1 exu_U22912(.A(bypass_rs1_data_btwn_mux[12]), .B(exu_n16312), .Y(exu_n24318));
INVX1 exu_U22913(.A(exu_n24318), .Y(exu_n6948));
AND2X1 exu_U22914(.A(alu_byp_rd_data_e[11]), .B(exu_n16316), .Y(exu_n24322));
INVX1 exu_U22915(.A(exu_n24322), .Y(exu_n6949));
AND2X1 exu_U22916(.A(bypass_rs1_data_btwn_mux[11]), .B(exu_n16312), .Y(exu_n24324));
INVX1 exu_U22917(.A(exu_n24324), .Y(exu_n6950));
AND2X1 exu_U22918(.A(alu_byp_rd_data_e[10]), .B(exu_n16316), .Y(exu_n24328));
INVX1 exu_U22919(.A(exu_n24328), .Y(exu_n6951));
AND2X1 exu_U22920(.A(bypass_rs1_data_btwn_mux[10]), .B(exu_n16312), .Y(exu_n24330));
INVX1 exu_U22921(.A(exu_n24330), .Y(exu_n6952));
AND2X1 exu_U22922(.A(alu_byp_rd_data_e[0]), .B(ecl_byp_rs1_mux2_sel_e), .Y(exu_n24334));
INVX1 exu_U22923(.A(exu_n24334), .Y(exu_n6953));
AND2X1 exu_U22924(.A(bypass_rs1_data_btwn_mux[0]), .B(exu_n16312), .Y(exu_n24336));
INVX1 exu_U22925(.A(exu_n24336), .Y(exu_n6954));
AND2X1 exu_U22926(.A(exu_n16302), .B(exu_tlu_wsr_data_m[9]), .Y(exu_n24340));
INVX1 exu_U22927(.A(exu_n24340), .Y(exu_n6955));
AND2X1 exu_U22928(.A(exu_tlu_wsr_data_m[8]), .B(exu_n16302), .Y(exu_n24344));
INVX1 exu_U22929(.A(exu_n24344), .Y(exu_n6956));
AND2X1 exu_U22930(.A(exu_tlu_wsr_data_m[7]), .B(exu_n16302), .Y(exu_n24348));
INVX1 exu_U22931(.A(exu_n24348), .Y(exu_n6957));
AND2X1 exu_U22932(.A(exu_tlu_wsr_data_m[6]), .B(exu_n16302), .Y(exu_n24352));
INVX1 exu_U22933(.A(exu_n24352), .Y(exu_n6958));
AND2X1 exu_U22934(.A(exu_tlu_wsr_data_m[63]), .B(exu_n16302), .Y(exu_n24356));
INVX1 exu_U22935(.A(exu_n24356), .Y(exu_n6959));
AND2X1 exu_U22936(.A(exu_tlu_wsr_data_m[62]), .B(exu_n16302), .Y(exu_n24360));
INVX1 exu_U22937(.A(exu_n24360), .Y(exu_n6960));
AND2X1 exu_U22938(.A(exu_tlu_wsr_data_m[61]), .B(exu_n16302), .Y(exu_n24364));
INVX1 exu_U22939(.A(exu_n24364), .Y(exu_n6961));
AND2X1 exu_U22940(.A(exu_tlu_wsr_data_m[60]), .B(exu_n16302), .Y(exu_n24368));
INVX1 exu_U22941(.A(exu_n24368), .Y(exu_n6962));
AND2X1 exu_U22942(.A(exu_tlu_wsr_data_m[5]), .B(exu_n16302), .Y(exu_n24372));
INVX1 exu_U22943(.A(exu_n24372), .Y(exu_n6963));
AND2X1 exu_U22944(.A(exu_tlu_wsr_data_m[59]), .B(exu_n16302), .Y(exu_n24376));
INVX1 exu_U22945(.A(exu_n24376), .Y(exu_n6964));
AND2X1 exu_U22946(.A(exu_tlu_wsr_data_m[58]), .B(exu_n16302), .Y(exu_n24380));
INVX1 exu_U22947(.A(exu_n24380), .Y(exu_n6965));
AND2X1 exu_U22948(.A(exu_tlu_wsr_data_m[57]), .B(exu_n16302), .Y(exu_n24384));
INVX1 exu_U22949(.A(exu_n24384), .Y(exu_n6966));
AND2X1 exu_U22950(.A(exu_tlu_wsr_data_m[56]), .B(exu_n16302), .Y(exu_n24388));
INVX1 exu_U22951(.A(exu_n24388), .Y(exu_n6967));
AND2X1 exu_U22952(.A(exu_tlu_wsr_data_m[55]), .B(exu_n16302), .Y(exu_n24392));
INVX1 exu_U22953(.A(exu_n24392), .Y(exu_n6968));
AND2X1 exu_U22954(.A(exu_tlu_wsr_data_m[54]), .B(exu_n16302), .Y(exu_n24396));
INVX1 exu_U22955(.A(exu_n24396), .Y(exu_n6969));
AND2X1 exu_U22956(.A(exu_tlu_wsr_data_m[53]), .B(exu_n16302), .Y(exu_n24400));
INVX1 exu_U22957(.A(exu_n24400), .Y(exu_n6970));
AND2X1 exu_U22958(.A(exu_tlu_wsr_data_m[52]), .B(exu_n16302), .Y(exu_n24404));
INVX1 exu_U22959(.A(exu_n24404), .Y(exu_n6971));
AND2X1 exu_U22960(.A(exu_tlu_wsr_data_m[51]), .B(exu_n16302), .Y(exu_n24408));
INVX1 exu_U22961(.A(exu_n24408), .Y(exu_n6972));
AND2X1 exu_U22962(.A(exu_tlu_wsr_data_m[50]), .B(exu_n16302), .Y(exu_n24412));
INVX1 exu_U22963(.A(exu_n24412), .Y(exu_n6973));
AND2X1 exu_U22964(.A(exu_tlu_wsr_data_m[4]), .B(exu_n16302), .Y(exu_n24416));
INVX1 exu_U22965(.A(exu_n24416), .Y(exu_n6974));
AND2X1 exu_U22966(.A(exu_tlu_wsr_data_m[49]), .B(exu_n16302), .Y(exu_n24420));
INVX1 exu_U22967(.A(exu_n24420), .Y(exu_n6975));
AND2X1 exu_U22968(.A(exu_tlu_wsr_data_m[48]), .B(exu_n16302), .Y(exu_n24424));
INVX1 exu_U22969(.A(exu_n24424), .Y(exu_n6976));
AND2X1 exu_U22970(.A(exu_tlu_wsr_data_m[47]), .B(exu_n16302), .Y(exu_n24428));
INVX1 exu_U22971(.A(exu_n24428), .Y(exu_n6977));
AND2X1 exu_U22972(.A(exu_tlu_wsr_data_m[46]), .B(exu_n16302), .Y(exu_n24432));
INVX1 exu_U22973(.A(exu_n24432), .Y(exu_n6978));
AND2X1 exu_U22974(.A(exu_tlu_wsr_data_m[45]), .B(exu_n16302), .Y(exu_n24436));
INVX1 exu_U22975(.A(exu_n24436), .Y(exu_n6979));
AND2X1 exu_U22976(.A(exu_tlu_wsr_data_m[44]), .B(exu_n16302), .Y(exu_n24440));
INVX1 exu_U22977(.A(exu_n24440), .Y(exu_n6980));
AND2X1 exu_U22978(.A(exu_tlu_wsr_data_m[43]), .B(exu_n16302), .Y(exu_n24444));
INVX1 exu_U22979(.A(exu_n24444), .Y(exu_n6981));
AND2X1 exu_U22980(.A(exu_tlu_wsr_data_m[42]), .B(exu_n16302), .Y(exu_n24448));
INVX1 exu_U22981(.A(exu_n24448), .Y(exu_n6982));
AND2X1 exu_U22982(.A(exu_tlu_wsr_data_m[41]), .B(exu_n16302), .Y(exu_n24452));
INVX1 exu_U22983(.A(exu_n24452), .Y(exu_n6983));
AND2X1 exu_U22984(.A(exu_tlu_wsr_data_m[40]), .B(exu_n16302), .Y(exu_n24456));
INVX1 exu_U22985(.A(exu_n24456), .Y(exu_n6984));
AND2X1 exu_U22986(.A(exu_tlu_wsr_data_m[3]), .B(exu_n16302), .Y(exu_n24460));
INVX1 exu_U22987(.A(exu_n24460), .Y(exu_n6985));
AND2X1 exu_U22988(.A(exu_tlu_wsr_data_m[39]), .B(exu_n16302), .Y(exu_n24464));
INVX1 exu_U22989(.A(exu_n24464), .Y(exu_n6986));
AND2X1 exu_U22990(.A(exu_tlu_wsr_data_m[38]), .B(exu_n16302), .Y(exu_n24468));
INVX1 exu_U22991(.A(exu_n24468), .Y(exu_n6987));
AND2X1 exu_U22992(.A(exu_tlu_wsr_data_m[37]), .B(exu_n16302), .Y(exu_n24472));
INVX1 exu_U22993(.A(exu_n24472), .Y(exu_n6988));
AND2X1 exu_U22994(.A(exu_tlu_wsr_data_m[36]), .B(exu_n16302), .Y(exu_n24476));
INVX1 exu_U22995(.A(exu_n24476), .Y(exu_n6989));
AND2X1 exu_U22996(.A(exu_tlu_wsr_data_m[35]), .B(exu_n16302), .Y(exu_n24480));
INVX1 exu_U22997(.A(exu_n24480), .Y(exu_n6990));
AND2X1 exu_U22998(.A(exu_tlu_wsr_data_m[34]), .B(exu_n16302), .Y(exu_n24484));
INVX1 exu_U22999(.A(exu_n24484), .Y(exu_n6991));
AND2X1 exu_U23000(.A(exu_tlu_wsr_data_m[33]), .B(exu_n16302), .Y(exu_n24488));
INVX1 exu_U23001(.A(exu_n24488), .Y(exu_n6992));
AND2X1 exu_U23002(.A(exu_tlu_wsr_data_m[32]), .B(exu_n16302), .Y(exu_n24492));
INVX1 exu_U23003(.A(exu_n24492), .Y(exu_n6993));
AND2X1 exu_U23004(.A(exu_tlu_wsr_data_m[31]), .B(exu_n16302), .Y(exu_n24496));
INVX1 exu_U23005(.A(exu_n24496), .Y(exu_n6994));
AND2X1 exu_U23006(.A(exu_tlu_wsr_data_m[30]), .B(exu_n16302), .Y(exu_n24500));
INVX1 exu_U23007(.A(exu_n24500), .Y(exu_n6995));
AND2X1 exu_U23008(.A(exu_tlu_wsr_data_m[2]), .B(exu_n16302), .Y(exu_n24504));
INVX1 exu_U23009(.A(exu_n24504), .Y(exu_n6996));
AND2X1 exu_U23010(.A(exu_tlu_wsr_data_m[29]), .B(exu_n16302), .Y(exu_n24508));
INVX1 exu_U23011(.A(exu_n24508), .Y(exu_n6997));
AND2X1 exu_U23012(.A(exu_tlu_wsr_data_m[28]), .B(exu_n16302), .Y(exu_n24512));
INVX1 exu_U23013(.A(exu_n24512), .Y(exu_n6998));
AND2X1 exu_U23014(.A(exu_tlu_wsr_data_m[27]), .B(exu_n16302), .Y(exu_n24516));
INVX1 exu_U23015(.A(exu_n24516), .Y(exu_n6999));
AND2X1 exu_U23016(.A(exu_tlu_wsr_data_m[26]), .B(exu_n16302), .Y(exu_n24520));
INVX1 exu_U23017(.A(exu_n24520), .Y(exu_n7000));
AND2X1 exu_U23018(.A(exu_tlu_wsr_data_m[25]), .B(exu_n16302), .Y(exu_n24524));
INVX1 exu_U23019(.A(exu_n24524), .Y(exu_n7001));
AND2X1 exu_U23020(.A(exu_tlu_wsr_data_m[24]), .B(exu_n16302), .Y(exu_n24528));
INVX1 exu_U23021(.A(exu_n24528), .Y(exu_n7002));
AND2X1 exu_U23022(.A(exu_tlu_wsr_data_m[23]), .B(exu_n16302), .Y(exu_n24532));
INVX1 exu_U23023(.A(exu_n24532), .Y(exu_n7003));
AND2X1 exu_U23024(.A(exu_tlu_wsr_data_m[22]), .B(exu_n16302), .Y(exu_n24536));
INVX1 exu_U23025(.A(exu_n24536), .Y(exu_n7004));
AND2X1 exu_U23026(.A(exu_tlu_wsr_data_m[21]), .B(exu_n16302), .Y(exu_n24540));
INVX1 exu_U23027(.A(exu_n24540), .Y(exu_n7005));
AND2X1 exu_U23028(.A(exu_tlu_wsr_data_m[20]), .B(exu_n16302), .Y(exu_n24544));
INVX1 exu_U23029(.A(exu_n24544), .Y(exu_n7006));
AND2X1 exu_U23030(.A(exu_tlu_wsr_data_m[1]), .B(exu_n16302), .Y(exu_n24548));
INVX1 exu_U23031(.A(exu_n24548), .Y(exu_n7007));
AND2X1 exu_U23032(.A(exu_tlu_wsr_data_m[19]), .B(exu_n16302), .Y(exu_n24552));
INVX1 exu_U23033(.A(exu_n24552), .Y(exu_n7008));
AND2X1 exu_U23034(.A(exu_tlu_wsr_data_m[18]), .B(exu_n16302), .Y(exu_n24556));
INVX1 exu_U23035(.A(exu_n24556), .Y(exu_n7009));
AND2X1 exu_U23036(.A(exu_tlu_wsr_data_m[17]), .B(exu_n16302), .Y(exu_n24560));
INVX1 exu_U23037(.A(exu_n24560), .Y(exu_n7010));
AND2X1 exu_U23038(.A(exu_tlu_wsr_data_m[16]), .B(exu_n16302), .Y(exu_n24564));
INVX1 exu_U23039(.A(exu_n24564), .Y(exu_n7011));
AND2X1 exu_U23040(.A(exu_tlu_wsr_data_m[15]), .B(exu_n16302), .Y(exu_n24568));
INVX1 exu_U23041(.A(exu_n24568), .Y(exu_n7012));
AND2X1 exu_U23042(.A(exu_tlu_wsr_data_m[14]), .B(exu_n16302), .Y(exu_n24572));
INVX1 exu_U23043(.A(exu_n24572), .Y(exu_n7013));
AND2X1 exu_U23044(.A(exu_tlu_wsr_data_m[13]), .B(exu_n16302), .Y(exu_n24576));
INVX1 exu_U23045(.A(exu_n24576), .Y(exu_n7014));
AND2X1 exu_U23046(.A(exu_tlu_wsr_data_m[12]), .B(exu_n16302), .Y(exu_n24580));
INVX1 exu_U23047(.A(exu_n24580), .Y(exu_n7015));
AND2X1 exu_U23048(.A(exu_tlu_wsr_data_m[11]), .B(exu_n16302), .Y(exu_n24584));
INVX1 exu_U23049(.A(exu_n24584), .Y(exu_n7016));
AND2X1 exu_U23050(.A(exu_tlu_wsr_data_m[10]), .B(exu_n16302), .Y(exu_n24588));
INVX1 exu_U23051(.A(exu_n24588), .Y(exu_n7017));
AND2X1 exu_U23052(.A(exu_tlu_wsr_data_m[0]), .B(exu_n16302), .Y(exu_n24592));
INVX1 exu_U23053(.A(exu_n24592), .Y(exu_n7018));
AND2X1 exu_U23054(.A(exu_n16306), .B(alu_byp_rd_data_e[9]), .Y(exu_n24596));
INVX1 exu_U23055(.A(exu_n24596), .Y(exu_n7019));
AND2X1 exu_U23056(.A(exu_n16303), .B(bypass_rcc_data_btwn_mux[9]), .Y(exu_n24598));
INVX1 exu_U23057(.A(exu_n24598), .Y(exu_n7020));
AND2X1 exu_U23058(.A(alu_byp_rd_data_e[8]), .B(exu_n16306), .Y(exu_n24602));
INVX1 exu_U23059(.A(exu_n24602), .Y(exu_n7021));
AND2X1 exu_U23060(.A(bypass_rcc_data_btwn_mux[8]), .B(exu_n16303), .Y(exu_n24604));
INVX1 exu_U23061(.A(exu_n24604), .Y(exu_n7022));
AND2X1 exu_U23062(.A(alu_byp_rd_data_e[7]), .B(exu_n16306), .Y(exu_n24608));
INVX1 exu_U23063(.A(exu_n24608), .Y(exu_n7023));
AND2X1 exu_U23064(.A(bypass_rcc_data_btwn_mux[7]), .B(exu_n16303), .Y(exu_n24610));
INVX1 exu_U23065(.A(exu_n24610), .Y(exu_n7024));
AND2X1 exu_U23066(.A(alu_byp_rd_data_e[6]), .B(exu_n16306), .Y(exu_n24614));
INVX1 exu_U23067(.A(exu_n24614), .Y(exu_n7025));
AND2X1 exu_U23068(.A(bypass_rcc_data_btwn_mux[6]), .B(exu_n16303), .Y(exu_n24616));
INVX1 exu_U23069(.A(exu_n24616), .Y(exu_n7026));
AND2X1 exu_U23070(.A(alu_byp_rd_data_e[63]), .B(exu_n16306), .Y(exu_n24620));
INVX1 exu_U23071(.A(exu_n24620), .Y(exu_n7027));
AND2X1 exu_U23072(.A(bypass_rcc_data_btwn_mux[63]), .B(exu_n16303), .Y(exu_n24622));
INVX1 exu_U23073(.A(exu_n24622), .Y(exu_n7028));
AND2X1 exu_U23074(.A(alu_byp_rd_data_e[62]), .B(exu_n16306), .Y(exu_n24626));
INVX1 exu_U23075(.A(exu_n24626), .Y(exu_n7029));
AND2X1 exu_U23076(.A(bypass_rcc_data_btwn_mux[62]), .B(exu_n16303), .Y(exu_n24628));
INVX1 exu_U23077(.A(exu_n24628), .Y(exu_n7030));
AND2X1 exu_U23078(.A(alu_byp_rd_data_e[61]), .B(exu_n16306), .Y(exu_n24632));
INVX1 exu_U23079(.A(exu_n24632), .Y(exu_n7031));
AND2X1 exu_U23080(.A(bypass_rcc_data_btwn_mux[61]), .B(exu_n16303), .Y(exu_n24634));
INVX1 exu_U23081(.A(exu_n24634), .Y(exu_n7032));
AND2X1 exu_U23082(.A(alu_byp_rd_data_e[60]), .B(exu_n16306), .Y(exu_n24638));
INVX1 exu_U23083(.A(exu_n24638), .Y(exu_n7033));
AND2X1 exu_U23084(.A(bypass_rcc_data_btwn_mux[60]), .B(exu_n16303), .Y(exu_n24640));
INVX1 exu_U23085(.A(exu_n24640), .Y(exu_n7034));
AND2X1 exu_U23086(.A(alu_byp_rd_data_e[5]), .B(exu_n16306), .Y(exu_n24644));
INVX1 exu_U23087(.A(exu_n24644), .Y(exu_n7035));
AND2X1 exu_U23088(.A(bypass_rcc_data_btwn_mux[5]), .B(exu_n16303), .Y(exu_n24646));
INVX1 exu_U23089(.A(exu_n24646), .Y(exu_n7036));
AND2X1 exu_U23090(.A(alu_byp_rd_data_e[59]), .B(exu_n16306), .Y(exu_n24650));
INVX1 exu_U23091(.A(exu_n24650), .Y(exu_n7037));
AND2X1 exu_U23092(.A(bypass_rcc_data_btwn_mux[59]), .B(exu_n16303), .Y(exu_n24652));
INVX1 exu_U23093(.A(exu_n24652), .Y(exu_n7038));
AND2X1 exu_U23094(.A(alu_byp_rd_data_e[58]), .B(exu_n16306), .Y(exu_n24656));
INVX1 exu_U23095(.A(exu_n24656), .Y(exu_n7039));
AND2X1 exu_U23096(.A(bypass_rcc_data_btwn_mux[58]), .B(exu_n16303), .Y(exu_n24658));
INVX1 exu_U23097(.A(exu_n24658), .Y(exu_n7040));
AND2X1 exu_U23098(.A(alu_byp_rd_data_e[57]), .B(exu_n16306), .Y(exu_n24662));
INVX1 exu_U23099(.A(exu_n24662), .Y(exu_n7041));
AND2X1 exu_U23100(.A(bypass_rcc_data_btwn_mux[57]), .B(exu_n16303), .Y(exu_n24664));
INVX1 exu_U23101(.A(exu_n24664), .Y(exu_n7042));
AND2X1 exu_U23102(.A(alu_byp_rd_data_e[56]), .B(exu_n16306), .Y(exu_n24668));
INVX1 exu_U23103(.A(exu_n24668), .Y(exu_n7043));
AND2X1 exu_U23104(.A(bypass_rcc_data_btwn_mux[56]), .B(exu_n16303), .Y(exu_n24670));
INVX1 exu_U23105(.A(exu_n24670), .Y(exu_n7044));
AND2X1 exu_U23106(.A(alu_byp_rd_data_e[55]), .B(exu_n16306), .Y(exu_n24674));
INVX1 exu_U23107(.A(exu_n24674), .Y(exu_n7045));
AND2X1 exu_U23108(.A(bypass_rcc_data_btwn_mux[55]), .B(exu_n16303), .Y(exu_n24676));
INVX1 exu_U23109(.A(exu_n24676), .Y(exu_n7046));
AND2X1 exu_U23110(.A(alu_byp_rd_data_e[54]), .B(exu_n16306), .Y(exu_n24680));
INVX1 exu_U23111(.A(exu_n24680), .Y(exu_n7047));
AND2X1 exu_U23112(.A(bypass_rcc_data_btwn_mux[54]), .B(exu_n16303), .Y(exu_n24682));
INVX1 exu_U23113(.A(exu_n24682), .Y(exu_n7048));
AND2X1 exu_U23114(.A(alu_byp_rd_data_e[53]), .B(exu_n16306), .Y(exu_n24686));
INVX1 exu_U23115(.A(exu_n24686), .Y(exu_n7049));
AND2X1 exu_U23116(.A(bypass_rcc_data_btwn_mux[53]), .B(exu_n16303), .Y(exu_n24688));
INVX1 exu_U23117(.A(exu_n24688), .Y(exu_n7050));
AND2X1 exu_U23118(.A(alu_byp_rd_data_e[52]), .B(exu_n16306), .Y(exu_n24692));
INVX1 exu_U23119(.A(exu_n24692), .Y(exu_n7051));
AND2X1 exu_U23120(.A(bypass_rcc_data_btwn_mux[52]), .B(exu_n16303), .Y(exu_n24694));
INVX1 exu_U23121(.A(exu_n24694), .Y(exu_n7052));
AND2X1 exu_U23122(.A(alu_byp_rd_data_e[51]), .B(exu_n16306), .Y(exu_n24698));
INVX1 exu_U23123(.A(exu_n24698), .Y(exu_n7053));
AND2X1 exu_U23124(.A(bypass_rcc_data_btwn_mux[51]), .B(exu_n16303), .Y(exu_n24700));
INVX1 exu_U23125(.A(exu_n24700), .Y(exu_n7054));
AND2X1 exu_U23126(.A(alu_byp_rd_data_e[50]), .B(exu_n16306), .Y(exu_n24704));
INVX1 exu_U23127(.A(exu_n24704), .Y(exu_n7055));
AND2X1 exu_U23128(.A(bypass_rcc_data_btwn_mux[50]), .B(exu_n16303), .Y(exu_n24706));
INVX1 exu_U23129(.A(exu_n24706), .Y(exu_n7056));
AND2X1 exu_U23130(.A(alu_byp_rd_data_e[4]), .B(exu_n16306), .Y(exu_n24710));
INVX1 exu_U23131(.A(exu_n24710), .Y(exu_n7057));
AND2X1 exu_U23132(.A(bypass_rcc_data_btwn_mux[4]), .B(exu_n16303), .Y(exu_n24712));
INVX1 exu_U23133(.A(exu_n24712), .Y(exu_n7058));
AND2X1 exu_U23134(.A(alu_byp_rd_data_e[49]), .B(exu_n16306), .Y(exu_n24716));
INVX1 exu_U23135(.A(exu_n24716), .Y(exu_n7059));
AND2X1 exu_U23136(.A(bypass_rcc_data_btwn_mux[49]), .B(exu_n16303), .Y(exu_n24718));
INVX1 exu_U23137(.A(exu_n24718), .Y(exu_n7060));
AND2X1 exu_U23138(.A(alu_byp_rd_data_e[48]), .B(exu_n16306), .Y(exu_n24722));
INVX1 exu_U23139(.A(exu_n24722), .Y(exu_n7061));
AND2X1 exu_U23140(.A(bypass_rcc_data_btwn_mux[48]), .B(exu_n16303), .Y(exu_n24724));
INVX1 exu_U23141(.A(exu_n24724), .Y(exu_n7062));
AND2X1 exu_U23142(.A(alu_byp_rd_data_e[47]), .B(exu_n16306), .Y(exu_n24728));
INVX1 exu_U23143(.A(exu_n24728), .Y(exu_n7063));
AND2X1 exu_U23144(.A(bypass_rcc_data_btwn_mux[47]), .B(exu_n16303), .Y(exu_n24730));
INVX1 exu_U23145(.A(exu_n24730), .Y(exu_n7064));
AND2X1 exu_U23146(.A(alu_byp_rd_data_e[46]), .B(exu_n16306), .Y(exu_n24734));
INVX1 exu_U23147(.A(exu_n24734), .Y(exu_n7065));
AND2X1 exu_U23148(.A(bypass_rcc_data_btwn_mux[46]), .B(exu_n16303), .Y(exu_n24736));
INVX1 exu_U23149(.A(exu_n24736), .Y(exu_n7066));
AND2X1 exu_U23150(.A(alu_byp_rd_data_e[45]), .B(exu_n16306), .Y(exu_n24740));
INVX1 exu_U23151(.A(exu_n24740), .Y(exu_n7067));
AND2X1 exu_U23152(.A(bypass_rcc_data_btwn_mux[45]), .B(exu_n16303), .Y(exu_n24742));
INVX1 exu_U23153(.A(exu_n24742), .Y(exu_n7068));
AND2X1 exu_U23154(.A(alu_byp_rd_data_e[44]), .B(exu_n16306), .Y(exu_n24746));
INVX1 exu_U23155(.A(exu_n24746), .Y(exu_n7069));
AND2X1 exu_U23156(.A(bypass_rcc_data_btwn_mux[44]), .B(exu_n16303), .Y(exu_n24748));
INVX1 exu_U23157(.A(exu_n24748), .Y(exu_n7070));
AND2X1 exu_U23158(.A(alu_byp_rd_data_e[43]), .B(exu_n16306), .Y(exu_n24752));
INVX1 exu_U23159(.A(exu_n24752), .Y(exu_n7071));
AND2X1 exu_U23160(.A(bypass_rcc_data_btwn_mux[43]), .B(exu_n16303), .Y(exu_n24754));
INVX1 exu_U23161(.A(exu_n24754), .Y(exu_n7072));
AND2X1 exu_U23162(.A(alu_byp_rd_data_e[42]), .B(exu_n16306), .Y(exu_n24758));
INVX1 exu_U23163(.A(exu_n24758), .Y(exu_n7073));
AND2X1 exu_U23164(.A(bypass_rcc_data_btwn_mux[42]), .B(exu_n16303), .Y(exu_n24760));
INVX1 exu_U23165(.A(exu_n24760), .Y(exu_n7074));
AND2X1 exu_U23166(.A(alu_byp_rd_data_e[41]), .B(exu_n16306), .Y(exu_n24764));
INVX1 exu_U23167(.A(exu_n24764), .Y(exu_n7075));
AND2X1 exu_U23168(.A(bypass_rcc_data_btwn_mux[41]), .B(exu_n16303), .Y(exu_n24766));
INVX1 exu_U23169(.A(exu_n24766), .Y(exu_n7076));
AND2X1 exu_U23170(.A(alu_byp_rd_data_e[40]), .B(exu_n16306), .Y(exu_n24770));
INVX1 exu_U23171(.A(exu_n24770), .Y(exu_n7077));
AND2X1 exu_U23172(.A(bypass_rcc_data_btwn_mux[40]), .B(exu_n16303), .Y(exu_n24772));
INVX1 exu_U23173(.A(exu_n24772), .Y(exu_n7078));
AND2X1 exu_U23174(.A(alu_byp_rd_data_e[3]), .B(exu_n16306), .Y(exu_n24776));
INVX1 exu_U23175(.A(exu_n24776), .Y(exu_n7079));
AND2X1 exu_U23176(.A(bypass_rcc_data_btwn_mux[3]), .B(exu_n16303), .Y(exu_n24778));
INVX1 exu_U23177(.A(exu_n24778), .Y(exu_n7080));
AND2X1 exu_U23178(.A(alu_byp_rd_data_e[39]), .B(exu_n16306), .Y(exu_n24782));
INVX1 exu_U23179(.A(exu_n24782), .Y(exu_n7081));
AND2X1 exu_U23180(.A(bypass_rcc_data_btwn_mux[39]), .B(exu_n16303), .Y(exu_n24784));
INVX1 exu_U23181(.A(exu_n24784), .Y(exu_n7082));
AND2X1 exu_U23182(.A(alu_byp_rd_data_e[38]), .B(exu_n16306), .Y(exu_n24788));
INVX1 exu_U23183(.A(exu_n24788), .Y(exu_n7083));
AND2X1 exu_U23184(.A(bypass_rcc_data_btwn_mux[38]), .B(exu_n16303), .Y(exu_n24790));
INVX1 exu_U23185(.A(exu_n24790), .Y(exu_n7084));
AND2X1 exu_U23186(.A(alu_byp_rd_data_e[37]), .B(exu_n16306), .Y(exu_n24794));
INVX1 exu_U23187(.A(exu_n24794), .Y(exu_n7085));
AND2X1 exu_U23188(.A(bypass_rcc_data_btwn_mux[37]), .B(exu_n16303), .Y(exu_n24796));
INVX1 exu_U23189(.A(exu_n24796), .Y(exu_n7086));
AND2X1 exu_U23190(.A(alu_byp_rd_data_e[36]), .B(exu_n16306), .Y(exu_n24800));
INVX1 exu_U23191(.A(exu_n24800), .Y(exu_n7087));
AND2X1 exu_U23192(.A(bypass_rcc_data_btwn_mux[36]), .B(exu_n16303), .Y(exu_n24802));
INVX1 exu_U23193(.A(exu_n24802), .Y(exu_n7088));
AND2X1 exu_U23194(.A(alu_byp_rd_data_e[35]), .B(exu_n16306), .Y(exu_n24806));
INVX1 exu_U23195(.A(exu_n24806), .Y(exu_n7089));
AND2X1 exu_U23196(.A(bypass_rcc_data_btwn_mux[35]), .B(exu_n16303), .Y(exu_n24808));
INVX1 exu_U23197(.A(exu_n24808), .Y(exu_n7090));
AND2X1 exu_U23198(.A(alu_byp_rd_data_e[34]), .B(exu_n16306), .Y(exu_n24812));
INVX1 exu_U23199(.A(exu_n24812), .Y(exu_n7091));
AND2X1 exu_U23200(.A(bypass_rcc_data_btwn_mux[34]), .B(exu_n16303), .Y(exu_n24814));
INVX1 exu_U23201(.A(exu_n24814), .Y(exu_n7092));
AND2X1 exu_U23202(.A(alu_byp_rd_data_e[33]), .B(exu_n16306), .Y(exu_n24818));
INVX1 exu_U23203(.A(exu_n24818), .Y(exu_n7093));
AND2X1 exu_U23204(.A(bypass_rcc_data_btwn_mux[33]), .B(exu_n16303), .Y(exu_n24820));
INVX1 exu_U23205(.A(exu_n24820), .Y(exu_n7094));
AND2X1 exu_U23206(.A(alu_byp_rd_data_e[32]), .B(exu_n16306), .Y(exu_n24824));
INVX1 exu_U23207(.A(exu_n24824), .Y(exu_n7095));
AND2X1 exu_U23208(.A(bypass_rcc_data_btwn_mux[32]), .B(exu_n16303), .Y(exu_n24826));
INVX1 exu_U23209(.A(exu_n24826), .Y(exu_n7096));
AND2X1 exu_U23210(.A(alu_byp_rd_data_e[31]), .B(exu_n16306), .Y(exu_n24830));
INVX1 exu_U23211(.A(exu_n24830), .Y(exu_n7097));
AND2X1 exu_U23212(.A(bypass_rcc_data_btwn_mux[31]), .B(exu_n16303), .Y(exu_n24832));
INVX1 exu_U23213(.A(exu_n24832), .Y(exu_n7098));
AND2X1 exu_U23214(.A(alu_byp_rd_data_e[30]), .B(exu_n16306), .Y(exu_n24836));
INVX1 exu_U23215(.A(exu_n24836), .Y(exu_n7099));
AND2X1 exu_U23216(.A(bypass_rcc_data_btwn_mux[30]), .B(exu_n16303), .Y(exu_n24838));
INVX1 exu_U23217(.A(exu_n24838), .Y(exu_n7100));
AND2X1 exu_U23218(.A(alu_byp_rd_data_e[2]), .B(exu_n16306), .Y(exu_n24842));
INVX1 exu_U23219(.A(exu_n24842), .Y(exu_n7101));
AND2X1 exu_U23220(.A(bypass_rcc_data_btwn_mux[2]), .B(exu_n16303), .Y(exu_n24844));
INVX1 exu_U23221(.A(exu_n24844), .Y(exu_n7102));
AND2X1 exu_U23222(.A(alu_byp_rd_data_e[29]), .B(exu_n16306), .Y(exu_n24848));
INVX1 exu_U23223(.A(exu_n24848), .Y(exu_n7103));
AND2X1 exu_U23224(.A(bypass_rcc_data_btwn_mux[29]), .B(exu_n16303), .Y(exu_n24850));
INVX1 exu_U23225(.A(exu_n24850), .Y(exu_n7104));
AND2X1 exu_U23226(.A(alu_byp_rd_data_e[28]), .B(exu_n16306), .Y(exu_n24854));
INVX1 exu_U23227(.A(exu_n24854), .Y(exu_n7105));
AND2X1 exu_U23228(.A(bypass_rcc_data_btwn_mux[28]), .B(exu_n16303), .Y(exu_n24856));
INVX1 exu_U23229(.A(exu_n24856), .Y(exu_n7106));
AND2X1 exu_U23230(.A(alu_byp_rd_data_e[27]), .B(exu_n16306), .Y(exu_n24860));
INVX1 exu_U23231(.A(exu_n24860), .Y(exu_n7107));
AND2X1 exu_U23232(.A(bypass_rcc_data_btwn_mux[27]), .B(exu_n16303), .Y(exu_n24862));
INVX1 exu_U23233(.A(exu_n24862), .Y(exu_n7108));
AND2X1 exu_U23234(.A(alu_byp_rd_data_e[26]), .B(exu_n16306), .Y(exu_n24866));
INVX1 exu_U23235(.A(exu_n24866), .Y(exu_n7109));
AND2X1 exu_U23236(.A(bypass_rcc_data_btwn_mux[26]), .B(exu_n16303), .Y(exu_n24868));
INVX1 exu_U23237(.A(exu_n24868), .Y(exu_n7110));
AND2X1 exu_U23238(.A(alu_byp_rd_data_e[25]), .B(exu_n16306), .Y(exu_n24872));
INVX1 exu_U23239(.A(exu_n24872), .Y(exu_n7111));
AND2X1 exu_U23240(.A(bypass_rcc_data_btwn_mux[25]), .B(exu_n16303), .Y(exu_n24874));
INVX1 exu_U23241(.A(exu_n24874), .Y(exu_n7112));
AND2X1 exu_U23242(.A(alu_byp_rd_data_e[24]), .B(exu_n16306), .Y(exu_n24878));
INVX1 exu_U23243(.A(exu_n24878), .Y(exu_n7113));
AND2X1 exu_U23244(.A(bypass_rcc_data_btwn_mux[24]), .B(exu_n16303), .Y(exu_n24880));
INVX1 exu_U23245(.A(exu_n24880), .Y(exu_n7114));
AND2X1 exu_U23246(.A(alu_byp_rd_data_e[23]), .B(exu_n16306), .Y(exu_n24884));
INVX1 exu_U23247(.A(exu_n24884), .Y(exu_n7115));
AND2X1 exu_U23248(.A(bypass_rcc_data_btwn_mux[23]), .B(exu_n16303), .Y(exu_n24886));
INVX1 exu_U23249(.A(exu_n24886), .Y(exu_n7116));
AND2X1 exu_U23250(.A(alu_byp_rd_data_e[22]), .B(exu_n16306), .Y(exu_n24890));
INVX1 exu_U23251(.A(exu_n24890), .Y(exu_n7117));
AND2X1 exu_U23252(.A(bypass_rcc_data_btwn_mux[22]), .B(exu_n16303), .Y(exu_n24892));
INVX1 exu_U23253(.A(exu_n24892), .Y(exu_n7118));
AND2X1 exu_U23254(.A(alu_byp_rd_data_e[21]), .B(exu_n16306), .Y(exu_n24896));
INVX1 exu_U23255(.A(exu_n24896), .Y(exu_n7119));
AND2X1 exu_U23256(.A(bypass_rcc_data_btwn_mux[21]), .B(exu_n16303), .Y(exu_n24898));
INVX1 exu_U23257(.A(exu_n24898), .Y(exu_n7120));
AND2X1 exu_U23258(.A(alu_byp_rd_data_e[20]), .B(exu_n16306), .Y(exu_n24902));
INVX1 exu_U23259(.A(exu_n24902), .Y(exu_n7121));
AND2X1 exu_U23260(.A(bypass_rcc_data_btwn_mux[20]), .B(exu_n16303), .Y(exu_n24904));
INVX1 exu_U23261(.A(exu_n24904), .Y(exu_n7122));
AND2X1 exu_U23262(.A(alu_byp_rd_data_e[1]), .B(exu_n16306), .Y(exu_n24908));
INVX1 exu_U23263(.A(exu_n24908), .Y(exu_n7123));
AND2X1 exu_U23264(.A(bypass_rcc_data_btwn_mux[1]), .B(exu_n16303), .Y(exu_n24910));
INVX1 exu_U23265(.A(exu_n24910), .Y(exu_n7124));
AND2X1 exu_U23266(.A(alu_byp_rd_data_e[19]), .B(exu_n16306), .Y(exu_n24914));
INVX1 exu_U23267(.A(exu_n24914), .Y(exu_n7125));
AND2X1 exu_U23268(.A(bypass_rcc_data_btwn_mux[19]), .B(exu_n16303), .Y(exu_n24916));
INVX1 exu_U23269(.A(exu_n24916), .Y(exu_n7126));
AND2X1 exu_U23270(.A(alu_byp_rd_data_e[18]), .B(exu_n16306), .Y(exu_n24920));
INVX1 exu_U23271(.A(exu_n24920), .Y(exu_n7127));
AND2X1 exu_U23272(.A(bypass_rcc_data_btwn_mux[18]), .B(exu_n16303), .Y(exu_n24922));
INVX1 exu_U23273(.A(exu_n24922), .Y(exu_n7128));
AND2X1 exu_U23274(.A(alu_byp_rd_data_e[17]), .B(exu_n16306), .Y(exu_n24926));
INVX1 exu_U23275(.A(exu_n24926), .Y(exu_n7129));
AND2X1 exu_U23276(.A(bypass_rcc_data_btwn_mux[17]), .B(exu_n16303), .Y(exu_n24928));
INVX1 exu_U23277(.A(exu_n24928), .Y(exu_n7130));
AND2X1 exu_U23278(.A(alu_byp_rd_data_e[16]), .B(exu_n16306), .Y(exu_n24932));
INVX1 exu_U23279(.A(exu_n24932), .Y(exu_n7131));
AND2X1 exu_U23280(.A(bypass_rcc_data_btwn_mux[16]), .B(exu_n16303), .Y(exu_n24934));
INVX1 exu_U23281(.A(exu_n24934), .Y(exu_n7132));
AND2X1 exu_U23282(.A(alu_byp_rd_data_e[15]), .B(exu_n16306), .Y(exu_n24938));
INVX1 exu_U23283(.A(exu_n24938), .Y(exu_n7133));
AND2X1 exu_U23284(.A(bypass_rcc_data_btwn_mux[15]), .B(exu_n16303), .Y(exu_n24940));
INVX1 exu_U23285(.A(exu_n24940), .Y(exu_n7134));
AND2X1 exu_U23286(.A(alu_byp_rd_data_e[14]), .B(exu_n16306), .Y(exu_n24944));
INVX1 exu_U23287(.A(exu_n24944), .Y(exu_n7135));
AND2X1 exu_U23288(.A(bypass_rcc_data_btwn_mux[14]), .B(exu_n16303), .Y(exu_n24946));
INVX1 exu_U23289(.A(exu_n24946), .Y(exu_n7136));
AND2X1 exu_U23290(.A(alu_byp_rd_data_e[13]), .B(exu_n16306), .Y(exu_n24950));
INVX1 exu_U23291(.A(exu_n24950), .Y(exu_n7137));
AND2X1 exu_U23292(.A(bypass_rcc_data_btwn_mux[13]), .B(exu_n16303), .Y(exu_n24952));
INVX1 exu_U23293(.A(exu_n24952), .Y(exu_n7138));
AND2X1 exu_U23294(.A(alu_byp_rd_data_e[12]), .B(exu_n16306), .Y(exu_n24956));
INVX1 exu_U23295(.A(exu_n24956), .Y(exu_n7139));
AND2X1 exu_U23296(.A(bypass_rcc_data_btwn_mux[12]), .B(exu_n16303), .Y(exu_n24958));
INVX1 exu_U23297(.A(exu_n24958), .Y(exu_n7140));
AND2X1 exu_U23298(.A(alu_byp_rd_data_e[11]), .B(exu_n16306), .Y(exu_n24962));
INVX1 exu_U23299(.A(exu_n24962), .Y(exu_n7141));
AND2X1 exu_U23300(.A(bypass_rcc_data_btwn_mux[11]), .B(exu_n16303), .Y(exu_n24964));
INVX1 exu_U23301(.A(exu_n24964), .Y(exu_n7142));
AND2X1 exu_U23302(.A(alu_byp_rd_data_e[10]), .B(exu_n16306), .Y(exu_n24968));
INVX1 exu_U23303(.A(exu_n24968), .Y(exu_n7143));
AND2X1 exu_U23304(.A(bypass_rcc_data_btwn_mux[10]), .B(exu_n16303), .Y(exu_n24970));
INVX1 exu_U23305(.A(exu_n24970), .Y(exu_n7144));
AND2X1 exu_U23306(.A(alu_byp_rd_data_e[0]), .B(exu_n16306), .Y(exu_n24974));
INVX1 exu_U23307(.A(exu_n24974), .Y(exu_n7145));
AND2X1 exu_U23308(.A(bypass_rcc_data_btwn_mux[0]), .B(exu_n16303), .Y(exu_n24976));
INVX1 exu_U23309(.A(exu_n24976), .Y(exu_n7146));
AND2X1 exu_U23310(.A(ecl_byplog_rs2_n30), .B(exu_n9999), .Y(exu_n24980));
INVX1 exu_U23311(.A(exu_n24980), .Y(exu_n7147));
AND2X1 exu_U23312(.A(exu_n16294), .B(exu_tlu_wsr_data_m[9]), .Y(exu_n24982));
INVX1 exu_U23313(.A(exu_n24982), .Y(exu_n7148));
AND2X1 exu_U23314(.A(exu_n10994), .B(ecl_byplog_rs2_n30), .Y(exu_n24986));
INVX1 exu_U23315(.A(exu_n24986), .Y(exu_n7149));
AND2X1 exu_U23316(.A(exu_tlu_wsr_data_m[8]), .B(exu_n16294), .Y(exu_n24988));
INVX1 exu_U23317(.A(exu_n24988), .Y(exu_n7150));
AND2X1 exu_U23318(.A(exu_n10995), .B(exu_n15963), .Y(exu_n24992));
INVX1 exu_U23319(.A(exu_n24992), .Y(exu_n7151));
AND2X1 exu_U23320(.A(exu_tlu_wsr_data_m[7]), .B(exu_n16294), .Y(exu_n24994));
INVX1 exu_U23321(.A(exu_n24994), .Y(exu_n7152));
AND2X1 exu_U23322(.A(exu_n10996), .B(ecl_byplog_rs2_n30), .Y(exu_n24998));
INVX1 exu_U23323(.A(exu_n24998), .Y(exu_n7153));
AND2X1 exu_U23324(.A(exu_tlu_wsr_data_m[6]), .B(exu_n16294), .Y(exu_n25000));
INVX1 exu_U23325(.A(exu_n25000), .Y(exu_n7154));
AND2X1 exu_U23326(.A(exu_n10997), .B(ecl_byplog_rs2_n30), .Y(exu_n25003));
INVX1 exu_U23327(.A(exu_n25003), .Y(exu_n7155));
AND2X1 exu_U23328(.A(exu_tlu_wsr_data_m[63]), .B(exu_n16294), .Y(exu_n25005));
INVX1 exu_U23329(.A(exu_n25005), .Y(exu_n7156));
AND2X1 exu_U23330(.A(exu_n10998), .B(ecl_byplog_rs2_n30), .Y(exu_n25008));
INVX1 exu_U23331(.A(exu_n25008), .Y(exu_n7157));
AND2X1 exu_U23332(.A(exu_tlu_wsr_data_m[62]), .B(exu_n16294), .Y(exu_n25010));
INVX1 exu_U23333(.A(exu_n25010), .Y(exu_n7158));
AND2X1 exu_U23334(.A(exu_n10999), .B(exu_n15963), .Y(exu_n25013));
INVX1 exu_U23335(.A(exu_n25013), .Y(exu_n7159));
AND2X1 exu_U23336(.A(exu_tlu_wsr_data_m[61]), .B(exu_n16294), .Y(exu_n25015));
INVX1 exu_U23337(.A(exu_n25015), .Y(exu_n7160));
AND2X1 exu_U23338(.A(exu_n11000), .B(ecl_byplog_rs2_n30), .Y(exu_n25018));
INVX1 exu_U23339(.A(exu_n25018), .Y(exu_n7161));
AND2X1 exu_U23340(.A(exu_tlu_wsr_data_m[60]), .B(exu_n16294), .Y(exu_n25020));
INVX1 exu_U23341(.A(exu_n25020), .Y(exu_n7162));
AND2X1 exu_U23342(.A(exu_n11001), .B(ecl_byplog_rs2_n30), .Y(exu_n25024));
INVX1 exu_U23343(.A(exu_n25024), .Y(exu_n7163));
AND2X1 exu_U23344(.A(exu_tlu_wsr_data_m[5]), .B(exu_n16294), .Y(exu_n25026));
INVX1 exu_U23345(.A(exu_n25026), .Y(exu_n7164));
AND2X1 exu_U23346(.A(exu_n11002), .B(ecl_byplog_rs2_n30), .Y(exu_n25029));
INVX1 exu_U23347(.A(exu_n25029), .Y(exu_n7165));
AND2X1 exu_U23348(.A(exu_tlu_wsr_data_m[59]), .B(exu_n16294), .Y(exu_n25031));
INVX1 exu_U23349(.A(exu_n25031), .Y(exu_n7166));
AND2X1 exu_U23350(.A(exu_n11003), .B(exu_n15963), .Y(exu_n25034));
INVX1 exu_U23351(.A(exu_n25034), .Y(exu_n7167));
AND2X1 exu_U23352(.A(exu_tlu_wsr_data_m[58]), .B(exu_n16294), .Y(exu_n25036));
INVX1 exu_U23353(.A(exu_n25036), .Y(exu_n7168));
AND2X1 exu_U23354(.A(exu_n11004), .B(ecl_byplog_rs2_n30), .Y(exu_n25039));
INVX1 exu_U23355(.A(exu_n25039), .Y(exu_n7169));
AND2X1 exu_U23356(.A(exu_tlu_wsr_data_m[57]), .B(exu_n16294), .Y(exu_n25041));
INVX1 exu_U23357(.A(exu_n25041), .Y(exu_n7170));
AND2X1 exu_U23358(.A(exu_n11005), .B(ecl_byplog_rs2_n30), .Y(exu_n25044));
INVX1 exu_U23359(.A(exu_n25044), .Y(exu_n7171));
AND2X1 exu_U23360(.A(exu_tlu_wsr_data_m[56]), .B(exu_n16294), .Y(exu_n25046));
INVX1 exu_U23361(.A(exu_n25046), .Y(exu_n7172));
AND2X1 exu_U23362(.A(exu_n11006), .B(exu_n15963), .Y(exu_n25049));
INVX1 exu_U23363(.A(exu_n25049), .Y(exu_n7173));
AND2X1 exu_U23364(.A(exu_tlu_wsr_data_m[55]), .B(exu_n16294), .Y(exu_n25051));
INVX1 exu_U23365(.A(exu_n25051), .Y(exu_n7174));
AND2X1 exu_U23366(.A(exu_n11007), .B(ecl_byplog_rs2_n30), .Y(exu_n25054));
INVX1 exu_U23367(.A(exu_n25054), .Y(exu_n7175));
AND2X1 exu_U23368(.A(exu_tlu_wsr_data_m[54]), .B(exu_n16294), .Y(exu_n25056));
INVX1 exu_U23369(.A(exu_n25056), .Y(exu_n7176));
AND2X1 exu_U23370(.A(exu_n11008), .B(ecl_byplog_rs2_n30), .Y(exu_n25059));
INVX1 exu_U23371(.A(exu_n25059), .Y(exu_n7177));
AND2X1 exu_U23372(.A(exu_tlu_wsr_data_m[53]), .B(exu_n16294), .Y(exu_n25061));
INVX1 exu_U23373(.A(exu_n25061), .Y(exu_n7178));
AND2X1 exu_U23374(.A(exu_n11009), .B(ecl_byplog_rs2_n30), .Y(exu_n25064));
INVX1 exu_U23375(.A(exu_n25064), .Y(exu_n7179));
AND2X1 exu_U23376(.A(exu_tlu_wsr_data_m[52]), .B(exu_n16294), .Y(exu_n25066));
INVX1 exu_U23377(.A(exu_n25066), .Y(exu_n7180));
AND2X1 exu_U23378(.A(exu_n11010), .B(exu_n15963), .Y(exu_n25069));
INVX1 exu_U23379(.A(exu_n25069), .Y(exu_n7181));
AND2X1 exu_U23380(.A(exu_tlu_wsr_data_m[51]), .B(exu_n16294), .Y(exu_n25071));
INVX1 exu_U23381(.A(exu_n25071), .Y(exu_n7182));
AND2X1 exu_U23382(.A(exu_n11011), .B(ecl_byplog_rs2_n30), .Y(exu_n25074));
INVX1 exu_U23383(.A(exu_n25074), .Y(exu_n7183));
AND2X1 exu_U23384(.A(exu_tlu_wsr_data_m[50]), .B(exu_n16294), .Y(exu_n25076));
INVX1 exu_U23385(.A(exu_n25076), .Y(exu_n7184));
AND2X1 exu_U23386(.A(exu_n11012), .B(exu_n15963), .Y(exu_n25080));
INVX1 exu_U23387(.A(exu_n25080), .Y(exu_n7185));
AND2X1 exu_U23388(.A(exu_tlu_wsr_data_m[4]), .B(exu_n16294), .Y(exu_n25082));
INVX1 exu_U23389(.A(exu_n25082), .Y(exu_n7186));
AND2X1 exu_U23390(.A(exu_n11013), .B(ecl_byplog_rs2_n30), .Y(exu_n25085));
INVX1 exu_U23391(.A(exu_n25085), .Y(exu_n7187));
AND2X1 exu_U23392(.A(exu_tlu_wsr_data_m[49]), .B(exu_n16294), .Y(exu_n25087));
INVX1 exu_U23393(.A(exu_n25087), .Y(exu_n7188));
AND2X1 exu_U23394(.A(exu_n11014), .B(exu_n15963), .Y(exu_n25090));
INVX1 exu_U23395(.A(exu_n25090), .Y(exu_n7189));
AND2X1 exu_U23396(.A(exu_tlu_wsr_data_m[48]), .B(exu_n16294), .Y(exu_n25092));
INVX1 exu_U23397(.A(exu_n25092), .Y(exu_n7190));
AND2X1 exu_U23398(.A(exu_n11015), .B(exu_n15963), .Y(exu_n25095));
INVX1 exu_U23399(.A(exu_n25095), .Y(exu_n7191));
AND2X1 exu_U23400(.A(exu_tlu_wsr_data_m[47]), .B(exu_n16294), .Y(exu_n25097));
INVX1 exu_U23401(.A(exu_n25097), .Y(exu_n7192));
AND2X1 exu_U23402(.A(exu_n11016), .B(ecl_byplog_rs2_n30), .Y(exu_n25100));
INVX1 exu_U23403(.A(exu_n25100), .Y(exu_n7193));
AND2X1 exu_U23404(.A(exu_tlu_wsr_data_m[46]), .B(exu_n16294), .Y(exu_n25102));
INVX1 exu_U23405(.A(exu_n25102), .Y(exu_n7194));
AND2X1 exu_U23406(.A(exu_n11017), .B(ecl_byplog_rs2_n30), .Y(exu_n25105));
INVX1 exu_U23407(.A(exu_n25105), .Y(exu_n7195));
AND2X1 exu_U23408(.A(exu_tlu_wsr_data_m[45]), .B(exu_n16294), .Y(exu_n25107));
INVX1 exu_U23409(.A(exu_n25107), .Y(exu_n7196));
AND2X1 exu_U23410(.A(exu_n11018), .B(exu_n15963), .Y(exu_n25110));
INVX1 exu_U23411(.A(exu_n25110), .Y(exu_n7197));
AND2X1 exu_U23412(.A(exu_tlu_wsr_data_m[44]), .B(exu_n16294), .Y(exu_n25112));
INVX1 exu_U23413(.A(exu_n25112), .Y(exu_n7198));
AND2X1 exu_U23414(.A(exu_n11019), .B(exu_n15963), .Y(exu_n25115));
INVX1 exu_U23415(.A(exu_n25115), .Y(exu_n7199));
AND2X1 exu_U23416(.A(exu_tlu_wsr_data_m[43]), .B(exu_n16294), .Y(exu_n25117));
INVX1 exu_U23417(.A(exu_n25117), .Y(exu_n7200));
AND2X1 exu_U23418(.A(exu_n11020), .B(exu_n15963), .Y(exu_n25120));
INVX1 exu_U23419(.A(exu_n25120), .Y(exu_n7201));
AND2X1 exu_U23420(.A(exu_tlu_wsr_data_m[42]), .B(exu_n16294), .Y(exu_n25122));
INVX1 exu_U23421(.A(exu_n25122), .Y(exu_n7202));
AND2X1 exu_U23422(.A(exu_n11021), .B(exu_n15963), .Y(exu_n25125));
INVX1 exu_U23423(.A(exu_n25125), .Y(exu_n7203));
AND2X1 exu_U23424(.A(exu_tlu_wsr_data_m[41]), .B(exu_n16294), .Y(exu_n25127));
INVX1 exu_U23425(.A(exu_n25127), .Y(exu_n7204));
AND2X1 exu_U23426(.A(exu_n11022), .B(exu_n15963), .Y(exu_n25130));
INVX1 exu_U23427(.A(exu_n25130), .Y(exu_n7205));
AND2X1 exu_U23428(.A(exu_tlu_wsr_data_m[40]), .B(exu_n16294), .Y(exu_n25132));
INVX1 exu_U23429(.A(exu_n25132), .Y(exu_n7206));
AND2X1 exu_U23430(.A(exu_n11023), .B(exu_n15963), .Y(exu_n25136));
INVX1 exu_U23431(.A(exu_n25136), .Y(exu_n7207));
AND2X1 exu_U23432(.A(exu_tlu_wsr_data_m[3]), .B(exu_n16294), .Y(exu_n25138));
INVX1 exu_U23433(.A(exu_n25138), .Y(exu_n7208));
AND2X1 exu_U23434(.A(exu_n11024), .B(exu_n15963), .Y(exu_n25141));
INVX1 exu_U23435(.A(exu_n25141), .Y(exu_n7209));
AND2X1 exu_U23436(.A(exu_tlu_wsr_data_m[39]), .B(exu_n16294), .Y(exu_n25143));
INVX1 exu_U23437(.A(exu_n25143), .Y(exu_n7210));
AND2X1 exu_U23438(.A(exu_n11025), .B(exu_n15963), .Y(exu_n25146));
INVX1 exu_U23439(.A(exu_n25146), .Y(exu_n7211));
AND2X1 exu_U23440(.A(exu_tlu_wsr_data_m[38]), .B(exu_n16294), .Y(exu_n25148));
INVX1 exu_U23441(.A(exu_n25148), .Y(exu_n7212));
AND2X1 exu_U23442(.A(exu_n11026), .B(exu_n15963), .Y(exu_n25151));
INVX1 exu_U23443(.A(exu_n25151), .Y(exu_n7213));
AND2X1 exu_U23444(.A(exu_tlu_wsr_data_m[37]), .B(exu_n16294), .Y(exu_n25153));
INVX1 exu_U23445(.A(exu_n25153), .Y(exu_n7214));
AND2X1 exu_U23446(.A(exu_n11027), .B(exu_n15963), .Y(exu_n25156));
INVX1 exu_U23447(.A(exu_n25156), .Y(exu_n7215));
AND2X1 exu_U23448(.A(exu_tlu_wsr_data_m[36]), .B(exu_n16294), .Y(exu_n25158));
INVX1 exu_U23449(.A(exu_n25158), .Y(exu_n7216));
AND2X1 exu_U23450(.A(exu_n11028), .B(exu_n15963), .Y(exu_n25161));
INVX1 exu_U23451(.A(exu_n25161), .Y(exu_n7217));
AND2X1 exu_U23452(.A(exu_tlu_wsr_data_m[35]), .B(exu_n16294), .Y(exu_n25163));
INVX1 exu_U23453(.A(exu_n25163), .Y(exu_n7218));
AND2X1 exu_U23454(.A(exu_n11029), .B(exu_n15963), .Y(exu_n25166));
INVX1 exu_U23455(.A(exu_n25166), .Y(exu_n7219));
AND2X1 exu_U23456(.A(exu_tlu_wsr_data_m[34]), .B(exu_n16294), .Y(exu_n25168));
INVX1 exu_U23457(.A(exu_n25168), .Y(exu_n7220));
AND2X1 exu_U23458(.A(exu_n11030), .B(exu_n15963), .Y(exu_n25171));
INVX1 exu_U23459(.A(exu_n25171), .Y(exu_n7221));
AND2X1 exu_U23460(.A(exu_tlu_wsr_data_m[33]), .B(exu_n16294), .Y(exu_n25173));
INVX1 exu_U23461(.A(exu_n25173), .Y(exu_n7222));
AND2X1 exu_U23462(.A(exu_n11031), .B(exu_n15963), .Y(exu_n25176));
INVX1 exu_U23463(.A(exu_n25176), .Y(exu_n7223));
AND2X1 exu_U23464(.A(exu_tlu_wsr_data_m[32]), .B(exu_n16294), .Y(exu_n25178));
INVX1 exu_U23465(.A(exu_n25178), .Y(exu_n7224));
AND2X1 exu_U23466(.A(exu_n11032), .B(exu_n15963), .Y(exu_n25182));
INVX1 exu_U23467(.A(exu_n25182), .Y(exu_n7225));
AND2X1 exu_U23468(.A(exu_tlu_wsr_data_m[31]), .B(exu_n16294), .Y(exu_n25184));
INVX1 exu_U23469(.A(exu_n25184), .Y(exu_n7226));
AND2X1 exu_U23470(.A(exu_n11033), .B(ecl_byplog_rs2_n30), .Y(exu_n25188));
INVX1 exu_U23471(.A(exu_n25188), .Y(exu_n7227));
AND2X1 exu_U23472(.A(exu_tlu_wsr_data_m[30]), .B(exu_n16294), .Y(exu_n25190));
INVX1 exu_U23473(.A(exu_n25190), .Y(exu_n7228));
AND2X1 exu_U23474(.A(exu_n11034), .B(ecl_byplog_rs2_n30), .Y(exu_n25194));
INVX1 exu_U23475(.A(exu_n25194), .Y(exu_n7229));
AND2X1 exu_U23476(.A(exu_tlu_wsr_data_m[2]), .B(exu_n16294), .Y(exu_n25196));
INVX1 exu_U23477(.A(exu_n25196), .Y(exu_n7230));
AND2X1 exu_U23478(.A(exu_n11035), .B(exu_n15963), .Y(exu_n25200));
INVX1 exu_U23479(.A(exu_n25200), .Y(exu_n7231));
AND2X1 exu_U23480(.A(exu_tlu_wsr_data_m[29]), .B(exu_n16294), .Y(exu_n25202));
INVX1 exu_U23481(.A(exu_n25202), .Y(exu_n7232));
AND2X1 exu_U23482(.A(exu_n11036), .B(ecl_byplog_rs2_n30), .Y(exu_n25206));
INVX1 exu_U23483(.A(exu_n25206), .Y(exu_n7233));
AND2X1 exu_U23484(.A(exu_tlu_wsr_data_m[28]), .B(exu_n16294), .Y(exu_n25208));
INVX1 exu_U23485(.A(exu_n25208), .Y(exu_n7234));
AND2X1 exu_U23486(.A(exu_n11037), .B(exu_n15963), .Y(exu_n25212));
INVX1 exu_U23487(.A(exu_n25212), .Y(exu_n7235));
AND2X1 exu_U23488(.A(exu_tlu_wsr_data_m[27]), .B(exu_n16294), .Y(exu_n25214));
INVX1 exu_U23489(.A(exu_n25214), .Y(exu_n7236));
AND2X1 exu_U23490(.A(exu_n11038), .B(exu_n15963), .Y(exu_n25218));
INVX1 exu_U23491(.A(exu_n25218), .Y(exu_n7237));
AND2X1 exu_U23492(.A(exu_tlu_wsr_data_m[26]), .B(exu_n16294), .Y(exu_n25220));
INVX1 exu_U23493(.A(exu_n25220), .Y(exu_n7238));
AND2X1 exu_U23494(.A(exu_n11039), .B(ecl_byplog_rs2_n30), .Y(exu_n25224));
INVX1 exu_U23495(.A(exu_n25224), .Y(exu_n7239));
AND2X1 exu_U23496(.A(exu_tlu_wsr_data_m[25]), .B(exu_n16294), .Y(exu_n25226));
INVX1 exu_U23497(.A(exu_n25226), .Y(exu_n7240));
AND2X1 exu_U23498(.A(exu_n11040), .B(ecl_byplog_rs2_n30), .Y(exu_n25230));
INVX1 exu_U23499(.A(exu_n25230), .Y(exu_n7241));
AND2X1 exu_U23500(.A(exu_tlu_wsr_data_m[24]), .B(exu_n16294), .Y(exu_n25232));
INVX1 exu_U23501(.A(exu_n25232), .Y(exu_n7242));
AND2X1 exu_U23502(.A(exu_n11041), .B(exu_n15963), .Y(exu_n25236));
INVX1 exu_U23503(.A(exu_n25236), .Y(exu_n7243));
AND2X1 exu_U23504(.A(exu_tlu_wsr_data_m[23]), .B(exu_n16294), .Y(exu_n25238));
INVX1 exu_U23505(.A(exu_n25238), .Y(exu_n7244));
AND2X1 exu_U23506(.A(exu_n11042), .B(ecl_byplog_rs2_n30), .Y(exu_n25242));
INVX1 exu_U23507(.A(exu_n25242), .Y(exu_n7245));
AND2X1 exu_U23508(.A(exu_tlu_wsr_data_m[22]), .B(exu_n16294), .Y(exu_n25244));
INVX1 exu_U23509(.A(exu_n25244), .Y(exu_n7246));
AND2X1 exu_U23510(.A(exu_n11043), .B(exu_n15963), .Y(exu_n25248));
INVX1 exu_U23511(.A(exu_n25248), .Y(exu_n7247));
AND2X1 exu_U23512(.A(exu_tlu_wsr_data_m[21]), .B(exu_n16294), .Y(exu_n25250));
INVX1 exu_U23513(.A(exu_n25250), .Y(exu_n7248));
AND2X1 exu_U23514(.A(exu_n11044), .B(exu_n15963), .Y(exu_n25254));
INVX1 exu_U23515(.A(exu_n25254), .Y(exu_n7249));
AND2X1 exu_U23516(.A(exu_tlu_wsr_data_m[20]), .B(exu_n16294), .Y(exu_n25256));
INVX1 exu_U23517(.A(exu_n25256), .Y(exu_n7250));
AND2X1 exu_U23518(.A(exu_n11045), .B(ecl_byplog_rs2_n30), .Y(exu_n25260));
INVX1 exu_U23519(.A(exu_n25260), .Y(exu_n7251));
AND2X1 exu_U23520(.A(exu_tlu_wsr_data_m[1]), .B(exu_n16294), .Y(exu_n25262));
INVX1 exu_U23521(.A(exu_n25262), .Y(exu_n7252));
AND2X1 exu_U23522(.A(exu_n11046), .B(ecl_byplog_rs2_n30), .Y(exu_n25266));
INVX1 exu_U23523(.A(exu_n25266), .Y(exu_n7253));
AND2X1 exu_U23524(.A(exu_tlu_wsr_data_m[19]), .B(exu_n16294), .Y(exu_n25268));
INVX1 exu_U23525(.A(exu_n25268), .Y(exu_n7254));
AND2X1 exu_U23526(.A(exu_n11047), .B(exu_n15963), .Y(exu_n25272));
INVX1 exu_U23527(.A(exu_n25272), .Y(exu_n7255));
AND2X1 exu_U23528(.A(exu_tlu_wsr_data_m[18]), .B(exu_n16294), .Y(exu_n25274));
INVX1 exu_U23529(.A(exu_n25274), .Y(exu_n7256));
AND2X1 exu_U23530(.A(exu_n11048), .B(ecl_byplog_rs2_n30), .Y(exu_n25278));
INVX1 exu_U23531(.A(exu_n25278), .Y(exu_n7257));
AND2X1 exu_U23532(.A(exu_tlu_wsr_data_m[17]), .B(exu_n16294), .Y(exu_n25280));
INVX1 exu_U23533(.A(exu_n25280), .Y(exu_n7258));
AND2X1 exu_U23534(.A(exu_n11049), .B(ecl_byplog_rs2_n30), .Y(exu_n25284));
INVX1 exu_U23535(.A(exu_n25284), .Y(exu_n7259));
AND2X1 exu_U23536(.A(exu_tlu_wsr_data_m[16]), .B(exu_n16294), .Y(exu_n25286));
INVX1 exu_U23537(.A(exu_n25286), .Y(exu_n7260));
AND2X1 exu_U23538(.A(exu_n11050), .B(ecl_byplog_rs2_n30), .Y(exu_n25290));
INVX1 exu_U23539(.A(exu_n25290), .Y(exu_n7261));
AND2X1 exu_U23540(.A(exu_tlu_wsr_data_m[15]), .B(exu_n16294), .Y(exu_n25292));
INVX1 exu_U23541(.A(exu_n25292), .Y(exu_n7262));
AND2X1 exu_U23542(.A(exu_n11051), .B(exu_n15963), .Y(exu_n25296));
INVX1 exu_U23543(.A(exu_n25296), .Y(exu_n7263));
AND2X1 exu_U23544(.A(exu_tlu_wsr_data_m[14]), .B(exu_n16294), .Y(exu_n25298));
INVX1 exu_U23545(.A(exu_n25298), .Y(exu_n7264));
AND2X1 exu_U23546(.A(exu_n11052), .B(ecl_byplog_rs2_n30), .Y(exu_n25302));
INVX1 exu_U23547(.A(exu_n25302), .Y(exu_n7265));
AND2X1 exu_U23548(.A(exu_tlu_wsr_data_m[13]), .B(exu_n16294), .Y(exu_n25304));
INVX1 exu_U23549(.A(exu_n25304), .Y(exu_n7266));
AND2X1 exu_U23550(.A(exu_n11053), .B(exu_n15963), .Y(exu_n25308));
INVX1 exu_U23551(.A(exu_n25308), .Y(exu_n7267));
AND2X1 exu_U23552(.A(exu_tlu_wsr_data_m[12]), .B(exu_n16294), .Y(exu_n25310));
INVX1 exu_U23553(.A(exu_n25310), .Y(exu_n7268));
AND2X1 exu_U23554(.A(exu_n11054), .B(ecl_byplog_rs2_n30), .Y(exu_n25314));
INVX1 exu_U23555(.A(exu_n25314), .Y(exu_n7269));
AND2X1 exu_U23556(.A(exu_tlu_wsr_data_m[11]), .B(exu_n16294), .Y(exu_n25316));
INVX1 exu_U23557(.A(exu_n25316), .Y(exu_n7270));
AND2X1 exu_U23558(.A(exu_n11055), .B(ecl_byplog_rs2_n30), .Y(exu_n25320));
INVX1 exu_U23559(.A(exu_n25320), .Y(exu_n7271));
AND2X1 exu_U23560(.A(exu_tlu_wsr_data_m[10]), .B(exu_n16294), .Y(exu_n25322));
INVX1 exu_U23561(.A(exu_n25322), .Y(exu_n7272));
AND2X1 exu_U23562(.A(exu_n11056), .B(ecl_byplog_rs2_n30), .Y(exu_n25326));
INVX1 exu_U23563(.A(exu_n25326), .Y(exu_n7273));
AND2X1 exu_U23564(.A(exu_tlu_wsr_data_m[0]), .B(exu_n16294), .Y(exu_n25328));
INVX1 exu_U23565(.A(exu_n25328), .Y(exu_n7274));
AND2X1 exu_U23566(.A(exu_n16299), .B(alu_byp_rd_data_e[9]), .Y(exu_n25332));
INVX1 exu_U23567(.A(exu_n25332), .Y(exu_n7275));
AND2X1 exu_U23568(.A(exu_n16295), .B(bypass_rs2_data_btwn_mux[9]), .Y(exu_n25334));
INVX1 exu_U23569(.A(exu_n25334), .Y(exu_n7276));
AND2X1 exu_U23570(.A(alu_byp_rd_data_e[8]), .B(exu_n16299), .Y(exu_n25338));
INVX1 exu_U23571(.A(exu_n25338), .Y(exu_n7277));
AND2X1 exu_U23572(.A(bypass_rs2_data_btwn_mux[8]), .B(exu_n16295), .Y(exu_n25340));
INVX1 exu_U23573(.A(exu_n25340), .Y(exu_n7278));
AND2X1 exu_U23574(.A(alu_byp_rd_data_e[7]), .B(exu_n16299), .Y(exu_n25344));
INVX1 exu_U23575(.A(exu_n25344), .Y(exu_n7279));
AND2X1 exu_U23576(.A(bypass_rs2_data_btwn_mux[7]), .B(exu_n16295), .Y(exu_n25346));
INVX1 exu_U23577(.A(exu_n25346), .Y(exu_n7280));
AND2X1 exu_U23578(.A(alu_byp_rd_data_e[6]), .B(exu_n16299), .Y(exu_n25350));
INVX1 exu_U23579(.A(exu_n25350), .Y(exu_n7281));
AND2X1 exu_U23580(.A(bypass_rs2_data_btwn_mux[6]), .B(exu_n16295), .Y(exu_n25352));
INVX1 exu_U23581(.A(exu_n25352), .Y(exu_n7282));
AND2X1 exu_U23582(.A(alu_byp_rd_data_e[63]), .B(exu_n16299), .Y(exu_n25356));
INVX1 exu_U23583(.A(exu_n25356), .Y(exu_n7283));
AND2X1 exu_U23584(.A(bypass_rs2_data_btwn_mux[63]), .B(exu_n16295), .Y(exu_n25358));
INVX1 exu_U23585(.A(exu_n25358), .Y(exu_n7284));
AND2X1 exu_U23586(.A(alu_byp_rd_data_e[62]), .B(exu_n16299), .Y(exu_n25362));
INVX1 exu_U23587(.A(exu_n25362), .Y(exu_n7285));
AND2X1 exu_U23588(.A(bypass_rs2_data_btwn_mux[62]), .B(exu_n16295), .Y(exu_n25364));
INVX1 exu_U23589(.A(exu_n25364), .Y(exu_n7286));
AND2X1 exu_U23590(.A(alu_byp_rd_data_e[61]), .B(exu_n16299), .Y(exu_n25368));
INVX1 exu_U23591(.A(exu_n25368), .Y(exu_n7287));
AND2X1 exu_U23592(.A(bypass_rs2_data_btwn_mux[61]), .B(exu_n16295), .Y(exu_n25370));
INVX1 exu_U23593(.A(exu_n25370), .Y(exu_n7288));
AND2X1 exu_U23594(.A(alu_byp_rd_data_e[60]), .B(exu_n16299), .Y(exu_n25374));
INVX1 exu_U23595(.A(exu_n25374), .Y(exu_n7289));
AND2X1 exu_U23596(.A(bypass_rs2_data_btwn_mux[60]), .B(exu_n16295), .Y(exu_n25376));
INVX1 exu_U23597(.A(exu_n25376), .Y(exu_n7290));
AND2X1 exu_U23598(.A(alu_byp_rd_data_e[5]), .B(exu_n16299), .Y(exu_n25380));
INVX1 exu_U23599(.A(exu_n25380), .Y(exu_n7291));
AND2X1 exu_U23600(.A(bypass_rs2_data_btwn_mux[5]), .B(exu_n16295), .Y(exu_n25382));
INVX1 exu_U23601(.A(exu_n25382), .Y(exu_n7292));
AND2X1 exu_U23602(.A(alu_byp_rd_data_e[59]), .B(exu_n16299), .Y(exu_n25386));
INVX1 exu_U23603(.A(exu_n25386), .Y(exu_n7293));
AND2X1 exu_U23604(.A(bypass_rs2_data_btwn_mux[59]), .B(exu_n16295), .Y(exu_n25388));
INVX1 exu_U23605(.A(exu_n25388), .Y(exu_n7294));
AND2X1 exu_U23606(.A(alu_byp_rd_data_e[58]), .B(exu_n16299), .Y(exu_n25392));
INVX1 exu_U23607(.A(exu_n25392), .Y(exu_n7295));
AND2X1 exu_U23608(.A(bypass_rs2_data_btwn_mux[58]), .B(exu_n16295), .Y(exu_n25394));
INVX1 exu_U23609(.A(exu_n25394), .Y(exu_n7296));
AND2X1 exu_U23610(.A(alu_byp_rd_data_e[57]), .B(exu_n16299), .Y(exu_n25398));
INVX1 exu_U23611(.A(exu_n25398), .Y(exu_n7297));
AND2X1 exu_U23612(.A(bypass_rs2_data_btwn_mux[57]), .B(exu_n16295), .Y(exu_n25400));
INVX1 exu_U23613(.A(exu_n25400), .Y(exu_n7298));
AND2X1 exu_U23614(.A(alu_byp_rd_data_e[56]), .B(exu_n16299), .Y(exu_n25404));
INVX1 exu_U23615(.A(exu_n25404), .Y(exu_n7299));
AND2X1 exu_U23616(.A(bypass_rs2_data_btwn_mux[56]), .B(exu_n16295), .Y(exu_n25406));
INVX1 exu_U23617(.A(exu_n25406), .Y(exu_n7300));
AND2X1 exu_U23618(.A(alu_byp_rd_data_e[55]), .B(exu_n16299), .Y(exu_n25410));
INVX1 exu_U23619(.A(exu_n25410), .Y(exu_n7301));
AND2X1 exu_U23620(.A(bypass_rs2_data_btwn_mux[55]), .B(exu_n16295), .Y(exu_n25412));
INVX1 exu_U23621(.A(exu_n25412), .Y(exu_n7302));
AND2X1 exu_U23622(.A(alu_byp_rd_data_e[54]), .B(exu_n16299), .Y(exu_n25416));
INVX1 exu_U23623(.A(exu_n25416), .Y(exu_n7303));
AND2X1 exu_U23624(.A(bypass_rs2_data_btwn_mux[54]), .B(exu_n16295), .Y(exu_n25418));
INVX1 exu_U23625(.A(exu_n25418), .Y(exu_n7304));
AND2X1 exu_U23626(.A(alu_byp_rd_data_e[53]), .B(exu_n16299), .Y(exu_n25422));
INVX1 exu_U23627(.A(exu_n25422), .Y(exu_n7305));
AND2X1 exu_U23628(.A(bypass_rs2_data_btwn_mux[53]), .B(exu_n16295), .Y(exu_n25424));
INVX1 exu_U23629(.A(exu_n25424), .Y(exu_n7306));
AND2X1 exu_U23630(.A(alu_byp_rd_data_e[52]), .B(exu_n16299), .Y(exu_n25428));
INVX1 exu_U23631(.A(exu_n25428), .Y(exu_n7307));
AND2X1 exu_U23632(.A(bypass_rs2_data_btwn_mux[52]), .B(exu_n16295), .Y(exu_n25430));
INVX1 exu_U23633(.A(exu_n25430), .Y(exu_n7308));
AND2X1 exu_U23634(.A(alu_byp_rd_data_e[51]), .B(exu_n16299), .Y(exu_n25434));
INVX1 exu_U23635(.A(exu_n25434), .Y(exu_n7309));
AND2X1 exu_U23636(.A(bypass_rs2_data_btwn_mux[51]), .B(exu_n16295), .Y(exu_n25436));
INVX1 exu_U23637(.A(exu_n25436), .Y(exu_n7310));
AND2X1 exu_U23638(.A(alu_byp_rd_data_e[50]), .B(exu_n16299), .Y(exu_n25440));
INVX1 exu_U23639(.A(exu_n25440), .Y(exu_n7311));
AND2X1 exu_U23640(.A(bypass_rs2_data_btwn_mux[50]), .B(exu_n16295), .Y(exu_n25442));
INVX1 exu_U23641(.A(exu_n25442), .Y(exu_n7312));
AND2X1 exu_U23642(.A(alu_byp_rd_data_e[4]), .B(exu_n16299), .Y(exu_n25446));
INVX1 exu_U23643(.A(exu_n25446), .Y(exu_n7313));
AND2X1 exu_U23644(.A(bypass_rs2_data_btwn_mux[4]), .B(exu_n16295), .Y(exu_n25448));
INVX1 exu_U23645(.A(exu_n25448), .Y(exu_n7314));
AND2X1 exu_U23646(.A(alu_byp_rd_data_e[49]), .B(exu_n16299), .Y(exu_n25452));
INVX1 exu_U23647(.A(exu_n25452), .Y(exu_n7315));
AND2X1 exu_U23648(.A(bypass_rs2_data_btwn_mux[49]), .B(exu_n16295), .Y(exu_n25454));
INVX1 exu_U23649(.A(exu_n25454), .Y(exu_n7316));
AND2X1 exu_U23650(.A(alu_byp_rd_data_e[48]), .B(exu_n16299), .Y(exu_n25458));
INVX1 exu_U23651(.A(exu_n25458), .Y(exu_n7317));
AND2X1 exu_U23652(.A(bypass_rs2_data_btwn_mux[48]), .B(exu_n16295), .Y(exu_n25460));
INVX1 exu_U23653(.A(exu_n25460), .Y(exu_n7318));
AND2X1 exu_U23654(.A(alu_byp_rd_data_e[47]), .B(exu_n16299), .Y(exu_n25464));
INVX1 exu_U23655(.A(exu_n25464), .Y(exu_n7319));
AND2X1 exu_U23656(.A(bypass_rs2_data_btwn_mux[47]), .B(exu_n16295), .Y(exu_n25466));
INVX1 exu_U23657(.A(exu_n25466), .Y(exu_n7320));
AND2X1 exu_U23658(.A(alu_byp_rd_data_e[46]), .B(exu_n16299), .Y(exu_n25470));
INVX1 exu_U23659(.A(exu_n25470), .Y(exu_n7321));
AND2X1 exu_U23660(.A(bypass_rs2_data_btwn_mux[46]), .B(exu_n16295), .Y(exu_n25472));
INVX1 exu_U23661(.A(exu_n25472), .Y(exu_n7322));
AND2X1 exu_U23662(.A(alu_byp_rd_data_e[45]), .B(exu_n16299), .Y(exu_n25476));
INVX1 exu_U23663(.A(exu_n25476), .Y(exu_n7323));
AND2X1 exu_U23664(.A(bypass_rs2_data_btwn_mux[45]), .B(exu_n16295), .Y(exu_n25478));
INVX1 exu_U23665(.A(exu_n25478), .Y(exu_n7324));
AND2X1 exu_U23666(.A(alu_byp_rd_data_e[44]), .B(exu_n16299), .Y(exu_n25482));
INVX1 exu_U23667(.A(exu_n25482), .Y(exu_n7325));
AND2X1 exu_U23668(.A(bypass_rs2_data_btwn_mux[44]), .B(exu_n16295), .Y(exu_n25484));
INVX1 exu_U23669(.A(exu_n25484), .Y(exu_n7326));
AND2X1 exu_U23670(.A(alu_byp_rd_data_e[43]), .B(exu_n16299), .Y(exu_n25488));
INVX1 exu_U23671(.A(exu_n25488), .Y(exu_n7327));
AND2X1 exu_U23672(.A(bypass_rs2_data_btwn_mux[43]), .B(exu_n16295), .Y(exu_n25490));
INVX1 exu_U23673(.A(exu_n25490), .Y(exu_n7328));
AND2X1 exu_U23674(.A(alu_byp_rd_data_e[42]), .B(exu_n16299), .Y(exu_n25494));
INVX1 exu_U23675(.A(exu_n25494), .Y(exu_n7329));
AND2X1 exu_U23676(.A(bypass_rs2_data_btwn_mux[42]), .B(exu_n16295), .Y(exu_n25496));
INVX1 exu_U23677(.A(exu_n25496), .Y(exu_n7330));
AND2X1 exu_U23678(.A(alu_byp_rd_data_e[41]), .B(exu_n16299), .Y(exu_n25500));
INVX1 exu_U23679(.A(exu_n25500), .Y(exu_n7331));
AND2X1 exu_U23680(.A(bypass_rs2_data_btwn_mux[41]), .B(exu_n16295), .Y(exu_n25502));
INVX1 exu_U23681(.A(exu_n25502), .Y(exu_n7332));
AND2X1 exu_U23682(.A(alu_byp_rd_data_e[40]), .B(exu_n16299), .Y(exu_n25506));
INVX1 exu_U23683(.A(exu_n25506), .Y(exu_n7333));
AND2X1 exu_U23684(.A(bypass_rs2_data_btwn_mux[40]), .B(exu_n16295), .Y(exu_n25508));
INVX1 exu_U23685(.A(exu_n25508), .Y(exu_n7334));
AND2X1 exu_U23686(.A(alu_byp_rd_data_e[3]), .B(exu_n16299), .Y(exu_n25512));
INVX1 exu_U23687(.A(exu_n25512), .Y(exu_n7335));
AND2X1 exu_U23688(.A(bypass_rs2_data_btwn_mux[3]), .B(exu_n16295), .Y(exu_n25514));
INVX1 exu_U23689(.A(exu_n25514), .Y(exu_n7336));
AND2X1 exu_U23690(.A(alu_byp_rd_data_e[39]), .B(exu_n16299), .Y(exu_n25518));
INVX1 exu_U23691(.A(exu_n25518), .Y(exu_n7337));
AND2X1 exu_U23692(.A(bypass_rs2_data_btwn_mux[39]), .B(exu_n16295), .Y(exu_n25520));
INVX1 exu_U23693(.A(exu_n25520), .Y(exu_n7338));
AND2X1 exu_U23694(.A(alu_byp_rd_data_e[38]), .B(exu_n16299), .Y(exu_n25524));
INVX1 exu_U23695(.A(exu_n25524), .Y(exu_n7339));
AND2X1 exu_U23696(.A(bypass_rs2_data_btwn_mux[38]), .B(exu_n16295), .Y(exu_n25526));
INVX1 exu_U23697(.A(exu_n25526), .Y(exu_n7340));
AND2X1 exu_U23698(.A(alu_byp_rd_data_e[37]), .B(exu_n16299), .Y(exu_n25530));
INVX1 exu_U23699(.A(exu_n25530), .Y(exu_n7341));
AND2X1 exu_U23700(.A(bypass_rs2_data_btwn_mux[37]), .B(exu_n16295), .Y(exu_n25532));
INVX1 exu_U23701(.A(exu_n25532), .Y(exu_n7342));
AND2X1 exu_U23702(.A(alu_byp_rd_data_e[36]), .B(exu_n16299), .Y(exu_n25536));
INVX1 exu_U23703(.A(exu_n25536), .Y(exu_n7343));
AND2X1 exu_U23704(.A(bypass_rs2_data_btwn_mux[36]), .B(exu_n16295), .Y(exu_n25538));
INVX1 exu_U23705(.A(exu_n25538), .Y(exu_n7344));
AND2X1 exu_U23706(.A(alu_byp_rd_data_e[35]), .B(exu_n16299), .Y(exu_n25542));
INVX1 exu_U23707(.A(exu_n25542), .Y(exu_n7345));
AND2X1 exu_U23708(.A(bypass_rs2_data_btwn_mux[35]), .B(exu_n16295), .Y(exu_n25544));
INVX1 exu_U23709(.A(exu_n25544), .Y(exu_n7346));
AND2X1 exu_U23710(.A(alu_byp_rd_data_e[34]), .B(exu_n16299), .Y(exu_n25548));
INVX1 exu_U23711(.A(exu_n25548), .Y(exu_n7347));
AND2X1 exu_U23712(.A(bypass_rs2_data_btwn_mux[34]), .B(exu_n16295), .Y(exu_n25550));
INVX1 exu_U23713(.A(exu_n25550), .Y(exu_n7348));
AND2X1 exu_U23714(.A(alu_byp_rd_data_e[33]), .B(exu_n16299), .Y(exu_n25554));
INVX1 exu_U23715(.A(exu_n25554), .Y(exu_n7349));
AND2X1 exu_U23716(.A(bypass_rs2_data_btwn_mux[33]), .B(exu_n16295), .Y(exu_n25556));
INVX1 exu_U23717(.A(exu_n25556), .Y(exu_n7350));
AND2X1 exu_U23718(.A(alu_byp_rd_data_e[32]), .B(exu_n16299), .Y(exu_n25560));
INVX1 exu_U23719(.A(exu_n25560), .Y(exu_n7351));
AND2X1 exu_U23720(.A(bypass_rs2_data_btwn_mux[32]), .B(exu_n16295), .Y(exu_n25562));
INVX1 exu_U23721(.A(exu_n25562), .Y(exu_n7352));
AND2X1 exu_U23722(.A(alu_byp_rd_data_e[31]), .B(exu_n16299), .Y(exu_n25566));
INVX1 exu_U23723(.A(exu_n25566), .Y(exu_n7353));
AND2X1 exu_U23724(.A(bypass_rs2_data_btwn_mux[31]), .B(exu_n16295), .Y(exu_n25568));
INVX1 exu_U23725(.A(exu_n25568), .Y(exu_n7354));
AND2X1 exu_U23726(.A(alu_byp_rd_data_e[30]), .B(exu_n16299), .Y(exu_n25572));
INVX1 exu_U23727(.A(exu_n25572), .Y(exu_n7355));
AND2X1 exu_U23728(.A(bypass_rs2_data_btwn_mux[30]), .B(exu_n16295), .Y(exu_n25574));
INVX1 exu_U23729(.A(exu_n25574), .Y(exu_n7356));
AND2X1 exu_U23730(.A(alu_byp_rd_data_e[2]), .B(exu_n16299), .Y(exu_n25578));
INVX1 exu_U23731(.A(exu_n25578), .Y(exu_n7357));
AND2X1 exu_U23732(.A(bypass_rs2_data_btwn_mux[2]), .B(exu_n16295), .Y(exu_n25580));
INVX1 exu_U23733(.A(exu_n25580), .Y(exu_n7358));
AND2X1 exu_U23734(.A(alu_byp_rd_data_e[29]), .B(exu_n16299), .Y(exu_n25584));
INVX1 exu_U23735(.A(exu_n25584), .Y(exu_n7359));
AND2X1 exu_U23736(.A(bypass_rs2_data_btwn_mux[29]), .B(exu_n16295), .Y(exu_n25586));
INVX1 exu_U23737(.A(exu_n25586), .Y(exu_n7360));
AND2X1 exu_U23738(.A(alu_byp_rd_data_e[28]), .B(exu_n16299), .Y(exu_n25590));
INVX1 exu_U23739(.A(exu_n25590), .Y(exu_n7361));
AND2X1 exu_U23740(.A(bypass_rs2_data_btwn_mux[28]), .B(exu_n16295), .Y(exu_n25592));
INVX1 exu_U23741(.A(exu_n25592), .Y(exu_n7362));
AND2X1 exu_U23742(.A(alu_byp_rd_data_e[27]), .B(exu_n16299), .Y(exu_n25596));
INVX1 exu_U23743(.A(exu_n25596), .Y(exu_n7363));
AND2X1 exu_U23744(.A(bypass_rs2_data_btwn_mux[27]), .B(exu_n16295), .Y(exu_n25598));
INVX1 exu_U23745(.A(exu_n25598), .Y(exu_n7364));
AND2X1 exu_U23746(.A(alu_byp_rd_data_e[26]), .B(exu_n16299), .Y(exu_n25602));
INVX1 exu_U23747(.A(exu_n25602), .Y(exu_n7365));
AND2X1 exu_U23748(.A(bypass_rs2_data_btwn_mux[26]), .B(exu_n16295), .Y(exu_n25604));
INVX1 exu_U23749(.A(exu_n25604), .Y(exu_n7366));
AND2X1 exu_U23750(.A(alu_byp_rd_data_e[25]), .B(exu_n16299), .Y(exu_n25608));
INVX1 exu_U23751(.A(exu_n25608), .Y(exu_n7367));
AND2X1 exu_U23752(.A(bypass_rs2_data_btwn_mux[25]), .B(exu_n16295), .Y(exu_n25610));
INVX1 exu_U23753(.A(exu_n25610), .Y(exu_n7368));
AND2X1 exu_U23754(.A(alu_byp_rd_data_e[24]), .B(exu_n16299), .Y(exu_n25614));
INVX1 exu_U23755(.A(exu_n25614), .Y(exu_n7369));
AND2X1 exu_U23756(.A(bypass_rs2_data_btwn_mux[24]), .B(exu_n16295), .Y(exu_n25616));
INVX1 exu_U23757(.A(exu_n25616), .Y(exu_n7370));
AND2X1 exu_U23758(.A(alu_byp_rd_data_e[23]), .B(exu_n16299), .Y(exu_n25620));
INVX1 exu_U23759(.A(exu_n25620), .Y(exu_n7371));
AND2X1 exu_U23760(.A(bypass_rs2_data_btwn_mux[23]), .B(exu_n16295), .Y(exu_n25622));
INVX1 exu_U23761(.A(exu_n25622), .Y(exu_n7372));
AND2X1 exu_U23762(.A(alu_byp_rd_data_e[22]), .B(exu_n16299), .Y(exu_n25626));
INVX1 exu_U23763(.A(exu_n25626), .Y(exu_n7373));
AND2X1 exu_U23764(.A(bypass_rs2_data_btwn_mux[22]), .B(exu_n16295), .Y(exu_n25628));
INVX1 exu_U23765(.A(exu_n25628), .Y(exu_n7374));
AND2X1 exu_U23766(.A(alu_byp_rd_data_e[21]), .B(exu_n16299), .Y(exu_n25632));
INVX1 exu_U23767(.A(exu_n25632), .Y(exu_n7375));
AND2X1 exu_U23768(.A(bypass_rs2_data_btwn_mux[21]), .B(exu_n16295), .Y(exu_n25634));
INVX1 exu_U23769(.A(exu_n25634), .Y(exu_n7376));
AND2X1 exu_U23770(.A(alu_byp_rd_data_e[20]), .B(exu_n16299), .Y(exu_n25638));
INVX1 exu_U23771(.A(exu_n25638), .Y(exu_n7377));
AND2X1 exu_U23772(.A(bypass_rs2_data_btwn_mux[20]), .B(exu_n16295), .Y(exu_n25640));
INVX1 exu_U23773(.A(exu_n25640), .Y(exu_n7378));
AND2X1 exu_U23774(.A(alu_byp_rd_data_e[1]), .B(exu_n16299), .Y(exu_n25644));
INVX1 exu_U23775(.A(exu_n25644), .Y(exu_n7379));
AND2X1 exu_U23776(.A(bypass_rs2_data_btwn_mux[1]), .B(exu_n16295), .Y(exu_n25646));
INVX1 exu_U23777(.A(exu_n25646), .Y(exu_n7380));
AND2X1 exu_U23778(.A(alu_byp_rd_data_e[19]), .B(exu_n16299), .Y(exu_n25650));
INVX1 exu_U23779(.A(exu_n25650), .Y(exu_n7381));
AND2X1 exu_U23780(.A(bypass_rs2_data_btwn_mux[19]), .B(exu_n16295), .Y(exu_n25652));
INVX1 exu_U23781(.A(exu_n25652), .Y(exu_n7382));
AND2X1 exu_U23782(.A(alu_byp_rd_data_e[18]), .B(exu_n16299), .Y(exu_n25656));
INVX1 exu_U23783(.A(exu_n25656), .Y(exu_n7383));
AND2X1 exu_U23784(.A(bypass_rs2_data_btwn_mux[18]), .B(exu_n16295), .Y(exu_n25658));
INVX1 exu_U23785(.A(exu_n25658), .Y(exu_n7384));
AND2X1 exu_U23786(.A(alu_byp_rd_data_e[17]), .B(exu_n16299), .Y(exu_n25662));
INVX1 exu_U23787(.A(exu_n25662), .Y(exu_n7385));
AND2X1 exu_U23788(.A(bypass_rs2_data_btwn_mux[17]), .B(exu_n16295), .Y(exu_n25664));
INVX1 exu_U23789(.A(exu_n25664), .Y(exu_n7386));
AND2X1 exu_U23790(.A(alu_byp_rd_data_e[16]), .B(exu_n16299), .Y(exu_n25668));
INVX1 exu_U23791(.A(exu_n25668), .Y(exu_n7387));
AND2X1 exu_U23792(.A(bypass_rs2_data_btwn_mux[16]), .B(exu_n16295), .Y(exu_n25670));
INVX1 exu_U23793(.A(exu_n25670), .Y(exu_n7388));
AND2X1 exu_U23794(.A(alu_byp_rd_data_e[15]), .B(exu_n16299), .Y(exu_n25674));
INVX1 exu_U23795(.A(exu_n25674), .Y(exu_n7389));
AND2X1 exu_U23796(.A(bypass_rs2_data_btwn_mux[15]), .B(exu_n16295), .Y(exu_n25676));
INVX1 exu_U23797(.A(exu_n25676), .Y(exu_n7390));
AND2X1 exu_U23798(.A(alu_byp_rd_data_e[14]), .B(exu_n16299), .Y(exu_n25680));
INVX1 exu_U23799(.A(exu_n25680), .Y(exu_n7391));
AND2X1 exu_U23800(.A(bypass_rs2_data_btwn_mux[14]), .B(exu_n16295), .Y(exu_n25682));
INVX1 exu_U23801(.A(exu_n25682), .Y(exu_n7392));
AND2X1 exu_U23802(.A(alu_byp_rd_data_e[13]), .B(exu_n16299), .Y(exu_n25686));
INVX1 exu_U23803(.A(exu_n25686), .Y(exu_n7393));
AND2X1 exu_U23804(.A(bypass_rs2_data_btwn_mux[13]), .B(exu_n16295), .Y(exu_n25688));
INVX1 exu_U23805(.A(exu_n25688), .Y(exu_n7394));
AND2X1 exu_U23806(.A(alu_byp_rd_data_e[12]), .B(exu_n16299), .Y(exu_n25692));
INVX1 exu_U23807(.A(exu_n25692), .Y(exu_n7395));
AND2X1 exu_U23808(.A(bypass_rs2_data_btwn_mux[12]), .B(exu_n16295), .Y(exu_n25694));
INVX1 exu_U23809(.A(exu_n25694), .Y(exu_n7396));
AND2X1 exu_U23810(.A(alu_byp_rd_data_e[11]), .B(exu_n16299), .Y(exu_n25698));
INVX1 exu_U23811(.A(exu_n25698), .Y(exu_n7397));
AND2X1 exu_U23812(.A(bypass_rs2_data_btwn_mux[11]), .B(exu_n16295), .Y(exu_n25700));
INVX1 exu_U23813(.A(exu_n25700), .Y(exu_n7398));
AND2X1 exu_U23814(.A(alu_byp_rd_data_e[10]), .B(exu_n16299), .Y(exu_n25704));
INVX1 exu_U23815(.A(exu_n25704), .Y(exu_n7399));
AND2X1 exu_U23816(.A(bypass_rs2_data_btwn_mux[10]), .B(exu_n16295), .Y(exu_n25706));
INVX1 exu_U23817(.A(exu_n25706), .Y(exu_n7400));
AND2X1 exu_U23818(.A(alu_byp_rd_data_e[0]), .B(exu_n16299), .Y(exu_n25710));
INVX1 exu_U23819(.A(exu_n25710), .Y(exu_n7401));
AND2X1 exu_U23820(.A(bypass_rs2_data_btwn_mux[0]), .B(exu_n16295), .Y(exu_n25712));
INVX1 exu_U23821(.A(exu_n25712), .Y(exu_n7402));
AND2X1 exu_U23822(.A(exu_n16290), .B(exu_tlu_wsr_data_m[9]), .Y(exu_n25716));
INVX1 exu_U23823(.A(exu_n25716), .Y(exu_n7403));
AND2X1 exu_U23824(.A(exu_tlu_wsr_data_m[8]), .B(exu_n16290), .Y(exu_n25720));
INVX1 exu_U23825(.A(exu_n25720), .Y(exu_n7404));
AND2X1 exu_U23826(.A(exu_tlu_wsr_data_m[7]), .B(exu_n16290), .Y(exu_n25724));
INVX1 exu_U23827(.A(exu_n25724), .Y(exu_n7405));
AND2X1 exu_U23828(.A(exu_tlu_wsr_data_m[6]), .B(exu_n16290), .Y(exu_n25728));
INVX1 exu_U23829(.A(exu_n25728), .Y(exu_n7406));
AND2X1 exu_U23830(.A(exu_tlu_wsr_data_m[63]), .B(exu_n16290), .Y(exu_n25732));
INVX1 exu_U23831(.A(exu_n25732), .Y(exu_n7407));
AND2X1 exu_U23832(.A(exu_tlu_wsr_data_m[62]), .B(exu_n16290), .Y(exu_n25736));
INVX1 exu_U23833(.A(exu_n25736), .Y(exu_n7408));
AND2X1 exu_U23834(.A(exu_tlu_wsr_data_m[61]), .B(exu_n16290), .Y(exu_n25740));
INVX1 exu_U23835(.A(exu_n25740), .Y(exu_n7409));
AND2X1 exu_U23836(.A(exu_tlu_wsr_data_m[60]), .B(exu_n16290), .Y(exu_n25744));
INVX1 exu_U23837(.A(exu_n25744), .Y(exu_n7410));
AND2X1 exu_U23838(.A(exu_tlu_wsr_data_m[5]), .B(exu_n16290), .Y(exu_n25748));
INVX1 exu_U23839(.A(exu_n25748), .Y(exu_n7411));
AND2X1 exu_U23840(.A(exu_tlu_wsr_data_m[59]), .B(exu_n16290), .Y(exu_n25752));
INVX1 exu_U23841(.A(exu_n25752), .Y(exu_n7412));
AND2X1 exu_U23842(.A(exu_tlu_wsr_data_m[58]), .B(exu_n16290), .Y(exu_n25756));
INVX1 exu_U23843(.A(exu_n25756), .Y(exu_n7413));
AND2X1 exu_U23844(.A(exu_tlu_wsr_data_m[57]), .B(exu_n16290), .Y(exu_n25760));
INVX1 exu_U23845(.A(exu_n25760), .Y(exu_n7414));
AND2X1 exu_U23846(.A(exu_tlu_wsr_data_m[56]), .B(exu_n16290), .Y(exu_n25764));
INVX1 exu_U23847(.A(exu_n25764), .Y(exu_n7415));
AND2X1 exu_U23848(.A(exu_tlu_wsr_data_m[55]), .B(exu_n16290), .Y(exu_n25768));
INVX1 exu_U23849(.A(exu_n25768), .Y(exu_n7416));
AND2X1 exu_U23850(.A(exu_tlu_wsr_data_m[54]), .B(exu_n16290), .Y(exu_n25772));
INVX1 exu_U23851(.A(exu_n25772), .Y(exu_n7417));
AND2X1 exu_U23852(.A(exu_tlu_wsr_data_m[53]), .B(exu_n16290), .Y(exu_n25776));
INVX1 exu_U23853(.A(exu_n25776), .Y(exu_n7418));
AND2X1 exu_U23854(.A(exu_tlu_wsr_data_m[52]), .B(exu_n16290), .Y(exu_n25780));
INVX1 exu_U23855(.A(exu_n25780), .Y(exu_n7419));
AND2X1 exu_U23856(.A(exu_tlu_wsr_data_m[51]), .B(exu_n16290), .Y(exu_n25784));
INVX1 exu_U23857(.A(exu_n25784), .Y(exu_n7420));
AND2X1 exu_U23858(.A(exu_tlu_wsr_data_m[50]), .B(exu_n16290), .Y(exu_n25788));
INVX1 exu_U23859(.A(exu_n25788), .Y(exu_n7421));
AND2X1 exu_U23860(.A(exu_tlu_wsr_data_m[4]), .B(exu_n16290), .Y(exu_n25792));
INVX1 exu_U23861(.A(exu_n25792), .Y(exu_n7422));
AND2X1 exu_U23862(.A(exu_tlu_wsr_data_m[49]), .B(exu_n16290), .Y(exu_n25796));
INVX1 exu_U23863(.A(exu_n25796), .Y(exu_n7423));
AND2X1 exu_U23864(.A(exu_tlu_wsr_data_m[48]), .B(exu_n16290), .Y(exu_n25800));
INVX1 exu_U23865(.A(exu_n25800), .Y(exu_n7424));
AND2X1 exu_U23866(.A(exu_tlu_wsr_data_m[47]), .B(exu_n16290), .Y(exu_n25804));
INVX1 exu_U23867(.A(exu_n25804), .Y(exu_n7425));
AND2X1 exu_U23868(.A(exu_tlu_wsr_data_m[46]), .B(exu_n16290), .Y(exu_n25808));
INVX1 exu_U23869(.A(exu_n25808), .Y(exu_n7426));
AND2X1 exu_U23870(.A(exu_tlu_wsr_data_m[45]), .B(exu_n16290), .Y(exu_n25812));
INVX1 exu_U23871(.A(exu_n25812), .Y(exu_n7427));
AND2X1 exu_U23872(.A(exu_tlu_wsr_data_m[44]), .B(exu_n16290), .Y(exu_n25816));
INVX1 exu_U23873(.A(exu_n25816), .Y(exu_n7428));
AND2X1 exu_U23874(.A(exu_tlu_wsr_data_m[43]), .B(exu_n16290), .Y(exu_n25820));
INVX1 exu_U23875(.A(exu_n25820), .Y(exu_n7429));
AND2X1 exu_U23876(.A(exu_tlu_wsr_data_m[42]), .B(exu_n16290), .Y(exu_n25824));
INVX1 exu_U23877(.A(exu_n25824), .Y(exu_n7430));
AND2X1 exu_U23878(.A(exu_tlu_wsr_data_m[41]), .B(exu_n16290), .Y(exu_n25828));
INVX1 exu_U23879(.A(exu_n25828), .Y(exu_n7431));
AND2X1 exu_U23880(.A(exu_tlu_wsr_data_m[40]), .B(exu_n16290), .Y(exu_n25832));
INVX1 exu_U23881(.A(exu_n25832), .Y(exu_n7432));
AND2X1 exu_U23882(.A(exu_tlu_wsr_data_m[3]), .B(exu_n16290), .Y(exu_n25836));
INVX1 exu_U23883(.A(exu_n25836), .Y(exu_n7433));
AND2X1 exu_U23884(.A(exu_tlu_wsr_data_m[39]), .B(exu_n16290), .Y(exu_n25840));
INVX1 exu_U23885(.A(exu_n25840), .Y(exu_n7434));
AND2X1 exu_U23886(.A(exu_tlu_wsr_data_m[38]), .B(exu_n16290), .Y(exu_n25844));
INVX1 exu_U23887(.A(exu_n25844), .Y(exu_n7435));
AND2X1 exu_U23888(.A(exu_tlu_wsr_data_m[37]), .B(exu_n16290), .Y(exu_n25848));
INVX1 exu_U23889(.A(exu_n25848), .Y(exu_n7436));
AND2X1 exu_U23890(.A(exu_tlu_wsr_data_m[36]), .B(exu_n16290), .Y(exu_n25852));
INVX1 exu_U23891(.A(exu_n25852), .Y(exu_n7437));
AND2X1 exu_U23892(.A(exu_tlu_wsr_data_m[35]), .B(exu_n16290), .Y(exu_n25856));
INVX1 exu_U23893(.A(exu_n25856), .Y(exu_n7438));
AND2X1 exu_U23894(.A(exu_tlu_wsr_data_m[34]), .B(exu_n16290), .Y(exu_n25860));
INVX1 exu_U23895(.A(exu_n25860), .Y(exu_n7439));
AND2X1 exu_U23896(.A(exu_tlu_wsr_data_m[33]), .B(exu_n16290), .Y(exu_n25864));
INVX1 exu_U23897(.A(exu_n25864), .Y(exu_n7440));
AND2X1 exu_U23898(.A(exu_tlu_wsr_data_m[32]), .B(exu_n16290), .Y(exu_n25868));
INVX1 exu_U23899(.A(exu_n25868), .Y(exu_n7441));
AND2X1 exu_U23900(.A(exu_tlu_wsr_data_m[31]), .B(exu_n16290), .Y(exu_n25872));
INVX1 exu_U23901(.A(exu_n25872), .Y(exu_n7442));
AND2X1 exu_U23902(.A(exu_tlu_wsr_data_m[30]), .B(exu_n16290), .Y(exu_n25876));
INVX1 exu_U23903(.A(exu_n25876), .Y(exu_n7443));
AND2X1 exu_U23904(.A(exu_tlu_wsr_data_m[2]), .B(exu_n16290), .Y(exu_n25880));
INVX1 exu_U23905(.A(exu_n25880), .Y(exu_n7444));
AND2X1 exu_U23906(.A(exu_tlu_wsr_data_m[29]), .B(exu_n16290), .Y(exu_n25884));
INVX1 exu_U23907(.A(exu_n25884), .Y(exu_n7445));
AND2X1 exu_U23908(.A(exu_tlu_wsr_data_m[28]), .B(exu_n16290), .Y(exu_n25888));
INVX1 exu_U23909(.A(exu_n25888), .Y(exu_n7446));
AND2X1 exu_U23910(.A(exu_tlu_wsr_data_m[27]), .B(exu_n16290), .Y(exu_n25892));
INVX1 exu_U23911(.A(exu_n25892), .Y(exu_n7447));
AND2X1 exu_U23912(.A(exu_tlu_wsr_data_m[26]), .B(exu_n16290), .Y(exu_n25896));
INVX1 exu_U23913(.A(exu_n25896), .Y(exu_n7448));
AND2X1 exu_U23914(.A(exu_tlu_wsr_data_m[25]), .B(exu_n16290), .Y(exu_n25900));
INVX1 exu_U23915(.A(exu_n25900), .Y(exu_n7449));
AND2X1 exu_U23916(.A(exu_tlu_wsr_data_m[24]), .B(exu_n16290), .Y(exu_n25904));
INVX1 exu_U23917(.A(exu_n25904), .Y(exu_n7450));
AND2X1 exu_U23918(.A(exu_tlu_wsr_data_m[23]), .B(exu_n16290), .Y(exu_n25908));
INVX1 exu_U23919(.A(exu_n25908), .Y(exu_n7451));
AND2X1 exu_U23920(.A(exu_tlu_wsr_data_m[22]), .B(exu_n16290), .Y(exu_n25912));
INVX1 exu_U23921(.A(exu_n25912), .Y(exu_n7452));
AND2X1 exu_U23922(.A(exu_tlu_wsr_data_m[21]), .B(exu_n16290), .Y(exu_n25916));
INVX1 exu_U23923(.A(exu_n25916), .Y(exu_n7453));
AND2X1 exu_U23924(.A(exu_tlu_wsr_data_m[20]), .B(exu_n16290), .Y(exu_n25920));
INVX1 exu_U23925(.A(exu_n25920), .Y(exu_n7454));
AND2X1 exu_U23926(.A(exu_tlu_wsr_data_m[1]), .B(exu_n16290), .Y(exu_n25924));
INVX1 exu_U23927(.A(exu_n25924), .Y(exu_n7455));
AND2X1 exu_U23928(.A(exu_tlu_wsr_data_m[19]), .B(exu_n16290), .Y(exu_n25928));
INVX1 exu_U23929(.A(exu_n25928), .Y(exu_n7456));
AND2X1 exu_U23930(.A(exu_tlu_wsr_data_m[18]), .B(exu_n16290), .Y(exu_n25932));
INVX1 exu_U23931(.A(exu_n25932), .Y(exu_n7457));
AND2X1 exu_U23932(.A(exu_tlu_wsr_data_m[17]), .B(exu_n16290), .Y(exu_n25936));
INVX1 exu_U23933(.A(exu_n25936), .Y(exu_n7458));
AND2X1 exu_U23934(.A(exu_tlu_wsr_data_m[16]), .B(exu_n16290), .Y(exu_n25940));
INVX1 exu_U23935(.A(exu_n25940), .Y(exu_n7459));
AND2X1 exu_U23936(.A(exu_tlu_wsr_data_m[15]), .B(exu_n16290), .Y(exu_n25944));
INVX1 exu_U23937(.A(exu_n25944), .Y(exu_n7460));
AND2X1 exu_U23938(.A(exu_tlu_wsr_data_m[14]), .B(exu_n16290), .Y(exu_n25948));
INVX1 exu_U23939(.A(exu_n25948), .Y(exu_n7461));
AND2X1 exu_U23940(.A(exu_tlu_wsr_data_m[13]), .B(exu_n16290), .Y(exu_n25952));
INVX1 exu_U23941(.A(exu_n25952), .Y(exu_n7462));
AND2X1 exu_U23942(.A(exu_tlu_wsr_data_m[12]), .B(exu_n16290), .Y(exu_n25956));
INVX1 exu_U23943(.A(exu_n25956), .Y(exu_n7463));
AND2X1 exu_U23944(.A(exu_tlu_wsr_data_m[11]), .B(exu_n16290), .Y(exu_n25960));
INVX1 exu_U23945(.A(exu_n25960), .Y(exu_n7464));
AND2X1 exu_U23946(.A(exu_tlu_wsr_data_m[10]), .B(exu_n16290), .Y(exu_n25964));
INVX1 exu_U23947(.A(exu_n25964), .Y(exu_n7465));
AND2X1 exu_U23948(.A(exu_tlu_wsr_data_m[0]), .B(exu_n16290), .Y(exu_n25968));
INVX1 exu_U23949(.A(exu_n25968), .Y(exu_n7466));
AND2X1 exu_U23950(.A(exu_n16292), .B(alu_byp_rd_data_e[9]), .Y(exu_n25972));
INVX1 exu_U23951(.A(exu_n25972), .Y(exu_n7467));
AND2X1 exu_U23952(.A(exu_n15961), .B(bypass_rs3_data_btwn_mux[9]), .Y(exu_n25974));
INVX1 exu_U23953(.A(exu_n25974), .Y(exu_n7468));
AND2X1 exu_U23954(.A(alu_byp_rd_data_e[8]), .B(exu_n16292), .Y(exu_n25978));
INVX1 exu_U23955(.A(exu_n25978), .Y(exu_n7469));
AND2X1 exu_U23956(.A(bypass_rs3_data_btwn_mux[8]), .B(exu_n15961), .Y(exu_n25980));
INVX1 exu_U23957(.A(exu_n25980), .Y(exu_n7470));
AND2X1 exu_U23958(.A(alu_byp_rd_data_e[7]), .B(exu_n16292), .Y(exu_n25984));
INVX1 exu_U23959(.A(exu_n25984), .Y(exu_n7471));
AND2X1 exu_U23960(.A(bypass_rs3_data_btwn_mux[7]), .B(exu_n15961), .Y(exu_n25986));
INVX1 exu_U23961(.A(exu_n25986), .Y(exu_n7472));
AND2X1 exu_U23962(.A(alu_byp_rd_data_e[6]), .B(exu_n16292), .Y(exu_n25990));
INVX1 exu_U23963(.A(exu_n25990), .Y(exu_n7473));
AND2X1 exu_U23964(.A(bypass_rs3_data_btwn_mux[6]), .B(exu_n15961), .Y(exu_n25992));
INVX1 exu_U23965(.A(exu_n25992), .Y(exu_n7474));
AND2X1 exu_U23966(.A(alu_byp_rd_data_e[63]), .B(exu_n16292), .Y(exu_n25996));
INVX1 exu_U23967(.A(exu_n25996), .Y(exu_n7475));
AND2X1 exu_U23968(.A(bypass_rs3_data_btwn_mux[63]), .B(exu_n15961), .Y(exu_n25998));
INVX1 exu_U23969(.A(exu_n25998), .Y(exu_n7476));
AND2X1 exu_U23970(.A(alu_byp_rd_data_e[62]), .B(exu_n16292), .Y(exu_n26002));
INVX1 exu_U23971(.A(exu_n26002), .Y(exu_n7477));
AND2X1 exu_U23972(.A(bypass_rs3_data_btwn_mux[62]), .B(exu_n15961), .Y(exu_n26004));
INVX1 exu_U23973(.A(exu_n26004), .Y(exu_n7478));
AND2X1 exu_U23974(.A(alu_byp_rd_data_e[61]), .B(exu_n16292), .Y(exu_n26008));
INVX1 exu_U23975(.A(exu_n26008), .Y(exu_n7479));
AND2X1 exu_U23976(.A(bypass_rs3_data_btwn_mux[61]), .B(exu_n15961), .Y(exu_n26010));
INVX1 exu_U23977(.A(exu_n26010), .Y(exu_n7480));
AND2X1 exu_U23978(.A(alu_byp_rd_data_e[60]), .B(exu_n16292), .Y(exu_n26014));
INVX1 exu_U23979(.A(exu_n26014), .Y(exu_n7481));
AND2X1 exu_U23980(.A(bypass_rs3_data_btwn_mux[60]), .B(exu_n15961), .Y(exu_n26016));
INVX1 exu_U23981(.A(exu_n26016), .Y(exu_n7482));
AND2X1 exu_U23982(.A(alu_byp_rd_data_e[5]), .B(exu_n16292), .Y(exu_n26020));
INVX1 exu_U23983(.A(exu_n26020), .Y(exu_n7483));
AND2X1 exu_U23984(.A(bypass_rs3_data_btwn_mux[5]), .B(exu_n15961), .Y(exu_n26022));
INVX1 exu_U23985(.A(exu_n26022), .Y(exu_n7484));
AND2X1 exu_U23986(.A(alu_byp_rd_data_e[59]), .B(exu_n16292), .Y(exu_n26026));
INVX1 exu_U23987(.A(exu_n26026), .Y(exu_n7485));
AND2X1 exu_U23988(.A(bypass_rs3_data_btwn_mux[59]), .B(exu_n15961), .Y(exu_n26028));
INVX1 exu_U23989(.A(exu_n26028), .Y(exu_n7486));
AND2X1 exu_U23990(.A(alu_byp_rd_data_e[58]), .B(exu_n16292), .Y(exu_n26032));
INVX1 exu_U23991(.A(exu_n26032), .Y(exu_n7487));
AND2X1 exu_U23992(.A(bypass_rs3_data_btwn_mux[58]), .B(exu_n15961), .Y(exu_n26034));
INVX1 exu_U23993(.A(exu_n26034), .Y(exu_n7488));
AND2X1 exu_U23994(.A(alu_byp_rd_data_e[57]), .B(exu_n16292), .Y(exu_n26038));
INVX1 exu_U23995(.A(exu_n26038), .Y(exu_n7489));
AND2X1 exu_U23996(.A(bypass_rs3_data_btwn_mux[57]), .B(exu_n15961), .Y(exu_n26040));
INVX1 exu_U23997(.A(exu_n26040), .Y(exu_n7490));
AND2X1 exu_U23998(.A(alu_byp_rd_data_e[56]), .B(exu_n16292), .Y(exu_n26044));
INVX1 exu_U23999(.A(exu_n26044), .Y(exu_n7491));
AND2X1 exu_U24000(.A(bypass_rs3_data_btwn_mux[56]), .B(exu_n15961), .Y(exu_n26046));
INVX1 exu_U24001(.A(exu_n26046), .Y(exu_n7492));
AND2X1 exu_U24002(.A(alu_byp_rd_data_e[55]), .B(exu_n16292), .Y(exu_n26050));
INVX1 exu_U24003(.A(exu_n26050), .Y(exu_n7493));
AND2X1 exu_U24004(.A(bypass_rs3_data_btwn_mux[55]), .B(exu_n19184), .Y(exu_n26052));
INVX1 exu_U24005(.A(exu_n26052), .Y(exu_n7494));
AND2X1 exu_U24006(.A(alu_byp_rd_data_e[54]), .B(exu_n16292), .Y(exu_n26056));
INVX1 exu_U24007(.A(exu_n26056), .Y(exu_n7495));
AND2X1 exu_U24008(.A(bypass_rs3_data_btwn_mux[54]), .B(exu_n15961), .Y(exu_n26058));
INVX1 exu_U24009(.A(exu_n26058), .Y(exu_n7496));
AND2X1 exu_U24010(.A(alu_byp_rd_data_e[53]), .B(exu_n16292), .Y(exu_n26062));
INVX1 exu_U24011(.A(exu_n26062), .Y(exu_n7497));
AND2X1 exu_U24012(.A(bypass_rs3_data_btwn_mux[53]), .B(exu_n19184), .Y(exu_n26064));
INVX1 exu_U24013(.A(exu_n26064), .Y(exu_n7498));
AND2X1 exu_U24014(.A(alu_byp_rd_data_e[52]), .B(exu_n16292), .Y(exu_n26068));
INVX1 exu_U24015(.A(exu_n26068), .Y(exu_n7499));
AND2X1 exu_U24016(.A(bypass_rs3_data_btwn_mux[52]), .B(exu_n15961), .Y(exu_n26070));
INVX1 exu_U24017(.A(exu_n26070), .Y(exu_n7500));
AND2X1 exu_U24018(.A(alu_byp_rd_data_e[51]), .B(exu_n16292), .Y(exu_n26074));
INVX1 exu_U24019(.A(exu_n26074), .Y(exu_n7501));
AND2X1 exu_U24020(.A(bypass_rs3_data_btwn_mux[51]), .B(exu_n19184), .Y(exu_n26076));
INVX1 exu_U24021(.A(exu_n26076), .Y(exu_n7502));
AND2X1 exu_U24022(.A(alu_byp_rd_data_e[50]), .B(exu_n16292), .Y(exu_n26080));
INVX1 exu_U24023(.A(exu_n26080), .Y(exu_n7503));
AND2X1 exu_U24024(.A(bypass_rs3_data_btwn_mux[50]), .B(exu_n15961), .Y(exu_n26082));
INVX1 exu_U24025(.A(exu_n26082), .Y(exu_n7504));
AND2X1 exu_U24026(.A(alu_byp_rd_data_e[4]), .B(exu_n16292), .Y(exu_n26086));
INVX1 exu_U24027(.A(exu_n26086), .Y(exu_n7505));
AND2X1 exu_U24028(.A(bypass_rs3_data_btwn_mux[4]), .B(exu_n19184), .Y(exu_n26088));
INVX1 exu_U24029(.A(exu_n26088), .Y(exu_n7506));
AND2X1 exu_U24030(.A(alu_byp_rd_data_e[49]), .B(exu_n16292), .Y(exu_n26092));
INVX1 exu_U24031(.A(exu_n26092), .Y(exu_n7507));
AND2X1 exu_U24032(.A(bypass_rs3_data_btwn_mux[49]), .B(exu_n15961), .Y(exu_n26094));
INVX1 exu_U24033(.A(exu_n26094), .Y(exu_n7508));
AND2X1 exu_U24034(.A(alu_byp_rd_data_e[48]), .B(exu_n16292), .Y(exu_n26098));
INVX1 exu_U24035(.A(exu_n26098), .Y(exu_n7509));
AND2X1 exu_U24036(.A(bypass_rs3_data_btwn_mux[48]), .B(exu_n19184), .Y(exu_n26100));
INVX1 exu_U24037(.A(exu_n26100), .Y(exu_n7510));
AND2X1 exu_U24038(.A(alu_byp_rd_data_e[47]), .B(exu_n16292), .Y(exu_n26104));
INVX1 exu_U24039(.A(exu_n26104), .Y(exu_n7511));
AND2X1 exu_U24040(.A(bypass_rs3_data_btwn_mux[47]), .B(exu_n15961), .Y(exu_n26106));
INVX1 exu_U24041(.A(exu_n26106), .Y(exu_n7512));
AND2X1 exu_U24042(.A(alu_byp_rd_data_e[46]), .B(exu_n16292), .Y(exu_n26110));
INVX1 exu_U24043(.A(exu_n26110), .Y(exu_n7513));
AND2X1 exu_U24044(.A(bypass_rs3_data_btwn_mux[46]), .B(exu_n19184), .Y(exu_n26112));
INVX1 exu_U24045(.A(exu_n26112), .Y(exu_n7514));
AND2X1 exu_U24046(.A(alu_byp_rd_data_e[45]), .B(exu_n16292), .Y(exu_n26116));
INVX1 exu_U24047(.A(exu_n26116), .Y(exu_n7515));
AND2X1 exu_U24048(.A(bypass_rs3_data_btwn_mux[45]), .B(exu_n15961), .Y(exu_n26118));
INVX1 exu_U24049(.A(exu_n26118), .Y(exu_n7516));
AND2X1 exu_U24050(.A(alu_byp_rd_data_e[44]), .B(exu_n16292), .Y(exu_n26122));
INVX1 exu_U24051(.A(exu_n26122), .Y(exu_n7517));
AND2X1 exu_U24052(.A(bypass_rs3_data_btwn_mux[44]), .B(exu_n19184), .Y(exu_n26124));
INVX1 exu_U24053(.A(exu_n26124), .Y(exu_n7518));
AND2X1 exu_U24054(.A(alu_byp_rd_data_e[43]), .B(exu_n16292), .Y(exu_n26128));
INVX1 exu_U24055(.A(exu_n26128), .Y(exu_n7519));
AND2X1 exu_U24056(.A(bypass_rs3_data_btwn_mux[43]), .B(exu_n15961), .Y(exu_n26130));
INVX1 exu_U24057(.A(exu_n26130), .Y(exu_n7520));
AND2X1 exu_U24058(.A(alu_byp_rd_data_e[42]), .B(exu_n16292), .Y(exu_n26134));
INVX1 exu_U24059(.A(exu_n26134), .Y(exu_n7521));
AND2X1 exu_U24060(.A(bypass_rs3_data_btwn_mux[42]), .B(exu_n15961), .Y(exu_n26136));
INVX1 exu_U24061(.A(exu_n26136), .Y(exu_n7522));
AND2X1 exu_U24062(.A(alu_byp_rd_data_e[41]), .B(exu_n16292), .Y(exu_n26140));
INVX1 exu_U24063(.A(exu_n26140), .Y(exu_n7523));
AND2X1 exu_U24064(.A(bypass_rs3_data_btwn_mux[41]), .B(exu_n19184), .Y(exu_n26142));
INVX1 exu_U24065(.A(exu_n26142), .Y(exu_n7524));
AND2X1 exu_U24066(.A(alu_byp_rd_data_e[40]), .B(exu_n16292), .Y(exu_n26146));
INVX1 exu_U24067(.A(exu_n26146), .Y(exu_n7525));
AND2X1 exu_U24068(.A(bypass_rs3_data_btwn_mux[40]), .B(exu_n15961), .Y(exu_n26148));
INVX1 exu_U24069(.A(exu_n26148), .Y(exu_n7526));
AND2X1 exu_U24070(.A(alu_byp_rd_data_e[3]), .B(exu_n16292), .Y(exu_n26152));
INVX1 exu_U24071(.A(exu_n26152), .Y(exu_n7527));
AND2X1 exu_U24072(.A(bypass_rs3_data_btwn_mux[3]), .B(exu_n19184), .Y(exu_n26154));
INVX1 exu_U24073(.A(exu_n26154), .Y(exu_n7528));
AND2X1 exu_U24074(.A(alu_byp_rd_data_e[39]), .B(exu_n16292), .Y(exu_n26158));
INVX1 exu_U24075(.A(exu_n26158), .Y(exu_n7529));
AND2X1 exu_U24076(.A(bypass_rs3_data_btwn_mux[39]), .B(exu_n19184), .Y(exu_n26160));
INVX1 exu_U24077(.A(exu_n26160), .Y(exu_n7530));
AND2X1 exu_U24078(.A(alu_byp_rd_data_e[38]), .B(exu_n16292), .Y(exu_n26164));
INVX1 exu_U24079(.A(exu_n26164), .Y(exu_n7531));
AND2X1 exu_U24080(.A(bypass_rs3_data_btwn_mux[38]), .B(exu_n15961), .Y(exu_n26166));
INVX1 exu_U24081(.A(exu_n26166), .Y(exu_n7532));
AND2X1 exu_U24082(.A(alu_byp_rd_data_e[37]), .B(exu_n16292), .Y(exu_n26170));
INVX1 exu_U24083(.A(exu_n26170), .Y(exu_n7533));
AND2X1 exu_U24084(.A(bypass_rs3_data_btwn_mux[37]), .B(exu_n15961), .Y(exu_n26172));
INVX1 exu_U24085(.A(exu_n26172), .Y(exu_n7534));
AND2X1 exu_U24086(.A(alu_byp_rd_data_e[36]), .B(exu_n16292), .Y(exu_n26176));
INVX1 exu_U24087(.A(exu_n26176), .Y(exu_n7535));
AND2X1 exu_U24088(.A(bypass_rs3_data_btwn_mux[36]), .B(exu_n19184), .Y(exu_n26178));
INVX1 exu_U24089(.A(exu_n26178), .Y(exu_n7536));
AND2X1 exu_U24090(.A(alu_byp_rd_data_e[35]), .B(exu_n16292), .Y(exu_n26182));
INVX1 exu_U24091(.A(exu_n26182), .Y(exu_n7537));
AND2X1 exu_U24092(.A(bypass_rs3_data_btwn_mux[35]), .B(exu_n15961), .Y(exu_n26184));
INVX1 exu_U24093(.A(exu_n26184), .Y(exu_n7538));
AND2X1 exu_U24094(.A(alu_byp_rd_data_e[34]), .B(exu_n16292), .Y(exu_n26188));
INVX1 exu_U24095(.A(exu_n26188), .Y(exu_n7539));
AND2X1 exu_U24096(.A(bypass_rs3_data_btwn_mux[34]), .B(exu_n19184), .Y(exu_n26190));
INVX1 exu_U24097(.A(exu_n26190), .Y(exu_n7540));
AND2X1 exu_U24098(.A(alu_byp_rd_data_e[33]), .B(exu_n16292), .Y(exu_n26194));
INVX1 exu_U24099(.A(exu_n26194), .Y(exu_n7541));
AND2X1 exu_U24100(.A(bypass_rs3_data_btwn_mux[33]), .B(exu_n19184), .Y(exu_n26196));
INVX1 exu_U24101(.A(exu_n26196), .Y(exu_n7542));
AND2X1 exu_U24102(.A(alu_byp_rd_data_e[32]), .B(exu_n16292), .Y(exu_n26200));
INVX1 exu_U24103(.A(exu_n26200), .Y(exu_n7543));
AND2X1 exu_U24104(.A(bypass_rs3_data_btwn_mux[32]), .B(exu_n15961), .Y(exu_n26202));
INVX1 exu_U24105(.A(exu_n26202), .Y(exu_n7544));
AND2X1 exu_U24106(.A(alu_byp_rd_data_e[31]), .B(exu_n16292), .Y(exu_n26206));
INVX1 exu_U24107(.A(exu_n26206), .Y(exu_n7545));
AND2X1 exu_U24108(.A(bypass_rs3_data_btwn_mux[31]), .B(exu_n15961), .Y(exu_n26208));
INVX1 exu_U24109(.A(exu_n26208), .Y(exu_n7546));
AND2X1 exu_U24110(.A(alu_byp_rd_data_e[30]), .B(exu_n16292), .Y(exu_n26212));
INVX1 exu_U24111(.A(exu_n26212), .Y(exu_n7547));
AND2X1 exu_U24112(.A(bypass_rs3_data_btwn_mux[30]), .B(exu_n15961), .Y(exu_n26214));
INVX1 exu_U24113(.A(exu_n26214), .Y(exu_n7548));
AND2X1 exu_U24114(.A(alu_byp_rd_data_e[2]), .B(exu_n16292), .Y(exu_n26218));
INVX1 exu_U24115(.A(exu_n26218), .Y(exu_n7549));
AND2X1 exu_U24116(.A(bypass_rs3_data_btwn_mux[2]), .B(exu_n19184), .Y(exu_n26220));
INVX1 exu_U24117(.A(exu_n26220), .Y(exu_n7550));
AND2X1 exu_U24118(.A(alu_byp_rd_data_e[29]), .B(exu_n16292), .Y(exu_n26224));
INVX1 exu_U24119(.A(exu_n26224), .Y(exu_n7551));
AND2X1 exu_U24120(.A(bypass_rs3_data_btwn_mux[29]), .B(exu_n19184), .Y(exu_n26226));
INVX1 exu_U24121(.A(exu_n26226), .Y(exu_n7552));
AND2X1 exu_U24122(.A(alu_byp_rd_data_e[28]), .B(exu_n16292), .Y(exu_n26230));
INVX1 exu_U24123(.A(exu_n26230), .Y(exu_n7553));
AND2X1 exu_U24124(.A(bypass_rs3_data_btwn_mux[28]), .B(exu_n15961), .Y(exu_n26232));
INVX1 exu_U24125(.A(exu_n26232), .Y(exu_n7554));
AND2X1 exu_U24126(.A(alu_byp_rd_data_e[27]), .B(exu_n16292), .Y(exu_n26236));
INVX1 exu_U24127(.A(exu_n26236), .Y(exu_n7555));
AND2X1 exu_U24128(.A(bypass_rs3_data_btwn_mux[27]), .B(exu_n19184), .Y(exu_n26238));
INVX1 exu_U24129(.A(exu_n26238), .Y(exu_n7556));
AND2X1 exu_U24130(.A(alu_byp_rd_data_e[26]), .B(exu_n16292), .Y(exu_n26242));
INVX1 exu_U24131(.A(exu_n26242), .Y(exu_n7557));
AND2X1 exu_U24132(.A(bypass_rs3_data_btwn_mux[26]), .B(exu_n19184), .Y(exu_n26244));
INVX1 exu_U24133(.A(exu_n26244), .Y(exu_n7558));
AND2X1 exu_U24134(.A(alu_byp_rd_data_e[25]), .B(exu_n16292), .Y(exu_n26248));
INVX1 exu_U24135(.A(exu_n26248), .Y(exu_n7559));
AND2X1 exu_U24136(.A(bypass_rs3_data_btwn_mux[25]), .B(exu_n19184), .Y(exu_n26250));
INVX1 exu_U24137(.A(exu_n26250), .Y(exu_n7560));
AND2X1 exu_U24138(.A(alu_byp_rd_data_e[24]), .B(exu_n16292), .Y(exu_n26254));
INVX1 exu_U24139(.A(exu_n26254), .Y(exu_n7561));
AND2X1 exu_U24140(.A(bypass_rs3_data_btwn_mux[24]), .B(exu_n15961), .Y(exu_n26256));
INVX1 exu_U24141(.A(exu_n26256), .Y(exu_n7562));
AND2X1 exu_U24142(.A(alu_byp_rd_data_e[23]), .B(exu_n16292), .Y(exu_n26260));
INVX1 exu_U24143(.A(exu_n26260), .Y(exu_n7563));
AND2X1 exu_U24144(.A(bypass_rs3_data_btwn_mux[23]), .B(exu_n15961), .Y(exu_n26262));
INVX1 exu_U24145(.A(exu_n26262), .Y(exu_n7564));
AND2X1 exu_U24146(.A(alu_byp_rd_data_e[22]), .B(exu_n16292), .Y(exu_n26266));
INVX1 exu_U24147(.A(exu_n26266), .Y(exu_n7565));
AND2X1 exu_U24148(.A(bypass_rs3_data_btwn_mux[22]), .B(exu_n19184), .Y(exu_n26268));
INVX1 exu_U24149(.A(exu_n26268), .Y(exu_n7566));
AND2X1 exu_U24150(.A(alu_byp_rd_data_e[21]), .B(exu_n16292), .Y(exu_n26272));
INVX1 exu_U24151(.A(exu_n26272), .Y(exu_n7567));
AND2X1 exu_U24152(.A(bypass_rs3_data_btwn_mux[21]), .B(exu_n19184), .Y(exu_n26274));
INVX1 exu_U24153(.A(exu_n26274), .Y(exu_n7568));
AND2X1 exu_U24154(.A(alu_byp_rd_data_e[20]), .B(exu_n16292), .Y(exu_n26278));
INVX1 exu_U24155(.A(exu_n26278), .Y(exu_n7569));
AND2X1 exu_U24156(.A(bypass_rs3_data_btwn_mux[20]), .B(exu_n15961), .Y(exu_n26280));
INVX1 exu_U24157(.A(exu_n26280), .Y(exu_n7570));
AND2X1 exu_U24158(.A(alu_byp_rd_data_e[1]), .B(exu_n16292), .Y(exu_n26284));
INVX1 exu_U24159(.A(exu_n26284), .Y(exu_n7571));
AND2X1 exu_U24160(.A(bypass_rs3_data_btwn_mux[1]), .B(exu_n19184), .Y(exu_n26286));
INVX1 exu_U24161(.A(exu_n26286), .Y(exu_n7572));
AND2X1 exu_U24162(.A(alu_byp_rd_data_e[19]), .B(exu_n16292), .Y(exu_n26290));
INVX1 exu_U24163(.A(exu_n26290), .Y(exu_n7573));
AND2X1 exu_U24164(.A(bypass_rs3_data_btwn_mux[19]), .B(exu_n19184), .Y(exu_n26292));
INVX1 exu_U24165(.A(exu_n26292), .Y(exu_n7574));
AND2X1 exu_U24166(.A(alu_byp_rd_data_e[18]), .B(exu_n16292), .Y(exu_n26296));
INVX1 exu_U24167(.A(exu_n26296), .Y(exu_n7575));
AND2X1 exu_U24168(.A(bypass_rs3_data_btwn_mux[18]), .B(exu_n19184), .Y(exu_n26298));
INVX1 exu_U24169(.A(exu_n26298), .Y(exu_n7576));
AND2X1 exu_U24170(.A(alu_byp_rd_data_e[17]), .B(exu_n16292), .Y(exu_n26302));
INVX1 exu_U24171(.A(exu_n26302), .Y(exu_n7577));
AND2X1 exu_U24172(.A(bypass_rs3_data_btwn_mux[17]), .B(exu_n19184), .Y(exu_n26304));
INVX1 exu_U24173(.A(exu_n26304), .Y(exu_n7578));
AND2X1 exu_U24174(.A(alu_byp_rd_data_e[16]), .B(exu_n16292), .Y(exu_n26308));
INVX1 exu_U24175(.A(exu_n26308), .Y(exu_n7579));
AND2X1 exu_U24176(.A(bypass_rs3_data_btwn_mux[16]), .B(exu_n19184), .Y(exu_n26310));
INVX1 exu_U24177(.A(exu_n26310), .Y(exu_n7580));
AND2X1 exu_U24178(.A(alu_byp_rd_data_e[15]), .B(exu_n16292), .Y(exu_n26314));
INVX1 exu_U24179(.A(exu_n26314), .Y(exu_n7581));
AND2X1 exu_U24180(.A(bypass_rs3_data_btwn_mux[15]), .B(exu_n19184), .Y(exu_n26316));
INVX1 exu_U24181(.A(exu_n26316), .Y(exu_n7582));
AND2X1 exu_U24182(.A(alu_byp_rd_data_e[14]), .B(exu_n16292), .Y(exu_n26320));
INVX1 exu_U24183(.A(exu_n26320), .Y(exu_n7583));
AND2X1 exu_U24184(.A(bypass_rs3_data_btwn_mux[14]), .B(exu_n19184), .Y(exu_n26322));
INVX1 exu_U24185(.A(exu_n26322), .Y(exu_n7584));
AND2X1 exu_U24186(.A(alu_byp_rd_data_e[13]), .B(exu_n16292), .Y(exu_n26326));
INVX1 exu_U24187(.A(exu_n26326), .Y(exu_n7585));
AND2X1 exu_U24188(.A(bypass_rs3_data_btwn_mux[13]), .B(exu_n19184), .Y(exu_n26328));
INVX1 exu_U24189(.A(exu_n26328), .Y(exu_n7586));
AND2X1 exu_U24190(.A(alu_byp_rd_data_e[12]), .B(exu_n16292), .Y(exu_n26332));
INVX1 exu_U24191(.A(exu_n26332), .Y(exu_n7587));
AND2X1 exu_U24192(.A(bypass_rs3_data_btwn_mux[12]), .B(exu_n19184), .Y(exu_n26334));
INVX1 exu_U24193(.A(exu_n26334), .Y(exu_n7588));
AND2X1 exu_U24194(.A(alu_byp_rd_data_e[11]), .B(exu_n16292), .Y(exu_n26338));
INVX1 exu_U24195(.A(exu_n26338), .Y(exu_n7589));
AND2X1 exu_U24196(.A(bypass_rs3_data_btwn_mux[11]), .B(exu_n19184), .Y(exu_n26340));
INVX1 exu_U24197(.A(exu_n26340), .Y(exu_n7590));
AND2X1 exu_U24198(.A(alu_byp_rd_data_e[10]), .B(exu_n16292), .Y(exu_n26344));
INVX1 exu_U24199(.A(exu_n26344), .Y(exu_n7591));
AND2X1 exu_U24200(.A(bypass_rs3_data_btwn_mux[10]), .B(exu_n19184), .Y(exu_n26346));
INVX1 exu_U24201(.A(exu_n26346), .Y(exu_n7592));
AND2X1 exu_U24202(.A(alu_byp_rd_data_e[0]), .B(exu_n16292), .Y(exu_n26350));
INVX1 exu_U24203(.A(exu_n26350), .Y(exu_n7593));
AND2X1 exu_U24204(.A(bypass_rs3_data_btwn_mux[0]), .B(exu_n19184), .Y(exu_n26352));
INVX1 exu_U24205(.A(exu_n26352), .Y(exu_n7594));
AND2X1 exu_U24206(.A(exu_n15977), .B(exu_n10240), .Y(exu_n26356));
INVX1 exu_U24207(.A(exu_n26356), .Y(exu_n7595));
AND2X1 exu_U24208(.A(ecl_sel_sum_e), .B(exu_ifu_brpc_e[9]), .Y(exu_n26358));
INVX1 exu_U24209(.A(exu_n26358), .Y(exu_n7596));
AND2X1 exu_U24210(.A(exu_n11235), .B(exu_n15977), .Y(exu_n26362));
INVX1 exu_U24211(.A(exu_n26362), .Y(exu_n7597));
AND2X1 exu_U24212(.A(exu_ifu_brpc_e[8]), .B(exu_n16157), .Y(exu_n26364));
INVX1 exu_U24213(.A(exu_n26364), .Y(exu_n7598));
AND2X1 exu_U24214(.A(exu_n11237), .B(exu_n15977), .Y(exu_n26368));
INVX1 exu_U24215(.A(exu_n26368), .Y(exu_n7599));
AND2X1 exu_U24216(.A(exu_ifu_brpc_e[7]), .B(ecl_sel_sum_e), .Y(exu_n26370));
INVX1 exu_U24217(.A(exu_n26370), .Y(exu_n7600));
AND2X1 exu_U24218(.A(exu_n11239), .B(exu_n15977), .Y(exu_n26374));
INVX1 exu_U24219(.A(exu_n26374), .Y(exu_n7601));
AND2X1 exu_U24220(.A(exu_ifu_brpc_e[6]), .B(exu_n16155), .Y(exu_n26376));
INVX1 exu_U24221(.A(exu_n26376), .Y(exu_n7602));
AND2X1 exu_U24222(.A(exu_n11241), .B(exu_n15977), .Y(exu_n26380));
INVX1 exu_U24223(.A(exu_n26380), .Y(exu_n7603));
AND2X1 exu_U24224(.A(exu_n11243), .B(exu_n15977), .Y(exu_n26385));
INVX1 exu_U24225(.A(exu_n26385), .Y(exu_n7604));
AND2X1 exu_U24226(.A(alu_adder_out[62]), .B(exu_n16157), .Y(exu_n26387));
INVX1 exu_U24227(.A(exu_n26387), .Y(exu_n7605));
AND2X1 exu_U24228(.A(exu_n11245), .B(exu_n15977), .Y(exu_n26391));
INVX1 exu_U24229(.A(exu_n26391), .Y(exu_n7606));
AND2X1 exu_U24230(.A(alu_adder_out[61]), .B(exu_n16158), .Y(exu_n26393));
INVX1 exu_U24231(.A(exu_n26393), .Y(exu_n7607));
AND2X1 exu_U24232(.A(exu_n11247), .B(exu_n15977), .Y(exu_n26397));
INVX1 exu_U24233(.A(exu_n26397), .Y(exu_n7608));
AND2X1 exu_U24234(.A(alu_adder_out[60]), .B(exu_n16157), .Y(exu_n26399));
INVX1 exu_U24235(.A(exu_n26399), .Y(exu_n7609));
AND2X1 exu_U24236(.A(exu_n11249), .B(exu_n15977), .Y(exu_n26403));
INVX1 exu_U24237(.A(exu_n26403), .Y(exu_n7610));
AND2X1 exu_U24238(.A(exu_ifu_brpc_e[5]), .B(exu_n16158), .Y(exu_n26405));
INVX1 exu_U24239(.A(exu_n26405), .Y(exu_n7611));
AND2X1 exu_U24240(.A(exu_n11251), .B(exu_n15977), .Y(exu_n26409));
INVX1 exu_U24241(.A(exu_n26409), .Y(exu_n7612));
AND2X1 exu_U24242(.A(alu_adder_out[59]), .B(exu_n16157), .Y(exu_n26411));
INVX1 exu_U24243(.A(exu_n26411), .Y(exu_n7613));
AND2X1 exu_U24244(.A(exu_n11253), .B(exu_n15977), .Y(exu_n26415));
INVX1 exu_U24245(.A(exu_n26415), .Y(exu_n7614));
AND2X1 exu_U24246(.A(alu_adder_out[58]), .B(exu_n16155), .Y(exu_n26417));
INVX1 exu_U24247(.A(exu_n26417), .Y(exu_n7615));
AND2X1 exu_U24248(.A(exu_n11255), .B(exu_n15977), .Y(exu_n26421));
INVX1 exu_U24249(.A(exu_n26421), .Y(exu_n7616));
AND2X1 exu_U24250(.A(alu_adder_out[57]), .B(exu_n16158), .Y(exu_n26423));
INVX1 exu_U24251(.A(exu_n26423), .Y(exu_n7617));
AND2X1 exu_U24252(.A(exu_n11257), .B(exu_n15977), .Y(exu_n26427));
INVX1 exu_U24253(.A(exu_n26427), .Y(exu_n7618));
AND2X1 exu_U24254(.A(alu_adder_out[56]), .B(ecl_sel_sum_e), .Y(exu_n26429));
INVX1 exu_U24255(.A(exu_n26429), .Y(exu_n7619));
AND2X1 exu_U24256(.A(exu_n11259), .B(exu_n15977), .Y(exu_n26433));
INVX1 exu_U24257(.A(exu_n26433), .Y(exu_n7620));
AND2X1 exu_U24258(.A(alu_adder_out[55]), .B(exu_n16155), .Y(exu_n26435));
INVX1 exu_U24259(.A(exu_n26435), .Y(exu_n7621));
AND2X1 exu_U24260(.A(exu_n11261), .B(exu_n15977), .Y(exu_n26439));
INVX1 exu_U24261(.A(exu_n26439), .Y(exu_n7622));
AND2X1 exu_U24262(.A(alu_adder_out[54]), .B(exu_n16158), .Y(exu_n26441));
INVX1 exu_U24263(.A(exu_n26441), .Y(exu_n7623));
AND2X1 exu_U24264(.A(exu_n11263), .B(exu_n15977), .Y(exu_n26445));
INVX1 exu_U24265(.A(exu_n26445), .Y(exu_n7624));
AND2X1 exu_U24266(.A(alu_adder_out[53]), .B(exu_n16158), .Y(exu_n26447));
INVX1 exu_U24267(.A(exu_n26447), .Y(exu_n7625));
AND2X1 exu_U24268(.A(exu_n11265), .B(exu_n15977), .Y(exu_n26451));
INVX1 exu_U24269(.A(exu_n26451), .Y(exu_n7626));
AND2X1 exu_U24270(.A(alu_adder_out[52]), .B(ecl_sel_sum_e), .Y(exu_n26453));
INVX1 exu_U24271(.A(exu_n26453), .Y(exu_n7627));
AND2X1 exu_U24272(.A(exu_n11267), .B(exu_n15977), .Y(exu_n26457));
INVX1 exu_U24273(.A(exu_n26457), .Y(exu_n7628));
AND2X1 exu_U24274(.A(alu_adder_out[51]), .B(exu_n16155), .Y(exu_n26459));
INVX1 exu_U24275(.A(exu_n26459), .Y(exu_n7629));
AND2X1 exu_U24276(.A(exu_n11269), .B(exu_n15977), .Y(exu_n26463));
INVX1 exu_U24277(.A(exu_n26463), .Y(exu_n7630));
AND2X1 exu_U24278(.A(alu_adder_out[50]), .B(exu_n16157), .Y(exu_n26465));
INVX1 exu_U24279(.A(exu_n26465), .Y(exu_n7631));
AND2X1 exu_U24280(.A(exu_n11271), .B(exu_n15977), .Y(exu_n26469));
INVX1 exu_U24281(.A(exu_n26469), .Y(exu_n7632));
AND2X1 exu_U24282(.A(exu_ifu_brpc_e[4]), .B(exu_n16158), .Y(exu_n26471));
INVX1 exu_U24283(.A(exu_n26471), .Y(exu_n7633));
AND2X1 exu_U24284(.A(exu_n11273), .B(exu_n15977), .Y(exu_n26475));
INVX1 exu_U24285(.A(exu_n26475), .Y(exu_n7634));
AND2X1 exu_U24286(.A(alu_adder_out[49]), .B(ecl_sel_sum_e), .Y(exu_n26477));
INVX1 exu_U24287(.A(exu_n26477), .Y(exu_n7635));
AND2X1 exu_U24288(.A(exu_n11275), .B(exu_n15977), .Y(exu_n26481));
INVX1 exu_U24289(.A(exu_n26481), .Y(exu_n7636));
AND2X1 exu_U24290(.A(alu_adder_out[48]), .B(ecl_sel_sum_e), .Y(exu_n26483));
INVX1 exu_U24291(.A(exu_n26483), .Y(exu_n7637));
AND2X1 exu_U24292(.A(exu_n11277), .B(exu_n15977), .Y(exu_n26487));
INVX1 exu_U24293(.A(exu_n26487), .Y(exu_n7638));
AND2X1 exu_U24294(.A(exu_ifu_brpc_e[47]), .B(exu_n16155), .Y(exu_n26489));
INVX1 exu_U24295(.A(exu_n26489), .Y(exu_n7639));
AND2X1 exu_U24296(.A(exu_n11279), .B(exu_n15977), .Y(exu_n26493));
INVX1 exu_U24297(.A(exu_n26493), .Y(exu_n7640));
AND2X1 exu_U24298(.A(exu_ifu_brpc_e[46]), .B(exu_n16157), .Y(exu_n26495));
INVX1 exu_U24299(.A(exu_n26495), .Y(exu_n7641));
AND2X1 exu_U24300(.A(exu_n11281), .B(exu_n15977), .Y(exu_n26499));
INVX1 exu_U24301(.A(exu_n26499), .Y(exu_n7642));
AND2X1 exu_U24302(.A(exu_ifu_brpc_e[45]), .B(exu_n16158), .Y(exu_n26501));
INVX1 exu_U24303(.A(exu_n26501), .Y(exu_n7643));
AND2X1 exu_U24304(.A(exu_n11283), .B(exu_n15977), .Y(exu_n26505));
INVX1 exu_U24305(.A(exu_n26505), .Y(exu_n7644));
AND2X1 exu_U24306(.A(exu_ifu_brpc_e[44]), .B(exu_n16155), .Y(exu_n26507));
INVX1 exu_U24307(.A(exu_n26507), .Y(exu_n7645));
AND2X1 exu_U24308(.A(exu_n11285), .B(exu_n15977), .Y(exu_n26511));
INVX1 exu_U24309(.A(exu_n26511), .Y(exu_n7646));
AND2X1 exu_U24310(.A(exu_ifu_brpc_e[43]), .B(ecl_sel_sum_e), .Y(exu_n26513));
INVX1 exu_U24311(.A(exu_n26513), .Y(exu_n7647));
AND2X1 exu_U24312(.A(exu_n11287), .B(exu_n15977), .Y(exu_n26517));
INVX1 exu_U24313(.A(exu_n26517), .Y(exu_n7648));
AND2X1 exu_U24314(.A(exu_ifu_brpc_e[42]), .B(exu_n16155), .Y(exu_n26519));
INVX1 exu_U24315(.A(exu_n26519), .Y(exu_n7649));
AND2X1 exu_U24316(.A(exu_n11289), .B(exu_n15977), .Y(exu_n26523));
INVX1 exu_U24317(.A(exu_n26523), .Y(exu_n7650));
AND2X1 exu_U24318(.A(exu_ifu_brpc_e[41]), .B(exu_n16157), .Y(exu_n26525));
INVX1 exu_U24319(.A(exu_n26525), .Y(exu_n7651));
AND2X1 exu_U24320(.A(exu_n11291), .B(exu_n15977), .Y(exu_n26529));
INVX1 exu_U24321(.A(exu_n26529), .Y(exu_n7652));
AND2X1 exu_U24322(.A(exu_ifu_brpc_e[40]), .B(exu_n16155), .Y(exu_n26531));
INVX1 exu_U24323(.A(exu_n26531), .Y(exu_n7653));
AND2X1 exu_U24324(.A(exu_n11293), .B(exu_n15977), .Y(exu_n26535));
INVX1 exu_U24325(.A(exu_n26535), .Y(exu_n7654));
AND2X1 exu_U24326(.A(exu_ifu_brpc_e[3]), .B(ecl_sel_sum_e), .Y(exu_n26537));
INVX1 exu_U24327(.A(exu_n26537), .Y(exu_n7655));
AND2X1 exu_U24328(.A(exu_n11295), .B(exu_n15977), .Y(exu_n26541));
INVX1 exu_U24329(.A(exu_n26541), .Y(exu_n7656));
AND2X1 exu_U24330(.A(exu_ifu_brpc_e[39]), .B(exu_n16155), .Y(exu_n26543));
INVX1 exu_U24331(.A(exu_n26543), .Y(exu_n7657));
AND2X1 exu_U24332(.A(exu_n11297), .B(exu_n15977), .Y(exu_n26547));
INVX1 exu_U24333(.A(exu_n26547), .Y(exu_n7658));
AND2X1 exu_U24334(.A(exu_ifu_brpc_e[38]), .B(exu_n16157), .Y(exu_n26549));
INVX1 exu_U24335(.A(exu_n26549), .Y(exu_n7659));
AND2X1 exu_U24336(.A(exu_n11299), .B(exu_n15977), .Y(exu_n26553));
INVX1 exu_U24337(.A(exu_n26553), .Y(exu_n7660));
AND2X1 exu_U24338(.A(exu_ifu_brpc_e[37]), .B(exu_n16158), .Y(exu_n26555));
INVX1 exu_U24339(.A(exu_n26555), .Y(exu_n7661));
AND2X1 exu_U24340(.A(exu_n11301), .B(exu_n15977), .Y(exu_n26559));
INVX1 exu_U24341(.A(exu_n26559), .Y(exu_n7662));
AND2X1 exu_U24342(.A(exu_ifu_brpc_e[36]), .B(exu_n16158), .Y(exu_n26561));
INVX1 exu_U24343(.A(exu_n26561), .Y(exu_n7663));
AND2X1 exu_U24344(.A(exu_n11303), .B(exu_n15977), .Y(exu_n26565));
INVX1 exu_U24345(.A(exu_n26565), .Y(exu_n7664));
AND2X1 exu_U24346(.A(exu_ifu_brpc_e[35]), .B(exu_n16157), .Y(exu_n26567));
INVX1 exu_U24347(.A(exu_n26567), .Y(exu_n7665));
AND2X1 exu_U24348(.A(exu_n11305), .B(exu_n15977), .Y(exu_n26571));
INVX1 exu_U24349(.A(exu_n26571), .Y(exu_n7666));
AND2X1 exu_U24350(.A(exu_ifu_brpc_e[34]), .B(ecl_sel_sum_e), .Y(exu_n26573));
INVX1 exu_U24351(.A(exu_n26573), .Y(exu_n7667));
AND2X1 exu_U24352(.A(exu_n11307), .B(exu_n15977), .Y(exu_n26577));
INVX1 exu_U24353(.A(exu_n26577), .Y(exu_n7668));
AND2X1 exu_U24354(.A(exu_ifu_brpc_e[33]), .B(exu_n16155), .Y(exu_n26579));
INVX1 exu_U24355(.A(exu_n26579), .Y(exu_n7669));
AND2X1 exu_U24356(.A(exu_n11309), .B(exu_n15977), .Y(exu_n26583));
INVX1 exu_U24357(.A(exu_n26583), .Y(exu_n7670));
AND2X1 exu_U24358(.A(exu_ifu_brpc_e[32]), .B(exu_n16157), .Y(exu_n26585));
INVX1 exu_U24359(.A(exu_n26585), .Y(exu_n7671));
AND2X1 exu_U24360(.A(exu_n11311), .B(exu_n15977), .Y(exu_n26589));
INVX1 exu_U24361(.A(exu_n26589), .Y(exu_n7672));
AND2X1 exu_U24362(.A(exu_n11313), .B(exu_n15977), .Y(exu_n26594));
INVX1 exu_U24363(.A(exu_n26594), .Y(exu_n7673));
AND2X1 exu_U24364(.A(exu_ifu_brpc_e[30]), .B(exu_n16158), .Y(exu_n26596));
INVX1 exu_U24365(.A(exu_n26596), .Y(exu_n7674));
AND2X1 exu_U24366(.A(exu_n11315), .B(exu_n15977), .Y(exu_n26600));
INVX1 exu_U24367(.A(exu_n26600), .Y(exu_n7675));
AND2X1 exu_U24368(.A(exu_ifu_brpc_e[2]), .B(ecl_sel_sum_e), .Y(exu_n26602));
INVX1 exu_U24369(.A(exu_n26602), .Y(exu_n7676));
AND2X1 exu_U24370(.A(exu_n11317), .B(exu_n15977), .Y(exu_n26606));
INVX1 exu_U24371(.A(exu_n26606), .Y(exu_n7677));
AND2X1 exu_U24372(.A(exu_ifu_brpc_e[29]), .B(exu_n16158), .Y(exu_n26608));
INVX1 exu_U24373(.A(exu_n26608), .Y(exu_n7678));
AND2X1 exu_U24374(.A(exu_n11319), .B(exu_n15977), .Y(exu_n26612));
INVX1 exu_U24375(.A(exu_n26612), .Y(exu_n7679));
AND2X1 exu_U24376(.A(exu_ifu_brpc_e[28]), .B(ecl_sel_sum_e), .Y(exu_n26614));
INVX1 exu_U24377(.A(exu_n26614), .Y(exu_n7680));
AND2X1 exu_U24378(.A(exu_n11321), .B(exu_n15977), .Y(exu_n26618));
INVX1 exu_U24379(.A(exu_n26618), .Y(exu_n7681));
AND2X1 exu_U24380(.A(exu_ifu_brpc_e[27]), .B(exu_n16155), .Y(exu_n26620));
INVX1 exu_U24381(.A(exu_n26620), .Y(exu_n7682));
AND2X1 exu_U24382(.A(exu_n11323), .B(exu_n15977), .Y(exu_n26624));
INVX1 exu_U24383(.A(exu_n26624), .Y(exu_n7683));
AND2X1 exu_U24384(.A(exu_ifu_brpc_e[26]), .B(exu_n16157), .Y(exu_n26626));
INVX1 exu_U24385(.A(exu_n26626), .Y(exu_n7684));
AND2X1 exu_U24386(.A(exu_n11325), .B(exu_n15977), .Y(exu_n26630));
INVX1 exu_U24387(.A(exu_n26630), .Y(exu_n7685));
AND2X1 exu_U24388(.A(exu_ifu_brpc_e[25]), .B(exu_n16158), .Y(exu_n26632));
INVX1 exu_U24389(.A(exu_n26632), .Y(exu_n7686));
AND2X1 exu_U24390(.A(exu_n11327), .B(exu_n15977), .Y(exu_n26636));
INVX1 exu_U24391(.A(exu_n26636), .Y(exu_n7687));
AND2X1 exu_U24392(.A(exu_ifu_brpc_e[24]), .B(ecl_sel_sum_e), .Y(exu_n26638));
INVX1 exu_U24393(.A(exu_n26638), .Y(exu_n7688));
AND2X1 exu_U24394(.A(exu_n11329), .B(exu_n15977), .Y(exu_n26642));
INVX1 exu_U24395(.A(exu_n26642), .Y(exu_n7689));
AND2X1 exu_U24396(.A(exu_ifu_brpc_e[23]), .B(exu_n16155), .Y(exu_n26644));
INVX1 exu_U24397(.A(exu_n26644), .Y(exu_n7690));
AND2X1 exu_U24398(.A(exu_n11331), .B(exu_n15977), .Y(exu_n26648));
INVX1 exu_U24399(.A(exu_n26648), .Y(exu_n7691));
AND2X1 exu_U24400(.A(exu_ifu_brpc_e[22]), .B(exu_n16157), .Y(exu_n26650));
INVX1 exu_U24401(.A(exu_n26650), .Y(exu_n7692));
AND2X1 exu_U24402(.A(exu_n11333), .B(exu_n15977), .Y(exu_n26654));
INVX1 exu_U24403(.A(exu_n26654), .Y(exu_n7693));
AND2X1 exu_U24404(.A(exu_ifu_brpc_e[21]), .B(exu_n16158), .Y(exu_n26656));
INVX1 exu_U24405(.A(exu_n26656), .Y(exu_n7694));
AND2X1 exu_U24406(.A(exu_n11335), .B(exu_n15977), .Y(exu_n26660));
INVX1 exu_U24407(.A(exu_n26660), .Y(exu_n7695));
AND2X1 exu_U24408(.A(exu_ifu_brpc_e[20]), .B(ecl_sel_sum_e), .Y(exu_n26662));
INVX1 exu_U24409(.A(exu_n26662), .Y(exu_n7696));
AND2X1 exu_U24410(.A(exu_n11337), .B(exu_n15977), .Y(exu_n26666));
INVX1 exu_U24411(.A(exu_n26666), .Y(exu_n7697));
AND2X1 exu_U24412(.A(exu_ifu_brpc_e[1]), .B(exu_n16155), .Y(exu_n26668));
INVX1 exu_U24413(.A(exu_n26668), .Y(exu_n7698));
AND2X1 exu_U24414(.A(exu_n11339), .B(exu_n15977), .Y(exu_n26672));
INVX1 exu_U24415(.A(exu_n26672), .Y(exu_n7699));
AND2X1 exu_U24416(.A(exu_ifu_brpc_e[19]), .B(exu_n16157), .Y(exu_n26674));
INVX1 exu_U24417(.A(exu_n26674), .Y(exu_n7700));
AND2X1 exu_U24418(.A(exu_n11341), .B(exu_n15977), .Y(exu_n26678));
INVX1 exu_U24419(.A(exu_n26678), .Y(exu_n7701));
AND2X1 exu_U24420(.A(exu_ifu_brpc_e[18]), .B(exu_n16158), .Y(exu_n26680));
INVX1 exu_U24421(.A(exu_n26680), .Y(exu_n7702));
AND2X1 exu_U24422(.A(exu_n11343), .B(exu_n15977), .Y(exu_n26684));
INVX1 exu_U24423(.A(exu_n26684), .Y(exu_n7703));
AND2X1 exu_U24424(.A(exu_ifu_brpc_e[17]), .B(ecl_sel_sum_e), .Y(exu_n26686));
INVX1 exu_U24425(.A(exu_n26686), .Y(exu_n7704));
AND2X1 exu_U24426(.A(exu_n11345), .B(exu_n15977), .Y(exu_n26690));
INVX1 exu_U24427(.A(exu_n26690), .Y(exu_n7705));
AND2X1 exu_U24428(.A(exu_ifu_brpc_e[16]), .B(exu_n16155), .Y(exu_n26692));
INVX1 exu_U24429(.A(exu_n26692), .Y(exu_n7706));
AND2X1 exu_U24430(.A(exu_n11347), .B(exu_n15977), .Y(exu_n26696));
INVX1 exu_U24431(.A(exu_n26696), .Y(exu_n7707));
AND2X1 exu_U24432(.A(exu_ifu_brpc_e[15]), .B(ecl_sel_sum_e), .Y(exu_n26698));
INVX1 exu_U24433(.A(exu_n26698), .Y(exu_n7708));
AND2X1 exu_U24434(.A(exu_n11349), .B(exu_n15977), .Y(exu_n26702));
INVX1 exu_U24435(.A(exu_n26702), .Y(exu_n7709));
AND2X1 exu_U24436(.A(exu_ifu_brpc_e[14]), .B(exu_n16155), .Y(exu_n26704));
INVX1 exu_U24437(.A(exu_n26704), .Y(exu_n7710));
AND2X1 exu_U24438(.A(exu_n11351), .B(exu_n15977), .Y(exu_n26708));
INVX1 exu_U24439(.A(exu_n26708), .Y(exu_n7711));
AND2X1 exu_U24440(.A(exu_ifu_brpc_e[13]), .B(ecl_sel_sum_e), .Y(exu_n26710));
INVX1 exu_U24441(.A(exu_n26710), .Y(exu_n7712));
AND2X1 exu_U24442(.A(exu_n11353), .B(exu_n15977), .Y(exu_n26714));
INVX1 exu_U24443(.A(exu_n26714), .Y(exu_n7713));
AND2X1 exu_U24444(.A(exu_ifu_brpc_e[12]), .B(ecl_sel_sum_e), .Y(exu_n26716));
INVX1 exu_U24445(.A(exu_n26716), .Y(exu_n7714));
AND2X1 exu_U24446(.A(exu_n11355), .B(exu_n15977), .Y(exu_n26720));
INVX1 exu_U24447(.A(exu_n26720), .Y(exu_n7715));
AND2X1 exu_U24448(.A(exu_ifu_brpc_e[11]), .B(exu_n16155), .Y(exu_n26722));
INVX1 exu_U24449(.A(exu_n26722), .Y(exu_n7716));
AND2X1 exu_U24450(.A(exu_n11357), .B(exu_n15977), .Y(exu_n26726));
INVX1 exu_U24451(.A(exu_n26726), .Y(exu_n7717));
AND2X1 exu_U24452(.A(exu_ifu_brpc_e[10]), .B(exu_n16155), .Y(exu_n26728));
INVX1 exu_U24453(.A(exu_n26728), .Y(exu_n7718));
AND2X1 exu_U24454(.A(exu_n11359), .B(exu_n15977), .Y(exu_n26732));
INVX1 exu_U24455(.A(exu_n26732), .Y(exu_n7719));
AND2X1 exu_U24456(.A(exu_ifu_brpc_e[0]), .B(ecl_sel_sum_e), .Y(exu_n26734));
INVX1 exu_U24457(.A(exu_n26734), .Y(exu_n7720));
AND2X1 exu_U24458(.A(exu_n16146), .B(shft_rshifterinput_b1[25]), .Y(exu_n26737));
INVX1 exu_U24459(.A(exu_n26737), .Y(exu_n7721));
AND2X1 exu_U24460(.A(exu_n16144), .B(exu_n15694), .Y(exu_n26739));
INVX1 exu_U24461(.A(exu_n26739), .Y(exu_n7722));
AND2X1 exu_U24462(.A(exu_n15727), .B(exu_n16144), .Y(exu_n26743));
INVX1 exu_U24463(.A(exu_n26743), .Y(exu_n7723));
AND2X1 exu_U24464(.A(exu_n15728), .B(exu_n16143), .Y(exu_n26747));
INVX1 exu_U24465(.A(exu_n26747), .Y(exu_n7724));
AND2X1 exu_U24466(.A(exu_n15729), .B(exu_n16144), .Y(exu_n26751));
INVX1 exu_U24467(.A(exu_n26751), .Y(exu_n7725));
INVX1 exu_U24468(.A(exu_n7728), .Y(exu_n7726));
INVX1 exu_U24469(.A(exu_n7726), .Y(exu_n7727));
AND2X1 exu_U24470(.A(exu_n16187), .B(exu_n16143), .Y(exu_n26755));
INVX1 exu_U24471(.A(exu_n26755), .Y(exu_n7728));
INVX1 exu_U24472(.A(exu_n7735), .Y(exu_n7729));
INVX1 exu_U24473(.A(exu_n7729), .Y(exu_n7730));
INVX1 exu_U24474(.A(exu_n7733), .Y(exu_n7731));
INVX1 exu_U24475(.A(exu_n7731), .Y(exu_n7732));
AND2X1 exu_U24476(.A(exu_n16187), .B(exu_n16144), .Y(exu_n26759));
INVX1 exu_U24477(.A(exu_n26759), .Y(exu_n7733));
INVX1 exu_U24478(.A(exu_n7777), .Y(exu_n7734));
INVX1 exu_U24479(.A(exu_n7734), .Y(exu_n7735));
INVX1 exu_U24480(.A(exu_n7738), .Y(exu_n7736));
INVX1 exu_U24481(.A(exu_n7736), .Y(exu_n7737));
AND2X1 exu_U24482(.A(exu_n16187), .B(exu_n16143), .Y(exu_n26763));
INVX1 exu_U24483(.A(exu_n26763), .Y(exu_n7738));
INVX1 exu_U24484(.A(exu_n7741), .Y(exu_n7739));
INVX1 exu_U24485(.A(exu_n7739), .Y(exu_n7740));
AND2X1 exu_U24486(.A(exu_n16187), .B(exu_n15399), .Y(exu_n26767));
INVX1 exu_U24487(.A(exu_n26767), .Y(exu_n7741));
AND2X1 exu_U24488(.A(exu_n15730), .B(exu_n16144), .Y(exu_n26771));
INVX1 exu_U24489(.A(exu_n26771), .Y(exu_n7742));
INVX1 exu_U24490(.A(exu_n7745), .Y(exu_n7743));
INVX1 exu_U24491(.A(exu_n7743), .Y(exu_n7744));
AND2X1 exu_U24492(.A(exu_n16187), .B(exu_n16143), .Y(exu_n26775));
INVX1 exu_U24493(.A(exu_n26775), .Y(exu_n7745));
INVX1 exu_U24494(.A(exu_n7748), .Y(exu_n7746));
INVX1 exu_U24495(.A(exu_n7746), .Y(exu_n7747));
AND2X1 exu_U24496(.A(exu_n16187), .B(exu_n16144), .Y(exu_n26779));
INVX1 exu_U24497(.A(exu_n26779), .Y(exu_n7748));
INVX1 exu_U24498(.A(exu_n7751), .Y(exu_n7749));
INVX1 exu_U24499(.A(exu_n7749), .Y(exu_n7750));
AND2X1 exu_U24500(.A(exu_n16187), .B(exu_n16142), .Y(exu_n26783));
INVX1 exu_U24501(.A(exu_n26783), .Y(exu_n7751));
INVX1 exu_U24502(.A(exu_n7754), .Y(exu_n7752));
INVX1 exu_U24503(.A(exu_n7752), .Y(exu_n7753));
AND2X1 exu_U24504(.A(exu_n16187), .B(exu_n16143), .Y(exu_n26787));
INVX1 exu_U24505(.A(exu_n26787), .Y(exu_n7754));
INVX1 exu_U24506(.A(exu_n7757), .Y(exu_n7755));
INVX1 exu_U24507(.A(exu_n7755), .Y(exu_n7756));
AND2X1 exu_U24508(.A(exu_n16187), .B(exu_n15399), .Y(exu_n26791));
INVX1 exu_U24509(.A(exu_n26791), .Y(exu_n7757));
INVX1 exu_U24510(.A(exu_n7760), .Y(exu_n7758));
INVX1 exu_U24511(.A(exu_n7758), .Y(exu_n7759));
AND2X1 exu_U24512(.A(exu_n16187), .B(exu_n16144), .Y(exu_n26795));
INVX1 exu_U24513(.A(exu_n26795), .Y(exu_n7760));
INVX1 exu_U24514(.A(exu_n7763), .Y(exu_n7761));
INVX1 exu_U24515(.A(exu_n7761), .Y(exu_n7762));
AND2X1 exu_U24516(.A(exu_n16187), .B(exu_n16142), .Y(exu_n26799));
INVX1 exu_U24517(.A(exu_n26799), .Y(exu_n7763));
INVX1 exu_U24518(.A(exu_n7766), .Y(exu_n7764));
INVX1 exu_U24519(.A(exu_n7764), .Y(exu_n7765));
AND2X1 exu_U24520(.A(exu_n16187), .B(exu_n16143), .Y(exu_n26803));
INVX1 exu_U24521(.A(exu_n26803), .Y(exu_n7766));
INVX1 exu_U24522(.A(exu_n7769), .Y(exu_n7767));
INVX1 exu_U24523(.A(exu_n7767), .Y(exu_n7768));
AND2X1 exu_U24524(.A(exu_n15403), .B(exu_n15399), .Y(exu_n26807));
INVX1 exu_U24525(.A(exu_n26807), .Y(exu_n7769));
INVX1 exu_U24526(.A(exu_n7772), .Y(exu_n7770));
INVX1 exu_U24527(.A(exu_n7770), .Y(exu_n7771));
AND2X1 exu_U24528(.A(exu_n16191), .B(exu_n16144), .Y(exu_n26811));
INVX1 exu_U24529(.A(exu_n26811), .Y(exu_n7772));
AND2X1 exu_U24530(.A(exu_n15731), .B(exu_n16142), .Y(exu_n26815));
INVX1 exu_U24531(.A(exu_n26815), .Y(exu_n7773));
INVX1 exu_U24532(.A(exu_n7776), .Y(exu_n7774));
INVX1 exu_U24533(.A(exu_n7774), .Y(exu_n7775));
AND2X1 exu_U24534(.A(exu_n16189), .B(exu_n16143), .Y(exu_n26819));
INVX1 exu_U24535(.A(exu_n26819), .Y(exu_n7776));
AND2X1 exu_U24536(.A(exu_n16189), .B(exu_n16146), .Y(exu_n26823));
INVX1 exu_U24537(.A(exu_n26823), .Y(exu_n7777));
INVX1 exu_U24538(.A(exu_n7780), .Y(exu_n7778));
INVX1 exu_U24539(.A(exu_n7778), .Y(exu_n7779));
AND2X1 exu_U24540(.A(exu_n15403), .B(exu_n15399), .Y(exu_n26824));
INVX1 exu_U24541(.A(exu_n26824), .Y(exu_n7780));
AND2X1 exu_U24542(.A(exu_n15721), .B(exu_n16146), .Y(exu_n26828));
INVX1 exu_U24543(.A(exu_n26828), .Y(exu_n7781));
INVX1 exu_U24544(.A(exu_n7784), .Y(exu_n7782));
INVX1 exu_U24545(.A(exu_n7782), .Y(exu_n7783));
AND2X1 exu_U24546(.A(exu_n16191), .B(exu_n16144), .Y(exu_n26829));
INVX1 exu_U24547(.A(exu_n26829), .Y(exu_n7784));
AND2X1 exu_U24548(.A(exu_n15722), .B(exu_n16146), .Y(exu_n26833));
INVX1 exu_U24549(.A(exu_n26833), .Y(exu_n7785));
INVX1 exu_U24550(.A(exu_n7788), .Y(exu_n7786));
INVX1 exu_U24551(.A(exu_n7786), .Y(exu_n7787));
AND2X1 exu_U24552(.A(exu_n16189), .B(exu_n16142), .Y(exu_n26834));
INVX1 exu_U24553(.A(exu_n26834), .Y(exu_n7788));
AND2X1 exu_U24554(.A(exu_n15723), .B(exu_n16146), .Y(exu_n26838));
INVX1 exu_U24555(.A(exu_n26838), .Y(exu_n7789));
INVX1 exu_U24556(.A(exu_n7792), .Y(exu_n7790));
INVX1 exu_U24557(.A(exu_n7790), .Y(exu_n7791));
AND2X1 exu_U24558(.A(exu_n15403), .B(exu_n16142), .Y(exu_n26839));
INVX1 exu_U24559(.A(exu_n26839), .Y(exu_n7792));
AND2X1 exu_U24560(.A(exu_n15724), .B(exu_n16146), .Y(exu_n26843));
INVX1 exu_U24561(.A(exu_n26843), .Y(exu_n7793));
INVX1 exu_U24562(.A(exu_n7796), .Y(exu_n7794));
INVX1 exu_U24563(.A(exu_n7794), .Y(exu_n7795));
AND2X1 exu_U24564(.A(exu_n16191), .B(exu_n16142), .Y(exu_n26844));
INVX1 exu_U24565(.A(exu_n26844), .Y(exu_n7796));
AND2X1 exu_U24566(.A(exu_n15725), .B(exu_n16146), .Y(exu_n26848));
INVX1 exu_U24567(.A(exu_n26848), .Y(exu_n7797));
INVX1 exu_U24568(.A(exu_n7800), .Y(exu_n7798));
INVX1 exu_U24569(.A(exu_n7798), .Y(exu_n7799));
AND2X1 exu_U24570(.A(exu_n16189), .B(exu_n16142), .Y(exu_n26849));
INVX1 exu_U24571(.A(exu_n26849), .Y(exu_n7800));
AND2X1 exu_U24572(.A(exu_n15726), .B(shft_shift16_e[1]), .Y(exu_n26853));
INVX1 exu_U24573(.A(exu_n26853), .Y(exu_n7801));
INVX1 exu_U24574(.A(exu_n7804), .Y(exu_n7802));
INVX1 exu_U24575(.A(exu_n7802), .Y(exu_n7803));
AND2X1 exu_U24576(.A(exu_n16190), .B(exu_n16142), .Y(exu_n26854));
INVX1 exu_U24577(.A(exu_n26854), .Y(exu_n7804));
AND2X1 exu_U24578(.A(exu_n15694), .B(exu_n16146), .Y(exu_n26858));
INVX1 exu_U24579(.A(exu_n26858), .Y(exu_n7805));
INVX1 exu_U24580(.A(exu_n7808), .Y(exu_n7806));
INVX1 exu_U24581(.A(exu_n7806), .Y(exu_n7807));
AND2X1 exu_U24582(.A(exu_n15403), .B(exu_n16142), .Y(exu_n26859));
INVX1 exu_U24583(.A(exu_n26859), .Y(exu_n7808));
AND2X1 exu_U24584(.A(exu_n15727), .B(shft_shift16_e[1]), .Y(exu_n26863));
INVX1 exu_U24585(.A(exu_n26863), .Y(exu_n7809));
INVX1 exu_U24586(.A(exu_n7812), .Y(exu_n7810));
INVX1 exu_U24587(.A(exu_n7810), .Y(exu_n7811));
AND2X1 exu_U24588(.A(exu_n16191), .B(exu_n16142), .Y(exu_n26864));
INVX1 exu_U24589(.A(exu_n26864), .Y(exu_n7812));
AND2X1 exu_U24590(.A(exu_n15732), .B(exu_n16142), .Y(exu_n26868));
INVX1 exu_U24591(.A(exu_n26868), .Y(exu_n7813));
AND2X1 exu_U24592(.A(exu_n15728), .B(exu_n16146), .Y(exu_n26872));
INVX1 exu_U24593(.A(exu_n26872), .Y(exu_n7814));
INVX1 exu_U24594(.A(exu_n7817), .Y(exu_n7815));
INVX1 exu_U24595(.A(exu_n7815), .Y(exu_n7816));
AND2X1 exu_U24596(.A(exu_n16188), .B(exu_n16142), .Y(exu_n26873));
INVX1 exu_U24597(.A(exu_n26873), .Y(exu_n7817));
AND2X1 exu_U24598(.A(exu_n15729), .B(shft_shift16_e[1]), .Y(exu_n26877));
INVX1 exu_U24599(.A(exu_n26877), .Y(exu_n7818));
INVX1 exu_U24600(.A(exu_n7821), .Y(exu_n7819));
INVX1 exu_U24601(.A(exu_n7819), .Y(exu_n7820));
AND2X1 exu_U24602(.A(exu_n16188), .B(exu_n16142), .Y(exu_n26878));
INVX1 exu_U24603(.A(exu_n26878), .Y(exu_n7821));
AND2X1 exu_U24604(.A(exu_n15730), .B(exu_n16146), .Y(exu_n26882));
INVX1 exu_U24605(.A(exu_n26882), .Y(exu_n7822));
INVX1 exu_U24606(.A(exu_n7825), .Y(exu_n7823));
INVX1 exu_U24607(.A(exu_n7823), .Y(exu_n7824));
AND2X1 exu_U24608(.A(exu_n16188), .B(exu_n16142), .Y(exu_n26883));
INVX1 exu_U24609(.A(exu_n26883), .Y(exu_n7825));
AND2X1 exu_U24610(.A(exu_n15731), .B(shft_shift16_e[1]), .Y(exu_n26887));
INVX1 exu_U24611(.A(exu_n26887), .Y(exu_n7826));
INVX1 exu_U24612(.A(exu_n7829), .Y(exu_n7827));
INVX1 exu_U24613(.A(exu_n7827), .Y(exu_n7828));
AND2X1 exu_U24614(.A(exu_n16188), .B(exu_n16142), .Y(exu_n26888));
INVX1 exu_U24615(.A(exu_n26888), .Y(exu_n7829));
AND2X1 exu_U24616(.A(exu_n15732), .B(exu_n16146), .Y(exu_n26892));
INVX1 exu_U24617(.A(exu_n26892), .Y(exu_n7830));
INVX1 exu_U24618(.A(exu_n7833), .Y(exu_n7831));
INVX1 exu_U24619(.A(exu_n7831), .Y(exu_n7832));
AND2X1 exu_U24620(.A(exu_n16188), .B(exu_n16143), .Y(exu_n26893));
INVX1 exu_U24621(.A(exu_n26893), .Y(exu_n7833));
AND2X1 exu_U24622(.A(exu_n15733), .B(shft_shift16_e[1]), .Y(exu_n26897));
INVX1 exu_U24623(.A(exu_n26897), .Y(exu_n7834));
INVX1 exu_U24624(.A(exu_n7837), .Y(exu_n7835));
INVX1 exu_U24625(.A(exu_n7835), .Y(exu_n7836));
AND2X1 exu_U24626(.A(exu_n16188), .B(exu_n16143), .Y(exu_n26898));
INVX1 exu_U24627(.A(exu_n26898), .Y(exu_n7837));
AND2X1 exu_U24628(.A(exu_n15734), .B(exu_n16146), .Y(exu_n26902));
INVX1 exu_U24629(.A(exu_n26902), .Y(exu_n7838));
INVX1 exu_U24630(.A(exu_n7841), .Y(exu_n7839));
INVX1 exu_U24631(.A(exu_n7839), .Y(exu_n7840));
AND2X1 exu_U24632(.A(exu_n16188), .B(exu_n16143), .Y(exu_n26903));
INVX1 exu_U24633(.A(exu_n26903), .Y(exu_n7841));
AND2X1 exu_U24634(.A(exu_n15735), .B(shft_shift16_e[1]), .Y(exu_n26907));
INVX1 exu_U24635(.A(exu_n26907), .Y(exu_n7842));
INVX1 exu_U24636(.A(exu_n7845), .Y(exu_n7843));
INVX1 exu_U24637(.A(exu_n7843), .Y(exu_n7844));
AND2X1 exu_U24638(.A(exu_n16188), .B(exu_n16143), .Y(exu_n26909));
INVX1 exu_U24639(.A(exu_n26909), .Y(exu_n7845));
AND2X1 exu_U24640(.A(exu_n15450), .B(exu_n16146), .Y(exu_n26912));
INVX1 exu_U24641(.A(exu_n26912), .Y(exu_n7846));
AND2X1 exu_U24642(.A(exu_n15451), .B(shft_shift16_e[1]), .Y(exu_n26916));
INVX1 exu_U24643(.A(exu_n26916), .Y(exu_n7847));
AND2X1 exu_U24644(.A(exu_n15733), .B(exu_n16143), .Y(exu_n26921));
INVX1 exu_U24645(.A(exu_n26921), .Y(exu_n7848));
AND2X1 exu_U24646(.A(exu_n15452), .B(exu_n16146), .Y(exu_n26924));
INVX1 exu_U24647(.A(exu_n26924), .Y(exu_n7849));
AND2X1 exu_U24648(.A(exu_n15453), .B(shft_shift16_e[1]), .Y(exu_n26928));
INVX1 exu_U24649(.A(exu_n26928), .Y(exu_n7850));
AND2X1 exu_U24650(.A(exu_n15454), .B(shft_shift16_e[1]), .Y(exu_n26932));
INVX1 exu_U24651(.A(exu_n26932), .Y(exu_n7851));
AND2X1 exu_U24652(.A(exu_n15455), .B(exu_n16146), .Y(exu_n26936));
INVX1 exu_U24653(.A(exu_n26936), .Y(exu_n7852));
AND2X1 exu_U24654(.A(exu_n15438), .B(shft_shift16_e[1]), .Y(exu_n26940));
INVX1 exu_U24655(.A(exu_n26940), .Y(exu_n7853));
AND2X1 exu_U24656(.A(exu_n15442), .B(shft_shift16_e[1]), .Y(exu_n26944));
INVX1 exu_U24657(.A(exu_n26944), .Y(exu_n7854));
AND2X1 exu_U24658(.A(exu_n15443), .B(exu_n16146), .Y(exu_n26948));
INVX1 exu_U24659(.A(exu_n26948), .Y(exu_n7855));
AND2X1 exu_U24660(.A(exu_n15444), .B(exu_n16146), .Y(exu_n26952));
INVX1 exu_U24661(.A(exu_n26952), .Y(exu_n7856));
AND2X1 exu_U24662(.A(exu_n15445), .B(shft_shift16_e[1]), .Y(exu_n26956));
INVX1 exu_U24663(.A(exu_n26956), .Y(exu_n7857));
AND2X1 exu_U24664(.A(exu_n15446), .B(shft_shift16_e[1]), .Y(exu_n26960));
INVX1 exu_U24665(.A(exu_n26960), .Y(exu_n7858));
AND2X1 exu_U24666(.A(exu_n15734), .B(exu_n16144), .Y(exu_n26965));
INVX1 exu_U24667(.A(exu_n26965), .Y(exu_n7859));
AND2X1 exu_U24668(.A(exu_n15447), .B(exu_n16146), .Y(exu_n26968));
INVX1 exu_U24669(.A(exu_n26968), .Y(exu_n7860));
INVX1 exu_U24670(.A(exu_n7865), .Y(exu_n7861));
INVX1 exu_U24671(.A(exu_n7861), .Y(exu_n7862));
AND2X1 exu_U24672(.A(exu_n15448), .B(exu_n16146), .Y(exu_n26972));
INVX1 exu_U24673(.A(exu_n26972), .Y(exu_n7863));
INVX1 exu_U24674(.A(exu_n7868), .Y(exu_n7864));
INVX1 exu_U24675(.A(exu_n7864), .Y(exu_n7865));
AND2X1 exu_U24676(.A(exu_n15449), .B(exu_n16146), .Y(exu_n26976));
INVX1 exu_U24677(.A(exu_n26976), .Y(exu_n7866));
INVX1 exu_U24678(.A(exu_n7870), .Y(exu_n7867));
INVX1 exu_U24679(.A(exu_n7867), .Y(exu_n7868));
AND2X1 exu_U24680(.A(exu_n15456), .B(exu_n16146), .Y(exu_n26980));
INVX1 exu_U24681(.A(exu_n26980), .Y(exu_n7869));
AND2X1 exu_U24682(.A(exu_n15403), .B(exu_n16144), .Y(exu_n26982));
INVX1 exu_U24683(.A(exu_n26982), .Y(exu_n7870));
AND2X1 exu_U24684(.A(exu_n15721), .B(exu_n16144), .Y(exu_n26986));
INVX1 exu_U24685(.A(exu_n26986), .Y(exu_n7871));
AND2X1 exu_U24686(.A(exu_n15722), .B(exu_n16144), .Y(exu_n26990));
INVX1 exu_U24687(.A(exu_n26990), .Y(exu_n7872));
AND2X1 exu_U24688(.A(exu_n15723), .B(exu_n16144), .Y(exu_n26994));
INVX1 exu_U24689(.A(exu_n26994), .Y(exu_n7873));
AND2X1 exu_U24690(.A(exu_n15724), .B(exu_n16144), .Y(exu_n26998));
INVX1 exu_U24691(.A(exu_n26998), .Y(exu_n7874));
AND2X1 exu_U24692(.A(exu_n15725), .B(exu_n15399), .Y(exu_n27002));
INVX1 exu_U24693(.A(exu_n27002), .Y(exu_n7875));
AND2X1 exu_U24694(.A(exu_n15726), .B(exu_n15399), .Y(exu_n27006));
INVX1 exu_U24695(.A(exu_n27006), .Y(exu_n7876));
AND2X1 exu_U24696(.A(exu_n15735), .B(exu_n15399), .Y(exu_n27010));
INVX1 exu_U24697(.A(exu_n27010), .Y(exu_n7877));
AND2X1 exu_U24698(.A(exu_n15400), .B(shft_rshift16_b1[13]), .Y(exu_n27014));
INVX1 exu_U24699(.A(exu_n27014), .Y(exu_n7878));
AND2X1 exu_U24700(.A(exu_n16234), .B(shft_rshift16_b1[21]), .Y(exu_n27016));
INVX1 exu_U24701(.A(exu_n27016), .Y(exu_n7879));
AND2X1 exu_U24702(.A(shft_rshift16_b1[12]), .B(exu_n15400), .Y(exu_n27020));
INVX1 exu_U24703(.A(exu_n27020), .Y(exu_n7880));
AND2X1 exu_U24704(.A(shft_rshift16_b1[20]), .B(exu_n16234), .Y(exu_n27022));
INVX1 exu_U24705(.A(exu_n27022), .Y(exu_n7881));
AND2X1 exu_U24706(.A(shft_rshift16_b1[11]), .B(exu_n15400), .Y(exu_n27026));
INVX1 exu_U24707(.A(exu_n27026), .Y(exu_n7882));
AND2X1 exu_U24708(.A(shft_rshift16_b1[19]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27028));
INVX1 exu_U24709(.A(exu_n27028), .Y(exu_n7883));
AND2X1 exu_U24710(.A(shft_rshift16_b1[10]), .B(exu_n16231), .Y(exu_n27032));
INVX1 exu_U24711(.A(exu_n27032), .Y(exu_n7884));
AND2X1 exu_U24712(.A(shft_rshift16_b1[18]), .B(exu_n16234), .Y(exu_n27034));
INVX1 exu_U24713(.A(exu_n27034), .Y(exu_n7885));
AND2X1 exu_U24714(.A(exu_n16189), .B(exu_n16231), .Y(exu_n27046));
INVX1 exu_U24715(.A(exu_n27046), .Y(exu_n7886));
AND2X1 exu_U24716(.A(exu_n16190), .B(exu_n16234), .Y(exu_n27047));
INVX1 exu_U24717(.A(exu_n27047), .Y(exu_n7887));
AND2X1 exu_U24718(.A(shft_rshift16_b1[9]), .B(exu_n16231), .Y(exu_n27051));
INVX1 exu_U24719(.A(exu_n27051), .Y(exu_n7888));
AND2X1 exu_U24720(.A(shft_rshift16_b1[17]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27053));
INVX1 exu_U24721(.A(exu_n27053), .Y(exu_n7889));
AND2X1 exu_U24722(.A(shft_rshift16_b1[63]), .B(exu_n16231), .Y(exu_n27057));
INVX1 exu_U24723(.A(exu_n27057), .Y(exu_n7890));
AND2X1 exu_U24724(.A(exu_n16190), .B(exu_n16234), .Y(exu_n27058));
INVX1 exu_U24725(.A(exu_n27058), .Y(exu_n7891));
AND2X1 exu_U24726(.A(shft_rshift16_b1[62]), .B(exu_n15400), .Y(exu_n27062));
INVX1 exu_U24727(.A(exu_n27062), .Y(exu_n7892));
AND2X1 exu_U24728(.A(exu_n16190), .B(ecl_shft_shift4_e[3]), .Y(exu_n27063));
INVX1 exu_U24729(.A(exu_n27063), .Y(exu_n7893));
AND2X1 exu_U24730(.A(shft_rshift16_b1[61]), .B(exu_n16231), .Y(exu_n27066));
INVX1 exu_U24731(.A(exu_n27066), .Y(exu_n7894));
AND2X1 exu_U24732(.A(shft_rshift16_b1[60]), .B(exu_n15400), .Y(exu_n27070));
INVX1 exu_U24733(.A(exu_n27070), .Y(exu_n7895));
AND2X1 exu_U24734(.A(shft_rshift16_b1[59]), .B(exu_n16231), .Y(exu_n27075));
INVX1 exu_U24735(.A(exu_n27075), .Y(exu_n7896));
AND2X1 exu_U24736(.A(shft_rshift16_b1[58]), .B(exu_n15400), .Y(exu_n27080));
INVX1 exu_U24737(.A(exu_n27080), .Y(exu_n7897));
AND2X1 exu_U24738(.A(shft_rshift16_b1[57]), .B(exu_n16231), .Y(exu_n27085));
INVX1 exu_U24739(.A(exu_n27085), .Y(exu_n7898));
AND2X1 exu_U24740(.A(shft_rshift16_b1[56]), .B(exu_n15400), .Y(exu_n27090));
INVX1 exu_U24741(.A(exu_n27090), .Y(exu_n7899));
AND2X1 exu_U24742(.A(shft_rshift16_b1[55]), .B(exu_n15400), .Y(exu_n27095));
INVX1 exu_U24743(.A(exu_n27095), .Y(exu_n7900));
AND2X1 exu_U24744(.A(shft_rshift16_b1[63]), .B(exu_n16234), .Y(exu_n27097));
INVX1 exu_U24745(.A(exu_n27097), .Y(exu_n7901));
AND2X1 exu_U24746(.A(shft_rshift16_b1[54]), .B(exu_n16231), .Y(exu_n27101));
INVX1 exu_U24747(.A(exu_n27101), .Y(exu_n7902));
AND2X1 exu_U24748(.A(shft_rshift16_b1[62]), .B(exu_n16234), .Y(exu_n27103));
INVX1 exu_U24749(.A(exu_n27103), .Y(exu_n7903));
AND2X1 exu_U24750(.A(shft_rshift16_b1[8]), .B(exu_n15400), .Y(exu_n27107));
INVX1 exu_U24751(.A(exu_n27107), .Y(exu_n7904));
AND2X1 exu_U24752(.A(shft_rshift16_b1[16]), .B(exu_n16234), .Y(exu_n27109));
INVX1 exu_U24753(.A(exu_n27109), .Y(exu_n7905));
AND2X1 exu_U24754(.A(shft_rshift16_b1[53]), .B(exu_n16231), .Y(exu_n27113));
INVX1 exu_U24755(.A(exu_n27113), .Y(exu_n7906));
AND2X1 exu_U24756(.A(shft_rshift16_b1[61]), .B(exu_n16234), .Y(exu_n27115));
INVX1 exu_U24757(.A(exu_n27115), .Y(exu_n7907));
AND2X1 exu_U24758(.A(shft_rshift16_b1[52]), .B(exu_n15400), .Y(exu_n27119));
INVX1 exu_U24759(.A(exu_n27119), .Y(exu_n7908));
AND2X1 exu_U24760(.A(shft_rshift16_b1[60]), .B(exu_n16234), .Y(exu_n27121));
INVX1 exu_U24761(.A(exu_n27121), .Y(exu_n7909));
AND2X1 exu_U24762(.A(shft_rshift16_b1[51]), .B(exu_n16231), .Y(exu_n27125));
INVX1 exu_U24763(.A(exu_n27125), .Y(exu_n7910));
AND2X1 exu_U24764(.A(shft_rshift16_b1[59]), .B(exu_n16234), .Y(exu_n27127));
INVX1 exu_U24765(.A(exu_n27127), .Y(exu_n7911));
AND2X1 exu_U24766(.A(shft_rshift16_b1[50]), .B(exu_n16231), .Y(exu_n27131));
INVX1 exu_U24767(.A(exu_n27131), .Y(exu_n7912));
AND2X1 exu_U24768(.A(shft_rshift16_b1[58]), .B(exu_n16234), .Y(exu_n27133));
INVX1 exu_U24769(.A(exu_n27133), .Y(exu_n7913));
AND2X1 exu_U24770(.A(shft_rshift16_b1[49]), .B(exu_n15400), .Y(exu_n27137));
INVX1 exu_U24771(.A(exu_n27137), .Y(exu_n7914));
AND2X1 exu_U24772(.A(shft_rshift16_b1[57]), .B(exu_n16234), .Y(exu_n27139));
INVX1 exu_U24773(.A(exu_n27139), .Y(exu_n7915));
AND2X1 exu_U24774(.A(shft_rshift16_b1[48]), .B(exu_n15400), .Y(exu_n27143));
INVX1 exu_U24775(.A(exu_n27143), .Y(exu_n7916));
AND2X1 exu_U24776(.A(shft_rshift16_b1[56]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27145));
INVX1 exu_U24777(.A(exu_n27145), .Y(exu_n7917));
AND2X1 exu_U24778(.A(shft_rshift16_b1[47]), .B(exu_n15400), .Y(exu_n27149));
INVX1 exu_U24779(.A(exu_n27149), .Y(exu_n7918));
AND2X1 exu_U24780(.A(shft_rshift16_b1[55]), .B(exu_n16234), .Y(exu_n27151));
INVX1 exu_U24781(.A(exu_n27151), .Y(exu_n7919));
AND2X1 exu_U24782(.A(shft_rshift16_b1[46]), .B(exu_n15400), .Y(exu_n27155));
INVX1 exu_U24783(.A(exu_n27155), .Y(exu_n7920));
AND2X1 exu_U24784(.A(shft_rshift16_b1[54]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27157));
INVX1 exu_U24785(.A(exu_n27157), .Y(exu_n7921));
AND2X1 exu_U24786(.A(shft_rshift16_b1[45]), .B(exu_n16231), .Y(exu_n27161));
INVX1 exu_U24787(.A(exu_n27161), .Y(exu_n7922));
AND2X1 exu_U24788(.A(shft_rshift16_b1[53]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27163));
INVX1 exu_U24789(.A(exu_n27163), .Y(exu_n7923));
AND2X1 exu_U24790(.A(shft_rshift16_b1[44]), .B(exu_n15400), .Y(exu_n27167));
INVX1 exu_U24791(.A(exu_n27167), .Y(exu_n7924));
AND2X1 exu_U24792(.A(shft_rshift16_b1[52]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27169));
INVX1 exu_U24793(.A(exu_n27169), .Y(exu_n7925));
AND2X1 exu_U24794(.A(shft_rshift16_b1[7]), .B(exu_n15400), .Y(exu_n27173));
INVX1 exu_U24795(.A(exu_n27173), .Y(exu_n7926));
AND2X1 exu_U24796(.A(shft_rshift16_b1[15]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27175));
INVX1 exu_U24797(.A(exu_n27175), .Y(exu_n7927));
AND2X1 exu_U24798(.A(shft_rshift16_b1[43]), .B(exu_n16231), .Y(exu_n27179));
INVX1 exu_U24799(.A(exu_n27179), .Y(exu_n7928));
AND2X1 exu_U24800(.A(shft_rshift16_b1[51]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27181));
INVX1 exu_U24801(.A(exu_n27181), .Y(exu_n7929));
AND2X1 exu_U24802(.A(shft_rshift16_b1[42]), .B(exu_n15400), .Y(exu_n27185));
INVX1 exu_U24803(.A(exu_n27185), .Y(exu_n7930));
AND2X1 exu_U24804(.A(shft_rshift16_b1[50]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27187));
INVX1 exu_U24805(.A(exu_n27187), .Y(exu_n7931));
AND2X1 exu_U24806(.A(shft_rshift16_b1[41]), .B(exu_n16231), .Y(exu_n27191));
INVX1 exu_U24807(.A(exu_n27191), .Y(exu_n7932));
AND2X1 exu_U24808(.A(shft_rshift16_b1[49]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27193));
INVX1 exu_U24809(.A(exu_n27193), .Y(exu_n7933));
AND2X1 exu_U24810(.A(shft_rshift16_b1[40]), .B(exu_n15400), .Y(exu_n27197));
INVX1 exu_U24811(.A(exu_n27197), .Y(exu_n7934));
AND2X1 exu_U24812(.A(shft_rshift16_b1[48]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27199));
INVX1 exu_U24813(.A(exu_n27199), .Y(exu_n7935));
AND2X1 exu_U24814(.A(shft_rshift16_b1[39]), .B(exu_n16231), .Y(exu_n27203));
INVX1 exu_U24815(.A(exu_n27203), .Y(exu_n7936));
AND2X1 exu_U24816(.A(shft_rshift16_b1[47]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27205));
INVX1 exu_U24817(.A(exu_n27205), .Y(exu_n7937));
AND2X1 exu_U24818(.A(shft_rshift16_b1[38]), .B(exu_n15400), .Y(exu_n27209));
INVX1 exu_U24819(.A(exu_n27209), .Y(exu_n7938));
AND2X1 exu_U24820(.A(shft_rshift16_b1[46]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27211));
INVX1 exu_U24821(.A(exu_n27211), .Y(exu_n7939));
AND2X1 exu_U24822(.A(shft_rshift16_b1[37]), .B(exu_n16231), .Y(exu_n27215));
INVX1 exu_U24823(.A(exu_n27215), .Y(exu_n7940));
AND2X1 exu_U24824(.A(shft_rshift16_b1[45]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27217));
INVX1 exu_U24825(.A(exu_n27217), .Y(exu_n7941));
AND2X1 exu_U24826(.A(shft_rshift16_b1[36]), .B(exu_n15400), .Y(exu_n27221));
INVX1 exu_U24827(.A(exu_n27221), .Y(exu_n7942));
AND2X1 exu_U24828(.A(shft_rshift16_b1[44]), .B(exu_n16234), .Y(exu_n27223));
INVX1 exu_U24829(.A(exu_n27223), .Y(exu_n7943));
AND2X1 exu_U24830(.A(shft_rshift16_b1[35]), .B(exu_n16231), .Y(exu_n27227));
INVX1 exu_U24831(.A(exu_n27227), .Y(exu_n7944));
AND2X1 exu_U24832(.A(shft_rshift16_b1[43]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27229));
INVX1 exu_U24833(.A(exu_n27229), .Y(exu_n7945));
AND2X1 exu_U24834(.A(shft_rshift16_b1[34]), .B(exu_n15400), .Y(exu_n27233));
INVX1 exu_U24835(.A(exu_n27233), .Y(exu_n7946));
AND2X1 exu_U24836(.A(shft_rshift16_b1[42]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27235));
INVX1 exu_U24837(.A(exu_n27235), .Y(exu_n7947));
AND2X1 exu_U24838(.A(shft_rshift16_b1[6]), .B(exu_n16231), .Y(exu_n27239));
INVX1 exu_U24839(.A(exu_n27239), .Y(exu_n7948));
AND2X1 exu_U24840(.A(shft_rshift16_b1[14]), .B(exu_n16234), .Y(exu_n27241));
INVX1 exu_U24841(.A(exu_n27241), .Y(exu_n7949));
AND2X1 exu_U24842(.A(shft_rshift16_b1[33]), .B(exu_n15400), .Y(exu_n27245));
INVX1 exu_U24843(.A(exu_n27245), .Y(exu_n7950));
AND2X1 exu_U24844(.A(shft_rshift16_b1[41]), .B(exu_n16234), .Y(exu_n27247));
INVX1 exu_U24845(.A(exu_n27247), .Y(exu_n7951));
AND2X1 exu_U24846(.A(shft_rshift16_b1[32]), .B(exu_n15400), .Y(exu_n27251));
INVX1 exu_U24847(.A(exu_n27251), .Y(exu_n7952));
AND2X1 exu_U24848(.A(shft_rshift16_b1[40]), .B(exu_n16234), .Y(exu_n27253));
INVX1 exu_U24849(.A(exu_n27253), .Y(exu_n7953));
AND2X1 exu_U24850(.A(shft_rshift16_b1[31]), .B(exu_n15400), .Y(exu_n27257));
INVX1 exu_U24851(.A(exu_n27257), .Y(exu_n7954));
AND2X1 exu_U24852(.A(shft_rshift16_b1[39]), .B(exu_n16234), .Y(exu_n27259));
INVX1 exu_U24853(.A(exu_n27259), .Y(exu_n7955));
AND2X1 exu_U24854(.A(shft_rshift16_b1[30]), .B(exu_n15400), .Y(exu_n27263));
INVX1 exu_U24855(.A(exu_n27263), .Y(exu_n7956));
AND2X1 exu_U24856(.A(shft_rshift16_b1[38]), .B(exu_n16234), .Y(exu_n27265));
INVX1 exu_U24857(.A(exu_n27265), .Y(exu_n7957));
AND2X1 exu_U24858(.A(shft_rshift16_b1[29]), .B(exu_n15400), .Y(exu_n27269));
INVX1 exu_U24859(.A(exu_n27269), .Y(exu_n7958));
AND2X1 exu_U24860(.A(shft_rshift16_b1[37]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27271));
INVX1 exu_U24861(.A(exu_n27271), .Y(exu_n7959));
AND2X1 exu_U24862(.A(shft_rshift16_b1[28]), .B(exu_n15400), .Y(exu_n27275));
INVX1 exu_U24863(.A(exu_n27275), .Y(exu_n7960));
AND2X1 exu_U24864(.A(shft_rshift16_b1[36]), .B(exu_n16234), .Y(exu_n27277));
INVX1 exu_U24865(.A(exu_n27277), .Y(exu_n7961));
AND2X1 exu_U24866(.A(shft_rshift16_b1[27]), .B(exu_n16231), .Y(exu_n27281));
INVX1 exu_U24867(.A(exu_n27281), .Y(exu_n7962));
AND2X1 exu_U24868(.A(shft_rshift16_b1[35]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27283));
INVX1 exu_U24869(.A(exu_n27283), .Y(exu_n7963));
AND2X1 exu_U24870(.A(shft_rshift16_b1[26]), .B(exu_n16231), .Y(exu_n27287));
INVX1 exu_U24871(.A(exu_n27287), .Y(exu_n7964));
AND2X1 exu_U24872(.A(shft_rshift16_b1[34]), .B(exu_n16234), .Y(exu_n27289));
INVX1 exu_U24873(.A(exu_n27289), .Y(exu_n7965));
AND2X1 exu_U24874(.A(shft_rshift16_b1[25]), .B(exu_n16231), .Y(exu_n27293));
INVX1 exu_U24875(.A(exu_n27293), .Y(exu_n7966));
AND2X1 exu_U24876(.A(shft_rshift16_b1[33]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27295));
INVX1 exu_U24877(.A(exu_n27295), .Y(exu_n7967));
AND2X1 exu_U24878(.A(shft_rshift16_b1[24]), .B(exu_n15400), .Y(exu_n27299));
INVX1 exu_U24879(.A(exu_n27299), .Y(exu_n7968));
AND2X1 exu_U24880(.A(shft_rshift16_b1[32]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27301));
INVX1 exu_U24881(.A(exu_n27301), .Y(exu_n7969));
AND2X1 exu_U24882(.A(shft_rshift16_b1[5]), .B(exu_n16231), .Y(exu_n27305));
INVX1 exu_U24883(.A(exu_n27305), .Y(exu_n7970));
AND2X1 exu_U24884(.A(shft_rshift16_b1[13]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27307));
INVX1 exu_U24885(.A(exu_n27307), .Y(exu_n7971));
AND2X1 exu_U24886(.A(shft_rshift16_b1[23]), .B(exu_n16231), .Y(exu_n27311));
INVX1 exu_U24887(.A(exu_n27311), .Y(exu_n7972));
AND2X1 exu_U24888(.A(shft_rshift16_b1[31]), .B(exu_n16234), .Y(exu_n27313));
INVX1 exu_U24889(.A(exu_n27313), .Y(exu_n7973));
AND2X1 exu_U24890(.A(shft_rshift16_b1[22]), .B(exu_n15400), .Y(exu_n27317));
INVX1 exu_U24891(.A(exu_n27317), .Y(exu_n7974));
AND2X1 exu_U24892(.A(shft_rshift16_b1[30]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27319));
INVX1 exu_U24893(.A(exu_n27319), .Y(exu_n7975));
AND2X1 exu_U24894(.A(shft_rshift16_b1[21]), .B(exu_n15400), .Y(exu_n27323));
INVX1 exu_U24895(.A(exu_n27323), .Y(exu_n7976));
AND2X1 exu_U24896(.A(shft_rshift16_b1[29]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27325));
INVX1 exu_U24897(.A(exu_n27325), .Y(exu_n7977));
AND2X1 exu_U24898(.A(shft_rshift16_b1[20]), .B(exu_n15400), .Y(exu_n27329));
INVX1 exu_U24899(.A(exu_n27329), .Y(exu_n7978));
AND2X1 exu_U24900(.A(shft_rshift16_b1[28]), .B(exu_n16234), .Y(exu_n27331));
INVX1 exu_U24901(.A(exu_n27331), .Y(exu_n7979));
AND2X1 exu_U24902(.A(shft_rshift16_b1[19]), .B(exu_n15400), .Y(exu_n27335));
INVX1 exu_U24903(.A(exu_n27335), .Y(exu_n7980));
AND2X1 exu_U24904(.A(shft_rshift16_b1[27]), .B(exu_n16234), .Y(exu_n27337));
INVX1 exu_U24905(.A(exu_n27337), .Y(exu_n7981));
AND2X1 exu_U24906(.A(shft_rshift16_b1[18]), .B(exu_n15400), .Y(exu_n27341));
INVX1 exu_U24907(.A(exu_n27341), .Y(exu_n7982));
AND2X1 exu_U24908(.A(shft_rshift16_b1[26]), .B(exu_n16234), .Y(exu_n27343));
INVX1 exu_U24909(.A(exu_n27343), .Y(exu_n7983));
AND2X1 exu_U24910(.A(shft_rshift16_b1[17]), .B(exu_n15400), .Y(exu_n27347));
INVX1 exu_U24911(.A(exu_n27347), .Y(exu_n7984));
AND2X1 exu_U24912(.A(shft_rshift16_b1[25]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27349));
INVX1 exu_U24913(.A(exu_n27349), .Y(exu_n7985));
AND2X1 exu_U24914(.A(shft_rshift16_b1[16]), .B(exu_n16231), .Y(exu_n27353));
INVX1 exu_U24915(.A(exu_n27353), .Y(exu_n7986));
AND2X1 exu_U24916(.A(shft_rshift16_b1[24]), .B(exu_n16234), .Y(exu_n27355));
INVX1 exu_U24917(.A(exu_n27355), .Y(exu_n7987));
AND2X1 exu_U24918(.A(shft_rshift16_b1[15]), .B(exu_n15400), .Y(exu_n27359));
INVX1 exu_U24919(.A(exu_n27359), .Y(exu_n7988));
AND2X1 exu_U24920(.A(shft_rshift16_b1[23]), .B(exu_n16234), .Y(exu_n27361));
INVX1 exu_U24921(.A(exu_n27361), .Y(exu_n7989));
AND2X1 exu_U24922(.A(shft_rshift16_b1[14]), .B(exu_n16231), .Y(exu_n27365));
INVX1 exu_U24923(.A(exu_n27365), .Y(exu_n7990));
AND2X1 exu_U24924(.A(shft_rshift16_b1[22]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27367));
INVX1 exu_U24925(.A(exu_n27367), .Y(exu_n7991));
AND2X1 exu_U24926(.A(shft_rshift16_b1[4]), .B(exu_n16231), .Y(exu_n27371));
INVX1 exu_U24927(.A(exu_n27371), .Y(exu_n7992));
AND2X1 exu_U24928(.A(shft_rshift16_b1[12]), .B(exu_n16234), .Y(exu_n27373));
INVX1 exu_U24929(.A(exu_n27373), .Y(exu_n7993));
AND2X1 exu_U24930(.A(exu_n16226), .B(shft_rshift4_b1[10]), .Y(exu_n27377));
INVX1 exu_U24931(.A(exu_n27377), .Y(exu_n7994));
AND2X1 exu_U24932(.A(exu_n16228), .B(shft_rshift4_b1[12]), .Y(exu_n27379));
INVX1 exu_U24933(.A(exu_n27379), .Y(exu_n7995));
AND2X1 exu_U24934(.A(shft_rshift4_b1[9]), .B(exu_n16225), .Y(exu_n27383));
INVX1 exu_U24935(.A(exu_n27383), .Y(exu_n7996));
AND2X1 exu_U24936(.A(shft_rshift4_b1[11]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27385));
INVX1 exu_U24937(.A(exu_n27385), .Y(exu_n7997));
AND2X1 exu_U24938(.A(shft_rshift4_b1[8]), .B(exu_n16225), .Y(exu_n27389));
INVX1 exu_U24939(.A(exu_n27389), .Y(exu_n7998));
AND2X1 exu_U24940(.A(shft_rshift4_b1[10]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27391));
INVX1 exu_U24941(.A(exu_n27391), .Y(exu_n7999));
AND2X1 exu_U24942(.A(shft_rshift4_b1[7]), .B(exu_n16225), .Y(exu_n27395));
INVX1 exu_U24943(.A(exu_n27395), .Y(exu_n8000));
AND2X1 exu_U24944(.A(shft_rshift4_b1[9]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27397));
INVX1 exu_U24945(.A(exu_n27397), .Y(exu_n8001));
AND2X1 exu_U24946(.A(exu_n16191), .B(exu_n16225), .Y(exu_n27401));
INVX1 exu_U24947(.A(exu_n27401), .Y(exu_n8002));
AND2X1 exu_U24948(.A(shft_rshift4_b1[63]), .B(exu_n16225), .Y(exu_n27404));
INVX1 exu_U24949(.A(exu_n27404), .Y(exu_n8003));
AND2X1 exu_U24950(.A(exu_n16191), .B(ecl_shft_shift1_e[3]), .Y(exu_n27406));
INVX1 exu_U24951(.A(exu_n27406), .Y(exu_n8004));
AND2X1 exu_U24952(.A(shft_rshift4_b1[62]), .B(exu_n16225), .Y(exu_n27410));
INVX1 exu_U24953(.A(exu_n27410), .Y(exu_n8005));
AND2X1 exu_U24954(.A(shft_rshift4_b1[61]), .B(exu_n16225), .Y(exu_n27415));
INVX1 exu_U24955(.A(exu_n27415), .Y(exu_n8006));
AND2X1 exu_U24956(.A(shft_rshift4_b1[63]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27417));
INVX1 exu_U24957(.A(exu_n27417), .Y(exu_n8007));
AND2X1 exu_U24958(.A(shft_rshift4_b1[6]), .B(exu_n16225), .Y(exu_n27421));
INVX1 exu_U24959(.A(exu_n27421), .Y(exu_n8008));
AND2X1 exu_U24960(.A(shft_rshift4_b1[8]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27423));
INVX1 exu_U24961(.A(exu_n27423), .Y(exu_n8009));
AND2X1 exu_U24962(.A(shft_rshift4_b1[60]), .B(exu_n16225), .Y(exu_n27427));
INVX1 exu_U24963(.A(exu_n27427), .Y(exu_n8010));
AND2X1 exu_U24964(.A(shft_rshift4_b1[62]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27429));
INVX1 exu_U24965(.A(exu_n27429), .Y(exu_n8011));
AND2X1 exu_U24966(.A(shft_rshift4_b1[59]), .B(exu_n16225), .Y(exu_n27433));
INVX1 exu_U24967(.A(exu_n27433), .Y(exu_n8012));
AND2X1 exu_U24968(.A(shft_rshift4_b1[61]), .B(exu_n16228), .Y(exu_n27435));
INVX1 exu_U24969(.A(exu_n27435), .Y(exu_n8013));
AND2X1 exu_U24970(.A(shft_rshift4_b1[58]), .B(exu_n16225), .Y(exu_n27439));
INVX1 exu_U24971(.A(exu_n27439), .Y(exu_n8014));
AND2X1 exu_U24972(.A(shft_rshift4_b1[60]), .B(exu_n16228), .Y(exu_n27441));
INVX1 exu_U24973(.A(exu_n27441), .Y(exu_n8015));
AND2X1 exu_U24974(.A(shft_rshift4_b1[57]), .B(exu_n16225), .Y(exu_n27445));
INVX1 exu_U24975(.A(exu_n27445), .Y(exu_n8016));
AND2X1 exu_U24976(.A(shft_rshift4_b1[59]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27447));
INVX1 exu_U24977(.A(exu_n27447), .Y(exu_n8017));
AND2X1 exu_U24978(.A(shft_rshift4_b1[56]), .B(exu_n16225), .Y(exu_n27451));
INVX1 exu_U24979(.A(exu_n27451), .Y(exu_n8018));
AND2X1 exu_U24980(.A(shft_rshift4_b1[58]), .B(exu_n16228), .Y(exu_n27453));
INVX1 exu_U24981(.A(exu_n27453), .Y(exu_n8019));
AND2X1 exu_U24982(.A(shft_rshift4_b1[55]), .B(exu_n16225), .Y(exu_n27457));
INVX1 exu_U24983(.A(exu_n27457), .Y(exu_n8020));
AND2X1 exu_U24984(.A(shft_rshift4_b1[57]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27459));
INVX1 exu_U24985(.A(exu_n27459), .Y(exu_n8021));
AND2X1 exu_U24986(.A(shft_rshift4_b1[54]), .B(exu_n16225), .Y(exu_n27463));
INVX1 exu_U24987(.A(exu_n27463), .Y(exu_n8022));
AND2X1 exu_U24988(.A(shft_rshift4_b1[56]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27465));
INVX1 exu_U24989(.A(exu_n27465), .Y(exu_n8023));
AND2X1 exu_U24990(.A(shft_rshift4_b1[53]), .B(exu_n16226), .Y(exu_n27469));
INVX1 exu_U24991(.A(exu_n27469), .Y(exu_n8024));
AND2X1 exu_U24992(.A(shft_rshift4_b1[55]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27471));
INVX1 exu_U24993(.A(exu_n27471), .Y(exu_n8025));
AND2X1 exu_U24994(.A(shft_rshift4_b1[52]), .B(exu_n16225), .Y(exu_n27475));
INVX1 exu_U24995(.A(exu_n27475), .Y(exu_n8026));
AND2X1 exu_U24996(.A(shft_rshift4_b1[54]), .B(exu_n16228), .Y(exu_n27477));
INVX1 exu_U24997(.A(exu_n27477), .Y(exu_n8027));
AND2X1 exu_U24998(.A(shft_rshift4_b1[51]), .B(exu_n16226), .Y(exu_n27481));
INVX1 exu_U24999(.A(exu_n27481), .Y(exu_n8028));
AND2X1 exu_U25000(.A(shft_rshift4_b1[53]), .B(exu_n16228), .Y(exu_n27483));
INVX1 exu_U25001(.A(exu_n27483), .Y(exu_n8029));
AND2X1 exu_U25002(.A(shft_rshift4_b1[5]), .B(exu_n16226), .Y(exu_n27487));
INVX1 exu_U25003(.A(exu_n27487), .Y(exu_n8030));
AND2X1 exu_U25004(.A(shft_rshift4_b1[7]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27489));
INVX1 exu_U25005(.A(exu_n27489), .Y(exu_n8031));
AND2X1 exu_U25006(.A(shft_rshift4_b1[50]), .B(exu_n16226), .Y(exu_n27493));
INVX1 exu_U25007(.A(exu_n27493), .Y(exu_n8032));
AND2X1 exu_U25008(.A(shft_rshift4_b1[52]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27495));
INVX1 exu_U25009(.A(exu_n27495), .Y(exu_n8033));
AND2X1 exu_U25010(.A(shft_rshift4_b1[49]), .B(exu_n16225), .Y(exu_n27499));
INVX1 exu_U25011(.A(exu_n27499), .Y(exu_n8034));
AND2X1 exu_U25012(.A(shft_rshift4_b1[51]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27501));
INVX1 exu_U25013(.A(exu_n27501), .Y(exu_n8035));
AND2X1 exu_U25014(.A(shft_rshift4_b1[48]), .B(exu_n16225), .Y(exu_n27505));
INVX1 exu_U25015(.A(exu_n27505), .Y(exu_n8036));
AND2X1 exu_U25016(.A(shft_rshift4_b1[50]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27507));
INVX1 exu_U25017(.A(exu_n27507), .Y(exu_n8037));
AND2X1 exu_U25018(.A(shft_rshift4_b1[47]), .B(exu_n16226), .Y(exu_n27511));
INVX1 exu_U25019(.A(exu_n27511), .Y(exu_n8038));
AND2X1 exu_U25020(.A(shft_rshift4_b1[49]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27513));
INVX1 exu_U25021(.A(exu_n27513), .Y(exu_n8039));
AND2X1 exu_U25022(.A(shft_rshift4_b1[46]), .B(exu_n16226), .Y(exu_n27517));
INVX1 exu_U25023(.A(exu_n27517), .Y(exu_n8040));
AND2X1 exu_U25024(.A(shft_rshift4_b1[48]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27519));
INVX1 exu_U25025(.A(exu_n27519), .Y(exu_n8041));
AND2X1 exu_U25026(.A(shft_rshift4_b1[45]), .B(exu_n16226), .Y(exu_n27523));
INVX1 exu_U25027(.A(exu_n27523), .Y(exu_n8042));
AND2X1 exu_U25028(.A(shft_rshift4_b1[47]), .B(exu_n16228), .Y(exu_n27525));
INVX1 exu_U25029(.A(exu_n27525), .Y(exu_n8043));
AND2X1 exu_U25030(.A(shft_rshift4_b1[44]), .B(exu_n16226), .Y(exu_n27529));
INVX1 exu_U25031(.A(exu_n27529), .Y(exu_n8044));
AND2X1 exu_U25032(.A(shft_rshift4_b1[46]), .B(exu_n16228), .Y(exu_n27531));
INVX1 exu_U25033(.A(exu_n27531), .Y(exu_n8045));
AND2X1 exu_U25034(.A(shft_rshift4_b1[43]), .B(exu_n16225), .Y(exu_n27535));
INVX1 exu_U25035(.A(exu_n27535), .Y(exu_n8046));
AND2X1 exu_U25036(.A(shft_rshift4_b1[45]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27537));
INVX1 exu_U25037(.A(exu_n27537), .Y(exu_n8047));
AND2X1 exu_U25038(.A(shft_rshift4_b1[42]), .B(exu_n16226), .Y(exu_n27541));
INVX1 exu_U25039(.A(exu_n27541), .Y(exu_n8048));
AND2X1 exu_U25040(.A(shft_rshift4_b1[44]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27543));
INVX1 exu_U25041(.A(exu_n27543), .Y(exu_n8049));
AND2X1 exu_U25042(.A(shft_rshift4_b1[41]), .B(exu_n16226), .Y(exu_n27547));
INVX1 exu_U25043(.A(exu_n27547), .Y(exu_n8050));
AND2X1 exu_U25044(.A(shft_rshift4_b1[43]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27549));
INVX1 exu_U25045(.A(exu_n27549), .Y(exu_n8051));
AND2X1 exu_U25046(.A(shft_rshift4_b1[4]), .B(exu_n16226), .Y(exu_n27553));
INVX1 exu_U25047(.A(exu_n27553), .Y(exu_n8052));
AND2X1 exu_U25048(.A(shft_rshift4_b1[6]), .B(exu_n16228), .Y(exu_n27555));
INVX1 exu_U25049(.A(exu_n27555), .Y(exu_n8053));
AND2X1 exu_U25050(.A(shft_rshift4_b1[40]), .B(exu_n16225), .Y(exu_n27559));
INVX1 exu_U25051(.A(exu_n27559), .Y(exu_n8054));
AND2X1 exu_U25052(.A(shft_rshift4_b1[42]), .B(exu_n16228), .Y(exu_n27561));
INVX1 exu_U25053(.A(exu_n27561), .Y(exu_n8055));
AND2X1 exu_U25054(.A(shft_rshift4_b1[39]), .B(exu_n16226), .Y(exu_n27565));
INVX1 exu_U25055(.A(exu_n27565), .Y(exu_n8056));
AND2X1 exu_U25056(.A(shft_rshift4_b1[41]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27567));
INVX1 exu_U25057(.A(exu_n27567), .Y(exu_n8057));
AND2X1 exu_U25058(.A(shft_rshift4_b1[38]), .B(exu_n16226), .Y(exu_n27571));
INVX1 exu_U25059(.A(exu_n27571), .Y(exu_n8058));
AND2X1 exu_U25060(.A(shft_rshift4_b1[40]), .B(exu_n16228), .Y(exu_n27573));
INVX1 exu_U25061(.A(exu_n27573), .Y(exu_n8059));
AND2X1 exu_U25062(.A(shft_rshift4_b1[37]), .B(exu_n16225), .Y(exu_n27577));
INVX1 exu_U25063(.A(exu_n27577), .Y(exu_n8060));
AND2X1 exu_U25064(.A(shft_rshift4_b1[39]), .B(exu_n16228), .Y(exu_n27579));
INVX1 exu_U25065(.A(exu_n27579), .Y(exu_n8061));
AND2X1 exu_U25066(.A(shft_rshift4_b1[36]), .B(exu_n16225), .Y(exu_n27583));
INVX1 exu_U25067(.A(exu_n27583), .Y(exu_n8062));
AND2X1 exu_U25068(.A(shft_rshift4_b1[38]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27585));
INVX1 exu_U25069(.A(exu_n27585), .Y(exu_n8063));
AND2X1 exu_U25070(.A(shft_rshift4_b1[35]), .B(exu_n16225), .Y(exu_n27589));
INVX1 exu_U25071(.A(exu_n27589), .Y(exu_n8064));
AND2X1 exu_U25072(.A(shft_rshift4_b1[37]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27591));
INVX1 exu_U25073(.A(exu_n27591), .Y(exu_n8065));
AND2X1 exu_U25074(.A(shft_rshift4_b1[34]), .B(exu_n16226), .Y(exu_n27595));
INVX1 exu_U25075(.A(exu_n27595), .Y(exu_n8066));
AND2X1 exu_U25076(.A(shft_rshift4_b1[36]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27597));
INVX1 exu_U25077(.A(exu_n27597), .Y(exu_n8067));
AND2X1 exu_U25078(.A(shft_rshift4_b1[33]), .B(exu_n16226), .Y(exu_n27601));
INVX1 exu_U25079(.A(exu_n27601), .Y(exu_n8068));
AND2X1 exu_U25080(.A(shft_rshift4_b1[35]), .B(exu_n16228), .Y(exu_n27603));
INVX1 exu_U25081(.A(exu_n27603), .Y(exu_n8069));
AND2X1 exu_U25082(.A(shft_rshift4_b1[32]), .B(exu_n16225), .Y(exu_n27607));
INVX1 exu_U25083(.A(exu_n27607), .Y(exu_n8070));
AND2X1 exu_U25084(.A(shft_rshift4_b1[34]), .B(exu_n16228), .Y(exu_n27609));
INVX1 exu_U25085(.A(exu_n27609), .Y(exu_n8071));
AND2X1 exu_U25086(.A(shft_rshift4_b1[31]), .B(exu_n16226), .Y(exu_n27613));
INVX1 exu_U25087(.A(exu_n27613), .Y(exu_n8072));
AND2X1 exu_U25088(.A(shft_rshift4_b1[33]), .B(exu_n16228), .Y(exu_n27615));
INVX1 exu_U25089(.A(exu_n27615), .Y(exu_n8073));
AND2X1 exu_U25090(.A(shft_rshift4_b1[3]), .B(exu_n16225), .Y(exu_n27619));
INVX1 exu_U25091(.A(exu_n27619), .Y(exu_n8074));
AND2X1 exu_U25092(.A(shft_rshift4_b1[5]), .B(exu_n16228), .Y(exu_n27621));
INVX1 exu_U25093(.A(exu_n27621), .Y(exu_n8075));
AND2X1 exu_U25094(.A(shft_rshift4_b1[30]), .B(exu_n16226), .Y(exu_n27625));
INVX1 exu_U25095(.A(exu_n27625), .Y(exu_n8076));
AND2X1 exu_U25096(.A(shft_rshift4_b1[32]), .B(exu_n16228), .Y(exu_n27627));
INVX1 exu_U25097(.A(exu_n27627), .Y(exu_n8077));
AND2X1 exu_U25098(.A(shft_rshift4_b1[29]), .B(exu_n16225), .Y(exu_n27631));
INVX1 exu_U25099(.A(exu_n27631), .Y(exu_n8078));
AND2X1 exu_U25100(.A(shft_rshift4_b1[31]), .B(exu_n16228), .Y(exu_n27633));
INVX1 exu_U25101(.A(exu_n27633), .Y(exu_n8079));
AND2X1 exu_U25102(.A(shft_rshift4_b1[28]), .B(exu_n16226), .Y(exu_n27637));
INVX1 exu_U25103(.A(exu_n27637), .Y(exu_n8080));
AND2X1 exu_U25104(.A(shft_rshift4_b1[30]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27639));
INVX1 exu_U25105(.A(exu_n27639), .Y(exu_n8081));
AND2X1 exu_U25106(.A(shft_rshift4_b1[27]), .B(exu_n16225), .Y(exu_n27643));
INVX1 exu_U25107(.A(exu_n27643), .Y(exu_n8082));
AND2X1 exu_U25108(.A(shft_rshift4_b1[29]), .B(exu_n16228), .Y(exu_n27645));
INVX1 exu_U25109(.A(exu_n27645), .Y(exu_n8083));
AND2X1 exu_U25110(.A(shft_rshift4_b1[26]), .B(exu_n16226), .Y(exu_n27649));
INVX1 exu_U25111(.A(exu_n27649), .Y(exu_n8084));
AND2X1 exu_U25112(.A(shft_rshift4_b1[28]), .B(exu_n16228), .Y(exu_n27651));
INVX1 exu_U25113(.A(exu_n27651), .Y(exu_n8085));
AND2X1 exu_U25114(.A(shft_rshift4_b1[25]), .B(exu_n16225), .Y(exu_n27655));
INVX1 exu_U25115(.A(exu_n27655), .Y(exu_n8086));
AND2X1 exu_U25116(.A(shft_rshift4_b1[27]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27657));
INVX1 exu_U25117(.A(exu_n27657), .Y(exu_n8087));
AND2X1 exu_U25118(.A(shft_rshift4_b1[24]), .B(exu_n16225), .Y(exu_n27661));
INVX1 exu_U25119(.A(exu_n27661), .Y(exu_n8088));
AND2X1 exu_U25120(.A(shft_rshift4_b1[26]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27663));
INVX1 exu_U25121(.A(exu_n27663), .Y(exu_n8089));
AND2X1 exu_U25122(.A(shft_rshift4_b1[23]), .B(exu_n16225), .Y(exu_n27667));
INVX1 exu_U25123(.A(exu_n27667), .Y(exu_n8090));
AND2X1 exu_U25124(.A(shft_rshift4_b1[25]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27669));
INVX1 exu_U25125(.A(exu_n27669), .Y(exu_n8091));
AND2X1 exu_U25126(.A(shft_rshift4_b1[22]), .B(exu_n16225), .Y(exu_n27673));
INVX1 exu_U25127(.A(exu_n27673), .Y(exu_n8092));
AND2X1 exu_U25128(.A(shft_rshift4_b1[24]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27675));
INVX1 exu_U25129(.A(exu_n27675), .Y(exu_n8093));
AND2X1 exu_U25130(.A(shft_rshift4_b1[21]), .B(exu_n16225), .Y(exu_n27679));
INVX1 exu_U25131(.A(exu_n27679), .Y(exu_n8094));
AND2X1 exu_U25132(.A(shft_rshift4_b1[23]), .B(exu_n16228), .Y(exu_n27681));
INVX1 exu_U25133(.A(exu_n27681), .Y(exu_n8095));
AND2X1 exu_U25134(.A(shft_rshift4_b1[2]), .B(exu_n16226), .Y(exu_n27685));
INVX1 exu_U25135(.A(exu_n27685), .Y(exu_n8096));
AND2X1 exu_U25136(.A(shft_rshift4_b1[4]), .B(exu_n16228), .Y(exu_n27687));
INVX1 exu_U25137(.A(exu_n27687), .Y(exu_n8097));
AND2X1 exu_U25138(.A(shft_rshift4_b1[20]), .B(exu_n16226), .Y(exu_n27691));
INVX1 exu_U25139(.A(exu_n27691), .Y(exu_n8098));
AND2X1 exu_U25140(.A(shft_rshift4_b1[22]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27693));
INVX1 exu_U25141(.A(exu_n27693), .Y(exu_n8099));
AND2X1 exu_U25142(.A(shft_rshift4_b1[19]), .B(exu_n16225), .Y(exu_n27697));
INVX1 exu_U25143(.A(exu_n27697), .Y(exu_n8100));
AND2X1 exu_U25144(.A(shft_rshift4_b1[21]), .B(exu_n16228), .Y(exu_n27699));
INVX1 exu_U25145(.A(exu_n27699), .Y(exu_n8101));
AND2X1 exu_U25146(.A(shft_rshift4_b1[18]), .B(exu_n16225), .Y(exu_n27703));
INVX1 exu_U25147(.A(exu_n27703), .Y(exu_n8102));
AND2X1 exu_U25148(.A(shft_rshift4_b1[20]), .B(exu_n16228), .Y(exu_n27705));
INVX1 exu_U25149(.A(exu_n27705), .Y(exu_n8103));
AND2X1 exu_U25150(.A(shft_rshift4_b1[17]), .B(exu_n16226), .Y(exu_n27709));
INVX1 exu_U25151(.A(exu_n27709), .Y(exu_n8104));
AND2X1 exu_U25152(.A(shft_rshift4_b1[19]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27711));
INVX1 exu_U25153(.A(exu_n27711), .Y(exu_n8105));
AND2X1 exu_U25154(.A(shft_rshift4_b1[16]), .B(exu_n16226), .Y(exu_n27715));
INVX1 exu_U25155(.A(exu_n27715), .Y(exu_n8106));
AND2X1 exu_U25156(.A(shft_rshift4_b1[18]), .B(exu_n16228), .Y(exu_n27717));
INVX1 exu_U25157(.A(exu_n27717), .Y(exu_n8107));
AND2X1 exu_U25158(.A(shft_rshift4_b1[15]), .B(exu_n16226), .Y(exu_n27721));
INVX1 exu_U25159(.A(exu_n27721), .Y(exu_n8108));
AND2X1 exu_U25160(.A(shft_rshift4_b1[17]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27723));
INVX1 exu_U25161(.A(exu_n27723), .Y(exu_n8109));
AND2X1 exu_U25162(.A(shft_rshift4_b1[14]), .B(exu_n16226), .Y(exu_n27727));
INVX1 exu_U25163(.A(exu_n27727), .Y(exu_n8110));
AND2X1 exu_U25164(.A(shft_rshift4_b1[16]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27729));
INVX1 exu_U25165(.A(exu_n27729), .Y(exu_n8111));
AND2X1 exu_U25166(.A(shft_rshift4_b1[13]), .B(exu_n16225), .Y(exu_n27733));
INVX1 exu_U25167(.A(exu_n27733), .Y(exu_n8112));
AND2X1 exu_U25168(.A(shft_rshift4_b1[15]), .B(exu_n16228), .Y(exu_n27735));
INVX1 exu_U25169(.A(exu_n27735), .Y(exu_n8113));
AND2X1 exu_U25170(.A(shft_rshift4_b1[12]), .B(exu_n16226), .Y(exu_n27739));
INVX1 exu_U25171(.A(exu_n27739), .Y(exu_n8114));
AND2X1 exu_U25172(.A(shft_rshift4_b1[14]), .B(exu_n16228), .Y(exu_n27741));
INVX1 exu_U25173(.A(exu_n27741), .Y(exu_n8115));
AND2X1 exu_U25174(.A(shft_rshift4_b1[11]), .B(exu_n16226), .Y(exu_n27745));
INVX1 exu_U25175(.A(exu_n27745), .Y(exu_n8116));
AND2X1 exu_U25176(.A(shft_rshift4_b1[13]), .B(ecl_shft_shift1_e[3]), .Y(exu_n27747));
INVX1 exu_U25177(.A(exu_n27747), .Y(exu_n8117));
AND2X1 exu_U25178(.A(shft_rshift4_b1[1]), .B(exu_n16226), .Y(exu_n27751));
INVX1 exu_U25179(.A(exu_n27751), .Y(exu_n8118));
AND2X1 exu_U25180(.A(shft_rshift4_b1[3]), .B(exu_n16228), .Y(exu_n27753));
INVX1 exu_U25181(.A(exu_n27753), .Y(exu_n8119));
AND2X1 exu_U25182(.A(shft_shifter_input_b1[47]), .B(exu_n16146), .Y(exu_n27761));
INVX1 exu_U25183(.A(exu_n27761), .Y(exu_n8120));
AND2X1 exu_U25184(.A(shft_rshifterinput_b1[15]), .B(exu_n16142), .Y(exu_n27763));
INVX1 exu_U25185(.A(exu_n27763), .Y(exu_n8121));
AND2X1 exu_U25186(.A(shft_shifter_input_b1[46]), .B(shft_shift16_e[1]), .Y(exu_n27767));
INVX1 exu_U25187(.A(exu_n27767), .Y(exu_n8122));
AND2X1 exu_U25188(.A(shft_rshifterinput_b1[14]), .B(exu_n15399), .Y(exu_n27769));
INVX1 exu_U25189(.A(exu_n27769), .Y(exu_n8123));
AND2X1 exu_U25190(.A(shft_shifter_input_b1[45]), .B(exu_n16146), .Y(exu_n27773));
INVX1 exu_U25191(.A(exu_n27773), .Y(exu_n8124));
AND2X1 exu_U25192(.A(shft_rshifterinput_b1[13]), .B(exu_n15399), .Y(exu_n27775));
INVX1 exu_U25193(.A(exu_n27775), .Y(exu_n8125));
AND2X1 exu_U25194(.A(shft_shifter_input_b1[44]), .B(shft_shift16_e[1]), .Y(exu_n27779));
INVX1 exu_U25195(.A(exu_n27779), .Y(exu_n8126));
AND2X1 exu_U25196(.A(shft_rshifterinput_b1[12]), .B(exu_n15399), .Y(exu_n27781));
INVX1 exu_U25197(.A(exu_n27781), .Y(exu_n8127));
AND2X1 exu_U25198(.A(shft_shifter_input_b1[43]), .B(shft_shift16_e[1]), .Y(exu_n27786));
INVX1 exu_U25199(.A(exu_n27786), .Y(exu_n8128));
AND2X1 exu_U25200(.A(shft_rshifterinput_b1[11]), .B(exu_n16143), .Y(exu_n27788));
INVX1 exu_U25201(.A(exu_n27788), .Y(exu_n8129));
AND2X1 exu_U25202(.A(shft_shifter_input_b1[42]), .B(exu_n16146), .Y(exu_n27792));
INVX1 exu_U25203(.A(exu_n27792), .Y(exu_n8130));
AND2X1 exu_U25204(.A(shft_rshifterinput_b1[10]), .B(exu_n15399), .Y(exu_n27794));
INVX1 exu_U25205(.A(exu_n27794), .Y(exu_n8131));
AND2X1 exu_U25206(.A(shft_shifter_input_b1[41]), .B(exu_n16146), .Y(exu_n27798));
INVX1 exu_U25207(.A(exu_n27798), .Y(exu_n8132));
AND2X1 exu_U25208(.A(shft_rshifterinput_b1[9]), .B(exu_n15399), .Y(exu_n27800));
INVX1 exu_U25209(.A(exu_n27800), .Y(exu_n8133));
AND2X1 exu_U25210(.A(shft_shifter_input_b1[40]), .B(shft_shift16_e[1]), .Y(exu_n27804));
INVX1 exu_U25211(.A(exu_n27804), .Y(exu_n8134));
AND2X1 exu_U25212(.A(shft_rshifterinput_b1[8]), .B(exu_n16143), .Y(exu_n27806));
INVX1 exu_U25213(.A(exu_n27806), .Y(exu_n8135));
AND2X1 exu_U25214(.A(shft_shifter_input_b1[39]), .B(exu_n16146), .Y(exu_n27810));
INVX1 exu_U25215(.A(exu_n27810), .Y(exu_n8136));
AND2X1 exu_U25216(.A(shft_rshifterinput_b1[7]), .B(exu_n16144), .Y(exu_n27812));
INVX1 exu_U25217(.A(exu_n27812), .Y(exu_n8137));
AND2X1 exu_U25218(.A(shft_shifter_input_b1[38]), .B(shft_shift16_e[1]), .Y(exu_n27816));
INVX1 exu_U25219(.A(exu_n27816), .Y(exu_n8138));
AND2X1 exu_U25220(.A(shft_rshifterinput_b1[6]), .B(exu_n15399), .Y(exu_n27818));
INVX1 exu_U25221(.A(exu_n27818), .Y(exu_n8139));
AND2X1 exu_U25222(.A(shft_shifter_input_b1[37]), .B(exu_n16146), .Y(exu_n27822));
INVX1 exu_U25223(.A(exu_n27822), .Y(exu_n8140));
AND2X1 exu_U25224(.A(shft_rshifterinput_b1[5]), .B(exu_n15399), .Y(exu_n27824));
INVX1 exu_U25225(.A(exu_n27824), .Y(exu_n8141));
AND2X1 exu_U25226(.A(shft_shifter_input_b1[36]), .B(shft_shift16_e[1]), .Y(exu_n27828));
INVX1 exu_U25227(.A(exu_n27828), .Y(exu_n8142));
AND2X1 exu_U25228(.A(shft_rshifterinput_b1[4]), .B(exu_n16143), .Y(exu_n27830));
INVX1 exu_U25229(.A(exu_n27830), .Y(exu_n8143));
AND2X1 exu_U25230(.A(shft_shifter_input_b1[35]), .B(exu_n16146), .Y(exu_n27834));
INVX1 exu_U25231(.A(exu_n27834), .Y(exu_n8144));
AND2X1 exu_U25232(.A(shft_rshifterinput_b1[3]), .B(exu_n15399), .Y(exu_n27836));
INVX1 exu_U25233(.A(exu_n27836), .Y(exu_n8145));
AND2X1 exu_U25234(.A(shft_shifter_input_b1[34]), .B(exu_n16146), .Y(exu_n27840));
INVX1 exu_U25235(.A(exu_n27840), .Y(exu_n8146));
AND2X1 exu_U25236(.A(shft_rshifterinput_b1[2]), .B(exu_n16144), .Y(exu_n27842));
INVX1 exu_U25237(.A(exu_n27842), .Y(exu_n8147));
AND2X1 exu_U25238(.A(shft_shifter_input_b1[33]), .B(shft_shift16_e[1]), .Y(exu_n27847));
INVX1 exu_U25239(.A(exu_n27847), .Y(exu_n8148));
AND2X1 exu_U25240(.A(shft_rshifterinput_b1[1]), .B(exu_n16143), .Y(exu_n27849));
INVX1 exu_U25241(.A(exu_n27849), .Y(exu_n8149));
AND2X1 exu_U25242(.A(shft_shifter_input_b1[32]), .B(shft_shift16_e[1]), .Y(exu_n27853));
INVX1 exu_U25243(.A(exu_n27853), .Y(exu_n8150));
AND2X1 exu_U25244(.A(shft_rshifterinput_b1[0]), .B(exu_n15399), .Y(exu_n27855));
INVX1 exu_U25245(.A(exu_n27855), .Y(exu_n8151));
AND2X1 exu_U25246(.A(shft_rshifterinput_b1[31]), .B(exu_n16146), .Y(exu_n27858));
INVX1 exu_U25247(.A(exu_n27858), .Y(exu_n8152));
AND2X1 exu_U25248(.A(shft_rshifterinput_b1[30]), .B(shft_shift16_e[1]), .Y(exu_n27862));
INVX1 exu_U25249(.A(exu_n27862), .Y(exu_n8153));
AND2X1 exu_U25250(.A(shft_rshifterinput_b1[29]), .B(shft_shift16_e[1]), .Y(exu_n27866));
INVX1 exu_U25251(.A(exu_n27866), .Y(exu_n8154));
AND2X1 exu_U25252(.A(shft_rshifterinput_b1[28]), .B(shft_shift16_e[1]), .Y(exu_n27870));
INVX1 exu_U25253(.A(exu_n27870), .Y(exu_n8155));
AND2X1 exu_U25254(.A(shft_rshifterinput_b1[27]), .B(exu_n16146), .Y(exu_n27874));
INVX1 exu_U25255(.A(exu_n27874), .Y(exu_n8156));
AND2X1 exu_U25256(.A(shft_rshifterinput_b1[26]), .B(exu_n16146), .Y(exu_n27878));
INVX1 exu_U25257(.A(exu_n27878), .Y(exu_n8157));
AND2X1 exu_U25258(.A(shft_rshifterinput_b1[25]), .B(shft_shift16_e[1]), .Y(exu_n27882));
INVX1 exu_U25259(.A(exu_n27882), .Y(exu_n8158));
AND2X1 exu_U25260(.A(shft_rshifterinput_b1[24]), .B(shft_shift16_e[1]), .Y(exu_n27886));
INVX1 exu_U25261(.A(exu_n27886), .Y(exu_n8159));
AND2X1 exu_U25262(.A(shft_rshifterinput_b1[23]), .B(shft_shift16_e[1]), .Y(exu_n27891));
INVX1 exu_U25263(.A(exu_n27891), .Y(exu_n8160));
AND2X1 exu_U25264(.A(shft_rshifterinput_b1[22]), .B(exu_n16146), .Y(exu_n27895));
INVX1 exu_U25265(.A(exu_n27895), .Y(exu_n8161));
AND2X1 exu_U25266(.A(shft_rshifterinput_b1[21]), .B(shft_shift16_e[1]), .Y(exu_n27899));
INVX1 exu_U25267(.A(exu_n27899), .Y(exu_n8162));
AND2X1 exu_U25268(.A(shft_rshifterinput_b1[20]), .B(shft_shift16_e[1]), .Y(exu_n27903));
INVX1 exu_U25269(.A(exu_n27903), .Y(exu_n8163));
AND2X1 exu_U25270(.A(shft_rshifterinput_b1[19]), .B(exu_n16146), .Y(exu_n27907));
INVX1 exu_U25271(.A(exu_n27907), .Y(exu_n8164));
AND2X1 exu_U25272(.A(shft_rshifterinput_b1[18]), .B(shft_shift16_e[1]), .Y(exu_n27911));
INVX1 exu_U25273(.A(exu_n27911), .Y(exu_n8165));
AND2X1 exu_U25274(.A(shft_rshifterinput_b1[17]), .B(exu_n16146), .Y(exu_n27915));
INVX1 exu_U25275(.A(exu_n27915), .Y(exu_n8166));
AND2X1 exu_U25276(.A(shft_rshifterinput_b1[16]), .B(shft_shift16_e[1]), .Y(exu_n27919));
INVX1 exu_U25277(.A(exu_n27919), .Y(exu_n8167));
AND2X1 exu_U25278(.A(shft_rshifterinput_b1[15]), .B(shft_shift16_e[1]), .Y(exu_n27923));
INVX1 exu_U25279(.A(exu_n27923), .Y(exu_n8168));
AND2X1 exu_U25280(.A(shft_rshifterinput_b1[14]), .B(exu_n16146), .Y(exu_n27926));
INVX1 exu_U25281(.A(exu_n27926), .Y(exu_n8169));
AND2X1 exu_U25282(.A(shft_rshifterinput_b1[13]), .B(exu_n16146), .Y(exu_n27930));
INVX1 exu_U25283(.A(exu_n27930), .Y(exu_n8170));
AND2X1 exu_U25284(.A(shft_rshifterinput_b1[12]), .B(shft_shift16_e[1]), .Y(exu_n27933));
INVX1 exu_U25285(.A(exu_n27933), .Y(exu_n8171));
AND2X1 exu_U25286(.A(shft_rshifterinput_b1[11]), .B(shft_shift16_e[1]), .Y(exu_n27936));
INVX1 exu_U25287(.A(exu_n27936), .Y(exu_n8172));
AND2X1 exu_U25288(.A(shft_rshifterinput_b1[10]), .B(shft_shift16_e[1]), .Y(exu_n27939));
INVX1 exu_U25289(.A(exu_n27939), .Y(exu_n8173));
AND2X1 exu_U25290(.A(shft_rshifterinput_b1[9]), .B(shft_shift16_e[1]), .Y(exu_n27942));
INVX1 exu_U25291(.A(exu_n27942), .Y(exu_n8174));
AND2X1 exu_U25292(.A(shft_rshifterinput_b1[8]), .B(shft_shift16_e[1]), .Y(exu_n27945));
INVX1 exu_U25293(.A(exu_n27945), .Y(exu_n8175));
AND2X1 exu_U25294(.A(shft_rshifterinput_b1[7]), .B(exu_n16146), .Y(exu_n27948));
INVX1 exu_U25295(.A(exu_n27948), .Y(exu_n8176));
AND2X1 exu_U25296(.A(shft_rshifterinput_b1[6]), .B(shft_shift16_e[1]), .Y(exu_n27951));
INVX1 exu_U25297(.A(exu_n27951), .Y(exu_n8177));
AND2X1 exu_U25298(.A(shft_rshifterinput_b1[5]), .B(shft_shift16_e[1]), .Y(exu_n27954));
INVX1 exu_U25299(.A(exu_n27954), .Y(exu_n8178));
AND2X1 exu_U25300(.A(shft_rshifterinput_b1[4]), .B(shft_shift16_e[1]), .Y(exu_n27957));
INVX1 exu_U25301(.A(exu_n27957), .Y(exu_n8179));
AND2X1 exu_U25302(.A(shft_rshifterinput_b1[3]), .B(exu_n16146), .Y(exu_n27961));
INVX1 exu_U25303(.A(exu_n27961), .Y(exu_n8180));
AND2X1 exu_U25304(.A(shft_rshifterinput_b1[2]), .B(shft_shift16_e[1]), .Y(exu_n27964));
INVX1 exu_U25305(.A(exu_n27964), .Y(exu_n8181));
AND2X1 exu_U25306(.A(shft_rshifterinput_b1[1]), .B(exu_n16146), .Y(exu_n27967));
INVX1 exu_U25307(.A(exu_n27967), .Y(exu_n8182));
AND2X1 exu_U25308(.A(shft_rshifterinput_b1[0]), .B(exu_n16146), .Y(exu_n27970));
INVX1 exu_U25309(.A(exu_n27970), .Y(exu_n8183));
AND2X1 exu_U25310(.A(exu_n15400), .B(exu_n27782), .Y(exu_n27980));
INVX1 exu_U25311(.A(exu_n27980), .Y(exu_n8184));
AND2X1 exu_U25312(.A(exu_n27843), .B(exu_n16231), .Y(exu_n27984));
INVX1 exu_U25313(.A(exu_n27984), .Y(exu_n8185));
AND2X1 exu_U25314(.A(exu_n27888), .B(exu_n15400), .Y(exu_n27988));
INVX1 exu_U25315(.A(exu_n27988), .Y(exu_n8186));
AND2X1 exu_U25316(.A(exu_n27927), .B(exu_n15400), .Y(exu_n27991));
INVX1 exu_U25317(.A(exu_n27991), .Y(exu_n8187));
AND2X1 exu_U25318(.A(shft_lshift16_b1[59]), .B(exu_n16231), .Y(exu_n27995));
INVX1 exu_U25319(.A(exu_n27995), .Y(exu_n8188));
AND2X1 exu_U25320(.A(shft_lshift16_b1[51]), .B(ecl_shft_shift4_e[3]), .Y(exu_n27997));
INVX1 exu_U25321(.A(exu_n27997), .Y(exu_n8189));
AND2X1 exu_U25322(.A(shft_lshift16_b1[58]), .B(exu_n15400), .Y(exu_n28001));
INVX1 exu_U25323(.A(exu_n28001), .Y(exu_n8190));
AND2X1 exu_U25324(.A(shft_lshift16_b1[50]), .B(exu_n16234), .Y(exu_n28003));
INVX1 exu_U25325(.A(exu_n28003), .Y(exu_n8191));
AND2X1 exu_U25326(.A(shft_lshift16_b1[57]), .B(exu_n15400), .Y(exu_n28007));
INVX1 exu_U25327(.A(exu_n28007), .Y(exu_n8192));
AND2X1 exu_U25328(.A(shft_lshift16_b1[49]), .B(exu_n16234), .Y(exu_n28009));
INVX1 exu_U25329(.A(exu_n28009), .Y(exu_n8193));
AND2X1 exu_U25330(.A(shft_lshift16_b1[56]), .B(exu_n16231), .Y(exu_n28013));
INVX1 exu_U25331(.A(exu_n28013), .Y(exu_n8194));
AND2X1 exu_U25332(.A(shft_lshift16_b1[48]), .B(exu_n16234), .Y(exu_n28015));
INVX1 exu_U25333(.A(exu_n28015), .Y(exu_n8195));
AND2X1 exu_U25334(.A(exu_n27958), .B(exu_n16231), .Y(exu_n28018));
INVX1 exu_U25335(.A(exu_n28018), .Y(exu_n8196));
AND2X1 exu_U25336(.A(shft_lshift16_b1[55]), .B(exu_n15400), .Y(exu_n28022));
INVX1 exu_U25337(.A(exu_n28022), .Y(exu_n8197));
AND2X1 exu_U25338(.A(shft_lshift16_b1[47]), .B(exu_n16234), .Y(exu_n28024));
INVX1 exu_U25339(.A(exu_n28024), .Y(exu_n8198));
AND2X1 exu_U25340(.A(shft_lshift16_b1[54]), .B(exu_n16231), .Y(exu_n28028));
INVX1 exu_U25341(.A(exu_n28028), .Y(exu_n8199));
AND2X1 exu_U25342(.A(shft_lshift16_b1[46]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28030));
INVX1 exu_U25343(.A(exu_n28030), .Y(exu_n8200));
AND2X1 exu_U25344(.A(shft_lshift16_b1[53]), .B(exu_n15400), .Y(exu_n28034));
INVX1 exu_U25345(.A(exu_n28034), .Y(exu_n8201));
AND2X1 exu_U25346(.A(shft_lshift16_b1[45]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28036));
INVX1 exu_U25347(.A(exu_n28036), .Y(exu_n8202));
AND2X1 exu_U25348(.A(shft_lshift16_b1[52]), .B(exu_n16231), .Y(exu_n28040));
INVX1 exu_U25349(.A(exu_n28040), .Y(exu_n8203));
AND2X1 exu_U25350(.A(shft_lshift16_b1[44]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28042));
INVX1 exu_U25351(.A(exu_n28042), .Y(exu_n8204));
AND2X1 exu_U25352(.A(shft_lshift16_b1[51]), .B(exu_n16231), .Y(exu_n28046));
INVX1 exu_U25353(.A(exu_n28046), .Y(exu_n8205));
AND2X1 exu_U25354(.A(shft_lshift16_b1[43]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28048));
INVX1 exu_U25355(.A(exu_n28048), .Y(exu_n8206));
AND2X1 exu_U25356(.A(shft_lshift16_b1[50]), .B(exu_n15400), .Y(exu_n28052));
INVX1 exu_U25357(.A(exu_n28052), .Y(exu_n8207));
AND2X1 exu_U25358(.A(shft_lshift16_b1[42]), .B(exu_n16234), .Y(exu_n28054));
INVX1 exu_U25359(.A(exu_n28054), .Y(exu_n8208));
AND2X1 exu_U25360(.A(shft_lshift16_b1[49]), .B(exu_n15400), .Y(exu_n28058));
INVX1 exu_U25361(.A(exu_n28058), .Y(exu_n8209));
AND2X1 exu_U25362(.A(shft_lshift16_b1[41]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28060));
INVX1 exu_U25363(.A(exu_n28060), .Y(exu_n8210));
AND2X1 exu_U25364(.A(shft_lshift16_b1[48]), .B(exu_n16231), .Y(exu_n28064));
INVX1 exu_U25365(.A(exu_n28064), .Y(exu_n8211));
AND2X1 exu_U25366(.A(shft_lshift16_b1[40]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28066));
INVX1 exu_U25367(.A(exu_n28066), .Y(exu_n8212));
AND2X1 exu_U25368(.A(shft_lshift16_b1[47]), .B(exu_n15400), .Y(exu_n28070));
INVX1 exu_U25369(.A(exu_n28070), .Y(exu_n8213));
AND2X1 exu_U25370(.A(shft_lshift16_b1[39]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28072));
INVX1 exu_U25371(.A(exu_n28072), .Y(exu_n8214));
AND2X1 exu_U25372(.A(shft_lshift16_b1[46]), .B(exu_n16231), .Y(exu_n28076));
INVX1 exu_U25373(.A(exu_n28076), .Y(exu_n8215));
AND2X1 exu_U25374(.A(shft_lshift16_b1[38]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28078));
INVX1 exu_U25375(.A(exu_n28078), .Y(exu_n8216));
AND2X1 exu_U25376(.A(exu_n27977), .B(exu_n16231), .Y(exu_n28081));
INVX1 exu_U25377(.A(exu_n28081), .Y(exu_n8217));
AND2X1 exu_U25378(.A(shft_lshift16_b1[45]), .B(exu_n15400), .Y(exu_n28085));
INVX1 exu_U25379(.A(exu_n28085), .Y(exu_n8218));
AND2X1 exu_U25380(.A(shft_lshift16_b1[37]), .B(exu_n16234), .Y(exu_n28087));
INVX1 exu_U25381(.A(exu_n28087), .Y(exu_n8219));
AND2X1 exu_U25382(.A(shft_lshift16_b1[44]), .B(exu_n15400), .Y(exu_n28091));
INVX1 exu_U25383(.A(exu_n28091), .Y(exu_n8220));
AND2X1 exu_U25384(.A(shft_lshift16_b1[36]), .B(exu_n16234), .Y(exu_n28093));
INVX1 exu_U25385(.A(exu_n28093), .Y(exu_n8221));
AND2X1 exu_U25386(.A(shft_lshift16_b1[43]), .B(exu_n16231), .Y(exu_n28097));
INVX1 exu_U25387(.A(exu_n28097), .Y(exu_n8222));
AND2X1 exu_U25388(.A(shft_lshift16_b1[35]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28099));
INVX1 exu_U25389(.A(exu_n28099), .Y(exu_n8223));
AND2X1 exu_U25390(.A(shft_lshift16_b1[42]), .B(exu_n15400), .Y(exu_n28103));
INVX1 exu_U25391(.A(exu_n28103), .Y(exu_n8224));
AND2X1 exu_U25392(.A(shft_lshift16_b1[34]), .B(exu_n16234), .Y(exu_n28105));
INVX1 exu_U25393(.A(exu_n28105), .Y(exu_n8225));
AND2X1 exu_U25394(.A(shft_lshift16_b1[41]), .B(exu_n16231), .Y(exu_n28109));
INVX1 exu_U25395(.A(exu_n28109), .Y(exu_n8226));
AND2X1 exu_U25396(.A(shft_lshift16_b1[33]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28111));
INVX1 exu_U25397(.A(exu_n28111), .Y(exu_n8227));
AND2X1 exu_U25398(.A(shft_lshift16_b1[40]), .B(exu_n16231), .Y(exu_n28115));
INVX1 exu_U25399(.A(exu_n28115), .Y(exu_n8228));
AND2X1 exu_U25400(.A(shft_lshift16_b1[32]), .B(ecl_shft_shift4_e[3]), .Y(exu_n28117));
INVX1 exu_U25401(.A(exu_n28117), .Y(exu_n8229));
AND2X1 exu_U25402(.A(shft_lshift16_b1[39]), .B(exu_n15400), .Y(exu_n28121));
INVX1 exu_U25403(.A(exu_n28121), .Y(exu_n8230));
AND2X1 exu_U25404(.A(exu_n15703), .B(exu_n16234), .Y(exu_n28123));
INVX1 exu_U25405(.A(exu_n28123), .Y(exu_n8231));
AND2X1 exu_U25406(.A(shft_lshift16_b1[38]), .B(exu_n15400), .Y(exu_n28127));
INVX1 exu_U25407(.A(exu_n28127), .Y(exu_n8232));
AND2X1 exu_U25408(.A(exu_n15704), .B(exu_n16234), .Y(exu_n28129));
INVX1 exu_U25409(.A(exu_n28129), .Y(exu_n8233));
AND2X1 exu_U25410(.A(shft_lshift16_b1[37]), .B(exu_n15400), .Y(exu_n28133));
INVX1 exu_U25411(.A(exu_n28133), .Y(exu_n8234));
AND2X1 exu_U25412(.A(exu_n15705), .B(ecl_shft_shift4_e[3]), .Y(exu_n28135));
INVX1 exu_U25413(.A(exu_n28135), .Y(exu_n8235));
AND2X1 exu_U25414(.A(shft_lshift16_b1[36]), .B(exu_n16231), .Y(exu_n28139));
INVX1 exu_U25415(.A(exu_n28139), .Y(exu_n8236));
AND2X1 exu_U25416(.A(exu_n15706), .B(exu_n16234), .Y(exu_n28141));
INVX1 exu_U25417(.A(exu_n28141), .Y(exu_n8237));
AND2X1 exu_U25418(.A(shft_lshift16_b1[35]), .B(exu_n16231), .Y(exu_n28146));
INVX1 exu_U25419(.A(exu_n28146), .Y(exu_n8238));
AND2X1 exu_U25420(.A(exu_n15707), .B(ecl_shft_shift4_e[3]), .Y(exu_n28148));
INVX1 exu_U25421(.A(exu_n28148), .Y(exu_n8239));
AND2X1 exu_U25422(.A(shft_lshift16_b1[34]), .B(exu_n16231), .Y(exu_n28152));
INVX1 exu_U25423(.A(exu_n28152), .Y(exu_n8240));
AND2X1 exu_U25424(.A(exu_n15708), .B(ecl_shft_shift4_e[3]), .Y(exu_n28154));
INVX1 exu_U25425(.A(exu_n28154), .Y(exu_n8241));
AND2X1 exu_U25426(.A(shft_lshift16_b1[33]), .B(exu_n15400), .Y(exu_n28158));
INVX1 exu_U25427(.A(exu_n28158), .Y(exu_n8242));
AND2X1 exu_U25428(.A(exu_n15709), .B(exu_n16234), .Y(exu_n28160));
INVX1 exu_U25429(.A(exu_n28160), .Y(exu_n8243));
AND2X1 exu_U25430(.A(shft_lshift16_b1[32]), .B(exu_n16231), .Y(exu_n28164));
INVX1 exu_U25431(.A(exu_n28164), .Y(exu_n8244));
AND2X1 exu_U25432(.A(exu_n15710), .B(exu_n16234), .Y(exu_n28166));
INVX1 exu_U25433(.A(exu_n28166), .Y(exu_n8245));
AND2X1 exu_U25434(.A(exu_n15703), .B(exu_n16231), .Y(exu_n28170));
INVX1 exu_U25435(.A(exu_n28170), .Y(exu_n8246));
AND2X1 exu_U25436(.A(exu_n15711), .B(exu_n16234), .Y(exu_n28172));
INVX1 exu_U25437(.A(exu_n28172), .Y(exu_n8247));
AND2X1 exu_U25438(.A(exu_n15704), .B(exu_n15400), .Y(exu_n28176));
INVX1 exu_U25439(.A(exu_n28176), .Y(exu_n8248));
AND2X1 exu_U25440(.A(exu_n15712), .B(ecl_shft_shift4_e[3]), .Y(exu_n28178));
INVX1 exu_U25441(.A(exu_n28178), .Y(exu_n8249));
AND2X1 exu_U25442(.A(exu_n15705), .B(exu_n16231), .Y(exu_n28182));
INVX1 exu_U25443(.A(exu_n28182), .Y(exu_n8250));
AND2X1 exu_U25444(.A(exu_n15713), .B(ecl_shft_shift4_e[3]), .Y(exu_n28184));
INVX1 exu_U25445(.A(exu_n28184), .Y(exu_n8251));
AND2X1 exu_U25446(.A(exu_n15706), .B(exu_n16231), .Y(exu_n28188));
INVX1 exu_U25447(.A(exu_n28188), .Y(exu_n8252));
AND2X1 exu_U25448(.A(exu_n15714), .B(ecl_shft_shift4_e[3]), .Y(exu_n28190));
INVX1 exu_U25449(.A(exu_n28190), .Y(exu_n8253));
AND2X1 exu_U25450(.A(exu_n15707), .B(exu_n16231), .Y(exu_n28194));
INVX1 exu_U25451(.A(exu_n28194), .Y(exu_n8254));
AND2X1 exu_U25452(.A(exu_n15715), .B(exu_n16234), .Y(exu_n28196));
INVX1 exu_U25453(.A(exu_n28196), .Y(exu_n8255));
AND2X1 exu_U25454(.A(exu_n15708), .B(exu_n15400), .Y(exu_n28200));
INVX1 exu_U25455(.A(exu_n28200), .Y(exu_n8256));
AND2X1 exu_U25456(.A(exu_n15716), .B(exu_n16234), .Y(exu_n28202));
INVX1 exu_U25457(.A(exu_n28202), .Y(exu_n8257));
AND2X1 exu_U25458(.A(exu_n15709), .B(exu_n15400), .Y(exu_n28207));
INVX1 exu_U25459(.A(exu_n28207), .Y(exu_n8258));
AND2X1 exu_U25460(.A(exu_n15717), .B(ecl_shft_shift4_e[3]), .Y(exu_n28209));
INVX1 exu_U25461(.A(exu_n28209), .Y(exu_n8259));
AND2X1 exu_U25462(.A(exu_n15710), .B(exu_n16231), .Y(exu_n28213));
INVX1 exu_U25463(.A(exu_n28213), .Y(exu_n8260));
AND2X1 exu_U25464(.A(exu_n15718), .B(ecl_shft_shift4_e[3]), .Y(exu_n28215));
INVX1 exu_U25465(.A(exu_n28215), .Y(exu_n8261));
AND2X1 exu_U25466(.A(exu_n15711), .B(exu_n16231), .Y(exu_n28219));
INVX1 exu_U25467(.A(exu_n28219), .Y(exu_n8262));
AND2X1 exu_U25468(.A(exu_n27971), .B(exu_n16234), .Y(exu_n28221));
INVX1 exu_U25469(.A(exu_n28221), .Y(exu_n8263));
AND2X1 exu_U25470(.A(exu_n15712), .B(exu_n15400), .Y(exu_n28225));
INVX1 exu_U25471(.A(exu_n28225), .Y(exu_n8264));
AND2X1 exu_U25472(.A(exu_n27972), .B(exu_n16234), .Y(exu_n28227));
INVX1 exu_U25473(.A(exu_n28227), .Y(exu_n8265));
AND2X1 exu_U25474(.A(exu_n15713), .B(exu_n16231), .Y(exu_n28231));
INVX1 exu_U25475(.A(exu_n28231), .Y(exu_n8266));
AND2X1 exu_U25476(.A(exu_n27973), .B(ecl_shft_shift4_e[3]), .Y(exu_n28233));
INVX1 exu_U25477(.A(exu_n28233), .Y(exu_n8267));
AND2X1 exu_U25478(.A(exu_n15714), .B(exu_n16231), .Y(exu_n28237));
INVX1 exu_U25479(.A(exu_n28237), .Y(exu_n8268));
AND2X1 exu_U25480(.A(exu_n27974), .B(ecl_shft_shift4_e[3]), .Y(exu_n28239));
INVX1 exu_U25481(.A(exu_n28239), .Y(exu_n8269));
AND2X1 exu_U25482(.A(exu_n15715), .B(exu_n15400), .Y(exu_n28243));
INVX1 exu_U25483(.A(exu_n28243), .Y(exu_n8270));
AND2X1 exu_U25484(.A(exu_n27975), .B(exu_n16234), .Y(exu_n28245));
INVX1 exu_U25485(.A(exu_n28245), .Y(exu_n8271));
AND2X1 exu_U25486(.A(exu_n15716), .B(exu_n16231), .Y(exu_n28249));
INVX1 exu_U25487(.A(exu_n28249), .Y(exu_n8272));
AND2X1 exu_U25488(.A(exu_n27976), .B(exu_n16234), .Y(exu_n28251));
INVX1 exu_U25489(.A(exu_n28251), .Y(exu_n8273));
AND2X1 exu_U25490(.A(exu_n15717), .B(exu_n16231), .Y(exu_n28255));
INVX1 exu_U25491(.A(exu_n28255), .Y(exu_n8274));
AND2X1 exu_U25492(.A(exu_n27754), .B(ecl_shft_shift4_e[3]), .Y(exu_n28257));
INVX1 exu_U25493(.A(exu_n28257), .Y(exu_n8275));
AND2X1 exu_U25494(.A(exu_n15718), .B(exu_n16231), .Y(exu_n28261));
INVX1 exu_U25495(.A(exu_n28261), .Y(exu_n8276));
AND2X1 exu_U25496(.A(exu_n27755), .B(ecl_shft_shift4_e[3]), .Y(exu_n28263));
INVX1 exu_U25497(.A(exu_n28263), .Y(exu_n8277));
AND2X1 exu_U25498(.A(exu_n27971), .B(exu_n16231), .Y(exu_n28268));
INVX1 exu_U25499(.A(exu_n28268), .Y(exu_n8278));
AND2X1 exu_U25500(.A(exu_n27756), .B(ecl_shft_shift4_e[3]), .Y(exu_n28270));
INVX1 exu_U25501(.A(exu_n28270), .Y(exu_n8279));
AND2X1 exu_U25502(.A(exu_n27972), .B(exu_n16231), .Y(exu_n28274));
INVX1 exu_U25503(.A(exu_n28274), .Y(exu_n8280));
AND2X1 exu_U25504(.A(exu_n27757), .B(exu_n16234), .Y(exu_n28276));
INVX1 exu_U25505(.A(exu_n28276), .Y(exu_n8281));
AND2X1 exu_U25506(.A(exu_n27973), .B(exu_n16231), .Y(exu_n28280));
INVX1 exu_U25507(.A(exu_n28280), .Y(exu_n8282));
AND2X1 exu_U25508(.A(exu_n27782), .B(exu_n16234), .Y(exu_n28282));
INVX1 exu_U25509(.A(exu_n28282), .Y(exu_n8283));
AND2X1 exu_U25510(.A(exu_n27974), .B(exu_n15400), .Y(exu_n28286));
INVX1 exu_U25511(.A(exu_n28286), .Y(exu_n8284));
AND2X1 exu_U25512(.A(exu_n27843), .B(exu_n16234), .Y(exu_n28288));
INVX1 exu_U25513(.A(exu_n28288), .Y(exu_n8285));
AND2X1 exu_U25514(.A(exu_n27975), .B(exu_n16231), .Y(exu_n28292));
INVX1 exu_U25515(.A(exu_n28292), .Y(exu_n8286));
AND2X1 exu_U25516(.A(exu_n27888), .B(exu_n16234), .Y(exu_n28294));
INVX1 exu_U25517(.A(exu_n28294), .Y(exu_n8287));
AND2X1 exu_U25518(.A(exu_n27976), .B(exu_n15400), .Y(exu_n28298));
INVX1 exu_U25519(.A(exu_n28298), .Y(exu_n8288));
AND2X1 exu_U25520(.A(exu_n27927), .B(ecl_shft_shift4_e[3]), .Y(exu_n28300));
INVX1 exu_U25521(.A(exu_n28300), .Y(exu_n8289));
AND2X1 exu_U25522(.A(exu_n27754), .B(exu_n16231), .Y(exu_n28304));
INVX1 exu_U25523(.A(exu_n28304), .Y(exu_n8290));
AND2X1 exu_U25524(.A(exu_n27958), .B(ecl_shft_shift4_e[3]), .Y(exu_n28306));
INVX1 exu_U25525(.A(exu_n28306), .Y(exu_n8291));
AND2X1 exu_U25526(.A(exu_n27755), .B(exu_n16231), .Y(exu_n28310));
INVX1 exu_U25527(.A(exu_n28310), .Y(exu_n8292));
AND2X1 exu_U25528(.A(exu_n27977), .B(exu_n16234), .Y(exu_n28312));
INVX1 exu_U25529(.A(exu_n28312), .Y(exu_n8293));
AND2X1 exu_U25530(.A(exu_n27756), .B(exu_n15400), .Y(exu_n28315));
INVX1 exu_U25531(.A(exu_n28315), .Y(exu_n8294));
AND2X1 exu_U25532(.A(exu_n27757), .B(exu_n15400), .Y(exu_n28319));
INVX1 exu_U25533(.A(exu_n28319), .Y(exu_n8295));
AND2X1 exu_U25534(.A(exu_n16226), .B(shft_lshift4_b1[8]), .Y(exu_n28325));
INVX1 exu_U25535(.A(exu_n28325), .Y(exu_n8296));
AND2X1 exu_U25536(.A(ecl_shft_shift1_e[3]), .B(exu_n15695), .Y(exu_n28327));
INVX1 exu_U25537(.A(exu_n28327), .Y(exu_n8297));
AND2X1 exu_U25538(.A(exu_n15693), .B(exu_n16226), .Y(exu_n28331));
INVX1 exu_U25539(.A(exu_n28331), .Y(exu_n8298));
AND2X1 exu_U25540(.A(exu_n15719), .B(exu_n16228), .Y(exu_n28333));
INVX1 exu_U25541(.A(exu_n28333), .Y(exu_n8299));
AND2X1 exu_U25542(.A(exu_n15695), .B(exu_n16226), .Y(exu_n28337));
INVX1 exu_U25543(.A(exu_n28337), .Y(exu_n8300));
AND2X1 exu_U25544(.A(exu_n15720), .B(ecl_shft_shift1_e[3]), .Y(exu_n28339));
INVX1 exu_U25545(.A(exu_n28339), .Y(exu_n8301));
AND2X1 exu_U25546(.A(exu_n15719), .B(exu_n16226), .Y(exu_n28343));
INVX1 exu_U25547(.A(exu_n28343), .Y(exu_n8302));
AND2X1 exu_U25548(.A(exu_n28142), .B(ecl_shft_shift1_e[3]), .Y(exu_n28345));
INVX1 exu_U25549(.A(exu_n28345), .Y(exu_n8303));
AND2X1 exu_U25550(.A(shft_lshift4_b1[62]), .B(exu_n16226), .Y(exu_n28349));
INVX1 exu_U25551(.A(exu_n28349), .Y(exu_n8304));
AND2X1 exu_U25552(.A(shft_lshift4_b1[60]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28351));
INVX1 exu_U25553(.A(exu_n28351), .Y(exu_n8305));
AND2X1 exu_U25554(.A(shft_lshift4_b1[61]), .B(exu_n16226), .Y(exu_n28355));
INVX1 exu_U25555(.A(exu_n28355), .Y(exu_n8306));
AND2X1 exu_U25556(.A(shft_lshift4_b1[59]), .B(exu_n16228), .Y(exu_n28357));
INVX1 exu_U25557(.A(exu_n28357), .Y(exu_n8307));
AND2X1 exu_U25558(.A(shft_lshift4_b1[60]), .B(exu_n16226), .Y(exu_n28361));
INVX1 exu_U25559(.A(exu_n28361), .Y(exu_n8308));
AND2X1 exu_U25560(.A(shft_lshift4_b1[58]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28363));
INVX1 exu_U25561(.A(exu_n28363), .Y(exu_n8309));
AND2X1 exu_U25562(.A(shft_lshift4_b1[59]), .B(exu_n16226), .Y(exu_n28367));
INVX1 exu_U25563(.A(exu_n28367), .Y(exu_n8310));
AND2X1 exu_U25564(.A(shft_lshift4_b1[57]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28369));
INVX1 exu_U25565(.A(exu_n28369), .Y(exu_n8311));
AND2X1 exu_U25566(.A(exu_n15720), .B(exu_n16226), .Y(exu_n28373));
INVX1 exu_U25567(.A(exu_n28373), .Y(exu_n8312));
AND2X1 exu_U25568(.A(exu_n28203), .B(exu_n16228), .Y(exu_n28375));
INVX1 exu_U25569(.A(exu_n28375), .Y(exu_n8313));
AND2X1 exu_U25570(.A(shft_lshift4_b1[58]), .B(exu_n16226), .Y(exu_n28379));
INVX1 exu_U25571(.A(exu_n28379), .Y(exu_n8314));
AND2X1 exu_U25572(.A(shft_lshift4_b1[56]), .B(exu_n16228), .Y(exu_n28381));
INVX1 exu_U25573(.A(exu_n28381), .Y(exu_n8315));
AND2X1 exu_U25574(.A(shft_lshift4_b1[57]), .B(exu_n16225), .Y(exu_n28385));
INVX1 exu_U25575(.A(exu_n28385), .Y(exu_n8316));
AND2X1 exu_U25576(.A(shft_lshift4_b1[55]), .B(exu_n16228), .Y(exu_n28387));
INVX1 exu_U25577(.A(exu_n28387), .Y(exu_n8317));
AND2X1 exu_U25578(.A(shft_lshift4_b1[56]), .B(exu_n16225), .Y(exu_n28391));
INVX1 exu_U25579(.A(exu_n28391), .Y(exu_n8318));
AND2X1 exu_U25580(.A(shft_lshift4_b1[54]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28393));
INVX1 exu_U25581(.A(exu_n28393), .Y(exu_n8319));
AND2X1 exu_U25582(.A(shft_lshift4_b1[55]), .B(exu_n16225), .Y(exu_n28397));
INVX1 exu_U25583(.A(exu_n28397), .Y(exu_n8320));
AND2X1 exu_U25584(.A(shft_lshift4_b1[53]), .B(exu_n16228), .Y(exu_n28399));
INVX1 exu_U25585(.A(exu_n28399), .Y(exu_n8321));
AND2X1 exu_U25586(.A(shft_lshift4_b1[54]), .B(exu_n16226), .Y(exu_n28403));
INVX1 exu_U25587(.A(exu_n28403), .Y(exu_n8322));
AND2X1 exu_U25588(.A(shft_lshift4_b1[52]), .B(exu_n16228), .Y(exu_n28405));
INVX1 exu_U25589(.A(exu_n28405), .Y(exu_n8323));
AND2X1 exu_U25590(.A(shft_lshift4_b1[53]), .B(exu_n16225), .Y(exu_n28409));
INVX1 exu_U25591(.A(exu_n28409), .Y(exu_n8324));
AND2X1 exu_U25592(.A(shft_lshift4_b1[51]), .B(exu_n16228), .Y(exu_n28411));
INVX1 exu_U25593(.A(exu_n28411), .Y(exu_n8325));
AND2X1 exu_U25594(.A(shft_lshift4_b1[52]), .B(exu_n16225), .Y(exu_n28415));
INVX1 exu_U25595(.A(exu_n28415), .Y(exu_n8326));
AND2X1 exu_U25596(.A(shft_lshift4_b1[50]), .B(exu_n16228), .Y(exu_n28417));
INVX1 exu_U25597(.A(exu_n28417), .Y(exu_n8327));
AND2X1 exu_U25598(.A(shft_lshift4_b1[51]), .B(exu_n16226), .Y(exu_n28421));
INVX1 exu_U25599(.A(exu_n28421), .Y(exu_n8328));
AND2X1 exu_U25600(.A(shft_lshift4_b1[49]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28423));
INVX1 exu_U25601(.A(exu_n28423), .Y(exu_n8329));
AND2X1 exu_U25602(.A(shft_lshift4_b1[50]), .B(exu_n16225), .Y(exu_n28427));
INVX1 exu_U25603(.A(exu_n28427), .Y(exu_n8330));
AND2X1 exu_U25604(.A(shft_lshift4_b1[48]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28429));
INVX1 exu_U25605(.A(exu_n28429), .Y(exu_n8331));
AND2X1 exu_U25606(.A(shft_lshift4_b1[49]), .B(exu_n16226), .Y(exu_n28433));
INVX1 exu_U25607(.A(exu_n28433), .Y(exu_n8332));
AND2X1 exu_U25608(.A(shft_lshift4_b1[47]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28435));
INVX1 exu_U25609(.A(exu_n28435), .Y(exu_n8333));
AND2X1 exu_U25610(.A(exu_n28142), .B(exu_n16226), .Y(exu_n28439));
INVX1 exu_U25611(.A(exu_n28439), .Y(exu_n8334));
AND2X1 exu_U25612(.A(exu_n28264), .B(exu_n16228), .Y(exu_n28441));
INVX1 exu_U25613(.A(exu_n28441), .Y(exu_n8335));
AND2X1 exu_U25614(.A(shft_lshift4_b1[48]), .B(exu_n16225), .Y(exu_n28445));
INVX1 exu_U25615(.A(exu_n28445), .Y(exu_n8336));
AND2X1 exu_U25616(.A(shft_lshift4_b1[46]), .B(exu_n16228), .Y(exu_n28447));
INVX1 exu_U25617(.A(exu_n28447), .Y(exu_n8337));
AND2X1 exu_U25618(.A(shft_lshift4_b1[47]), .B(exu_n16225), .Y(exu_n28451));
INVX1 exu_U25619(.A(exu_n28451), .Y(exu_n8338));
AND2X1 exu_U25620(.A(shft_lshift4_b1[45]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28453));
INVX1 exu_U25621(.A(exu_n28453), .Y(exu_n8339));
AND2X1 exu_U25622(.A(shft_lshift4_b1[46]), .B(exu_n16226), .Y(exu_n28457));
INVX1 exu_U25623(.A(exu_n28457), .Y(exu_n8340));
AND2X1 exu_U25624(.A(shft_lshift4_b1[44]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28459));
INVX1 exu_U25625(.A(exu_n28459), .Y(exu_n8341));
AND2X1 exu_U25626(.A(shft_lshift4_b1[45]), .B(exu_n16226), .Y(exu_n28463));
INVX1 exu_U25627(.A(exu_n28463), .Y(exu_n8342));
AND2X1 exu_U25628(.A(shft_lshift4_b1[43]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28465));
INVX1 exu_U25629(.A(exu_n28465), .Y(exu_n8343));
AND2X1 exu_U25630(.A(shft_lshift4_b1[44]), .B(exu_n16225), .Y(exu_n28469));
INVX1 exu_U25631(.A(exu_n28469), .Y(exu_n8344));
AND2X1 exu_U25632(.A(shft_lshift4_b1[42]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28471));
INVX1 exu_U25633(.A(exu_n28471), .Y(exu_n8345));
AND2X1 exu_U25634(.A(shft_lshift4_b1[43]), .B(exu_n16225), .Y(exu_n28475));
INVX1 exu_U25635(.A(exu_n28475), .Y(exu_n8346));
AND2X1 exu_U25636(.A(shft_lshift4_b1[41]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28477));
INVX1 exu_U25637(.A(exu_n28477), .Y(exu_n8347));
AND2X1 exu_U25638(.A(shft_lshift4_b1[42]), .B(exu_n16225), .Y(exu_n28481));
INVX1 exu_U25639(.A(exu_n28481), .Y(exu_n8348));
AND2X1 exu_U25640(.A(shft_lshift4_b1[40]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28483));
INVX1 exu_U25641(.A(exu_n28483), .Y(exu_n8349));
AND2X1 exu_U25642(.A(shft_lshift4_b1[41]), .B(exu_n16226), .Y(exu_n28487));
INVX1 exu_U25643(.A(exu_n28487), .Y(exu_n8350));
AND2X1 exu_U25644(.A(shft_lshift4_b1[39]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28489));
INVX1 exu_U25645(.A(exu_n28489), .Y(exu_n8351));
AND2X1 exu_U25646(.A(shft_lshift4_b1[40]), .B(exu_n16225), .Y(exu_n28493));
INVX1 exu_U25647(.A(exu_n28493), .Y(exu_n8352));
AND2X1 exu_U25648(.A(shft_lshift4_b1[38]), .B(exu_n16228), .Y(exu_n28495));
INVX1 exu_U25649(.A(exu_n28495), .Y(exu_n8353));
AND2X1 exu_U25650(.A(shft_lshift4_b1[39]), .B(exu_n16225), .Y(exu_n28499));
INVX1 exu_U25651(.A(exu_n28499), .Y(exu_n8354));
AND2X1 exu_U25652(.A(shft_lshift4_b1[37]), .B(exu_n16228), .Y(exu_n28501));
INVX1 exu_U25653(.A(exu_n28501), .Y(exu_n8355));
AND2X1 exu_U25654(.A(exu_n28203), .B(exu_n16225), .Y(exu_n28505));
INVX1 exu_U25655(.A(exu_n28505), .Y(exu_n8356));
AND2X1 exu_U25656(.A(exu_n28321), .B(exu_n16228), .Y(exu_n28507));
INVX1 exu_U25657(.A(exu_n28507), .Y(exu_n8357));
AND2X1 exu_U25658(.A(shft_lshift4_b1[38]), .B(exu_n16226), .Y(exu_n28511));
INVX1 exu_U25659(.A(exu_n28511), .Y(exu_n8358));
AND2X1 exu_U25660(.A(shft_lshift4_b1[36]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28513));
INVX1 exu_U25661(.A(exu_n28513), .Y(exu_n8359));
AND2X1 exu_U25662(.A(shft_lshift4_b1[37]), .B(exu_n16225), .Y(exu_n28517));
INVX1 exu_U25663(.A(exu_n28517), .Y(exu_n8360));
AND2X1 exu_U25664(.A(shft_lshift4_b1[35]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28519));
INVX1 exu_U25665(.A(exu_n28519), .Y(exu_n8361));
AND2X1 exu_U25666(.A(shft_lshift4_b1[36]), .B(exu_n16225), .Y(exu_n28523));
INVX1 exu_U25667(.A(exu_n28523), .Y(exu_n8362));
AND2X1 exu_U25668(.A(shft_lshift4_b1[34]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28525));
INVX1 exu_U25669(.A(exu_n28525), .Y(exu_n8363));
AND2X1 exu_U25670(.A(shft_lshift4_b1[35]), .B(exu_n16225), .Y(exu_n28529));
INVX1 exu_U25671(.A(exu_n28529), .Y(exu_n8364));
AND2X1 exu_U25672(.A(shft_lshift4_b1[33]), .B(exu_n16228), .Y(exu_n28531));
INVX1 exu_U25673(.A(exu_n28531), .Y(exu_n8365));
AND2X1 exu_U25674(.A(shft_lshift4_b1[34]), .B(exu_n16226), .Y(exu_n28535));
INVX1 exu_U25675(.A(exu_n28535), .Y(exu_n8366));
AND2X1 exu_U25676(.A(shft_lshift4_b1[32]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28537));
INVX1 exu_U25677(.A(exu_n28537), .Y(exu_n8367));
AND2X1 exu_U25678(.A(shft_lshift4_b1[33]), .B(exu_n16225), .Y(exu_n28541));
INVX1 exu_U25679(.A(exu_n28541), .Y(exu_n8368));
AND2X1 exu_U25680(.A(shft_lshift4_b1[31]), .B(exu_n16228), .Y(exu_n28543));
INVX1 exu_U25681(.A(exu_n28543), .Y(exu_n8369));
AND2X1 exu_U25682(.A(shft_lshift4_b1[32]), .B(exu_n16226), .Y(exu_n28547));
INVX1 exu_U25683(.A(exu_n28547), .Y(exu_n8370));
AND2X1 exu_U25684(.A(shft_lshift4_b1[30]), .B(exu_n16228), .Y(exu_n28549));
INVX1 exu_U25685(.A(exu_n28549), .Y(exu_n8371));
AND2X1 exu_U25686(.A(shft_lshift4_b1[31]), .B(exu_n16226), .Y(exu_n28553));
INVX1 exu_U25687(.A(exu_n28553), .Y(exu_n8372));
AND2X1 exu_U25688(.A(shft_lshift4_b1[29]), .B(exu_n16228), .Y(exu_n28555));
INVX1 exu_U25689(.A(exu_n28555), .Y(exu_n8373));
AND2X1 exu_U25690(.A(shft_lshift4_b1[30]), .B(exu_n16225), .Y(exu_n28559));
INVX1 exu_U25691(.A(exu_n28559), .Y(exu_n8374));
AND2X1 exu_U25692(.A(shft_lshift4_b1[28]), .B(exu_n16228), .Y(exu_n28561));
INVX1 exu_U25693(.A(exu_n28561), .Y(exu_n8375));
AND2X1 exu_U25694(.A(shft_lshift4_b1[29]), .B(exu_n16226), .Y(exu_n28565));
INVX1 exu_U25695(.A(exu_n28565), .Y(exu_n8376));
AND2X1 exu_U25696(.A(shft_lshift4_b1[27]), .B(exu_n16228), .Y(exu_n28567));
INVX1 exu_U25697(.A(exu_n28567), .Y(exu_n8377));
AND2X1 exu_U25698(.A(exu_n28264), .B(exu_n16225), .Y(exu_n28570));
INVX1 exu_U25699(.A(exu_n28570), .Y(exu_n8378));
AND2X1 exu_U25700(.A(shft_lshift4_b1[28]), .B(exu_n16226), .Y(exu_n28575));
INVX1 exu_U25701(.A(exu_n28575), .Y(exu_n8379));
AND2X1 exu_U25702(.A(shft_lshift4_b1[26]), .B(exu_n16228), .Y(exu_n28577));
INVX1 exu_U25703(.A(exu_n28577), .Y(exu_n8380));
AND2X1 exu_U25704(.A(shft_lshift4_b1[27]), .B(exu_n16226), .Y(exu_n28581));
INVX1 exu_U25705(.A(exu_n28581), .Y(exu_n8381));
AND2X1 exu_U25706(.A(shft_lshift4_b1[25]), .B(exu_n16228), .Y(exu_n28583));
INVX1 exu_U25707(.A(exu_n28583), .Y(exu_n8382));
AND2X1 exu_U25708(.A(shft_lshift4_b1[26]), .B(exu_n16226), .Y(exu_n28587));
INVX1 exu_U25709(.A(exu_n28587), .Y(exu_n8383));
AND2X1 exu_U25710(.A(shft_lshift4_b1[24]), .B(exu_n16228), .Y(exu_n28589));
INVX1 exu_U25711(.A(exu_n28589), .Y(exu_n8384));
AND2X1 exu_U25712(.A(shft_lshift4_b1[25]), .B(exu_n16225), .Y(exu_n28593));
INVX1 exu_U25713(.A(exu_n28593), .Y(exu_n8385));
AND2X1 exu_U25714(.A(shft_lshift4_b1[23]), .B(exu_n16228), .Y(exu_n28595));
INVX1 exu_U25715(.A(exu_n28595), .Y(exu_n8386));
AND2X1 exu_U25716(.A(shft_lshift4_b1[24]), .B(exu_n16226), .Y(exu_n28599));
INVX1 exu_U25717(.A(exu_n28599), .Y(exu_n8387));
AND2X1 exu_U25718(.A(shft_lshift4_b1[22]), .B(exu_n16228), .Y(exu_n28601));
INVX1 exu_U25719(.A(exu_n28601), .Y(exu_n8388));
AND2X1 exu_U25720(.A(shft_lshift4_b1[23]), .B(exu_n16226), .Y(exu_n28605));
INVX1 exu_U25721(.A(exu_n28605), .Y(exu_n8389));
AND2X1 exu_U25722(.A(shft_lshift4_b1[21]), .B(exu_n16228), .Y(exu_n28607));
INVX1 exu_U25723(.A(exu_n28607), .Y(exu_n8390));
AND2X1 exu_U25724(.A(shft_lshift4_b1[22]), .B(exu_n16225), .Y(exu_n28611));
INVX1 exu_U25725(.A(exu_n28611), .Y(exu_n8391));
AND2X1 exu_U25726(.A(shft_lshift4_b1[20]), .B(exu_n16228), .Y(exu_n28613));
INVX1 exu_U25727(.A(exu_n28613), .Y(exu_n8392));
AND2X1 exu_U25728(.A(shft_lshift4_b1[21]), .B(exu_n16226), .Y(exu_n28617));
INVX1 exu_U25729(.A(exu_n28617), .Y(exu_n8393));
AND2X1 exu_U25730(.A(shft_lshift4_b1[19]), .B(exu_n16228), .Y(exu_n28619));
INVX1 exu_U25731(.A(exu_n28619), .Y(exu_n8394));
AND2X1 exu_U25732(.A(shft_lshift4_b1[20]), .B(exu_n16225), .Y(exu_n28623));
INVX1 exu_U25733(.A(exu_n28623), .Y(exu_n8395));
AND2X1 exu_U25734(.A(shft_lshift4_b1[18]), .B(exu_n16228), .Y(exu_n28625));
INVX1 exu_U25735(.A(exu_n28625), .Y(exu_n8396));
AND2X1 exu_U25736(.A(shft_lshift4_b1[19]), .B(exu_n16226), .Y(exu_n28629));
INVX1 exu_U25737(.A(exu_n28629), .Y(exu_n8397));
AND2X1 exu_U25738(.A(shft_lshift4_b1[17]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28631));
INVX1 exu_U25739(.A(exu_n28631), .Y(exu_n8398));
AND2X1 exu_U25740(.A(exu_n28321), .B(exu_n16226), .Y(exu_n28634));
INVX1 exu_U25741(.A(exu_n28634), .Y(exu_n8399));
AND2X1 exu_U25742(.A(shft_lshift4_b1[18]), .B(exu_n16226), .Y(exu_n28638));
INVX1 exu_U25743(.A(exu_n28638), .Y(exu_n8400));
AND2X1 exu_U25744(.A(shft_lshift4_b1[16]), .B(exu_n16228), .Y(exu_n28640));
INVX1 exu_U25745(.A(exu_n28640), .Y(exu_n8401));
AND2X1 exu_U25746(.A(shft_lshift4_b1[17]), .B(exu_n16226), .Y(exu_n28644));
INVX1 exu_U25747(.A(exu_n28644), .Y(exu_n8402));
AND2X1 exu_U25748(.A(shft_lshift4_b1[15]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28646));
INVX1 exu_U25749(.A(exu_n28646), .Y(exu_n8403));
AND2X1 exu_U25750(.A(shft_lshift4_b1[16]), .B(exu_n16225), .Y(exu_n28650));
INVX1 exu_U25751(.A(exu_n28650), .Y(exu_n8404));
AND2X1 exu_U25752(.A(shft_lshift4_b1[14]), .B(exu_n16228), .Y(exu_n28652));
INVX1 exu_U25753(.A(exu_n28652), .Y(exu_n8405));
AND2X1 exu_U25754(.A(shft_lshift4_b1[15]), .B(exu_n16225), .Y(exu_n28656));
INVX1 exu_U25755(.A(exu_n28656), .Y(exu_n8406));
AND2X1 exu_U25756(.A(shft_lshift4_b1[13]), .B(ecl_shft_shift1_e[3]), .Y(exu_n28658));
INVX1 exu_U25757(.A(exu_n28658), .Y(exu_n8407));
AND2X1 exu_U25758(.A(shft_lshift4_b1[14]), .B(exu_n16226), .Y(exu_n28662));
INVX1 exu_U25759(.A(exu_n28662), .Y(exu_n8408));
AND2X1 exu_U25760(.A(shft_lshift4_b1[12]), .B(exu_n16228), .Y(exu_n28664));
INVX1 exu_U25761(.A(exu_n28664), .Y(exu_n8409));
AND2X1 exu_U25762(.A(shft_lshift4_b1[13]), .B(exu_n16225), .Y(exu_n28668));
INVX1 exu_U25763(.A(exu_n28668), .Y(exu_n8410));
AND2X1 exu_U25764(.A(shft_lshift4_b1[11]), .B(exu_n16228), .Y(exu_n28670));
INVX1 exu_U25765(.A(exu_n28670), .Y(exu_n8411));
AND2X1 exu_U25766(.A(shft_lshift4_b1[12]), .B(exu_n16225), .Y(exu_n28674));
INVX1 exu_U25767(.A(exu_n28674), .Y(exu_n8412));
AND2X1 exu_U25768(.A(shft_lshift4_b1[10]), .B(exu_n16228), .Y(exu_n28676));
INVX1 exu_U25769(.A(exu_n28676), .Y(exu_n8413));
AND2X1 exu_U25770(.A(shft_lshift4_b1[11]), .B(exu_n16225), .Y(exu_n28680));
INVX1 exu_U25771(.A(exu_n28680), .Y(exu_n8414));
AND2X1 exu_U25772(.A(shft_lshift4_b1[9]), .B(exu_n16228), .Y(exu_n28682));
INVX1 exu_U25773(.A(exu_n28682), .Y(exu_n8415));
AND2X1 exu_U25774(.A(shft_lshift4_b1[10]), .B(exu_n16226), .Y(exu_n28686));
INVX1 exu_U25775(.A(exu_n28686), .Y(exu_n8416));
AND2X1 exu_U25776(.A(shft_lshift4_b1[8]), .B(exu_n16228), .Y(exu_n28688));
INVX1 exu_U25777(.A(exu_n28688), .Y(exu_n8417));
AND2X1 exu_U25778(.A(shft_lshift4_b1[9]), .B(exu_n16226), .Y(exu_n28692));
INVX1 exu_U25779(.A(exu_n28692), .Y(exu_n8418));
AND2X1 exu_U25780(.A(exu_n15693), .B(exu_n16228), .Y(exu_n28694));
INVX1 exu_U25781(.A(exu_n28694), .Y(exu_n8419));
AND2X1 exu_U25782(.A(ecl_divcntl_n61), .B(exu_n10696), .Y(exu_n28699));
INVX1 exu_U25783(.A(exu_n28699), .Y(exu_n8420));
AND2X1 exu_U25784(.A(exu_n16252), .B(div_curr_q[9]), .Y(exu_n28701));
INVX1 exu_U25785(.A(exu_n28701), .Y(exu_n8421));
AND2X1 exu_U25786(.A(exu_n11892), .B(ecl_divcntl_n61), .Y(exu_n28705));
INVX1 exu_U25787(.A(exu_n28705), .Y(exu_n8422));
AND2X1 exu_U25788(.A(div_curr_q[8]), .B(exu_n16252), .Y(exu_n28707));
INVX1 exu_U25789(.A(exu_n28707), .Y(exu_n8423));
AND2X1 exu_U25790(.A(exu_n11893), .B(ecl_divcntl_n61), .Y(exu_n28711));
INVX1 exu_U25791(.A(exu_n28711), .Y(exu_n8424));
AND2X1 exu_U25792(.A(div_curr_q[7]), .B(ecl_div_sel_64b), .Y(exu_n28713));
INVX1 exu_U25793(.A(exu_n28713), .Y(exu_n8425));
AND2X1 exu_U25794(.A(exu_n11894), .B(ecl_divcntl_n61), .Y(exu_n28717));
INVX1 exu_U25795(.A(exu_n28717), .Y(exu_n8426));
AND2X1 exu_U25796(.A(div_curr_q[6]), .B(ecl_div_sel_64b), .Y(exu_n28719));
INVX1 exu_U25797(.A(exu_n28719), .Y(exu_n8427));
AND2X1 exu_U25798(.A(exu_n11895), .B(ecl_divcntl_n61), .Y(exu_n28727));
INVX1 exu_U25799(.A(exu_n28727), .Y(exu_n8428));
AND2X1 exu_U25800(.A(div_curr_q[5]), .B(ecl_div_sel_64b), .Y(exu_n28729));
INVX1 exu_U25801(.A(exu_n28729), .Y(exu_n8429));
AND2X1 exu_U25802(.A(exu_n11896), .B(ecl_divcntl_n61), .Y(exu_n28743));
INVX1 exu_U25803(.A(exu_n28743), .Y(exu_n8430));
AND2X1 exu_U25804(.A(div_curr_q[4]), .B(exu_n16252), .Y(exu_n28745));
INVX1 exu_U25805(.A(exu_n28745), .Y(exu_n8431));
AND2X1 exu_U25806(.A(exu_n11897), .B(ecl_divcntl_n61), .Y(exu_n28759));
INVX1 exu_U25807(.A(exu_n28759), .Y(exu_n8432));
AND2X1 exu_U25808(.A(div_curr_q[3]), .B(ecl_div_sel_64b), .Y(exu_n28761));
INVX1 exu_U25809(.A(exu_n28761), .Y(exu_n8433));
AND2X1 exu_U25810(.A(div_curr_q[31]), .B(exu_n16252), .Y(exu_n28772));
INVX1 exu_U25811(.A(exu_n28772), .Y(exu_n8434));
AND2X1 exu_U25812(.A(exu_n11898), .B(ecl_divcntl_n61), .Y(exu_n28776));
INVX1 exu_U25813(.A(exu_n28776), .Y(exu_n8435));
AND2X1 exu_U25814(.A(div_curr_q[30]), .B(ecl_div_sel_64b), .Y(exu_n28778));
INVX1 exu_U25815(.A(exu_n28778), .Y(exu_n8436));
AND2X1 exu_U25816(.A(exu_n11899), .B(ecl_divcntl_n61), .Y(exu_n28782));
INVX1 exu_U25817(.A(exu_n28782), .Y(exu_n8437));
AND2X1 exu_U25818(.A(div_curr_q[2]), .B(ecl_div_sel_64b), .Y(exu_n28784));
INVX1 exu_U25819(.A(exu_n28784), .Y(exu_n8438));
AND2X1 exu_U25820(.A(exu_n11900), .B(ecl_divcntl_n61), .Y(exu_n28788));
INVX1 exu_U25821(.A(exu_n28788), .Y(exu_n8439));
AND2X1 exu_U25822(.A(div_curr_q[29]), .B(ecl_div_sel_64b), .Y(exu_n28790));
INVX1 exu_U25823(.A(exu_n28790), .Y(exu_n8440));
AND2X1 exu_U25824(.A(exu_n11901), .B(ecl_divcntl_n61), .Y(exu_n28794));
INVX1 exu_U25825(.A(exu_n28794), .Y(exu_n8441));
AND2X1 exu_U25826(.A(div_curr_q[28]), .B(ecl_div_sel_64b), .Y(exu_n28796));
INVX1 exu_U25827(.A(exu_n28796), .Y(exu_n8442));
AND2X1 exu_U25828(.A(exu_n11902), .B(ecl_divcntl_n61), .Y(exu_n28800));
INVX1 exu_U25829(.A(exu_n28800), .Y(exu_n8443));
AND2X1 exu_U25830(.A(div_curr_q[27]), .B(ecl_div_sel_64b), .Y(exu_n28802));
INVX1 exu_U25831(.A(exu_n28802), .Y(exu_n8444));
AND2X1 exu_U25832(.A(exu_n11903), .B(ecl_divcntl_n61), .Y(exu_n28806));
INVX1 exu_U25833(.A(exu_n28806), .Y(exu_n8445));
AND2X1 exu_U25834(.A(div_curr_q[26]), .B(ecl_div_sel_64b), .Y(exu_n28808));
INVX1 exu_U25835(.A(exu_n28808), .Y(exu_n8446));
AND2X1 exu_U25836(.A(exu_n11904), .B(ecl_divcntl_n61), .Y(exu_n28812));
INVX1 exu_U25837(.A(exu_n28812), .Y(exu_n8447));
AND2X1 exu_U25838(.A(div_curr_q[25]), .B(ecl_div_sel_64b), .Y(exu_n28814));
INVX1 exu_U25839(.A(exu_n28814), .Y(exu_n8448));
AND2X1 exu_U25840(.A(exu_n11905), .B(ecl_divcntl_n61), .Y(exu_n28818));
INVX1 exu_U25841(.A(exu_n28818), .Y(exu_n8449));
AND2X1 exu_U25842(.A(div_curr_q[24]), .B(ecl_div_sel_64b), .Y(exu_n28820));
INVX1 exu_U25843(.A(exu_n28820), .Y(exu_n8450));
AND2X1 exu_U25844(.A(exu_n11906), .B(ecl_divcntl_n61), .Y(exu_n28824));
INVX1 exu_U25845(.A(exu_n28824), .Y(exu_n8451));
AND2X1 exu_U25846(.A(div_curr_q[23]), .B(ecl_div_sel_64b), .Y(exu_n28826));
INVX1 exu_U25847(.A(exu_n28826), .Y(exu_n8452));
AND2X1 exu_U25848(.A(exu_n11907), .B(ecl_divcntl_n61), .Y(exu_n28830));
INVX1 exu_U25849(.A(exu_n28830), .Y(exu_n8453));
AND2X1 exu_U25850(.A(div_curr_q[22]), .B(exu_n16252), .Y(exu_n28832));
INVX1 exu_U25851(.A(exu_n28832), .Y(exu_n8454));
AND2X1 exu_U25852(.A(exu_n11908), .B(ecl_divcntl_n61), .Y(exu_n28836));
INVX1 exu_U25853(.A(exu_n28836), .Y(exu_n8455));
AND2X1 exu_U25854(.A(div_curr_q[21]), .B(exu_n16252), .Y(exu_n28838));
INVX1 exu_U25855(.A(exu_n28838), .Y(exu_n8456));
AND2X1 exu_U25856(.A(exu_n11909), .B(ecl_divcntl_n61), .Y(exu_n28842));
INVX1 exu_U25857(.A(exu_n28842), .Y(exu_n8457));
AND2X1 exu_U25858(.A(div_curr_q[20]), .B(ecl_div_sel_64b), .Y(exu_n28844));
INVX1 exu_U25859(.A(exu_n28844), .Y(exu_n8458));
AND2X1 exu_U25860(.A(exu_n11910), .B(ecl_divcntl_n61), .Y(exu_n28848));
INVX1 exu_U25861(.A(exu_n28848), .Y(exu_n8459));
AND2X1 exu_U25862(.A(div_curr_q[1]), .B(ecl_div_sel_64b), .Y(exu_n28850));
INVX1 exu_U25863(.A(exu_n28850), .Y(exu_n8460));
AND2X1 exu_U25864(.A(exu_n11911), .B(ecl_divcntl_n61), .Y(exu_n28854));
INVX1 exu_U25865(.A(exu_n28854), .Y(exu_n8461));
AND2X1 exu_U25866(.A(div_curr_q[19]), .B(ecl_div_sel_64b), .Y(exu_n28856));
INVX1 exu_U25867(.A(exu_n28856), .Y(exu_n8462));
AND2X1 exu_U25868(.A(exu_n11912), .B(ecl_divcntl_n61), .Y(exu_n28860));
INVX1 exu_U25869(.A(exu_n28860), .Y(exu_n8463));
AND2X1 exu_U25870(.A(div_curr_q[18]), .B(ecl_div_sel_64b), .Y(exu_n28862));
INVX1 exu_U25871(.A(exu_n28862), .Y(exu_n8464));
AND2X1 exu_U25872(.A(exu_n11913), .B(ecl_divcntl_n61), .Y(exu_n28866));
INVX1 exu_U25873(.A(exu_n28866), .Y(exu_n8465));
AND2X1 exu_U25874(.A(div_curr_q[17]), .B(exu_n16252), .Y(exu_n28868));
INVX1 exu_U25875(.A(exu_n28868), .Y(exu_n8466));
AND2X1 exu_U25876(.A(exu_n11914), .B(ecl_divcntl_n61), .Y(exu_n28872));
INVX1 exu_U25877(.A(exu_n28872), .Y(exu_n8467));
AND2X1 exu_U25878(.A(div_curr_q[16]), .B(exu_n16252), .Y(exu_n28874));
INVX1 exu_U25879(.A(exu_n28874), .Y(exu_n8468));
AND2X1 exu_U25880(.A(exu_n11915), .B(ecl_divcntl_n61), .Y(exu_n28878));
INVX1 exu_U25881(.A(exu_n28878), .Y(exu_n8469));
AND2X1 exu_U25882(.A(div_curr_q[15]), .B(exu_n16252), .Y(exu_n28880));
INVX1 exu_U25883(.A(exu_n28880), .Y(exu_n8470));
AND2X1 exu_U25884(.A(exu_n11916), .B(ecl_divcntl_n61), .Y(exu_n28884));
INVX1 exu_U25885(.A(exu_n28884), .Y(exu_n8471));
AND2X1 exu_U25886(.A(div_curr_q[14]), .B(exu_n16252), .Y(exu_n28886));
INVX1 exu_U25887(.A(exu_n28886), .Y(exu_n8472));
AND2X1 exu_U25888(.A(exu_n11917), .B(ecl_divcntl_n61), .Y(exu_n28890));
INVX1 exu_U25889(.A(exu_n28890), .Y(exu_n8473));
AND2X1 exu_U25890(.A(div_curr_q[13]), .B(exu_n16252), .Y(exu_n28892));
INVX1 exu_U25891(.A(exu_n28892), .Y(exu_n8474));
AND2X1 exu_U25892(.A(exu_n11918), .B(ecl_divcntl_n61), .Y(exu_n28896));
INVX1 exu_U25893(.A(exu_n28896), .Y(exu_n8475));
AND2X1 exu_U25894(.A(div_curr_q[12]), .B(exu_n16252), .Y(exu_n28898));
INVX1 exu_U25895(.A(exu_n28898), .Y(exu_n8476));
AND2X1 exu_U25896(.A(exu_n11919), .B(ecl_divcntl_n61), .Y(exu_n28902));
INVX1 exu_U25897(.A(exu_n28902), .Y(exu_n8477));
AND2X1 exu_U25898(.A(div_curr_q[11]), .B(exu_n16252), .Y(exu_n28904));
INVX1 exu_U25899(.A(exu_n28904), .Y(exu_n8478));
AND2X1 exu_U25900(.A(exu_n11920), .B(ecl_divcntl_n61), .Y(exu_n28908));
INVX1 exu_U25901(.A(exu_n28908), .Y(exu_n8479));
AND2X1 exu_U25902(.A(div_curr_q[10]), .B(exu_n16252), .Y(exu_n28910));
INVX1 exu_U25903(.A(exu_n28910), .Y(exu_n8480));
AND2X1 exu_U25904(.A(exu_n11921), .B(ecl_divcntl_n61), .Y(exu_n28914));
INVX1 exu_U25905(.A(exu_n28914), .Y(exu_n8481));
AND2X1 exu_U25906(.A(div_curr_q[0]), .B(ecl_div_sel_64b), .Y(exu_n28916));
INVX1 exu_U25907(.A(exu_n28916), .Y(exu_n8482));
AND2X1 exu_U25908(.A(exu_n16238), .B(alu_logic_result_xor[9]), .Y(exu_n28920));
INVX1 exu_U25909(.A(exu_n28920), .Y(exu_n8483));
AND2X1 exu_U25910(.A(exu_n16240), .B(alu_logic_result_and[9]), .Y(exu_n28922));
INVX1 exu_U25911(.A(exu_n28922), .Y(exu_n8484));
AND2X1 exu_U25912(.A(alu_logic_result_xor[8]), .B(exu_n16238), .Y(exu_n28926));
INVX1 exu_U25913(.A(exu_n28926), .Y(exu_n8485));
AND2X1 exu_U25914(.A(alu_logic_result_and[8]), .B(exu_n16240), .Y(exu_n28928));
INVX1 exu_U25915(.A(exu_n28928), .Y(exu_n8486));
AND2X1 exu_U25916(.A(alu_logic_result_xor[7]), .B(exu_n16238), .Y(exu_n28932));
INVX1 exu_U25917(.A(exu_n28932), .Y(exu_n8487));
AND2X1 exu_U25918(.A(alu_logic_result_and[7]), .B(exu_n16240), .Y(exu_n28934));
INVX1 exu_U25919(.A(exu_n28934), .Y(exu_n8488));
AND2X1 exu_U25920(.A(alu_logic_result_xor[6]), .B(exu_n16238), .Y(exu_n28938));
INVX1 exu_U25921(.A(exu_n28938), .Y(exu_n8489));
AND2X1 exu_U25922(.A(alu_logic_result_and[6]), .B(exu_n16240), .Y(exu_n28940));
INVX1 exu_U25923(.A(exu_n28940), .Y(exu_n8490));
AND2X1 exu_U25924(.A(alu_logic_result_xor[63]), .B(exu_n16238), .Y(exu_n28944));
INVX1 exu_U25925(.A(exu_n28944), .Y(exu_n8491));
AND2X1 exu_U25926(.A(alu_logic_result_and[63]), .B(exu_n16240), .Y(exu_n28946));
INVX1 exu_U25927(.A(exu_n28946), .Y(exu_n8492));
AND2X1 exu_U25928(.A(alu_logic_result_xor[62]), .B(exu_n16238), .Y(exu_n28950));
INVX1 exu_U25929(.A(exu_n28950), .Y(exu_n8493));
AND2X1 exu_U25930(.A(alu_logic_result_and[62]), .B(exu_n16240), .Y(exu_n28952));
INVX1 exu_U25931(.A(exu_n28952), .Y(exu_n8494));
AND2X1 exu_U25932(.A(alu_logic_result_xor[61]), .B(exu_n16238), .Y(exu_n28956));
INVX1 exu_U25933(.A(exu_n28956), .Y(exu_n8495));
AND2X1 exu_U25934(.A(alu_logic_result_and[61]), .B(exu_n16240), .Y(exu_n28958));
INVX1 exu_U25935(.A(exu_n28958), .Y(exu_n8496));
AND2X1 exu_U25936(.A(alu_logic_result_xor[60]), .B(exu_n16238), .Y(exu_n28962));
INVX1 exu_U25937(.A(exu_n28962), .Y(exu_n8497));
AND2X1 exu_U25938(.A(alu_logic_result_and[60]), .B(exu_n16240), .Y(exu_n28964));
INVX1 exu_U25939(.A(exu_n28964), .Y(exu_n8498));
AND2X1 exu_U25940(.A(alu_logic_result_xor[5]), .B(exu_n16238), .Y(exu_n28968));
INVX1 exu_U25941(.A(exu_n28968), .Y(exu_n8499));
AND2X1 exu_U25942(.A(alu_logic_result_and[5]), .B(exu_n16240), .Y(exu_n28970));
INVX1 exu_U25943(.A(exu_n28970), .Y(exu_n8500));
AND2X1 exu_U25944(.A(alu_logic_result_xor[59]), .B(exu_n16238), .Y(exu_n28974));
INVX1 exu_U25945(.A(exu_n28974), .Y(exu_n8501));
AND2X1 exu_U25946(.A(alu_logic_result_and[59]), .B(exu_n16240), .Y(exu_n28976));
INVX1 exu_U25947(.A(exu_n28976), .Y(exu_n8502));
AND2X1 exu_U25948(.A(alu_logic_result_xor[58]), .B(exu_n16238), .Y(exu_n28980));
INVX1 exu_U25949(.A(exu_n28980), .Y(exu_n8503));
AND2X1 exu_U25950(.A(alu_logic_result_and[58]), .B(exu_n16240), .Y(exu_n28982));
INVX1 exu_U25951(.A(exu_n28982), .Y(exu_n8504));
AND2X1 exu_U25952(.A(alu_logic_result_xor[57]), .B(exu_n16238), .Y(exu_n28986));
INVX1 exu_U25953(.A(exu_n28986), .Y(exu_n8505));
AND2X1 exu_U25954(.A(alu_logic_result_and[57]), .B(exu_n16240), .Y(exu_n28988));
INVX1 exu_U25955(.A(exu_n28988), .Y(exu_n8506));
AND2X1 exu_U25956(.A(alu_logic_result_xor[56]), .B(exu_n16238), .Y(exu_n28992));
INVX1 exu_U25957(.A(exu_n28992), .Y(exu_n8507));
AND2X1 exu_U25958(.A(alu_logic_result_and[56]), .B(exu_n16240), .Y(exu_n28994));
INVX1 exu_U25959(.A(exu_n28994), .Y(exu_n8508));
AND2X1 exu_U25960(.A(alu_logic_result_xor[55]), .B(exu_n16238), .Y(exu_n28998));
INVX1 exu_U25961(.A(exu_n28998), .Y(exu_n8509));
AND2X1 exu_U25962(.A(alu_logic_result_and[55]), .B(exu_n16240), .Y(exu_n29000));
INVX1 exu_U25963(.A(exu_n29000), .Y(exu_n8510));
AND2X1 exu_U25964(.A(alu_logic_result_xor[54]), .B(exu_n16238), .Y(exu_n29004));
INVX1 exu_U25965(.A(exu_n29004), .Y(exu_n8511));
AND2X1 exu_U25966(.A(alu_logic_result_and[54]), .B(exu_n16240), .Y(exu_n29006));
INVX1 exu_U25967(.A(exu_n29006), .Y(exu_n8512));
AND2X1 exu_U25968(.A(alu_logic_result_xor[53]), .B(exu_n16238), .Y(exu_n29010));
INVX1 exu_U25969(.A(exu_n29010), .Y(exu_n8513));
AND2X1 exu_U25970(.A(alu_logic_result_and[53]), .B(exu_n16240), .Y(exu_n29012));
INVX1 exu_U25971(.A(exu_n29012), .Y(exu_n8514));
AND2X1 exu_U25972(.A(alu_logic_result_xor[52]), .B(exu_n16238), .Y(exu_n29016));
INVX1 exu_U25973(.A(exu_n29016), .Y(exu_n8515));
AND2X1 exu_U25974(.A(alu_logic_result_and[52]), .B(exu_n16240), .Y(exu_n29018));
INVX1 exu_U25975(.A(exu_n29018), .Y(exu_n8516));
AND2X1 exu_U25976(.A(alu_logic_result_xor[51]), .B(exu_n16238), .Y(exu_n29022));
INVX1 exu_U25977(.A(exu_n29022), .Y(exu_n8517));
AND2X1 exu_U25978(.A(alu_logic_result_and[51]), .B(exu_n16240), .Y(exu_n29024));
INVX1 exu_U25979(.A(exu_n29024), .Y(exu_n8518));
AND2X1 exu_U25980(.A(alu_logic_result_xor[50]), .B(exu_n16238), .Y(exu_n29028));
INVX1 exu_U25981(.A(exu_n29028), .Y(exu_n8519));
AND2X1 exu_U25982(.A(alu_logic_result_and[50]), .B(exu_n16240), .Y(exu_n29030));
INVX1 exu_U25983(.A(exu_n29030), .Y(exu_n8520));
AND2X1 exu_U25984(.A(alu_logic_result_xor[4]), .B(exu_n16238), .Y(exu_n29034));
INVX1 exu_U25985(.A(exu_n29034), .Y(exu_n8521));
AND2X1 exu_U25986(.A(alu_logic_result_and[4]), .B(exu_n16240), .Y(exu_n29036));
INVX1 exu_U25987(.A(exu_n29036), .Y(exu_n8522));
AND2X1 exu_U25988(.A(alu_logic_result_xor[49]), .B(exu_n16238), .Y(exu_n29040));
INVX1 exu_U25989(.A(exu_n29040), .Y(exu_n8523));
AND2X1 exu_U25990(.A(alu_logic_result_and[49]), .B(exu_n16240), .Y(exu_n29042));
INVX1 exu_U25991(.A(exu_n29042), .Y(exu_n8524));
AND2X1 exu_U25992(.A(alu_logic_result_xor[48]), .B(exu_n16238), .Y(exu_n29046));
INVX1 exu_U25993(.A(exu_n29046), .Y(exu_n8525));
AND2X1 exu_U25994(.A(alu_logic_result_and[48]), .B(exu_n16240), .Y(exu_n29048));
INVX1 exu_U25995(.A(exu_n29048), .Y(exu_n8526));
AND2X1 exu_U25996(.A(alu_logic_result_xor[47]), .B(exu_n16238), .Y(exu_n29052));
INVX1 exu_U25997(.A(exu_n29052), .Y(exu_n8527));
AND2X1 exu_U25998(.A(alu_logic_result_and[47]), .B(exu_n16240), .Y(exu_n29054));
INVX1 exu_U25999(.A(exu_n29054), .Y(exu_n8528));
AND2X1 exu_U26000(.A(alu_logic_result_xor[46]), .B(exu_n16238), .Y(exu_n29058));
INVX1 exu_U26001(.A(exu_n29058), .Y(exu_n8529));
AND2X1 exu_U26002(.A(alu_logic_result_and[46]), .B(exu_n16240), .Y(exu_n29060));
INVX1 exu_U26003(.A(exu_n29060), .Y(exu_n8530));
AND2X1 exu_U26004(.A(alu_logic_result_xor[45]), .B(exu_n16238), .Y(exu_n29064));
INVX1 exu_U26005(.A(exu_n29064), .Y(exu_n8531));
AND2X1 exu_U26006(.A(alu_logic_result_and[45]), .B(exu_n16240), .Y(exu_n29066));
INVX1 exu_U26007(.A(exu_n29066), .Y(exu_n8532));
AND2X1 exu_U26008(.A(alu_logic_result_xor[44]), .B(exu_n16238), .Y(exu_n29070));
INVX1 exu_U26009(.A(exu_n29070), .Y(exu_n8533));
AND2X1 exu_U26010(.A(alu_logic_result_and[44]), .B(exu_n16240), .Y(exu_n29072));
INVX1 exu_U26011(.A(exu_n29072), .Y(exu_n8534));
AND2X1 exu_U26012(.A(alu_logic_result_xor[43]), .B(exu_n16238), .Y(exu_n29076));
INVX1 exu_U26013(.A(exu_n29076), .Y(exu_n8535));
AND2X1 exu_U26014(.A(alu_logic_result_and[43]), .B(exu_n16240), .Y(exu_n29078));
INVX1 exu_U26015(.A(exu_n29078), .Y(exu_n8536));
AND2X1 exu_U26016(.A(alu_logic_result_xor[42]), .B(exu_n16238), .Y(exu_n29082));
INVX1 exu_U26017(.A(exu_n29082), .Y(exu_n8537));
AND2X1 exu_U26018(.A(alu_logic_result_and[42]), .B(exu_n16240), .Y(exu_n29084));
INVX1 exu_U26019(.A(exu_n29084), .Y(exu_n8538));
AND2X1 exu_U26020(.A(alu_logic_result_xor[41]), .B(exu_n16238), .Y(exu_n29088));
INVX1 exu_U26021(.A(exu_n29088), .Y(exu_n8539));
AND2X1 exu_U26022(.A(alu_logic_result_and[41]), .B(exu_n16240), .Y(exu_n29090));
INVX1 exu_U26023(.A(exu_n29090), .Y(exu_n8540));
AND2X1 exu_U26024(.A(alu_logic_result_xor[40]), .B(exu_n16238), .Y(exu_n29094));
INVX1 exu_U26025(.A(exu_n29094), .Y(exu_n8541));
AND2X1 exu_U26026(.A(alu_logic_result_and[40]), .B(exu_n16240), .Y(exu_n29096));
INVX1 exu_U26027(.A(exu_n29096), .Y(exu_n8542));
AND2X1 exu_U26028(.A(alu_logic_result_xor[3]), .B(exu_n16238), .Y(exu_n29100));
INVX1 exu_U26029(.A(exu_n29100), .Y(exu_n8543));
AND2X1 exu_U26030(.A(alu_logic_result_and[3]), .B(exu_n16240), .Y(exu_n29102));
INVX1 exu_U26031(.A(exu_n29102), .Y(exu_n8544));
AND2X1 exu_U26032(.A(alu_logic_result_xor[39]), .B(exu_n16238), .Y(exu_n29106));
INVX1 exu_U26033(.A(exu_n29106), .Y(exu_n8545));
AND2X1 exu_U26034(.A(alu_logic_result_and[39]), .B(exu_n16240), .Y(exu_n29108));
INVX1 exu_U26035(.A(exu_n29108), .Y(exu_n8546));
AND2X1 exu_U26036(.A(alu_logic_result_xor[38]), .B(exu_n16238), .Y(exu_n29112));
INVX1 exu_U26037(.A(exu_n29112), .Y(exu_n8547));
AND2X1 exu_U26038(.A(alu_logic_result_and[38]), .B(exu_n16240), .Y(exu_n29114));
INVX1 exu_U26039(.A(exu_n29114), .Y(exu_n8548));
AND2X1 exu_U26040(.A(alu_logic_result_xor[37]), .B(exu_n16238), .Y(exu_n29118));
INVX1 exu_U26041(.A(exu_n29118), .Y(exu_n8549));
AND2X1 exu_U26042(.A(alu_logic_result_and[37]), .B(exu_n16240), .Y(exu_n29120));
INVX1 exu_U26043(.A(exu_n29120), .Y(exu_n8550));
AND2X1 exu_U26044(.A(alu_logic_result_xor[36]), .B(exu_n16238), .Y(exu_n29124));
INVX1 exu_U26045(.A(exu_n29124), .Y(exu_n8551));
AND2X1 exu_U26046(.A(alu_logic_result_and[36]), .B(exu_n16240), .Y(exu_n29126));
INVX1 exu_U26047(.A(exu_n29126), .Y(exu_n8552));
AND2X1 exu_U26048(.A(alu_logic_result_xor[35]), .B(exu_n16238), .Y(exu_n29130));
INVX1 exu_U26049(.A(exu_n29130), .Y(exu_n8553));
AND2X1 exu_U26050(.A(alu_logic_result_and[35]), .B(exu_n16240), .Y(exu_n29132));
INVX1 exu_U26051(.A(exu_n29132), .Y(exu_n8554));
AND2X1 exu_U26052(.A(alu_logic_result_xor[34]), .B(exu_n16238), .Y(exu_n29136));
INVX1 exu_U26053(.A(exu_n29136), .Y(exu_n8555));
AND2X1 exu_U26054(.A(alu_logic_result_and[34]), .B(exu_n16240), .Y(exu_n29138));
INVX1 exu_U26055(.A(exu_n29138), .Y(exu_n8556));
AND2X1 exu_U26056(.A(alu_logic_result_xor[33]), .B(exu_n16238), .Y(exu_n29142));
INVX1 exu_U26057(.A(exu_n29142), .Y(exu_n8557));
AND2X1 exu_U26058(.A(alu_logic_result_and[33]), .B(exu_n16240), .Y(exu_n29144));
INVX1 exu_U26059(.A(exu_n29144), .Y(exu_n8558));
AND2X1 exu_U26060(.A(alu_logic_result_xor[32]), .B(exu_n16238), .Y(exu_n29148));
INVX1 exu_U26061(.A(exu_n29148), .Y(exu_n8559));
AND2X1 exu_U26062(.A(alu_logic_result_and[32]), .B(exu_n16240), .Y(exu_n29150));
INVX1 exu_U26063(.A(exu_n29150), .Y(exu_n8560));
AND2X1 exu_U26064(.A(alu_logic_result_xor[31]), .B(exu_n16238), .Y(exu_n29154));
INVX1 exu_U26065(.A(exu_n29154), .Y(exu_n8561));
AND2X1 exu_U26066(.A(alu_logic_result_and[31]), .B(exu_n16240), .Y(exu_n29156));
INVX1 exu_U26067(.A(exu_n29156), .Y(exu_n8562));
AND2X1 exu_U26068(.A(alu_logic_result_xor[30]), .B(exu_n16238), .Y(exu_n29160));
INVX1 exu_U26069(.A(exu_n29160), .Y(exu_n8563));
AND2X1 exu_U26070(.A(alu_logic_result_and[30]), .B(exu_n16240), .Y(exu_n29162));
INVX1 exu_U26071(.A(exu_n29162), .Y(exu_n8564));
AND2X1 exu_U26072(.A(alu_logic_result_xor[2]), .B(exu_n16238), .Y(exu_n29166));
INVX1 exu_U26073(.A(exu_n29166), .Y(exu_n8565));
AND2X1 exu_U26074(.A(alu_logic_result_and[2]), .B(exu_n16240), .Y(exu_n29168));
INVX1 exu_U26075(.A(exu_n29168), .Y(exu_n8566));
AND2X1 exu_U26076(.A(alu_logic_result_xor[29]), .B(exu_n16238), .Y(exu_n29172));
INVX1 exu_U26077(.A(exu_n29172), .Y(exu_n8567));
AND2X1 exu_U26078(.A(alu_logic_result_and[29]), .B(exu_n16240), .Y(exu_n29174));
INVX1 exu_U26079(.A(exu_n29174), .Y(exu_n8568));
AND2X1 exu_U26080(.A(alu_logic_result_xor[28]), .B(exu_n16238), .Y(exu_n29178));
INVX1 exu_U26081(.A(exu_n29178), .Y(exu_n8569));
AND2X1 exu_U26082(.A(alu_logic_result_and[28]), .B(exu_n16240), .Y(exu_n29180));
INVX1 exu_U26083(.A(exu_n29180), .Y(exu_n8570));
AND2X1 exu_U26084(.A(alu_logic_result_xor[27]), .B(exu_n16238), .Y(exu_n29184));
INVX1 exu_U26085(.A(exu_n29184), .Y(exu_n8571));
AND2X1 exu_U26086(.A(alu_logic_result_and[27]), .B(exu_n16240), .Y(exu_n29186));
INVX1 exu_U26087(.A(exu_n29186), .Y(exu_n8572));
AND2X1 exu_U26088(.A(alu_logic_result_xor[26]), .B(exu_n16238), .Y(exu_n29190));
INVX1 exu_U26089(.A(exu_n29190), .Y(exu_n8573));
AND2X1 exu_U26090(.A(alu_logic_result_and[26]), .B(exu_n16240), .Y(exu_n29192));
INVX1 exu_U26091(.A(exu_n29192), .Y(exu_n8574));
AND2X1 exu_U26092(.A(alu_logic_result_xor[25]), .B(exu_n16238), .Y(exu_n29196));
INVX1 exu_U26093(.A(exu_n29196), .Y(exu_n8575));
AND2X1 exu_U26094(.A(alu_logic_result_and[25]), .B(exu_n16240), .Y(exu_n29198));
INVX1 exu_U26095(.A(exu_n29198), .Y(exu_n8576));
AND2X1 exu_U26096(.A(alu_logic_result_xor[24]), .B(exu_n16238), .Y(exu_n29202));
INVX1 exu_U26097(.A(exu_n29202), .Y(exu_n8577));
AND2X1 exu_U26098(.A(alu_logic_result_and[24]), .B(exu_n16240), .Y(exu_n29204));
INVX1 exu_U26099(.A(exu_n29204), .Y(exu_n8578));
AND2X1 exu_U26100(.A(alu_logic_result_xor[23]), .B(exu_n16238), .Y(exu_n29208));
INVX1 exu_U26101(.A(exu_n29208), .Y(exu_n8579));
AND2X1 exu_U26102(.A(alu_logic_result_and[23]), .B(exu_n16240), .Y(exu_n29210));
INVX1 exu_U26103(.A(exu_n29210), .Y(exu_n8580));
AND2X1 exu_U26104(.A(alu_logic_result_xor[22]), .B(exu_n16238), .Y(exu_n29214));
INVX1 exu_U26105(.A(exu_n29214), .Y(exu_n8581));
AND2X1 exu_U26106(.A(alu_logic_result_and[22]), .B(exu_n16240), .Y(exu_n29216));
INVX1 exu_U26107(.A(exu_n29216), .Y(exu_n8582));
AND2X1 exu_U26108(.A(alu_logic_result_xor[21]), .B(exu_n16238), .Y(exu_n29220));
INVX1 exu_U26109(.A(exu_n29220), .Y(exu_n8583));
AND2X1 exu_U26110(.A(alu_logic_result_and[21]), .B(exu_n16240), .Y(exu_n29222));
INVX1 exu_U26111(.A(exu_n29222), .Y(exu_n8584));
AND2X1 exu_U26112(.A(alu_logic_result_xor[20]), .B(exu_n16238), .Y(exu_n29226));
INVX1 exu_U26113(.A(exu_n29226), .Y(exu_n8585));
AND2X1 exu_U26114(.A(alu_logic_result_and[20]), .B(exu_n16240), .Y(exu_n29228));
INVX1 exu_U26115(.A(exu_n29228), .Y(exu_n8586));
AND2X1 exu_U26116(.A(alu_logic_result_xor[1]), .B(exu_n16238), .Y(exu_n29232));
INVX1 exu_U26117(.A(exu_n29232), .Y(exu_n8587));
AND2X1 exu_U26118(.A(alu_logic_result_and[1]), .B(exu_n16240), .Y(exu_n29234));
INVX1 exu_U26119(.A(exu_n29234), .Y(exu_n8588));
AND2X1 exu_U26120(.A(alu_logic_result_xor[19]), .B(exu_n16238), .Y(exu_n29238));
INVX1 exu_U26121(.A(exu_n29238), .Y(exu_n8589));
AND2X1 exu_U26122(.A(alu_logic_result_and[19]), .B(exu_n16240), .Y(exu_n29240));
INVX1 exu_U26123(.A(exu_n29240), .Y(exu_n8590));
AND2X1 exu_U26124(.A(alu_logic_result_xor[18]), .B(exu_n16238), .Y(exu_n29244));
INVX1 exu_U26125(.A(exu_n29244), .Y(exu_n8591));
AND2X1 exu_U26126(.A(alu_logic_result_and[18]), .B(exu_n16240), .Y(exu_n29246));
INVX1 exu_U26127(.A(exu_n29246), .Y(exu_n8592));
AND2X1 exu_U26128(.A(alu_logic_result_xor[17]), .B(exu_n16238), .Y(exu_n29250));
INVX1 exu_U26129(.A(exu_n29250), .Y(exu_n8593));
AND2X1 exu_U26130(.A(alu_logic_result_and[17]), .B(exu_n16240), .Y(exu_n29252));
INVX1 exu_U26131(.A(exu_n29252), .Y(exu_n8594));
AND2X1 exu_U26132(.A(alu_logic_result_xor[16]), .B(exu_n16238), .Y(exu_n29256));
INVX1 exu_U26133(.A(exu_n29256), .Y(exu_n8595));
AND2X1 exu_U26134(.A(alu_logic_result_and[16]), .B(exu_n16240), .Y(exu_n29258));
INVX1 exu_U26135(.A(exu_n29258), .Y(exu_n8596));
AND2X1 exu_U26136(.A(alu_logic_result_xor[15]), .B(exu_n16238), .Y(exu_n29262));
INVX1 exu_U26137(.A(exu_n29262), .Y(exu_n8597));
AND2X1 exu_U26138(.A(alu_logic_result_and[15]), .B(exu_n16240), .Y(exu_n29264));
INVX1 exu_U26139(.A(exu_n29264), .Y(exu_n8598));
AND2X1 exu_U26140(.A(alu_logic_result_xor[14]), .B(exu_n16238), .Y(exu_n29268));
INVX1 exu_U26141(.A(exu_n29268), .Y(exu_n8599));
AND2X1 exu_U26142(.A(alu_logic_result_and[14]), .B(exu_n16240), .Y(exu_n29270));
INVX1 exu_U26143(.A(exu_n29270), .Y(exu_n8600));
AND2X1 exu_U26144(.A(alu_logic_result_xor[13]), .B(exu_n16238), .Y(exu_n29274));
INVX1 exu_U26145(.A(exu_n29274), .Y(exu_n8601));
AND2X1 exu_U26146(.A(alu_logic_result_and[13]), .B(exu_n16240), .Y(exu_n29276));
INVX1 exu_U26147(.A(exu_n29276), .Y(exu_n8602));
AND2X1 exu_U26148(.A(alu_logic_result_xor[12]), .B(exu_n16238), .Y(exu_n29280));
INVX1 exu_U26149(.A(exu_n29280), .Y(exu_n8603));
AND2X1 exu_U26150(.A(alu_logic_result_and[12]), .B(exu_n16240), .Y(exu_n29282));
INVX1 exu_U26151(.A(exu_n29282), .Y(exu_n8604));
AND2X1 exu_U26152(.A(alu_logic_result_xor[11]), .B(exu_n16238), .Y(exu_n29286));
INVX1 exu_U26153(.A(exu_n29286), .Y(exu_n8605));
AND2X1 exu_U26154(.A(alu_logic_result_and[11]), .B(exu_n16240), .Y(exu_n29288));
INVX1 exu_U26155(.A(exu_n29288), .Y(exu_n8606));
AND2X1 exu_U26156(.A(alu_logic_result_xor[10]), .B(exu_n16238), .Y(exu_n29292));
INVX1 exu_U26157(.A(exu_n29292), .Y(exu_n8607));
AND2X1 exu_U26158(.A(alu_logic_result_and[10]), .B(exu_n16240), .Y(exu_n29294));
INVX1 exu_U26159(.A(exu_n29294), .Y(exu_n8608));
AND2X1 exu_U26160(.A(alu_logic_result_xor[0]), .B(exu_n16238), .Y(exu_n29298));
INVX1 exu_U26161(.A(exu_n29298), .Y(exu_n8609));
AND2X1 exu_U26162(.A(alu_logic_result_and[0]), .B(exu_n16240), .Y(exu_n29300));
INVX1 exu_U26163(.A(exu_n29300), .Y(exu_n8610));
AND2X1 exu_U26164(.A(exu_spu_rs3_data_e[9]), .B(exu_n16170), .Y(exu_n30402));
INVX1 exu_U26165(.A(exu_n30402), .Y(exu_n8611));
AND2X1 exu_U26166(.A(exu_spu_rs3_data_e[8]), .B(exu_n16168), .Y(exu_n30404));
INVX1 exu_U26167(.A(exu_n30404), .Y(exu_n8612));
AND2X1 exu_U26168(.A(exu_spu_rs3_data_e[7]), .B(exu_n16168), .Y(exu_n30406));
INVX1 exu_U26169(.A(exu_n30406), .Y(exu_n8613));
AND2X1 exu_U26170(.A(exu_spu_rs3_data_e[6]), .B(exu_n16169), .Y(exu_n30408));
INVX1 exu_U26171(.A(exu_n30408), .Y(exu_n8614));
AND2X1 exu_U26172(.A(exu_spu_rs3_data_e[5]), .B(exu_n16168), .Y(exu_n30414));
INVX1 exu_U26173(.A(exu_n30414), .Y(exu_n8615));
AND2X1 exu_U26174(.A(exu_spu_rs3_data_e[4]), .B(exu_n16168), .Y(exu_n30426));
INVX1 exu_U26175(.A(exu_n30426), .Y(exu_n8616));
AND2X1 exu_U26176(.A(exu_spu_rs3_data_e[3]), .B(exu_n16168), .Y(exu_n30438));
INVX1 exu_U26177(.A(exu_n30438), .Y(exu_n8617));
AND2X1 exu_U26178(.A(exu_spu_rs3_data_e[31]), .B(exu_n16170), .Y(exu_n30448));
INVX1 exu_U26179(.A(exu_n30448), .Y(exu_n8618));
AND2X1 exu_U26180(.A(exu_spu_rs3_data_e[30]), .B(exu_n16168), .Y(exu_n30450));
INVX1 exu_U26181(.A(exu_n30450), .Y(exu_n8619));
AND2X1 exu_U26182(.A(exu_spu_rs3_data_e[2]), .B(exu_n16167), .Y(exu_n30452));
INVX1 exu_U26183(.A(exu_n30452), .Y(exu_n8620));
AND2X1 exu_U26184(.A(exu_spu_rs3_data_e[29]), .B(exu_n16169), .Y(exu_n30454));
INVX1 exu_U26185(.A(exu_n30454), .Y(exu_n8621));
AND2X1 exu_U26186(.A(exu_spu_rs3_data_e[28]), .B(exu_n16167), .Y(exu_n30456));
INVX1 exu_U26187(.A(exu_n30456), .Y(exu_n8622));
AND2X1 exu_U26188(.A(exu_spu_rs3_data_e[27]), .B(exu_n16168), .Y(exu_n30458));
INVX1 exu_U26189(.A(exu_n30458), .Y(exu_n8623));
AND2X1 exu_U26190(.A(exu_spu_rs3_data_e[26]), .B(exu_n16168), .Y(exu_n30460));
INVX1 exu_U26191(.A(exu_n30460), .Y(exu_n8624));
AND2X1 exu_U26192(.A(exu_spu_rs3_data_e[25]), .B(exu_n16167), .Y(exu_n30462));
INVX1 exu_U26193(.A(exu_n30462), .Y(exu_n8625));
AND2X1 exu_U26194(.A(exu_spu_rs3_data_e[24]), .B(exu_n16170), .Y(exu_n30464));
INVX1 exu_U26195(.A(exu_n30464), .Y(exu_n8626));
AND2X1 exu_U26196(.A(exu_spu_rs3_data_e[23]), .B(exu_n16169), .Y(exu_n30466));
INVX1 exu_U26197(.A(exu_n30466), .Y(exu_n8627));
AND2X1 exu_U26198(.A(exu_spu_rs3_data_e[22]), .B(exu_n16170), .Y(exu_n30468));
INVX1 exu_U26199(.A(exu_n30468), .Y(exu_n8628));
AND2X1 exu_U26200(.A(exu_spu_rs3_data_e[21]), .B(exu_n16167), .Y(exu_n30470));
INVX1 exu_U26201(.A(exu_n30470), .Y(exu_n8629));
AND2X1 exu_U26202(.A(exu_spu_rs3_data_e[20]), .B(exu_n16169), .Y(exu_n30472));
INVX1 exu_U26203(.A(exu_n30472), .Y(exu_n8630));
AND2X1 exu_U26204(.A(exu_spu_rs3_data_e[1]), .B(exu_n16168), .Y(exu_n30474));
INVX1 exu_U26205(.A(exu_n30474), .Y(exu_n8631));
AND2X1 exu_U26206(.A(exu_spu_rs3_data_e[19]), .B(exu_n16168), .Y(exu_n30476));
INVX1 exu_U26207(.A(exu_n30476), .Y(exu_n8632));
AND2X1 exu_U26208(.A(exu_spu_rs3_data_e[18]), .B(exu_n16168), .Y(exu_n30478));
INVX1 exu_U26209(.A(exu_n30478), .Y(exu_n8633));
AND2X1 exu_U26210(.A(exu_spu_rs3_data_e[17]), .B(exu_n16168), .Y(exu_n30480));
INVX1 exu_U26211(.A(exu_n30480), .Y(exu_n8634));
AND2X1 exu_U26212(.A(exu_spu_rs3_data_e[16]), .B(exu_n16168), .Y(exu_n30482));
INVX1 exu_U26213(.A(exu_n30482), .Y(exu_n8635));
AND2X1 exu_U26214(.A(exu_spu_rs3_data_e[15]), .B(exu_n16168), .Y(exu_n30484));
INVX1 exu_U26215(.A(exu_n30484), .Y(exu_n8636));
AND2X1 exu_U26216(.A(exu_spu_rs3_data_e[14]), .B(exu_n16168), .Y(exu_n30486));
INVX1 exu_U26217(.A(exu_n30486), .Y(exu_n8637));
AND2X1 exu_U26218(.A(exu_spu_rs3_data_e[13]), .B(exu_n16168), .Y(exu_n30488));
INVX1 exu_U26219(.A(exu_n30488), .Y(exu_n8638));
AND2X1 exu_U26220(.A(exu_spu_rs3_data_e[12]), .B(exu_n16168), .Y(exu_n30490));
INVX1 exu_U26221(.A(exu_n30490), .Y(exu_n8639));
AND2X1 exu_U26222(.A(exu_spu_rs3_data_e[11]), .B(exu_n16168), .Y(exu_n30492));
INVX1 exu_U26223(.A(exu_n30492), .Y(exu_n8640));
AND2X1 exu_U26224(.A(exu_spu_rs3_data_e[10]), .B(exu_n16168), .Y(exu_n30494));
INVX1 exu_U26225(.A(exu_n30494), .Y(exu_n8641));
AND2X1 exu_U26226(.A(exu_spu_rs3_data_e[0]), .B(exu_n16168), .Y(exu_n30496));
INVX1 exu_U26227(.A(exu_n30496), .Y(exu_n8642));
AND2X1 exu_U26228(.A(alu_ecl_add_n64_e), .B(exu_n16262), .Y(exu_n30506));
INVX1 exu_U26229(.A(exu_n30506), .Y(exu_n8643));
AND2X1 exu_U26230(.A(alu_adder_out[62]), .B(exu_n16262), .Y(exu_n30508));
INVX1 exu_U26231(.A(exu_n30508), .Y(exu_n8644));
AND2X1 exu_U26232(.A(alu_adder_out[61]), .B(exu_n16262), .Y(exu_n30510));
INVX1 exu_U26233(.A(exu_n30510), .Y(exu_n8645));
AND2X1 exu_U26234(.A(alu_adder_out[60]), .B(exu_n16262), .Y(exu_n30512));
INVX1 exu_U26235(.A(exu_n30512), .Y(exu_n8646));
AND2X1 exu_U26236(.A(alu_adder_out[59]), .B(exu_n16262), .Y(exu_n30516));
INVX1 exu_U26237(.A(exu_n30516), .Y(exu_n8647));
AND2X1 exu_U26238(.A(alu_adder_out[58]), .B(exu_n16262), .Y(exu_n30518));
INVX1 exu_U26239(.A(exu_n30518), .Y(exu_n8648));
AND2X1 exu_U26240(.A(alu_adder_out[57]), .B(exu_n16262), .Y(exu_n30520));
INVX1 exu_U26241(.A(exu_n30520), .Y(exu_n8649));
AND2X1 exu_U26242(.A(alu_adder_out[56]), .B(exu_n16262), .Y(exu_n30522));
INVX1 exu_U26243(.A(exu_n30522), .Y(exu_n8650));
AND2X1 exu_U26244(.A(alu_adder_out[55]), .B(exu_n16262), .Y(exu_n30524));
INVX1 exu_U26245(.A(exu_n30524), .Y(exu_n8651));
AND2X1 exu_U26246(.A(alu_adder_out[54]), .B(exu_n16262), .Y(exu_n30526));
INVX1 exu_U26247(.A(exu_n30526), .Y(exu_n8652));
AND2X1 exu_U26248(.A(alu_adder_out[53]), .B(exu_n16262), .Y(exu_n30528));
INVX1 exu_U26249(.A(exu_n30528), .Y(exu_n8653));
AND2X1 exu_U26250(.A(alu_adder_out[52]), .B(exu_n16262), .Y(exu_n30530));
INVX1 exu_U26251(.A(exu_n30530), .Y(exu_n8654));
AND2X1 exu_U26252(.A(alu_adder_out[51]), .B(exu_n16262), .Y(exu_n30532));
INVX1 exu_U26253(.A(exu_n30532), .Y(exu_n8655));
AND2X1 exu_U26254(.A(alu_adder_out[50]), .B(exu_n16262), .Y(exu_n30534));
INVX1 exu_U26255(.A(exu_n30534), .Y(exu_n8656));
AND2X1 exu_U26256(.A(alu_adder_out[49]), .B(exu_n16262), .Y(exu_n30538));
INVX1 exu_U26257(.A(exu_n30538), .Y(exu_n8657));
AND2X1 exu_U26258(.A(alu_adder_out[48]), .B(exu_n16262), .Y(exu_n30540));
INVX1 exu_U26259(.A(exu_n30540), .Y(exu_n8658));
AND2X1 exu_U26260(.A(exu_ifu_brpc_e[47]), .B(exu_n16262), .Y(exu_n30542));
INVX1 exu_U26261(.A(exu_n30542), .Y(exu_n8659));
AND2X1 exu_U26262(.A(alu_logic_out_9), .B(exu_n16161), .Y(exu_n30626));
INVX1 exu_U26263(.A(exu_n30626), .Y(exu_n8660));
AND2X1 exu_U26264(.A(alu_logic_out_8), .B(exu_n16161), .Y(exu_n30628));
INVX1 exu_U26265(.A(exu_n30628), .Y(exu_n8661));
AND2X1 exu_U26266(.A(alu_logic_out_7), .B(exu_n16161), .Y(exu_n30630));
INVX1 exu_U26267(.A(exu_n30630), .Y(exu_n8662));
AND2X1 exu_U26268(.A(alu_logic_out_6), .B(exu_n16161), .Y(exu_n30632));
INVX1 exu_U26269(.A(exu_n30632), .Y(exu_n8663));
AND2X1 exu_U26270(.A(alu_ecl_log_n64_e), .B(exu_n16161), .Y(exu_n30634));
INVX1 exu_U26271(.A(exu_n30634), .Y(exu_n8664));
AND2X1 exu_U26272(.A(alu_logic_out[62]), .B(exu_n16161), .Y(exu_n30636));
INVX1 exu_U26273(.A(exu_n30636), .Y(exu_n8665));
AND2X1 exu_U26274(.A(alu_logic_out[61]), .B(exu_n16161), .Y(exu_n30638));
INVX1 exu_U26275(.A(exu_n30638), .Y(exu_n8666));
AND2X1 exu_U26276(.A(alu_logic_out[60]), .B(exu_n16161), .Y(exu_n30640));
INVX1 exu_U26277(.A(exu_n30640), .Y(exu_n8667));
AND2X1 exu_U26278(.A(alu_logic_out_5), .B(exu_n16161), .Y(exu_n30642));
INVX1 exu_U26279(.A(exu_n30642), .Y(exu_n8668));
AND2X1 exu_U26280(.A(alu_logic_out[59]), .B(exu_n16161), .Y(exu_n30644));
INVX1 exu_U26281(.A(exu_n30644), .Y(exu_n8669));
AND2X1 exu_U26282(.A(alu_logic_out[58]), .B(exu_n16156), .Y(exu_n30646));
INVX1 exu_U26283(.A(exu_n30646), .Y(exu_n8670));
AND2X1 exu_U26284(.A(alu_logic_out[57]), .B(exu_n16156), .Y(exu_n30648));
INVX1 exu_U26285(.A(exu_n30648), .Y(exu_n8671));
AND2X1 exu_U26286(.A(alu_logic_out[56]), .B(exu_n16156), .Y(exu_n30650));
INVX1 exu_U26287(.A(exu_n30650), .Y(exu_n8672));
AND2X1 exu_U26288(.A(alu_logic_out[55]), .B(exu_n16156), .Y(exu_n30652));
INVX1 exu_U26289(.A(exu_n30652), .Y(exu_n8673));
AND2X1 exu_U26290(.A(alu_logic_out[54]), .B(exu_n16156), .Y(exu_n30654));
INVX1 exu_U26291(.A(exu_n30654), .Y(exu_n8674));
AND2X1 exu_U26292(.A(alu_logic_out[53]), .B(exu_n16160), .Y(exu_n30656));
INVX1 exu_U26293(.A(exu_n30656), .Y(exu_n8675));
AND2X1 exu_U26294(.A(alu_logic_out[52]), .B(exu_n16156), .Y(exu_n30658));
INVX1 exu_U26295(.A(exu_n30658), .Y(exu_n8676));
AND2X1 exu_U26296(.A(alu_logic_out[51]), .B(exu_n16156), .Y(exu_n30660));
INVX1 exu_U26297(.A(exu_n30660), .Y(exu_n8677));
AND2X1 exu_U26298(.A(alu_logic_out[50]), .B(exu_n16161), .Y(exu_n30662));
INVX1 exu_U26299(.A(exu_n30662), .Y(exu_n8678));
AND2X1 exu_U26300(.A(alu_logic_out_4), .B(exu_n16159), .Y(exu_n30664));
INVX1 exu_U26301(.A(exu_n30664), .Y(exu_n8679));
AND2X1 exu_U26302(.A(alu_logic_out[49]), .B(exu_n16160), .Y(exu_n30666));
INVX1 exu_U26303(.A(exu_n30666), .Y(exu_n8680));
AND2X1 exu_U26304(.A(alu_logic_out[48]), .B(exu_n16160), .Y(exu_n30668));
INVX1 exu_U26305(.A(exu_n30668), .Y(exu_n8681));
AND2X1 exu_U26306(.A(alu_logic_out[47]), .B(exu_n16156), .Y(exu_n30670));
INVX1 exu_U26307(.A(exu_n30670), .Y(exu_n8682));
AND2X1 exu_U26308(.A(alu_logic_out[46]), .B(exu_n16159), .Y(exu_n30672));
INVX1 exu_U26309(.A(exu_n30672), .Y(exu_n8683));
AND2X1 exu_U26310(.A(alu_logic_out[45]), .B(exu_n16161), .Y(exu_n30674));
INVX1 exu_U26311(.A(exu_n30674), .Y(exu_n8684));
AND2X1 exu_U26312(.A(alu_logic_out[44]), .B(exu_n16156), .Y(exu_n30676));
INVX1 exu_U26313(.A(exu_n30676), .Y(exu_n8685));
AND2X1 exu_U26314(.A(alu_logic_out[43]), .B(exu_n16156), .Y(exu_n30678));
INVX1 exu_U26315(.A(exu_n30678), .Y(exu_n8686));
AND2X1 exu_U26316(.A(alu_logic_out[42]), .B(exu_n16159), .Y(exu_n30680));
INVX1 exu_U26317(.A(exu_n30680), .Y(exu_n8687));
AND2X1 exu_U26318(.A(alu_logic_out[41]), .B(exu_n16156), .Y(exu_n30682));
INVX1 exu_U26319(.A(exu_n30682), .Y(exu_n8688));
AND2X1 exu_U26320(.A(alu_logic_out[40]), .B(exu_n16161), .Y(exu_n30684));
INVX1 exu_U26321(.A(exu_n30684), .Y(exu_n8689));
AND2X1 exu_U26322(.A(alu_logic_out_3), .B(exu_n16159), .Y(exu_n30686));
INVX1 exu_U26323(.A(exu_n30686), .Y(exu_n8690));
AND2X1 exu_U26324(.A(alu_logic_out[39]), .B(exu_n16156), .Y(exu_n30688));
INVX1 exu_U26325(.A(exu_n30688), .Y(exu_n8691));
AND2X1 exu_U26326(.A(alu_logic_out[38]), .B(exu_n16161), .Y(exu_n30690));
INVX1 exu_U26327(.A(exu_n30690), .Y(exu_n8692));
AND2X1 exu_U26328(.A(alu_logic_out[37]), .B(exu_n16159), .Y(exu_n30692));
INVX1 exu_U26329(.A(exu_n30692), .Y(exu_n8693));
AND2X1 exu_U26330(.A(alu_logic_out[36]), .B(exu_n16156), .Y(exu_n30694));
INVX1 exu_U26331(.A(exu_n30694), .Y(exu_n8694));
AND2X1 exu_U26332(.A(alu_logic_out[35]), .B(exu_n16161), .Y(exu_n30696));
INVX1 exu_U26333(.A(exu_n30696), .Y(exu_n8695));
AND2X1 exu_U26334(.A(alu_logic_out[34]), .B(exu_n16159), .Y(exu_n30698));
INVX1 exu_U26335(.A(exu_n30698), .Y(exu_n8696));
AND2X1 exu_U26336(.A(alu_logic_out[33]), .B(exu_n16156), .Y(exu_n30700));
INVX1 exu_U26337(.A(exu_n30700), .Y(exu_n8697));
AND2X1 exu_U26338(.A(alu_logic_out[32]), .B(exu_n16161), .Y(exu_n30702));
INVX1 exu_U26339(.A(exu_n30702), .Y(exu_n8698));
AND2X1 exu_U26340(.A(alu_ecl_log_n32_e), .B(exu_n16159), .Y(exu_n30704));
INVX1 exu_U26341(.A(exu_n30704), .Y(exu_n8699));
AND2X1 exu_U26342(.A(alu_logic_out_30), .B(exu_n16159), .Y(exu_n30706));
INVX1 exu_U26343(.A(exu_n30706), .Y(exu_n8700));
AND2X1 exu_U26344(.A(alu_logic_out_2), .B(exu_n16160), .Y(exu_n30708));
INVX1 exu_U26345(.A(exu_n30708), .Y(exu_n8701));
AND2X1 exu_U26346(.A(alu_logic_out_29), .B(exu_n16161), .Y(exu_n30710));
INVX1 exu_U26347(.A(exu_n30710), .Y(exu_n8702));
AND2X1 exu_U26348(.A(alu_logic_out_28), .B(exu_n16156), .Y(exu_n30712));
INVX1 exu_U26349(.A(exu_n30712), .Y(exu_n8703));
AND2X1 exu_U26350(.A(alu_logic_out_27), .B(exu_n16159), .Y(exu_n30714));
INVX1 exu_U26351(.A(exu_n30714), .Y(exu_n8704));
AND2X1 exu_U26352(.A(alu_logic_out_26), .B(exu_n16159), .Y(exu_n30716));
INVX1 exu_U26353(.A(exu_n30716), .Y(exu_n8705));
AND2X1 exu_U26354(.A(alu_logic_out_25), .B(exu_n16160), .Y(exu_n30718));
INVX1 exu_U26355(.A(exu_n30718), .Y(exu_n8706));
AND2X1 exu_U26356(.A(alu_logic_out_24), .B(exu_n16161), .Y(exu_n30720));
INVX1 exu_U26357(.A(exu_n30720), .Y(exu_n8707));
AND2X1 exu_U26358(.A(alu_logic_out_23), .B(exu_n16156), .Y(exu_n30722));
INVX1 exu_U26359(.A(exu_n30722), .Y(exu_n8708));
AND2X1 exu_U26360(.A(alu_logic_out_22), .B(exu_n16159), .Y(exu_n30724));
INVX1 exu_U26361(.A(exu_n30724), .Y(exu_n8709));
AND2X1 exu_U26362(.A(alu_logic_out_21), .B(exu_n16159), .Y(exu_n30726));
INVX1 exu_U26363(.A(exu_n30726), .Y(exu_n8710));
AND2X1 exu_U26364(.A(alu_logic_out_20), .B(exu_n16160), .Y(exu_n30728));
INVX1 exu_U26365(.A(exu_n30728), .Y(exu_n8711));
AND2X1 exu_U26366(.A(alu_logic_out_1), .B(exu_n16161), .Y(exu_n30730));
INVX1 exu_U26367(.A(exu_n30730), .Y(exu_n8712));
AND2X1 exu_U26368(.A(alu_logic_out_19), .B(exu_n16156), .Y(exu_n30732));
INVX1 exu_U26369(.A(exu_n30732), .Y(exu_n8713));
AND2X1 exu_U26370(.A(alu_logic_out_18), .B(exu_n16159), .Y(exu_n30734));
INVX1 exu_U26371(.A(exu_n30734), .Y(exu_n8714));
AND2X1 exu_U26372(.A(alu_logic_out_17), .B(exu_n16156), .Y(exu_n30736));
INVX1 exu_U26373(.A(exu_n30736), .Y(exu_n8715));
AND2X1 exu_U26374(.A(alu_logic_out_16), .B(exu_n16160), .Y(exu_n30738));
INVX1 exu_U26375(.A(exu_n30738), .Y(exu_n8716));
AND2X1 exu_U26376(.A(alu_logic_out_15), .B(exu_n16159), .Y(exu_n30740));
INVX1 exu_U26377(.A(exu_n30740), .Y(exu_n8717));
AND2X1 exu_U26378(.A(alu_logic_out_14), .B(exu_n16156), .Y(exu_n30742));
INVX1 exu_U26379(.A(exu_n30742), .Y(exu_n8718));
AND2X1 exu_U26380(.A(alu_logic_out_13), .B(exu_n16160), .Y(exu_n30744));
INVX1 exu_U26381(.A(exu_n30744), .Y(exu_n8719));
AND2X1 exu_U26382(.A(alu_logic_out_12), .B(exu_n16161), .Y(exu_n30746));
INVX1 exu_U26383(.A(exu_n30746), .Y(exu_n8720));
AND2X1 exu_U26384(.A(alu_logic_out_11), .B(exu_n16159), .Y(exu_n30748));
INVX1 exu_U26385(.A(exu_n30748), .Y(exu_n8721));
AND2X1 exu_U26386(.A(alu_logic_out_10), .B(exu_n16161), .Y(exu_n30750));
INVX1 exu_U26387(.A(exu_n30750), .Y(exu_n8722));
AND2X1 exu_U26388(.A(alu_logic_out_0), .B(exu_n16156), .Y(exu_n30752));
INVX1 exu_U26389(.A(exu_n30752), .Y(exu_n8723));
AND2X1 exu_U26390(.A(shft_lshift1[8]), .B(exu_n16236), .Y(exu_n30756));
INVX1 exu_U26391(.A(exu_n30756), .Y(exu_n8724));
AND2X1 exu_U26392(.A(shft_lshift1[7]), .B(exu_n16236), .Y(exu_n30758));
INVX1 exu_U26393(.A(exu_n30758), .Y(exu_n8725));
AND2X1 exu_U26394(.A(shft_lshift1[6]), .B(exu_n16236), .Y(exu_n30760));
INVX1 exu_U26395(.A(exu_n30760), .Y(exu_n8726));
AND2X1 exu_U26396(.A(shft_lshift1[63]), .B(exu_n16236), .Y(exu_n30762));
INVX1 exu_U26397(.A(exu_n30762), .Y(exu_n8727));
AND2X1 exu_U26398(.A(shft_lshift1[62]), .B(exu_n16236), .Y(exu_n30764));
INVX1 exu_U26399(.A(exu_n30764), .Y(exu_n8728));
AND2X1 exu_U26400(.A(shft_lshift1[61]), .B(exu_n16236), .Y(exu_n30766));
INVX1 exu_U26401(.A(exu_n30766), .Y(exu_n8729));
AND2X1 exu_U26402(.A(shft_lshift1[60]), .B(exu_n16236), .Y(exu_n30768));
INVX1 exu_U26403(.A(exu_n30768), .Y(exu_n8730));
AND2X1 exu_U26404(.A(shft_lshift1[5]), .B(exu_n16236), .Y(exu_n30770));
INVX1 exu_U26405(.A(exu_n30770), .Y(exu_n8731));
AND2X1 exu_U26406(.A(shft_lshift1[59]), .B(exu_n16236), .Y(exu_n30772));
INVX1 exu_U26407(.A(exu_n30772), .Y(exu_n8732));
AND2X1 exu_U26408(.A(shft_lshift1[58]), .B(exu_n16236), .Y(exu_n30774));
INVX1 exu_U26409(.A(exu_n30774), .Y(exu_n8733));
AND2X1 exu_U26410(.A(shft_lshift1[57]), .B(exu_n16236), .Y(exu_n30776));
INVX1 exu_U26411(.A(exu_n30776), .Y(exu_n8734));
AND2X1 exu_U26412(.A(shft_lshift1[56]), .B(exu_n16236), .Y(exu_n30778));
INVX1 exu_U26413(.A(exu_n30778), .Y(exu_n8735));
AND2X1 exu_U26414(.A(shft_lshift1[55]), .B(exu_n16236), .Y(exu_n30780));
INVX1 exu_U26415(.A(exu_n30780), .Y(exu_n8736));
AND2X1 exu_U26416(.A(shft_lshift1[54]), .B(exu_n16236), .Y(exu_n30782));
INVX1 exu_U26417(.A(exu_n30782), .Y(exu_n8737));
AND2X1 exu_U26418(.A(shft_lshift1[53]), .B(exu_n16236), .Y(exu_n30784));
INVX1 exu_U26419(.A(exu_n30784), .Y(exu_n8738));
AND2X1 exu_U26420(.A(shft_lshift1[52]), .B(exu_n16236), .Y(exu_n30786));
INVX1 exu_U26421(.A(exu_n30786), .Y(exu_n8739));
AND2X1 exu_U26422(.A(shft_lshift1[51]), .B(exu_n16236), .Y(exu_n30788));
INVX1 exu_U26423(.A(exu_n30788), .Y(exu_n8740));
AND2X1 exu_U26424(.A(shft_lshift1[50]), .B(exu_n16236), .Y(exu_n30790));
INVX1 exu_U26425(.A(exu_n30790), .Y(exu_n8741));
AND2X1 exu_U26426(.A(shft_lshift1[4]), .B(exu_n16236), .Y(exu_n30792));
INVX1 exu_U26427(.A(exu_n30792), .Y(exu_n8742));
AND2X1 exu_U26428(.A(shft_lshift1[49]), .B(exu_n16236), .Y(exu_n30794));
INVX1 exu_U26429(.A(exu_n30794), .Y(exu_n8743));
AND2X1 exu_U26430(.A(shft_lshift1[48]), .B(exu_n16236), .Y(exu_n30796));
INVX1 exu_U26431(.A(exu_n30796), .Y(exu_n8744));
AND2X1 exu_U26432(.A(shft_lshift1[47]), .B(exu_n16236), .Y(exu_n30798));
INVX1 exu_U26433(.A(exu_n30798), .Y(exu_n8745));
AND2X1 exu_U26434(.A(shft_lshift1[46]), .B(exu_n16236), .Y(exu_n30800));
INVX1 exu_U26435(.A(exu_n30800), .Y(exu_n8746));
AND2X1 exu_U26436(.A(shft_lshift1[45]), .B(exu_n16236), .Y(exu_n30802));
INVX1 exu_U26437(.A(exu_n30802), .Y(exu_n8747));
AND2X1 exu_U26438(.A(shft_lshift1[44]), .B(exu_n16236), .Y(exu_n30804));
INVX1 exu_U26439(.A(exu_n30804), .Y(exu_n8748));
AND2X1 exu_U26440(.A(shft_lshift1[43]), .B(exu_n16236), .Y(exu_n30806));
INVX1 exu_U26441(.A(exu_n30806), .Y(exu_n8749));
AND2X1 exu_U26442(.A(shft_lshift1[42]), .B(exu_n16236), .Y(exu_n30808));
INVX1 exu_U26443(.A(exu_n30808), .Y(exu_n8750));
AND2X1 exu_U26444(.A(shft_lshift1[41]), .B(exu_n16236), .Y(exu_n30810));
INVX1 exu_U26445(.A(exu_n30810), .Y(exu_n8751));
AND2X1 exu_U26446(.A(shft_lshift1[40]), .B(exu_n16236), .Y(exu_n30812));
INVX1 exu_U26447(.A(exu_n30812), .Y(exu_n8752));
AND2X1 exu_U26448(.A(shft_lshift1[3]), .B(exu_n16236), .Y(exu_n30814));
INVX1 exu_U26449(.A(exu_n30814), .Y(exu_n8753));
AND2X1 exu_U26450(.A(shft_lshift1[39]), .B(exu_n16236), .Y(exu_n30816));
INVX1 exu_U26451(.A(exu_n30816), .Y(exu_n8754));
AND2X1 exu_U26452(.A(shft_lshift1[38]), .B(exu_n16236), .Y(exu_n30818));
INVX1 exu_U26453(.A(exu_n30818), .Y(exu_n8755));
AND2X1 exu_U26454(.A(shft_lshift1[37]), .B(exu_n16236), .Y(exu_n30820));
INVX1 exu_U26455(.A(exu_n30820), .Y(exu_n8756));
AND2X1 exu_U26456(.A(shft_lshift1[36]), .B(exu_n16236), .Y(exu_n30822));
INVX1 exu_U26457(.A(exu_n30822), .Y(exu_n8757));
AND2X1 exu_U26458(.A(shft_lshift1[35]), .B(exu_n16236), .Y(exu_n30824));
INVX1 exu_U26459(.A(exu_n30824), .Y(exu_n8758));
AND2X1 exu_U26460(.A(shft_lshift1[34]), .B(exu_n16236), .Y(exu_n30826));
INVX1 exu_U26461(.A(exu_n30826), .Y(exu_n8759));
AND2X1 exu_U26462(.A(shft_lshift1[33]), .B(exu_n16236), .Y(exu_n30828));
INVX1 exu_U26463(.A(exu_n30828), .Y(exu_n8760));
AND2X1 exu_U26464(.A(shft_lshift1[32]), .B(exu_n16236), .Y(exu_n30830));
INVX1 exu_U26465(.A(exu_n30830), .Y(exu_n8761));
AND2X1 exu_U26466(.A(shft_lshift1[31]), .B(exu_n16236), .Y(exu_n30832));
INVX1 exu_U26467(.A(exu_n30832), .Y(exu_n8762));
AND2X1 exu_U26468(.A(shft_lshift1[30]), .B(exu_n16236), .Y(exu_n30834));
INVX1 exu_U26469(.A(exu_n30834), .Y(exu_n8763));
AND2X1 exu_U26470(.A(shft_lshift1[2]), .B(exu_n16236), .Y(exu_n30836));
INVX1 exu_U26471(.A(exu_n30836), .Y(exu_n8764));
AND2X1 exu_U26472(.A(shft_lshift1[29]), .B(exu_n16236), .Y(exu_n30838));
INVX1 exu_U26473(.A(exu_n30838), .Y(exu_n8765));
AND2X1 exu_U26474(.A(shft_lshift1[28]), .B(exu_n16236), .Y(exu_n30840));
INVX1 exu_U26475(.A(exu_n30840), .Y(exu_n8766));
AND2X1 exu_U26476(.A(shft_lshift1[27]), .B(exu_n16236), .Y(exu_n30842));
INVX1 exu_U26477(.A(exu_n30842), .Y(exu_n8767));
AND2X1 exu_U26478(.A(shft_lshift1[26]), .B(exu_n16236), .Y(exu_n30844));
INVX1 exu_U26479(.A(exu_n30844), .Y(exu_n8768));
AND2X1 exu_U26480(.A(shft_lshift1[25]), .B(exu_n16236), .Y(exu_n30846));
INVX1 exu_U26481(.A(exu_n30846), .Y(exu_n8769));
AND2X1 exu_U26482(.A(shft_lshift1[24]), .B(exu_n16236), .Y(exu_n30848));
INVX1 exu_U26483(.A(exu_n30848), .Y(exu_n8770));
AND2X1 exu_U26484(.A(shft_lshift1[23]), .B(exu_n16236), .Y(exu_n30850));
INVX1 exu_U26485(.A(exu_n30850), .Y(exu_n8771));
AND2X1 exu_U26486(.A(shft_lshift1[22]), .B(exu_n16236), .Y(exu_n30852));
INVX1 exu_U26487(.A(exu_n30852), .Y(exu_n8772));
AND2X1 exu_U26488(.A(shft_lshift1[21]), .B(exu_n16236), .Y(exu_n30854));
INVX1 exu_U26489(.A(exu_n30854), .Y(exu_n8773));
AND2X1 exu_U26490(.A(shft_lshift1[20]), .B(exu_n16236), .Y(exu_n30856));
INVX1 exu_U26491(.A(exu_n30856), .Y(exu_n8774));
AND2X1 exu_U26492(.A(exu_n11057), .B(exu_n16236), .Y(exu_n30858));
INVX1 exu_U26493(.A(exu_n30858), .Y(exu_n8775));
AND2X1 exu_U26494(.A(shft_lshift1[19]), .B(exu_n16236), .Y(exu_n30860));
INVX1 exu_U26495(.A(exu_n30860), .Y(exu_n8776));
AND2X1 exu_U26496(.A(shft_lshift1[18]), .B(exu_n16236), .Y(exu_n30862));
INVX1 exu_U26497(.A(exu_n30862), .Y(exu_n8777));
AND2X1 exu_U26498(.A(shft_lshift1[17]), .B(exu_n16236), .Y(exu_n30864));
INVX1 exu_U26499(.A(exu_n30864), .Y(exu_n8778));
AND2X1 exu_U26500(.A(shft_lshift1[16]), .B(exu_n16236), .Y(exu_n30866));
INVX1 exu_U26501(.A(exu_n30866), .Y(exu_n8779));
AND2X1 exu_U26502(.A(shft_lshift1[15]), .B(exu_n16236), .Y(exu_n30868));
INVX1 exu_U26503(.A(exu_n30868), .Y(exu_n8780));
AND2X1 exu_U26504(.A(shft_lshift1[14]), .B(exu_n16236), .Y(exu_n30870));
INVX1 exu_U26505(.A(exu_n30870), .Y(exu_n8781));
AND2X1 exu_U26506(.A(shft_lshift1[13]), .B(exu_n16236), .Y(exu_n30872));
INVX1 exu_U26507(.A(exu_n30872), .Y(exu_n8782));
AND2X1 exu_U26508(.A(shft_lshift1[12]), .B(exu_n16236), .Y(exu_n30874));
INVX1 exu_U26509(.A(exu_n30874), .Y(exu_n8783));
AND2X1 exu_U26510(.A(shft_lshift1[11]), .B(exu_n16236), .Y(exu_n30876));
INVX1 exu_U26511(.A(exu_n30876), .Y(exu_n8784));
AND2X1 exu_U26512(.A(shft_lshift1[10]), .B(exu_n16236), .Y(exu_n30878));
INVX1 exu_U26513(.A(exu_n30878), .Y(exu_n8785));
AND2X1 exu_U26514(.A(exu_n28695), .B(exu_n16236), .Y(exu_n30880));
INVX1 exu_U26515(.A(exu_n30880), .Y(exu_n8786));
AND2X1 exu_U26516(.A(div_mul_result[8]), .B(exu_n16196), .Y(exu_n30948));
INVX1 exu_U26517(.A(exu_n30948), .Y(exu_n8787));
AND2X1 exu_U26518(.A(div_mul_result[7]), .B(exu_n16196), .Y(exu_n30950));
INVX1 exu_U26519(.A(exu_n30950), .Y(exu_n8788));
AND2X1 exu_U26520(.A(div_mul_result[6]), .B(exu_n16196), .Y(exu_n30952));
INVX1 exu_U26521(.A(exu_n30952), .Y(exu_n8789));
AND2X1 exu_U26522(.A(div_mul_result[63]), .B(exu_n16198), .Y(exu_n30954));
INVX1 exu_U26523(.A(exu_n30954), .Y(exu_n8790));
AND2X1 exu_U26524(.A(div_mul_result[62]), .B(exu_n16196), .Y(exu_n30956));
INVX1 exu_U26525(.A(exu_n30956), .Y(exu_n8791));
AND2X1 exu_U26526(.A(div_mul_result[61]), .B(exu_n16196), .Y(exu_n30958));
INVX1 exu_U26527(.A(exu_n30958), .Y(exu_n8792));
AND2X1 exu_U26528(.A(div_mul_result[60]), .B(exu_n16199), .Y(exu_n30960));
INVX1 exu_U26529(.A(exu_n30960), .Y(exu_n8793));
AND2X1 exu_U26530(.A(div_mul_result[5]), .B(exu_n16196), .Y(exu_n30962));
INVX1 exu_U26531(.A(exu_n30962), .Y(exu_n8794));
AND2X1 exu_U26532(.A(div_mul_result[59]), .B(exu_n16198), .Y(exu_n30964));
INVX1 exu_U26533(.A(exu_n30964), .Y(exu_n8795));
AND2X1 exu_U26534(.A(div_mul_result[58]), .B(exu_n16196), .Y(exu_n30966));
INVX1 exu_U26535(.A(exu_n30966), .Y(exu_n8796));
AND2X1 exu_U26536(.A(div_mul_result[57]), .B(exu_n16196), .Y(exu_n30968));
INVX1 exu_U26537(.A(exu_n30968), .Y(exu_n8797));
AND2X1 exu_U26538(.A(div_mul_result[56]), .B(exu_n16199), .Y(exu_n30970));
INVX1 exu_U26539(.A(exu_n30970), .Y(exu_n8798));
AND2X1 exu_U26540(.A(div_mul_result[55]), .B(exu_n16196), .Y(exu_n30972));
INVX1 exu_U26541(.A(exu_n30972), .Y(exu_n8799));
AND2X1 exu_U26542(.A(div_mul_result[54]), .B(exu_n16198), .Y(exu_n30974));
INVX1 exu_U26543(.A(exu_n30974), .Y(exu_n8800));
AND2X1 exu_U26544(.A(div_mul_result[53]), .B(exu_n16202), .Y(exu_n30976));
INVX1 exu_U26545(.A(exu_n30976), .Y(exu_n8801));
AND2X1 exu_U26546(.A(div_mul_result[52]), .B(exu_n16202), .Y(exu_n30978));
INVX1 exu_U26547(.A(exu_n30978), .Y(exu_n8802));
AND2X1 exu_U26548(.A(div_mul_result[51]), .B(exu_n16202), .Y(exu_n30980));
INVX1 exu_U26549(.A(exu_n30980), .Y(exu_n8803));
AND2X1 exu_U26550(.A(div_mul_result[50]), .B(exu_n16202), .Y(exu_n30982));
INVX1 exu_U26551(.A(exu_n30982), .Y(exu_n8804));
AND2X1 exu_U26552(.A(div_mul_result[4]), .B(exu_n16202), .Y(exu_n30984));
INVX1 exu_U26553(.A(exu_n30984), .Y(exu_n8805));
AND2X1 exu_U26554(.A(div_mul_result[49]), .B(exu_n16202), .Y(exu_n30986));
INVX1 exu_U26555(.A(exu_n30986), .Y(exu_n8806));
AND2X1 exu_U26556(.A(div_mul_result[48]), .B(exu_n16202), .Y(exu_n30988));
INVX1 exu_U26557(.A(exu_n30988), .Y(exu_n8807));
AND2X1 exu_U26558(.A(div_mul_result[47]), .B(exu_n16202), .Y(exu_n30990));
INVX1 exu_U26559(.A(exu_n30990), .Y(exu_n8808));
AND2X1 exu_U26560(.A(div_mul_result[46]), .B(exu_n16202), .Y(exu_n30992));
INVX1 exu_U26561(.A(exu_n30992), .Y(exu_n8809));
AND2X1 exu_U26562(.A(div_mul_result[45]), .B(exu_n16202), .Y(exu_n30994));
INVX1 exu_U26563(.A(exu_n30994), .Y(exu_n8810));
AND2X1 exu_U26564(.A(div_mul_result[44]), .B(exu_n16202), .Y(exu_n30996));
INVX1 exu_U26565(.A(exu_n30996), .Y(exu_n8811));
AND2X1 exu_U26566(.A(div_mul_result[43]), .B(exu_n16202), .Y(exu_n30998));
INVX1 exu_U26567(.A(exu_n30998), .Y(exu_n8812));
AND2X1 exu_U26568(.A(div_mul_result[42]), .B(exu_n16202), .Y(exu_n31000));
INVX1 exu_U26569(.A(exu_n31000), .Y(exu_n8813));
AND2X1 exu_U26570(.A(div_mul_result[41]), .B(exu_n16202), .Y(exu_n31002));
INVX1 exu_U26571(.A(exu_n31002), .Y(exu_n8814));
AND2X1 exu_U26572(.A(div_mul_result[40]), .B(exu_n16202), .Y(exu_n31004));
INVX1 exu_U26573(.A(exu_n31004), .Y(exu_n8815));
AND2X1 exu_U26574(.A(div_mul_result[3]), .B(exu_n16201), .Y(exu_n31006));
INVX1 exu_U26575(.A(exu_n31006), .Y(exu_n8816));
AND2X1 exu_U26576(.A(div_mul_result[39]), .B(exu_n16201), .Y(exu_n31008));
INVX1 exu_U26577(.A(exu_n31008), .Y(exu_n8817));
AND2X1 exu_U26578(.A(div_mul_result[38]), .B(exu_n16201), .Y(exu_n31010));
INVX1 exu_U26579(.A(exu_n31010), .Y(exu_n8818));
AND2X1 exu_U26580(.A(div_mul_result[37]), .B(exu_n16201), .Y(exu_n31012));
INVX1 exu_U26581(.A(exu_n31012), .Y(exu_n8819));
AND2X1 exu_U26582(.A(div_mul_result[36]), .B(exu_n16201), .Y(exu_n31014));
INVX1 exu_U26583(.A(exu_n31014), .Y(exu_n8820));
AND2X1 exu_U26584(.A(div_mul_result[35]), .B(exu_n16201), .Y(exu_n31016));
INVX1 exu_U26585(.A(exu_n31016), .Y(exu_n8821));
AND2X1 exu_U26586(.A(div_mul_result[34]), .B(exu_n16201), .Y(exu_n31018));
INVX1 exu_U26587(.A(exu_n31018), .Y(exu_n8822));
AND2X1 exu_U26588(.A(div_mul_result[33]), .B(exu_n16201), .Y(exu_n31020));
INVX1 exu_U26589(.A(exu_n31020), .Y(exu_n8823));
AND2X1 exu_U26590(.A(div_mul_result[32]), .B(exu_n16201), .Y(exu_n31022));
INVX1 exu_U26591(.A(exu_n31022), .Y(exu_n8824));
AND2X1 exu_U26592(.A(div_mul_result[31]), .B(exu_n16201), .Y(exu_n31024));
INVX1 exu_U26593(.A(exu_n31024), .Y(exu_n8825));
AND2X1 exu_U26594(.A(div_mul_result[30]), .B(exu_n16201), .Y(exu_n31026));
INVX1 exu_U26595(.A(exu_n31026), .Y(exu_n8826));
AND2X1 exu_U26596(.A(div_mul_result[2]), .B(exu_n16201), .Y(exu_n31028));
INVX1 exu_U26597(.A(exu_n31028), .Y(exu_n8827));
AND2X1 exu_U26598(.A(div_mul_result[29]), .B(exu_n16201), .Y(exu_n31030));
INVX1 exu_U26599(.A(exu_n31030), .Y(exu_n8828));
AND2X1 exu_U26600(.A(div_mul_result[28]), .B(exu_n16201), .Y(exu_n31032));
INVX1 exu_U26601(.A(exu_n31032), .Y(exu_n8829));
AND2X1 exu_U26602(.A(div_mul_result[27]), .B(exu_n16201), .Y(exu_n31034));
INVX1 exu_U26603(.A(exu_n31034), .Y(exu_n8830));
AND2X1 exu_U26604(.A(div_mul_result[26]), .B(exu_n16200), .Y(exu_n31036));
INVX1 exu_U26605(.A(exu_n31036), .Y(exu_n8831));
AND2X1 exu_U26606(.A(div_mul_result[25]), .B(exu_n16200), .Y(exu_n31038));
INVX1 exu_U26607(.A(exu_n31038), .Y(exu_n8832));
AND2X1 exu_U26608(.A(div_mul_result[24]), .B(exu_n16200), .Y(exu_n31040));
INVX1 exu_U26609(.A(exu_n31040), .Y(exu_n8833));
AND2X1 exu_U26610(.A(div_mul_result[23]), .B(exu_n16200), .Y(exu_n31042));
INVX1 exu_U26611(.A(exu_n31042), .Y(exu_n8834));
AND2X1 exu_U26612(.A(div_mul_result[22]), .B(exu_n16200), .Y(exu_n31044));
INVX1 exu_U26613(.A(exu_n31044), .Y(exu_n8835));
AND2X1 exu_U26614(.A(div_mul_result[21]), .B(exu_n16200), .Y(exu_n31046));
INVX1 exu_U26615(.A(exu_n31046), .Y(exu_n8836));
AND2X1 exu_U26616(.A(div_mul_result[20]), .B(exu_n16200), .Y(exu_n31048));
INVX1 exu_U26617(.A(exu_n31048), .Y(exu_n8837));
AND2X1 exu_U26618(.A(div_mul_result[1]), .B(exu_n16200), .Y(exu_n31050));
INVX1 exu_U26619(.A(exu_n31050), .Y(exu_n8838));
AND2X1 exu_U26620(.A(div_mul_result[19]), .B(exu_n16200), .Y(exu_n31052));
INVX1 exu_U26621(.A(exu_n31052), .Y(exu_n8839));
AND2X1 exu_U26622(.A(div_mul_result[18]), .B(exu_n16200), .Y(exu_n31054));
INVX1 exu_U26623(.A(exu_n31054), .Y(exu_n8840));
AND2X1 exu_U26624(.A(div_mul_result[17]), .B(exu_n16200), .Y(exu_n31056));
INVX1 exu_U26625(.A(exu_n31056), .Y(exu_n8841));
AND2X1 exu_U26626(.A(div_mul_result[16]), .B(exu_n16200), .Y(exu_n31058));
INVX1 exu_U26627(.A(exu_n31058), .Y(exu_n8842));
AND2X1 exu_U26628(.A(div_mul_result[15]), .B(exu_n16200), .Y(exu_n31060));
INVX1 exu_U26629(.A(exu_n31060), .Y(exu_n8843));
AND2X1 exu_U26630(.A(div_mul_result[14]), .B(exu_n16200), .Y(exu_n31062));
INVX1 exu_U26631(.A(exu_n31062), .Y(exu_n8844));
AND2X1 exu_U26632(.A(div_mul_result[13]), .B(exu_n16200), .Y(exu_n31064));
INVX1 exu_U26633(.A(exu_n31064), .Y(exu_n8845));
AND2X1 exu_U26634(.A(div_mul_result[12]), .B(exu_n16199), .Y(exu_n31066));
INVX1 exu_U26635(.A(exu_n31066), .Y(exu_n8846));
AND2X1 exu_U26636(.A(div_mul_result[11]), .B(exu_n16199), .Y(exu_n31068));
INVX1 exu_U26637(.A(exu_n31068), .Y(exu_n8847));
AND2X1 exu_U26638(.A(div_mul_result[10]), .B(exu_n16199), .Y(exu_n31070));
INVX1 exu_U26639(.A(exu_n31070), .Y(exu_n8848));
AND2X1 exu_U26640(.A(div_mul_result[0]), .B(exu_n16199), .Y(exu_n31072));
INVX1 exu_U26641(.A(exu_n31072), .Y(exu_n8849));
AND2X1 exu_U26642(.A(div_curr_q[8]), .B(exu_n16257), .Y(exu_n31074));
INVX1 exu_U26643(.A(exu_n31074), .Y(exu_n8850));
AND2X1 exu_U26644(.A(div_curr_q[7]), .B(exu_n16257), .Y(exu_n31076));
INVX1 exu_U26645(.A(exu_n31076), .Y(exu_n8851));
AND2X1 exu_U26646(.A(div_curr_q[6]), .B(exu_n16257), .Y(exu_n31078));
INVX1 exu_U26647(.A(exu_n31078), .Y(exu_n8852));
AND2X1 exu_U26648(.A(div_curr_q[5]), .B(exu_n16257), .Y(exu_n31080));
INVX1 exu_U26649(.A(exu_n31080), .Y(exu_n8853));
AND2X1 exu_U26650(.A(div_curr_q[62]), .B(exu_n16257), .Y(exu_n31082));
INVX1 exu_U26651(.A(exu_n31082), .Y(exu_n8854));
AND2X1 exu_U26652(.A(div_curr_q[61]), .B(exu_n16257), .Y(exu_n31084));
INVX1 exu_U26653(.A(exu_n31084), .Y(exu_n8855));
AND2X1 exu_U26654(.A(div_curr_q[60]), .B(exu_n16257), .Y(exu_n31086));
INVX1 exu_U26655(.A(exu_n31086), .Y(exu_n8856));
AND2X1 exu_U26656(.A(div_curr_q[59]), .B(exu_n16257), .Y(exu_n31088));
INVX1 exu_U26657(.A(exu_n31088), .Y(exu_n8857));
AND2X1 exu_U26658(.A(div_curr_q[4]), .B(exu_n16257), .Y(exu_n31090));
INVX1 exu_U26659(.A(exu_n31090), .Y(exu_n8858));
AND2X1 exu_U26660(.A(div_curr_q[58]), .B(exu_n16257), .Y(exu_n31092));
INVX1 exu_U26661(.A(exu_n31092), .Y(exu_n8859));
AND2X1 exu_U26662(.A(div_curr_q[57]), .B(exu_n16257), .Y(exu_n31094));
INVX1 exu_U26663(.A(exu_n31094), .Y(exu_n8860));
AND2X1 exu_U26664(.A(div_curr_q[56]), .B(exu_n16257), .Y(exu_n31096));
INVX1 exu_U26665(.A(exu_n31096), .Y(exu_n8861));
AND2X1 exu_U26666(.A(div_curr_q[55]), .B(exu_n16257), .Y(exu_n31098));
INVX1 exu_U26667(.A(exu_n31098), .Y(exu_n8862));
AND2X1 exu_U26668(.A(div_curr_q[54]), .B(exu_n16257), .Y(exu_n31100));
INVX1 exu_U26669(.A(exu_n31100), .Y(exu_n8863));
AND2X1 exu_U26670(.A(div_curr_q[53]), .B(exu_n16257), .Y(exu_n31102));
INVX1 exu_U26671(.A(exu_n31102), .Y(exu_n8864));
AND2X1 exu_U26672(.A(div_curr_q[52]), .B(exu_n16257), .Y(exu_n31104));
INVX1 exu_U26673(.A(exu_n31104), .Y(exu_n8865));
AND2X1 exu_U26674(.A(div_curr_q[51]), .B(exu_n16257), .Y(exu_n31106));
INVX1 exu_U26675(.A(exu_n31106), .Y(exu_n8866));
AND2X1 exu_U26676(.A(div_curr_q[50]), .B(exu_n16257), .Y(exu_n31108));
INVX1 exu_U26677(.A(exu_n31108), .Y(exu_n8867));
AND2X1 exu_U26678(.A(div_curr_q[49]), .B(exu_n16257), .Y(exu_n31110));
INVX1 exu_U26679(.A(exu_n31110), .Y(exu_n8868));
AND2X1 exu_U26680(.A(div_curr_q[3]), .B(exu_n16257), .Y(exu_n31112));
INVX1 exu_U26681(.A(exu_n31112), .Y(exu_n8869));
AND2X1 exu_U26682(.A(div_curr_q[48]), .B(exu_n16257), .Y(exu_n31114));
INVX1 exu_U26683(.A(exu_n31114), .Y(exu_n8870));
AND2X1 exu_U26684(.A(div_curr_q[47]), .B(exu_n16257), .Y(exu_n31116));
INVX1 exu_U26685(.A(exu_n31116), .Y(exu_n8871));
AND2X1 exu_U26686(.A(div_curr_q[46]), .B(exu_n16257), .Y(exu_n31118));
INVX1 exu_U26687(.A(exu_n31118), .Y(exu_n8872));
AND2X1 exu_U26688(.A(div_curr_q[45]), .B(exu_n16257), .Y(exu_n31120));
INVX1 exu_U26689(.A(exu_n31120), .Y(exu_n8873));
AND2X1 exu_U26690(.A(div_curr_q[44]), .B(exu_n16257), .Y(exu_n31122));
INVX1 exu_U26691(.A(exu_n31122), .Y(exu_n8874));
AND2X1 exu_U26692(.A(div_curr_q[43]), .B(exu_n16257), .Y(exu_n31124));
INVX1 exu_U26693(.A(exu_n31124), .Y(exu_n8875));
AND2X1 exu_U26694(.A(div_curr_q[42]), .B(exu_n16257), .Y(exu_n31126));
INVX1 exu_U26695(.A(exu_n31126), .Y(exu_n8876));
AND2X1 exu_U26696(.A(div_curr_q[41]), .B(exu_n16257), .Y(exu_n31128));
INVX1 exu_U26697(.A(exu_n31128), .Y(exu_n8877));
AND2X1 exu_U26698(.A(div_curr_q[40]), .B(exu_n16257), .Y(exu_n31130));
INVX1 exu_U26699(.A(exu_n31130), .Y(exu_n8878));
AND2X1 exu_U26700(.A(div_curr_q[39]), .B(exu_n16257), .Y(exu_n31132));
INVX1 exu_U26701(.A(exu_n31132), .Y(exu_n8879));
AND2X1 exu_U26702(.A(div_curr_q[2]), .B(exu_n16257), .Y(exu_n31134));
INVX1 exu_U26703(.A(exu_n31134), .Y(exu_n8880));
AND2X1 exu_U26704(.A(div_curr_q[38]), .B(exu_n16257), .Y(exu_n31136));
INVX1 exu_U26705(.A(exu_n31136), .Y(exu_n8881));
AND2X1 exu_U26706(.A(div_curr_q[37]), .B(exu_n16257), .Y(exu_n31138));
INVX1 exu_U26707(.A(exu_n31138), .Y(exu_n8882));
AND2X1 exu_U26708(.A(div_curr_q[36]), .B(exu_n16257), .Y(exu_n31140));
INVX1 exu_U26709(.A(exu_n31140), .Y(exu_n8883));
AND2X1 exu_U26710(.A(div_curr_q[35]), .B(exu_n16257), .Y(exu_n31142));
INVX1 exu_U26711(.A(exu_n31142), .Y(exu_n8884));
AND2X1 exu_U26712(.A(div_curr_q[34]), .B(exu_n16257), .Y(exu_n31144));
INVX1 exu_U26713(.A(exu_n31144), .Y(exu_n8885));
AND2X1 exu_U26714(.A(div_curr_q[33]), .B(exu_n16257), .Y(exu_n31146));
INVX1 exu_U26715(.A(exu_n31146), .Y(exu_n8886));
AND2X1 exu_U26716(.A(div_curr_q[32]), .B(exu_n16257), .Y(exu_n31148));
INVX1 exu_U26717(.A(exu_n31148), .Y(exu_n8887));
AND2X1 exu_U26718(.A(div_curr_q[31]), .B(exu_n16257), .Y(exu_n31150));
INVX1 exu_U26719(.A(exu_n31150), .Y(exu_n8888));
AND2X1 exu_U26720(.A(div_curr_q[30]), .B(exu_n16257), .Y(exu_n31152));
INVX1 exu_U26721(.A(exu_n31152), .Y(exu_n8889));
AND2X1 exu_U26722(.A(div_curr_q[29]), .B(exu_n16257), .Y(exu_n31154));
INVX1 exu_U26723(.A(exu_n31154), .Y(exu_n8890));
AND2X1 exu_U26724(.A(div_curr_q[1]), .B(exu_n16257), .Y(exu_n31156));
INVX1 exu_U26725(.A(exu_n31156), .Y(exu_n8891));
AND2X1 exu_U26726(.A(div_curr_q[28]), .B(exu_n16257), .Y(exu_n31158));
INVX1 exu_U26727(.A(exu_n31158), .Y(exu_n8892));
AND2X1 exu_U26728(.A(div_curr_q[27]), .B(exu_n16257), .Y(exu_n31160));
INVX1 exu_U26729(.A(exu_n31160), .Y(exu_n8893));
AND2X1 exu_U26730(.A(div_curr_q[26]), .B(exu_n16257), .Y(exu_n31162));
INVX1 exu_U26731(.A(exu_n31162), .Y(exu_n8894));
AND2X1 exu_U26732(.A(div_curr_q[25]), .B(exu_n16257), .Y(exu_n31164));
INVX1 exu_U26733(.A(exu_n31164), .Y(exu_n8895));
AND2X1 exu_U26734(.A(div_curr_q[24]), .B(exu_n16257), .Y(exu_n31166));
INVX1 exu_U26735(.A(exu_n31166), .Y(exu_n8896));
AND2X1 exu_U26736(.A(div_curr_q[23]), .B(exu_n16257), .Y(exu_n31168));
INVX1 exu_U26737(.A(exu_n31168), .Y(exu_n8897));
AND2X1 exu_U26738(.A(div_curr_q[22]), .B(exu_n16257), .Y(exu_n31170));
INVX1 exu_U26739(.A(exu_n31170), .Y(exu_n8898));
AND2X1 exu_U26740(.A(div_curr_q[21]), .B(exu_n16257), .Y(exu_n31172));
INVX1 exu_U26741(.A(exu_n31172), .Y(exu_n8899));
AND2X1 exu_U26742(.A(div_curr_q[20]), .B(exu_n16257), .Y(exu_n31174));
INVX1 exu_U26743(.A(exu_n31174), .Y(exu_n8900));
AND2X1 exu_U26744(.A(div_curr_q[19]), .B(exu_n16257), .Y(exu_n31176));
INVX1 exu_U26745(.A(exu_n31176), .Y(exu_n8901));
AND2X1 exu_U26746(.A(div_curr_q[0]), .B(exu_n16257), .Y(exu_n31178));
INVX1 exu_U26747(.A(exu_n31178), .Y(exu_n8902));
AND2X1 exu_U26748(.A(div_curr_q[18]), .B(exu_n16257), .Y(exu_n31180));
INVX1 exu_U26749(.A(exu_n31180), .Y(exu_n8903));
AND2X1 exu_U26750(.A(div_curr_q[17]), .B(exu_n16257), .Y(exu_n31182));
INVX1 exu_U26751(.A(exu_n31182), .Y(exu_n8904));
AND2X1 exu_U26752(.A(div_curr_q[16]), .B(exu_n16257), .Y(exu_n31184));
INVX1 exu_U26753(.A(exu_n31184), .Y(exu_n8905));
AND2X1 exu_U26754(.A(div_curr_q[15]), .B(exu_n16257), .Y(exu_n31186));
INVX1 exu_U26755(.A(exu_n31186), .Y(exu_n8906));
AND2X1 exu_U26756(.A(div_curr_q[14]), .B(exu_n16257), .Y(exu_n31188));
INVX1 exu_U26757(.A(exu_n31188), .Y(exu_n8907));
AND2X1 exu_U26758(.A(div_curr_q[13]), .B(exu_n16257), .Y(exu_n31190));
INVX1 exu_U26759(.A(exu_n31190), .Y(exu_n8908));
AND2X1 exu_U26760(.A(div_curr_q[12]), .B(exu_n16257), .Y(exu_n31192));
INVX1 exu_U26761(.A(exu_n31192), .Y(exu_n8909));
AND2X1 exu_U26762(.A(div_curr_q[11]), .B(exu_n16257), .Y(exu_n31194));
INVX1 exu_U26763(.A(exu_n31194), .Y(exu_n8910));
AND2X1 exu_U26764(.A(div_curr_q[10]), .B(exu_n16257), .Y(exu_n31196));
INVX1 exu_U26765(.A(exu_n31196), .Y(exu_n8911));
AND2X1 exu_U26766(.A(div_curr_q[9]), .B(exu_n16257), .Y(exu_n31198));
INVX1 exu_U26767(.A(exu_n31198), .Y(exu_n8912));
AND2X1 exu_U26768(.A(div_d_63), .B(exu_n16257), .Y(exu_n31200));
INVX1 exu_U26769(.A(exu_n31200), .Y(exu_n8913));
AND2X1 exu_U26770(.A(div_spr_out[9]), .B(exu_n16205), .Y(exu_n31202));
INVX1 exu_U26771(.A(exu_n31202), .Y(exu_n8914));
AND2X1 exu_U26772(.A(div_spr_out[8]), .B(exu_n16206), .Y(exu_n31204));
INVX1 exu_U26773(.A(exu_n31204), .Y(exu_n8915));
AND2X1 exu_U26774(.A(div_spr_out[7]), .B(exu_n16216), .Y(exu_n31206));
INVX1 exu_U26775(.A(exu_n31206), .Y(exu_n8916));
AND2X1 exu_U26776(.A(div_spr_out[6]), .B(exu_n16219), .Y(exu_n31208));
INVX1 exu_U26777(.A(exu_n31208), .Y(exu_n8917));
AND2X1 exu_U26778(.A(div_spr_out[63]), .B(exu_n16218), .Y(exu_n31210));
INVX1 exu_U26779(.A(exu_n31210), .Y(exu_n8918));
AND2X1 exu_U26780(.A(div_spr_out[62]), .B(exu_n16218), .Y(exu_n31212));
INVX1 exu_U26781(.A(exu_n31212), .Y(exu_n8919));
AND2X1 exu_U26782(.A(div_spr_out[61]), .B(exu_n16205), .Y(exu_n31214));
INVX1 exu_U26783(.A(exu_n31214), .Y(exu_n8920));
AND2X1 exu_U26784(.A(div_spr_out[60]), .B(exu_n16216), .Y(exu_n31216));
INVX1 exu_U26785(.A(exu_n31216), .Y(exu_n8921));
AND2X1 exu_U26786(.A(div_spr_out[5]), .B(exu_n16215), .Y(exu_n31218));
INVX1 exu_U26787(.A(exu_n31218), .Y(exu_n8922));
AND2X1 exu_U26788(.A(div_spr_out[59]), .B(exu_n16217), .Y(exu_n31220));
INVX1 exu_U26789(.A(exu_n31220), .Y(exu_n8923));
AND2X1 exu_U26790(.A(div_spr_out[58]), .B(exu_n16219), .Y(exu_n31222));
INVX1 exu_U26791(.A(exu_n31222), .Y(exu_n8924));
AND2X1 exu_U26792(.A(div_spr_out[57]), .B(exu_n16206), .Y(exu_n31224));
INVX1 exu_U26793(.A(exu_n31224), .Y(exu_n8925));
AND2X1 exu_U26794(.A(div_spr_out[56]), .B(exu_n16218), .Y(exu_n31226));
INVX1 exu_U26795(.A(exu_n31226), .Y(exu_n8926));
AND2X1 exu_U26796(.A(div_spr_out[55]), .B(exu_n16205), .Y(exu_n31228));
INVX1 exu_U26797(.A(exu_n31228), .Y(exu_n8927));
AND2X1 exu_U26798(.A(div_spr_out[54]), .B(exu_n16216), .Y(exu_n31230));
INVX1 exu_U26799(.A(exu_n31230), .Y(exu_n8928));
AND2X1 exu_U26800(.A(div_spr_out[53]), .B(exu_n16215), .Y(exu_n31232));
INVX1 exu_U26801(.A(exu_n31232), .Y(exu_n8929));
AND2X1 exu_U26802(.A(div_spr_out[52]), .B(exu_n16217), .Y(exu_n31234));
INVX1 exu_U26803(.A(exu_n31234), .Y(exu_n8930));
AND2X1 exu_U26804(.A(div_spr_out[51]), .B(exu_n16219), .Y(exu_n31236));
INVX1 exu_U26805(.A(exu_n31236), .Y(exu_n8931));
AND2X1 exu_U26806(.A(div_spr_out[50]), .B(exu_n16206), .Y(exu_n31238));
INVX1 exu_U26807(.A(exu_n31238), .Y(exu_n8932));
AND2X1 exu_U26808(.A(div_spr_out[4]), .B(exu_n16218), .Y(exu_n31240));
INVX1 exu_U26809(.A(exu_n31240), .Y(exu_n8933));
AND2X1 exu_U26810(.A(div_spr_out[49]), .B(exu_n16205), .Y(exu_n31242));
INVX1 exu_U26811(.A(exu_n31242), .Y(exu_n8934));
AND2X1 exu_U26812(.A(div_spr_out[48]), .B(exu_n16215), .Y(exu_n31244));
INVX1 exu_U26813(.A(exu_n31244), .Y(exu_n8935));
AND2X1 exu_U26814(.A(div_spr_out[47]), .B(exu_n16217), .Y(exu_n31246));
INVX1 exu_U26815(.A(exu_n31246), .Y(exu_n8936));
AND2X1 exu_U26816(.A(div_spr_out[46]), .B(exu_n16205), .Y(exu_n31248));
INVX1 exu_U26817(.A(exu_n31248), .Y(exu_n8937));
AND2X1 exu_U26818(.A(div_spr_out[45]), .B(exu_n16215), .Y(exu_n31250));
INVX1 exu_U26819(.A(exu_n31250), .Y(exu_n8938));
AND2X1 exu_U26820(.A(div_spr_out[44]), .B(exu_n16217), .Y(exu_n31252));
INVX1 exu_U26821(.A(exu_n31252), .Y(exu_n8939));
AND2X1 exu_U26822(.A(div_spr_out[43]), .B(exu_n16205), .Y(exu_n31254));
INVX1 exu_U26823(.A(exu_n31254), .Y(exu_n8940));
AND2X1 exu_U26824(.A(div_spr_out[42]), .B(exu_n16215), .Y(exu_n31256));
INVX1 exu_U26825(.A(exu_n31256), .Y(exu_n8941));
AND2X1 exu_U26826(.A(div_spr_out[41]), .B(exu_n16217), .Y(exu_n31258));
INVX1 exu_U26827(.A(exu_n31258), .Y(exu_n8942));
AND2X1 exu_U26828(.A(div_spr_out[40]), .B(exu_n16205), .Y(exu_n31260));
INVX1 exu_U26829(.A(exu_n31260), .Y(exu_n8943));
AND2X1 exu_U26830(.A(div_spr_out[3]), .B(exu_n16219), .Y(exu_n31262));
INVX1 exu_U26831(.A(exu_n31262), .Y(exu_n8944));
AND2X1 exu_U26832(.A(div_spr_out[39]), .B(exu_n16206), .Y(exu_n31264));
INVX1 exu_U26833(.A(exu_n31264), .Y(exu_n8945));
AND2X1 exu_U26834(.A(div_spr_out[38]), .B(exu_n16218), .Y(exu_n31266));
INVX1 exu_U26835(.A(exu_n31266), .Y(exu_n8946));
AND2X1 exu_U26836(.A(div_spr_out[37]), .B(exu_n16216), .Y(exu_n31268));
INVX1 exu_U26837(.A(exu_n31268), .Y(exu_n8947));
AND2X1 exu_U26838(.A(div_spr_out[36]), .B(exu_n16205), .Y(exu_n31270));
INVX1 exu_U26839(.A(exu_n31270), .Y(exu_n8948));
AND2X1 exu_U26840(.A(div_spr_out[35]), .B(exu_n16205), .Y(exu_n31272));
INVX1 exu_U26841(.A(exu_n31272), .Y(exu_n8949));
AND2X1 exu_U26842(.A(div_spr_out[34]), .B(exu_n16205), .Y(exu_n31274));
INVX1 exu_U26843(.A(exu_n31274), .Y(exu_n8950));
AND2X1 exu_U26844(.A(div_spr_out[33]), .B(exu_n16205), .Y(exu_n31276));
INVX1 exu_U26845(.A(exu_n31276), .Y(exu_n8951));
AND2X1 exu_U26846(.A(div_spr_out[32]), .B(exu_n16217), .Y(exu_n31278));
INVX1 exu_U26847(.A(exu_n31278), .Y(exu_n8952));
AND2X1 exu_U26848(.A(div_spr_out[31]), .B(exu_n16205), .Y(exu_n31280));
INVX1 exu_U26849(.A(exu_n31280), .Y(exu_n8953));
AND2X1 exu_U26850(.A(div_spr_out[30]), .B(exu_n16219), .Y(exu_n31282));
INVX1 exu_U26851(.A(exu_n31282), .Y(exu_n8954));
AND2X1 exu_U26852(.A(div_spr_out[2]), .B(exu_n16206), .Y(exu_n31284));
INVX1 exu_U26853(.A(exu_n31284), .Y(exu_n8955));
AND2X1 exu_U26854(.A(div_spr_out[29]), .B(exu_n16218), .Y(exu_n31286));
INVX1 exu_U26855(.A(exu_n31286), .Y(exu_n8956));
AND2X1 exu_U26856(.A(div_spr_out[28]), .B(exu_n16216), .Y(exu_n31288));
INVX1 exu_U26857(.A(exu_n31288), .Y(exu_n8957));
AND2X1 exu_U26858(.A(div_spr_out[27]), .B(exu_n16215), .Y(exu_n31290));
INVX1 exu_U26859(.A(exu_n31290), .Y(exu_n8958));
AND2X1 exu_U26860(.A(div_spr_out[26]), .B(exu_n16217), .Y(exu_n31292));
INVX1 exu_U26861(.A(exu_n31292), .Y(exu_n8959));
AND2X1 exu_U26862(.A(div_spr_out[25]), .B(exu_n16205), .Y(exu_n31294));
INVX1 exu_U26863(.A(exu_n31294), .Y(exu_n8960));
AND2X1 exu_U26864(.A(div_spr_out[24]), .B(exu_n16219), .Y(exu_n31296));
INVX1 exu_U26865(.A(exu_n31296), .Y(exu_n8961));
AND2X1 exu_U26866(.A(div_spr_out[23]), .B(exu_n16206), .Y(exu_n31298));
INVX1 exu_U26867(.A(exu_n31298), .Y(exu_n8962));
AND2X1 exu_U26868(.A(div_spr_out[22]), .B(exu_n16219), .Y(exu_n31300));
INVX1 exu_U26869(.A(exu_n31300), .Y(exu_n8963));
AND2X1 exu_U26870(.A(div_spr_out[21]), .B(exu_n16219), .Y(exu_n31302));
INVX1 exu_U26871(.A(exu_n31302), .Y(exu_n8964));
AND2X1 exu_U26872(.A(div_spr_out[20]), .B(exu_n16219), .Y(exu_n31304));
INVX1 exu_U26873(.A(exu_n31304), .Y(exu_n8965));
AND2X1 exu_U26874(.A(div_spr_out[1]), .B(exu_n16219), .Y(exu_n31306));
INVX1 exu_U26875(.A(exu_n31306), .Y(exu_n8966));
AND2X1 exu_U26876(.A(div_spr_out[19]), .B(exu_n16219), .Y(exu_n31308));
INVX1 exu_U26877(.A(exu_n31308), .Y(exu_n8967));
AND2X1 exu_U26878(.A(div_spr_out[18]), .B(exu_n16219), .Y(exu_n31310));
INVX1 exu_U26879(.A(exu_n31310), .Y(exu_n8968));
AND2X1 exu_U26880(.A(div_spr_out[17]), .B(exu_n16219), .Y(exu_n31312));
INVX1 exu_U26881(.A(exu_n31312), .Y(exu_n8969));
AND2X1 exu_U26882(.A(div_spr_out[16]), .B(exu_n16219), .Y(exu_n31314));
INVX1 exu_U26883(.A(exu_n31314), .Y(exu_n8970));
AND2X1 exu_U26884(.A(div_spr_out[15]), .B(exu_n16219), .Y(exu_n31316));
INVX1 exu_U26885(.A(exu_n31316), .Y(exu_n8971));
AND2X1 exu_U26886(.A(div_spr_out[14]), .B(exu_n16219), .Y(exu_n31318));
INVX1 exu_U26887(.A(exu_n31318), .Y(exu_n8972));
AND2X1 exu_U26888(.A(div_spr_out[13]), .B(exu_n16218), .Y(exu_n31320));
INVX1 exu_U26889(.A(exu_n31320), .Y(exu_n8973));
AND2X1 exu_U26890(.A(div_spr_out[12]), .B(exu_n16217), .Y(exu_n31322));
INVX1 exu_U26891(.A(exu_n31322), .Y(exu_n8974));
AND2X1 exu_U26892(.A(div_spr_out[11]), .B(exu_n16216), .Y(exu_n31324));
INVX1 exu_U26893(.A(exu_n31324), .Y(exu_n8975));
AND2X1 exu_U26894(.A(div_spr_out[10]), .B(exu_n16206), .Y(exu_n31326));
INVX1 exu_U26895(.A(exu_n31326), .Y(exu_n8976));
AND2X1 exu_U26896(.A(div_spr_out[0]), .B(exu_n16216), .Y(exu_n31328));
INVX1 exu_U26897(.A(exu_n31328), .Y(exu_n8977));
AND2X1 exu_U26898(.A(ecl_writeback_ecl_sel_mul_g), .B(ecl_mdqctl_wb_multhr_g[1]), .Y(exu_n31460));
INVX1 exu_U26899(.A(exu_n31460), .Y(exu_n8978));
AND2X1 exu_U26900(.A(exu_n16271), .B(ecl_writeback_dfill_tid_g2[1]), .Y(exu_n31462));
INVX1 exu_U26901(.A(exu_n31462), .Y(exu_n8979));
AND2X1 exu_U26902(.A(ecl_mdqctl_wb_multhr_g[0]), .B(ecl_writeback_ecl_sel_mul_g), .Y(exu_n31466));
INVX1 exu_U26903(.A(exu_n31466), .Y(exu_n8980));
AND2X1 exu_U26904(.A(ecl_writeback_dfill_tid_g2[0]), .B(exu_n16271), .Y(exu_n31468));
INVX1 exu_U26905(.A(exu_n31468), .Y(exu_n8981));
AND2X1 exu_U26906(.A(rml_cwp_swap_keep_state[0]), .B(rml_cwp_swap_slot0_state_valid[1]), .Y(exu_n31471));
INVX1 exu_U26907(.A(exu_n31471), .Y(exu_n8982));
AND2X1 exu_U26908(.A(rml_cwp_swap_keep_state[1]), .B(rml_cwp_swap_slot1_state_valid[1]), .Y(exu_n31476));
INVX1 exu_U26909(.A(exu_n31476), .Y(exu_n8983));
AND2X1 exu_U26910(.A(rml_cwp_swap_keep_state[2]), .B(rml_cwp_swap_slot2_state_valid[1]), .Y(exu_n31481));
INVX1 exu_U26911(.A(exu_n31481), .Y(exu_n8984));
AND2X1 exu_U26912(.A(rml_cwp_swap_keep_state[3]), .B(rml_cwp_swap_slot3_state_valid[1]), .Y(exu_n31486));
INVX1 exu_U26913(.A(exu_n31486), .Y(exu_n8985));
OR2X1 exu_U26914(.A(exu_n12039), .B(exu_n14927), .Y(exu_n31619));
INVX1 exu_U26915(.A(exu_n31619), .Y(exu_n8986));
OR2X1 exu_U26916(.A(byp_alu_rcc_data_e[1]), .B(byp_alu_rcc_data_e[19]), .Y(exu_n31623));
INVX1 exu_U26917(.A(exu_n31623), .Y(exu_n8987));
OR2X1 exu_U26918(.A(byp_alu_rcc_data_e[23]), .B(byp_alu_rcc_data_e[22]), .Y(exu_n31625));
INVX1 exu_U26919(.A(exu_n31625), .Y(exu_n8988));
OR2X1 exu_U26920(.A(byp_alu_rcc_data_e[12]), .B(byp_alu_rcc_data_e[11]), .Y(exu_n31629));
INVX1 exu_U26921(.A(exu_n31629), .Y(exu_n8989));
OR2X1 exu_U26922(.A(byp_alu_rcc_data_e[16]), .B(byp_alu_rcc_data_e[15]), .Y(exu_n31631));
INVX1 exu_U26923(.A(exu_n31631), .Y(exu_n8990));
OR2X1 exu_U26924(.A(exu_n12041), .B(exu_n14929), .Y(exu_n31633));
INVX1 exu_U26925(.A(exu_n31633), .Y(exu_n8991));
OR2X1 exu_U26926(.A(byp_alu_rcc_data_e[5]), .B(byp_alu_rcc_data_e[4]), .Y(exu_n31637));
INVX1 exu_U26927(.A(exu_n31637), .Y(exu_n8992));
OR2X1 exu_U26928(.A(byp_alu_rcc_data_e[9]), .B(byp_alu_rcc_data_e[8]), .Y(exu_n31639));
INVX1 exu_U26929(.A(exu_n31639), .Y(exu_n8993));
OR2X1 exu_U26930(.A(byp_alu_rcc_data_e[27]), .B(byp_alu_rcc_data_e[26]), .Y(exu_n31643));
INVX1 exu_U26931(.A(exu_n31643), .Y(exu_n8994));
OR2X1 exu_U26932(.A(byp_alu_rcc_data_e[30]), .B(byp_alu_rcc_data_e[2]), .Y(exu_n31645));
INVX1 exu_U26933(.A(exu_n31645), .Y(exu_n8995));
OR2X1 exu_U26934(.A(exu_n12043), .B(exu_n14931), .Y(exu_n31649));
INVX1 exu_U26935(.A(exu_n31649), .Y(exu_n8996));
OR2X1 exu_U26936(.A(byp_alu_rcc_data_e[33]), .B(byp_alu_rcc_data_e[51]), .Y(exu_n31653));
INVX1 exu_U26937(.A(exu_n31653), .Y(exu_n8997));
OR2X1 exu_U26938(.A(byp_alu_rcc_data_e[55]), .B(byp_alu_rcc_data_e[54]), .Y(exu_n31655));
INVX1 exu_U26939(.A(exu_n31655), .Y(exu_n8998));
OR2X1 exu_U26940(.A(byp_alu_rcc_data_e[44]), .B(byp_alu_rcc_data_e[43]), .Y(exu_n31659));
INVX1 exu_U26941(.A(exu_n31659), .Y(exu_n8999));
OR2X1 exu_U26942(.A(byp_alu_rcc_data_e[48]), .B(byp_alu_rcc_data_e[47]), .Y(exu_n31661));
INVX1 exu_U26943(.A(exu_n31661), .Y(exu_n9000));
OR2X1 exu_U26944(.A(exu_n12045), .B(exu_n14933), .Y(exu_n31663));
INVX1 exu_U26945(.A(exu_n31663), .Y(exu_n9001));
OR2X1 exu_U26946(.A(byp_alu_rcc_data_e[37]), .B(byp_alu_rcc_data_e[36]), .Y(exu_n31667));
INVX1 exu_U26947(.A(exu_n31667), .Y(exu_n9002));
OR2X1 exu_U26948(.A(byp_alu_rcc_data_e[41]), .B(byp_alu_rcc_data_e[40]), .Y(exu_n31669));
INVX1 exu_U26949(.A(exu_n31669), .Y(exu_n9003));
OR2X1 exu_U26950(.A(byp_alu_rcc_data_e[59]), .B(byp_alu_rcc_data_e[58]), .Y(exu_n31673));
INVX1 exu_U26951(.A(exu_n31673), .Y(exu_n9004));
OR2X1 exu_U26952(.A(byp_alu_rcc_data_e[62]), .B(byp_alu_rcc_data_e[34]), .Y(exu_n31675));
INVX1 exu_U26953(.A(exu_n31675), .Y(exu_n9005));
OR2X1 exu_U26954(.A(exu_n12047), .B(exu_n14935), .Y(exu_n31679));
INVX1 exu_U26955(.A(exu_n31679), .Y(exu_n9006));
OR2X1 exu_U26956(.A(div_u32eql_inxor[1]), .B(div_u32eql_inxor[19]), .Y(exu_n31683));
INVX1 exu_U26957(.A(exu_n31683), .Y(exu_n9007));
OR2X1 exu_U26958(.A(div_u32eql_inxor[23]), .B(div_u32eql_inxor[22]), .Y(exu_n31685));
INVX1 exu_U26959(.A(exu_n31685), .Y(exu_n9008));
OR2X1 exu_U26960(.A(div_u32eql_inxor[12]), .B(div_u32eql_inxor[11]), .Y(exu_n31688));
INVX1 exu_U26961(.A(exu_n31688), .Y(exu_n9009));
OR2X1 exu_U26962(.A(div_u32eql_inxor[16]), .B(div_u32eql_inxor[15]), .Y(exu_n31690));
INVX1 exu_U26963(.A(exu_n31690), .Y(exu_n9010));
OR2X1 exu_U26964(.A(exu_n12049), .B(exu_n14937), .Y(exu_n31692));
INVX1 exu_U26965(.A(exu_n31692), .Y(exu_n9011));
OR2X1 exu_U26966(.A(div_u32eql_inxor[5]), .B(div_u32eql_inxor[4]), .Y(exu_n31696));
INVX1 exu_U26967(.A(exu_n31696), .Y(exu_n9012));
OR2X1 exu_U26968(.A(div_u32eql_inxor[9]), .B(div_u32eql_inxor[8]), .Y(exu_n31698));
INVX1 exu_U26969(.A(exu_n31698), .Y(exu_n9013));
OR2X1 exu_U26970(.A(div_u32eql_inxor[27]), .B(div_u32eql_inxor[26]), .Y(exu_n31702));
INVX1 exu_U26971(.A(exu_n31702), .Y(exu_n9014));
OR2X1 exu_U26972(.A(div_u32eql_inxor[30]), .B(div_u32eql_inxor[2]), .Y(exu_n31704));
INVX1 exu_U26973(.A(exu_n31704), .Y(exu_n9015));
AND2X1 exu_U26974(.A(rml_cwp_swap_sel[2]), .B(rml_cwp_swap_slot2_data[9]), .Y(rml_cwp_cwp_output_mux_n4));
INVX1 exu_U26975(.A(rml_cwp_cwp_output_mux_n4), .Y(exu_n9016));
AND2X1 exu_U26976(.A(exu_n15025), .B(rml_cwp_swap_slot0_data[9]), .Y(rml_cwp_cwp_output_mux_n6));
INVX1 exu_U26977(.A(rml_cwp_cwp_output_mux_n6), .Y(exu_n9017));
AND2X1 exu_U26978(.A(rml_cwp_swap_slot2_data[8]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n10));
INVX1 exu_U26979(.A(rml_cwp_cwp_output_mux_n10), .Y(exu_n9018));
AND2X1 exu_U26980(.A(rml_cwp_swap_slot0_data[8]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n12));
INVX1 exu_U26981(.A(rml_cwp_cwp_output_mux_n12), .Y(exu_n9019));
AND2X1 exu_U26982(.A(rml_cwp_swap_slot2_data[7]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n16));
INVX1 exu_U26983(.A(rml_cwp_cwp_output_mux_n16), .Y(exu_n9020));
AND2X1 exu_U26984(.A(rml_cwp_swap_slot0_data[7]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n18));
INVX1 exu_U26985(.A(rml_cwp_cwp_output_mux_n18), .Y(exu_n9021));
AND2X1 exu_U26986(.A(rml_cwp_swap_slot2_data[6]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n22));
INVX1 exu_U26987(.A(rml_cwp_cwp_output_mux_n22), .Y(exu_n9022));
AND2X1 exu_U26988(.A(rml_cwp_swap_slot0_data[6]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n24));
INVX1 exu_U26989(.A(rml_cwp_cwp_output_mux_n24), .Y(exu_n9023));
AND2X1 exu_U26990(.A(rml_cwp_swap_slot2_data[5]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n28));
INVX1 exu_U26991(.A(rml_cwp_cwp_output_mux_n28), .Y(exu_n9024));
AND2X1 exu_U26992(.A(rml_cwp_swap_slot0_data[5]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n30));
INVX1 exu_U26993(.A(rml_cwp_cwp_output_mux_n30), .Y(exu_n9025));
AND2X1 exu_U26994(.A(rml_cwp_swap_slot2_data[4]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n34));
INVX1 exu_U26995(.A(rml_cwp_cwp_output_mux_n34), .Y(exu_n9026));
AND2X1 exu_U26996(.A(rml_cwp_swap_slot0_data[4]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n36));
INVX1 exu_U26997(.A(rml_cwp_cwp_output_mux_n36), .Y(exu_n9027));
AND2X1 exu_U26998(.A(rml_cwp_swap_slot2_data[3]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n40));
INVX1 exu_U26999(.A(rml_cwp_cwp_output_mux_n40), .Y(exu_n9028));
AND2X1 exu_U27000(.A(rml_cwp_swap_slot0_data[3]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n42));
INVX1 exu_U27001(.A(rml_cwp_cwp_output_mux_n42), .Y(exu_n9029));
AND2X1 exu_U27002(.A(rml_cwp_swap_slot2_data[2]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n46));
INVX1 exu_U27003(.A(rml_cwp_cwp_output_mux_n46), .Y(exu_n9030));
AND2X1 exu_U27004(.A(rml_cwp_swap_slot0_data[2]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n48));
INVX1 exu_U27005(.A(rml_cwp_cwp_output_mux_n48), .Y(exu_n9031));
AND2X1 exu_U27006(.A(rml_cwp_swap_slot2_data[1]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n52));
INVX1 exu_U27007(.A(rml_cwp_cwp_output_mux_n52), .Y(exu_n9032));
AND2X1 exu_U27008(.A(rml_cwp_swap_slot0_data[1]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n54));
INVX1 exu_U27009(.A(rml_cwp_cwp_output_mux_n54), .Y(exu_n9033));
AND2X1 exu_U27010(.A(rml_cwp_swap_slot2_state[1]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n58));
INVX1 exu_U27011(.A(rml_cwp_cwp_output_mux_n58), .Y(exu_n9034));
AND2X1 exu_U27012(.A(rml_cwp_swap_slot0_state[1]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n60));
INVX1 exu_U27013(.A(rml_cwp_cwp_output_mux_n60), .Y(exu_n9035));
AND2X1 exu_U27014(.A(rml_cwp_swap_slot2_state_valid[0]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n64));
INVX1 exu_U27015(.A(rml_cwp_cwp_output_mux_n64), .Y(exu_n9036));
AND2X1 exu_U27016(.A(rml_cwp_swap_slot0_state_valid[0]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n66));
INVX1 exu_U27017(.A(rml_cwp_cwp_output_mux_n66), .Y(exu_n9037));
AND2X1 exu_U27018(.A(rml_cwp_swap_slot2_data[12]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n70));
INVX1 exu_U27019(.A(rml_cwp_cwp_output_mux_n70), .Y(exu_n9038));
AND2X1 exu_U27020(.A(rml_cwp_swap_slot0_data[12]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n72));
INVX1 exu_U27021(.A(rml_cwp_cwp_output_mux_n72), .Y(exu_n9039));
AND2X1 exu_U27022(.A(rml_cwp_swap_slot2_data[11]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n76));
INVX1 exu_U27023(.A(rml_cwp_cwp_output_mux_n76), .Y(exu_n9040));
AND2X1 exu_U27024(.A(rml_cwp_swap_slot0_data[11]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n78));
INVX1 exu_U27025(.A(rml_cwp_cwp_output_mux_n78), .Y(exu_n9041));
AND2X1 exu_U27026(.A(rml_cwp_swap_slot2_data[10]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n82));
INVX1 exu_U27027(.A(rml_cwp_cwp_output_mux_n82), .Y(exu_n9042));
AND2X1 exu_U27028(.A(rml_cwp_swap_slot0_data[10]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n84));
INVX1 exu_U27029(.A(rml_cwp_cwp_output_mux_n84), .Y(exu_n9043));
AND2X1 exu_U27030(.A(rml_cwp_swap_slot2_data[0]), .B(rml_cwp_swap_sel[2]), .Y(rml_cwp_cwp_output_mux_n88));
INVX1 exu_U27031(.A(rml_cwp_cwp_output_mux_n88), .Y(exu_n9044));
AND2X1 exu_U27032(.A(rml_cwp_swap_slot0_data[0]), .B(exu_n15025), .Y(rml_cwp_cwp_output_mux_n90));
INVX1 exu_U27033(.A(rml_cwp_cwp_output_mux_n90), .Y(exu_n9045));
AND2X1 exu_U27034(.A(rml_cwp_cwp_output_queue_n22), .B(exu_n10312), .Y(rml_cwp_cwp_output_queue_n18));
INVX1 exu_U27035(.A(rml_cwp_cwp_output_queue_n18), .Y(exu_n9046));
AND2X1 exu_U27036(.A(exu_n16617), .B(exu_n10314), .Y(rml_cwp_cwp_output_queue_n23));
INVX1 exu_U27037(.A(rml_cwp_cwp_output_queue_n23), .Y(exu_n9047));
AND2X1 exu_U27038(.A(exu_n16511), .B(exu_n16624), .Y(rml_cwp_cwp_output_queue_n27));
INVX1 exu_U27039(.A(rml_cwp_cwp_output_queue_n27), .Y(exu_n9048));
AND2X1 exu_U27040(.A(rml_cwp_cwp_output_queue_n26), .B(exu_n10315), .Y(rml_cwp_cwp_output_queue_n28));
INVX1 exu_U27041(.A(rml_cwp_cwp_output_queue_n28), .Y(exu_n9049));
AND2X1 exu_U27042(.A(rml_cwp_cwp_output_queue_pv[3]), .B(exu_n16511), .Y(rml_cwp_cwp_output_queue_n32));
INVX1 exu_U27043(.A(rml_cwp_cwp_output_queue_n32), .Y(exu_n9050));
AND2X1 exu_U27044(.A(exu_n11557), .B(exu_n16624), .Y(rml_cwp_cwp_output_queue_n34));
INVX1 exu_U27045(.A(rml_cwp_cwp_output_queue_n34), .Y(exu_n9051));
AND2X1 exu_U27046(.A(rml_cwp_swap_req_vec[0]), .B(exu_n15365), .Y(rml_cwp_cwp_output_queue_n37));
INVX1 exu_U27047(.A(rml_cwp_cwp_output_queue_n37), .Y(exu_n9052));
AND2X1 exu_U27048(.A(rml_cwp_cwp_output_queue_pv[1]), .B(exu_n16625), .Y(rml_cwp_cwp_output_queue_n38));
INVX1 exu_U27049(.A(rml_cwp_cwp_output_queue_n38), .Y(exu_n9053));
AND2X1 exu_U27050(.A(exu_n15851), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n20));
INVX1 exu_U27051(.A(rml_cwp_slot0_data_mux_n20), .Y(exu_n9054));
AND2X1 exu_U27052(.A(exu_n15852), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n24));
INVX1 exu_U27053(.A(rml_cwp_slot0_data_mux_n24), .Y(exu_n9055));
AND2X1 exu_U27054(.A(exu_n15853), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n28));
INVX1 exu_U27055(.A(rml_cwp_slot0_data_mux_n28), .Y(exu_n9056));
AND2X1 exu_U27056(.A(rml_rml_ecl_cwp_e[2]), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n32));
INVX1 exu_U27057(.A(rml_cwp_slot0_data_mux_n32), .Y(exu_n9057));
AND2X1 exu_U27058(.A(rml_rml_ecl_cwp_e[1]), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n36));
INVX1 exu_U27059(.A(rml_cwp_slot0_data_mux_n36), .Y(exu_n9058));
AND2X1 exu_U27060(.A(rml_rml_ecl_cwp_e[0]), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n52));
INVX1 exu_U27061(.A(rml_cwp_slot0_data_mux_n52), .Y(exu_n9059));
OR2X1 exu_U27062(.A(exu_n16622), .B(exu_n14939), .Y(ecl_divcntl_cnt6_n12));
INVX1 exu_U27063(.A(ecl_divcntl_cnt6_n12), .Y(exu_n9060));
AND2X1 exu_U27064(.A(ecl_divcntl_cnt6_n20), .B(exu_n10344), .Y(ecl_divcntl_cnt6_n18));
INVX1 exu_U27065(.A(ecl_divcntl_cnt6_n18), .Y(exu_n9061));
AND2X1 exu_U27066(.A(exu_n16622), .B(ecl_divcntl_div_state_1), .Y(ecl_divcntl_cnt6_n25));
INVX1 exu_U27067(.A(ecl_divcntl_cnt6_n25), .Y(exu_n9062));
OR2X1 exu_U27068(.A(exu_n12051), .B(exu_n14940), .Y(ecl_byplog_rs1_w_comp7_n2));
INVX1 exu_U27069(.A(ecl_byplog_rs1_w_comp7_n2), .Y(exu_n9063));
AND2X1 exu_U27070(.A(exu_n15028), .B(ecl_eccctl_rs1_ce_m), .Y(ecl_eccctl_ecc_synd7_mux_n4));
INVX1 exu_U27071(.A(ecl_eccctl_ecc_synd7_mux_n4), .Y(exu_n9064));
AND2X1 exu_U27072(.A(exu_n15975), .B(ecl_ifu_exu_rs1_m[4]), .Y(ecl_eccctl_ecc_rd_mux_n4));
INVX1 exu_U27073(.A(ecl_eccctl_ecc_rd_mux_n4), .Y(exu_n9065));
AND2X1 exu_U27074(.A(ecl_ifu_exu_rs3_m[3]), .B(ecl_ecc_sel_rs3_m_l), .Y(ecl_eccctl_ecc_rd_mux_n6));
INVX1 exu_U27075(.A(ecl_eccctl_ecc_rd_mux_n6), .Y(exu_n9066));
AND2X1 exu_U27076(.A(ecl_ifu_exu_rs1_m[3]), .B(ecl_ecc_sel_rs1_m_l), .Y(ecl_eccctl_ecc_rd_mux_n8));
INVX1 exu_U27077(.A(ecl_eccctl_ecc_rd_mux_n8), .Y(exu_n9067));
AND2X1 exu_U27078(.A(ecl_ifu_exu_rs3_m[2]), .B(ecl_ecc_sel_rs3_m_l), .Y(ecl_eccctl_ecc_rd_mux_n10));
INVX1 exu_U27079(.A(ecl_eccctl_ecc_rd_mux_n10), .Y(exu_n9068));
AND2X1 exu_U27080(.A(ecl_ifu_exu_rs1_m[2]), .B(ecl_ecc_sel_rs1_m_l), .Y(ecl_eccctl_ecc_rd_mux_n12));
INVX1 exu_U27081(.A(ecl_eccctl_ecc_rd_mux_n12), .Y(exu_n9069));
AND2X1 exu_U27082(.A(ecl_ifu_exu_rs3_m[1]), .B(ecl_ecc_sel_rs3_m_l), .Y(ecl_eccctl_ecc_rd_mux_n14));
INVX1 exu_U27083(.A(ecl_eccctl_ecc_rd_mux_n14), .Y(exu_n9070));
AND2X1 exu_U27084(.A(ecl_ifu_exu_rs1_m[1]), .B(ecl_ecc_sel_rs1_m_l), .Y(ecl_eccctl_ecc_rd_mux_n16));
INVX1 exu_U27085(.A(ecl_eccctl_ecc_rd_mux_n16), .Y(exu_n9071));
AND2X1 exu_U27086(.A(ecl_ifu_exu_rs3_m[0]), .B(exu_n15973), .Y(ecl_eccctl_ecc_rd_mux_n18));
INVX1 exu_U27087(.A(ecl_eccctl_ecc_rd_mux_n18), .Y(exu_n9072));
AND2X1 exu_U27088(.A(ecl_ifu_exu_rs1_m[0]), .B(exu_n15975), .Y(ecl_eccctl_ecc_rd_mux_n20));
INVX1 exu_U27089(.A(ecl_eccctl_ecc_rd_mux_n20), .Y(exu_n9073));
AND2X1 exu_U27090(.A(exu_n15692), .B(rml_ecl_cansave_d[2]), .Y(ecl_writeback_rdpr_mux1_n4));
INVX1 exu_U27091(.A(ecl_writeback_rdpr_mux1_n4), .Y(exu_n9074));
AND2X1 exu_U27092(.A(ecl_writeback_n72), .B(rml_ecl_canrestore_d[2]), .Y(ecl_writeback_rdpr_mux1_n6));
INVX1 exu_U27093(.A(ecl_writeback_rdpr_mux1_n6), .Y(exu_n9075));
AND2X1 exu_U27094(.A(rml_ecl_cansave_d[1]), .B(exu_n15692), .Y(ecl_writeback_rdpr_mux1_n10));
INVX1 exu_U27095(.A(ecl_writeback_rdpr_mux1_n10), .Y(exu_n9076));
AND2X1 exu_U27096(.A(rml_ecl_canrestore_d[1]), .B(ecl_writeback_n72), .Y(ecl_writeback_rdpr_mux1_n12));
INVX1 exu_U27097(.A(ecl_writeback_rdpr_mux1_n12), .Y(exu_n9077));
AND2X1 exu_U27098(.A(rml_ecl_cansave_d[0]), .B(exu_n15692), .Y(ecl_writeback_rdpr_mux1_n16));
INVX1 exu_U27099(.A(ecl_writeback_rdpr_mux1_n16), .Y(exu_n9078));
AND2X1 exu_U27100(.A(rml_ecl_canrestore_d[0]), .B(ecl_writeback_n72), .Y(ecl_writeback_rdpr_mux1_n18));
INVX1 exu_U27101(.A(ecl_writeback_rdpr_mux1_n18), .Y(exu_n9079));
AND2X1 exu_U27102(.A(ecl_writeback_ecl_sel_mul_g), .B(ecl_mdqctl_wb_mulrd_g[4]), .Y(ecl_writeback_rd_g_mux_n4));
INVX1 exu_U27103(.A(ecl_writeback_rd_g_mux_n4), .Y(exu_n9080));
AND2X1 exu_U27104(.A(ecl_byp_sel_load_g), .B(ecl_wb_byplog_rd_g2[4]), .Y(ecl_writeback_rd_g_mux_n6));
INVX1 exu_U27105(.A(ecl_writeback_rd_g_mux_n6), .Y(exu_n9081));
AND2X1 exu_U27106(.A(ecl_mdqctl_wb_mulrd_g[3]), .B(ecl_writeback_ecl_sel_mul_g), .Y(ecl_writeback_rd_g_mux_n10));
INVX1 exu_U27107(.A(ecl_writeback_rd_g_mux_n10), .Y(exu_n9082));
AND2X1 exu_U27108(.A(ecl_wb_byplog_rd_g2[3]), .B(ecl_byp_sel_load_g), .Y(ecl_writeback_rd_g_mux_n12));
INVX1 exu_U27109(.A(ecl_writeback_rd_g_mux_n12), .Y(exu_n9083));
AND2X1 exu_U27110(.A(ecl_mdqctl_wb_mulrd_g[2]), .B(ecl_writeback_ecl_sel_mul_g), .Y(ecl_writeback_rd_g_mux_n16));
INVX1 exu_U27111(.A(ecl_writeback_rd_g_mux_n16), .Y(exu_n9084));
AND2X1 exu_U27112(.A(ecl_wb_byplog_rd_g2[2]), .B(ecl_byp_sel_load_g), .Y(ecl_writeback_rd_g_mux_n18));
INVX1 exu_U27113(.A(ecl_writeback_rd_g_mux_n18), .Y(exu_n9085));
AND2X1 exu_U27114(.A(ecl_mdqctl_wb_mulrd_g[1]), .B(ecl_writeback_ecl_sel_mul_g), .Y(ecl_writeback_rd_g_mux_n22));
INVX1 exu_U27115(.A(ecl_writeback_rd_g_mux_n22), .Y(exu_n9086));
AND2X1 exu_U27116(.A(ecl_wb_byplog_rd_g2[1]), .B(ecl_byp_sel_load_g), .Y(ecl_writeback_rd_g_mux_n24));
INVX1 exu_U27117(.A(ecl_writeback_rd_g_mux_n24), .Y(exu_n9087));
AND2X1 exu_U27118(.A(ecl_mdqctl_wb_mulrd_g[0]), .B(ecl_writeback_ecl_sel_mul_g), .Y(ecl_writeback_rd_g_mux_n28));
INVX1 exu_U27119(.A(ecl_writeback_rd_g_mux_n28), .Y(exu_n9088));
AND2X1 exu_U27120(.A(ecl_wb_byplog_rd_g2[0]), .B(ecl_byp_sel_load_g), .Y(ecl_writeback_rd_g_mux_n30));
INVX1 exu_U27121(.A(ecl_writeback_rd_g_mux_n30), .Y(exu_n9089));
AND2X1 exu_U27122(.A(exu_n15933), .B(exu_tlu_ccr2_w[7]), .Y(ecl_ccr_mux_ccr_out_n4));
INVX1 exu_U27123(.A(ecl_ccr_mux_ccr_out_n4), .Y(exu_n9090));
AND2X1 exu_U27124(.A(exu_n15935), .B(exu_tlu_ccr0_w[7]), .Y(ecl_ccr_mux_ccr_out_n6));
INVX1 exu_U27125(.A(ecl_ccr_mux_ccr_out_n6), .Y(exu_n9091));
AND2X1 exu_U27126(.A(exu_tlu_ccr2_w[6]), .B(exu_n15933), .Y(ecl_ccr_mux_ccr_out_n10));
INVX1 exu_U27127(.A(ecl_ccr_mux_ccr_out_n10), .Y(exu_n9092));
AND2X1 exu_U27128(.A(exu_tlu_ccr0_w[6]), .B(exu_n15935), .Y(ecl_ccr_mux_ccr_out_n12));
INVX1 exu_U27129(.A(ecl_ccr_mux_ccr_out_n12), .Y(exu_n9093));
AND2X1 exu_U27130(.A(exu_tlu_ccr2_w[5]), .B(exu_n15933), .Y(ecl_ccr_mux_ccr_out_n16));
INVX1 exu_U27131(.A(ecl_ccr_mux_ccr_out_n16), .Y(exu_n9094));
AND2X1 exu_U27132(.A(exu_tlu_ccr0_w[5]), .B(exu_n15935), .Y(ecl_ccr_mux_ccr_out_n18));
INVX1 exu_U27133(.A(ecl_ccr_mux_ccr_out_n18), .Y(exu_n9095));
AND2X1 exu_U27134(.A(exu_tlu_ccr2_w[4]), .B(exu_n15933), .Y(ecl_ccr_mux_ccr_out_n22));
INVX1 exu_U27135(.A(ecl_ccr_mux_ccr_out_n22), .Y(exu_n9096));
AND2X1 exu_U27136(.A(exu_tlu_ccr0_w[4]), .B(exu_n15935), .Y(ecl_ccr_mux_ccr_out_n24));
INVX1 exu_U27137(.A(ecl_ccr_mux_ccr_out_n24), .Y(exu_n9097));
AND2X1 exu_U27138(.A(exu_tlu_ccr2_w[3]), .B(exu_n15933), .Y(ecl_ccr_mux_ccr_out_n28));
INVX1 exu_U27139(.A(ecl_ccr_mux_ccr_out_n28), .Y(exu_n9098));
AND2X1 exu_U27140(.A(exu_tlu_ccr0_w[3]), .B(exu_n15935), .Y(ecl_ccr_mux_ccr_out_n30));
INVX1 exu_U27141(.A(ecl_ccr_mux_ccr_out_n30), .Y(exu_n9099));
AND2X1 exu_U27142(.A(exu_tlu_ccr2_w[2]), .B(exu_n15933), .Y(ecl_ccr_mux_ccr_out_n34));
INVX1 exu_U27143(.A(ecl_ccr_mux_ccr_out_n34), .Y(exu_n9100));
AND2X1 exu_U27144(.A(exu_tlu_ccr0_w[2]), .B(exu_n15935), .Y(ecl_ccr_mux_ccr_out_n36));
INVX1 exu_U27145(.A(ecl_ccr_mux_ccr_out_n36), .Y(exu_n9101));
AND2X1 exu_U27146(.A(exu_tlu_ccr2_w[1]), .B(exu_n15933), .Y(ecl_ccr_mux_ccr_out_n40));
INVX1 exu_U27147(.A(ecl_ccr_mux_ccr_out_n40), .Y(exu_n9102));
AND2X1 exu_U27148(.A(exu_tlu_ccr0_w[1]), .B(exu_n15935), .Y(ecl_ccr_mux_ccr_out_n42));
INVX1 exu_U27149(.A(ecl_ccr_mux_ccr_out_n42), .Y(exu_n9103));
AND2X1 exu_U27150(.A(exu_tlu_ccr2_w[0]), .B(exu_n15933), .Y(ecl_ccr_mux_ccr_out_n46));
INVX1 exu_U27151(.A(ecl_ccr_mux_ccr_out_n46), .Y(exu_n9104));
AND2X1 exu_U27152(.A(exu_tlu_ccr0_w[0]), .B(exu_n15935), .Y(ecl_ccr_mux_ccr_out_n48));
INVX1 exu_U27153(.A(ecl_ccr_mux_ccr_out_n48), .Y(exu_n9105));
AND2X1 exu_U27154(.A(ecl_ccr_wen_thr0_w), .B(exu_n15686), .Y(ecl_ccr_mux_ccrin0_n4));
INVX1 exu_U27155(.A(ecl_ccr_mux_ccrin0_n4), .Y(exu_n9106));
AND2X1 exu_U27156(.A(exu_n15702), .B(ecl_ccr_wen_thr0_w), .Y(ecl_ccr_mux_ccrin0_n8));
INVX1 exu_U27157(.A(ecl_ccr_mux_ccrin0_n8), .Y(exu_n9107));
AND2X1 exu_U27158(.A(exu_n15699), .B(ecl_ccr_wen_thr0_w), .Y(ecl_ccr_mux_ccrin0_n20));
INVX1 exu_U27159(.A(ecl_ccr_mux_ccrin0_n20), .Y(exu_n9108));
AND2X1 exu_U27160(.A(exu_n15698), .B(ecl_ccr_wen_thr0_w), .Y(ecl_ccr_mux_ccrin0_n24));
INVX1 exu_U27161(.A(ecl_ccr_mux_ccrin0_n24), .Y(exu_n9109));
AND2X1 exu_U27162(.A(exu_n15697), .B(ecl_ccr_wen_thr0_w), .Y(ecl_ccr_mux_ccrin0_n28));
INVX1 exu_U27163(.A(ecl_ccr_mux_ccrin0_n28), .Y(exu_n9110));
AND2X1 exu_U27164(.A(exu_n15696), .B(ecl_ccr_wen_thr0_w), .Y(ecl_ccr_mux_ccrin0_n32));
INVX1 exu_U27165(.A(ecl_ccr_mux_ccrin0_n32), .Y(exu_n9111));
AND2X1 exu_U27166(.A(rml_agp_thr[2]), .B(rml_agp_thr2[1]), .Y(rml_mux_agp_out1_n4));
INVX1 exu_U27167(.A(rml_mux_agp_out1_n4), .Y(exu_n9112));
AND2X1 exu_U27168(.A(exu_n15440), .B(rml_agp_thr0[1]), .Y(rml_mux_agp_out1_n6));
INVX1 exu_U27169(.A(rml_mux_agp_out1_n6), .Y(exu_n9113));
AND2X1 exu_U27170(.A(rml_agp_thr2[0]), .B(rml_agp_thr[2]), .Y(rml_mux_agp_out1_n10));
INVX1 exu_U27171(.A(rml_mux_agp_out1_n10), .Y(exu_n9114));
AND2X1 exu_U27172(.A(rml_agp_thr0[0]), .B(exu_n15440), .Y(rml_mux_agp_out1_n12));
INVX1 exu_U27173(.A(rml_mux_agp_out1_n12), .Y(exu_n9115));
AND2X1 exu_U27174(.A(exu_n11608), .B(exu_n10378), .Y(rml_cwp_swapping));
INVX1 exu_U27175(.A(rml_cwp_swapping), .Y(exu_n9116));
AND2X1 exu_U27176(.A(ecl_rml_thr_w[3]), .B(rml_cwp_n28), .Y(rml_cwp_n27));
INVX1 exu_U27177(.A(rml_cwp_n27), .Y(exu_n9117));
AND2X1 exu_U27178(.A(ecl_rml_thr_w[2]), .B(rml_cwp_n28), .Y(rml_cwp_n29));
INVX1 exu_U27179(.A(rml_cwp_n29), .Y(exu_n9118));
AND2X1 exu_U27180(.A(exu_n15957), .B(rml_cwp_n28), .Y(rml_cwp_n30));
INVX1 exu_U27181(.A(rml_cwp_n30), .Y(exu_n9119));
AND2X1 exu_U27182(.A(exu_n15959), .B(rml_cwp_n28), .Y(rml_cwp_n31));
INVX1 exu_U27183(.A(rml_cwp_n31), .Y(exu_n9120));
AND2X1 exu_U27184(.A(rml_cwp_swap_thr[0]), .B(rml_cwp_N99), .Y(rml_cwp_n46));
INVX1 exu_U27185(.A(rml_cwp_n46), .Y(exu_n9121));
OR2X1 exu_U27186(.A(rml_cwp_n88), .B(rml_cwp_n89), .Y(rml_cwp_n66));
INVX1 exu_U27187(.A(rml_cwp_n66), .Y(exu_n9122));
OR2X1 exu_U27188(.A(rml_cwp_n85), .B(rml_cwp_n86), .Y(rml_cwp_n68));
INVX1 exu_U27189(.A(rml_cwp_n68), .Y(exu_n9123));
OR2X1 exu_U27190(.A(rml_cwp_n82), .B(rml_cwp_n83), .Y(rml_cwp_n70));
INVX1 exu_U27191(.A(rml_cwp_n70), .Y(exu_n9124));
OR2X1 exu_U27192(.A(rml_cwp_n79), .B(rml_cwp_n80), .Y(rml_cwp_n72));
INVX1 exu_U27193(.A(rml_cwp_n72), .Y(exu_n9125));
OR2X1 exu_U27194(.A(rml_cwp_just_swapped), .B(rml_cwp_n104), .Y(rml_cwp_n103));
INVX1 exu_U27195(.A(rml_cwp_n103), .Y(exu_n9126));
AND2X1 exu_U27196(.A(exu_n15940), .B(rml_spill_cwp_e[2]), .Y(rml_next_cwp_mux_n2));
INVX1 exu_U27197(.A(rml_next_cwp_mux_n2), .Y(exu_n9127));
AND2X1 exu_U27198(.A(rml_full_swap_e), .B(rml_rml_next_cwp_e[2]), .Y(rml_next_cwp_mux_n4));
INVX1 exu_U27199(.A(rml_next_cwp_mux_n4), .Y(exu_n9128));
AND2X1 exu_U27200(.A(rml_spill_cwp_e[1]), .B(exu_n15940), .Y(rml_next_cwp_mux_n6));
INVX1 exu_U27201(.A(rml_next_cwp_mux_n6), .Y(exu_n9129));
AND2X1 exu_U27202(.A(rml_rml_next_cwp_e[1]), .B(rml_full_swap_e), .Y(rml_next_cwp_mux_n8));
INVX1 exu_U27203(.A(rml_next_cwp_mux_n8), .Y(exu_n9130));
AND2X1 exu_U27204(.A(rml_spill_cwp_e[0]), .B(exu_n15940), .Y(rml_next_cwp_mux_n10));
INVX1 exu_U27205(.A(rml_next_cwp_mux_n10), .Y(exu_n9131));
AND2X1 exu_U27206(.A(exu_n16569), .B(rml_full_swap_e), .Y(rml_next_cwp_mux_n12));
INVX1 exu_U27207(.A(rml_next_cwp_mux_n12), .Y(exu_n9132));
AND2X1 exu_U27208(.A(rml_save_e), .B(rml_cwp_inc_n6), .Y(rml_cwp_inc_n5));
INVX1 exu_U27209(.A(rml_cwp_inc_n5), .Y(exu_n9133));
AND2X1 exu_U27210(.A(exu_n16259), .B(div_out64[9]), .Y(div_d_mux_n4));
INVX1 exu_U27211(.A(div_d_mux_n4), .Y(exu_n9134));
AND2X1 exu_U27212(.A(div_curr_q[35]), .B(exu_n16259), .Y(div_d_mux_n8));
INVX1 exu_U27213(.A(div_d_mux_n8), .Y(exu_n9135));
AND2X1 exu_U27214(.A(div_curr_q[34]), .B(exu_n16258), .Y(div_d_mux_n12));
INVX1 exu_U27215(.A(div_d_mux_n12), .Y(exu_n9136));
AND2X1 exu_U27216(.A(div_curr_q[33]), .B(exu_n16259), .Y(div_d_mux_n16));
INVX1 exu_U27217(.A(div_d_mux_n16), .Y(exu_n9137));
AND2X1 exu_U27218(.A(div_curr_q[32]), .B(exu_n16258), .Y(div_d_mux_n20));
INVX1 exu_U27219(.A(div_d_mux_n20), .Y(exu_n9138));
AND2X1 exu_U27220(.A(div_curr_q[31]), .B(exu_n16258), .Y(div_d_mux_n24));
INVX1 exu_U27221(.A(div_d_mux_n24), .Y(exu_n9139));
AND2X1 exu_U27222(.A(div_curr_q[30]), .B(exu_n16259), .Y(div_d_mux_n28));
INVX1 exu_U27223(.A(div_d_mux_n28), .Y(exu_n9140));
AND2X1 exu_U27224(.A(div_curr_q[29]), .B(exu_n16259), .Y(div_d_mux_n32));
INVX1 exu_U27225(.A(div_d_mux_n32), .Y(exu_n9141));
AND2X1 exu_U27226(.A(div_curr_q[28]), .B(exu_n16259), .Y(div_d_mux_n36));
INVX1 exu_U27227(.A(div_d_mux_n36), .Y(exu_n9142));
AND2X1 exu_U27228(.A(div_curr_q[27]), .B(exu_n16259), .Y(div_d_mux_n40));
INVX1 exu_U27229(.A(div_d_mux_n40), .Y(exu_n9143));
AND2X1 exu_U27230(.A(div_curr_q[26]), .B(exu_n16258), .Y(div_d_mux_n44));
INVX1 exu_U27231(.A(div_d_mux_n44), .Y(exu_n9144));
AND2X1 exu_U27232(.A(div_out64[8]), .B(exu_n16258), .Y(div_d_mux_n48));
INVX1 exu_U27233(.A(div_d_mux_n48), .Y(exu_n9145));
AND2X1 exu_U27234(.A(div_curr_q[25]), .B(exu_n16259), .Y(div_d_mux_n52));
INVX1 exu_U27235(.A(div_d_mux_n52), .Y(exu_n9146));
AND2X1 exu_U27236(.A(div_curr_q[24]), .B(exu_n16259), .Y(div_d_mux_n56));
INVX1 exu_U27237(.A(div_d_mux_n56), .Y(exu_n9147));
AND2X1 exu_U27238(.A(div_curr_q[23]), .B(exu_n16259), .Y(div_d_mux_n60));
INVX1 exu_U27239(.A(div_d_mux_n60), .Y(exu_n9148));
AND2X1 exu_U27240(.A(div_curr_q[22]), .B(exu_n16258), .Y(div_d_mux_n64));
INVX1 exu_U27241(.A(div_d_mux_n64), .Y(exu_n9149));
AND2X1 exu_U27242(.A(div_curr_q[21]), .B(exu_n16258), .Y(div_d_mux_n68));
INVX1 exu_U27243(.A(div_d_mux_n68), .Y(exu_n9150));
AND2X1 exu_U27244(.A(div_curr_q[20]), .B(exu_n16258), .Y(div_d_mux_n72));
INVX1 exu_U27245(.A(div_d_mux_n72), .Y(exu_n9151));
AND2X1 exu_U27246(.A(div_curr_q[19]), .B(exu_n16259), .Y(div_d_mux_n76));
INVX1 exu_U27247(.A(div_d_mux_n76), .Y(exu_n9152));
AND2X1 exu_U27248(.A(div_curr_q[18]), .B(exu_n16259), .Y(div_d_mux_n80));
INVX1 exu_U27249(.A(div_d_mux_n80), .Y(exu_n9153));
AND2X1 exu_U27250(.A(div_curr_q[17]), .B(exu_n16258), .Y(div_d_mux_n84));
INVX1 exu_U27251(.A(div_d_mux_n84), .Y(exu_n9154));
AND2X1 exu_U27252(.A(div_curr_q[16]), .B(exu_n16259), .Y(div_d_mux_n88));
INVX1 exu_U27253(.A(div_d_mux_n88), .Y(exu_n9155));
AND2X1 exu_U27254(.A(div_out64[7]), .B(exu_n16259), .Y(div_d_mux_n92));
INVX1 exu_U27255(.A(div_d_mux_n92), .Y(exu_n9156));
AND2X1 exu_U27256(.A(div_curr_q[15]), .B(exu_n16258), .Y(div_d_mux_n96));
INVX1 exu_U27257(.A(div_d_mux_n96), .Y(exu_n9157));
AND2X1 exu_U27258(.A(div_curr_q[14]), .B(exu_n16259), .Y(div_d_mux_n100));
INVX1 exu_U27259(.A(div_d_mux_n100), .Y(exu_n9158));
AND2X1 exu_U27260(.A(div_curr_q[13]), .B(exu_n16258), .Y(div_d_mux_n104));
INVX1 exu_U27261(.A(div_d_mux_n104), .Y(exu_n9159));
AND2X1 exu_U27262(.A(div_curr_q[12]), .B(exu_n16258), .Y(div_d_mux_n108));
INVX1 exu_U27263(.A(div_d_mux_n108), .Y(exu_n9160));
AND2X1 exu_U27264(.A(div_curr_q[11]), .B(exu_n16258), .Y(div_d_mux_n112));
INVX1 exu_U27265(.A(div_d_mux_n112), .Y(exu_n9161));
AND2X1 exu_U27266(.A(div_curr_q[10]), .B(exu_n16258), .Y(div_d_mux_n116));
INVX1 exu_U27267(.A(div_d_mux_n116), .Y(exu_n9162));
AND2X1 exu_U27268(.A(div_curr_q[9]), .B(exu_n16259), .Y(div_d_mux_n120));
INVX1 exu_U27269(.A(div_d_mux_n120), .Y(exu_n9163));
AND2X1 exu_U27270(.A(div_curr_q[8]), .B(exu_n16259), .Y(div_d_mux_n124));
INVX1 exu_U27271(.A(div_d_mux_n124), .Y(exu_n9164));
AND2X1 exu_U27272(.A(div_curr_q[7]), .B(exu_n16258), .Y(div_d_mux_n128));
INVX1 exu_U27273(.A(div_d_mux_n128), .Y(exu_n9165));
AND2X1 exu_U27274(.A(div_curr_q[6]), .B(exu_n16258), .Y(div_d_mux_n132));
INVX1 exu_U27275(.A(div_d_mux_n132), .Y(exu_n9166));
AND2X1 exu_U27276(.A(div_out64[6]), .B(exu_n16259), .Y(div_d_mux_n136));
INVX1 exu_U27277(.A(div_d_mux_n136), .Y(exu_n9167));
AND2X1 exu_U27278(.A(div_curr_q[5]), .B(exu_n16259), .Y(div_d_mux_n140));
INVX1 exu_U27279(.A(div_d_mux_n140), .Y(exu_n9168));
AND2X1 exu_U27280(.A(div_curr_q[4]), .B(exu_n16259), .Y(div_d_mux_n144));
INVX1 exu_U27281(.A(div_d_mux_n144), .Y(exu_n9169));
AND2X1 exu_U27282(.A(div_curr_q[3]), .B(exu_n16259), .Y(div_d_mux_n148));
INVX1 exu_U27283(.A(div_d_mux_n148), .Y(exu_n9170));
AND2X1 exu_U27284(.A(div_curr_q[2]), .B(exu_n16258), .Y(div_d_mux_n152));
INVX1 exu_U27285(.A(div_d_mux_n152), .Y(exu_n9171));
AND2X1 exu_U27286(.A(div_curr_q[1]), .B(exu_n16258), .Y(div_d_mux_n156));
INVX1 exu_U27287(.A(div_d_mux_n156), .Y(exu_n9172));
AND2X1 exu_U27288(.A(div_curr_q[0]), .B(exu_n16259), .Y(div_d_mux_n160));
INVX1 exu_U27289(.A(div_d_mux_n160), .Y(exu_n9173));
AND2X1 exu_U27290(.A(div_out64[63]), .B(exu_n16258), .Y(div_d_mux_n164));
INVX1 exu_U27291(.A(div_d_mux_n164), .Y(exu_n9174));
AND2X1 exu_U27292(.A(div_out64[62]), .B(exu_n16258), .Y(div_d_mux_n168));
INVX1 exu_U27293(.A(div_d_mux_n168), .Y(exu_n9175));
AND2X1 exu_U27294(.A(div_out64[61]), .B(exu_n16258), .Y(div_d_mux_n172));
INVX1 exu_U27295(.A(div_d_mux_n172), .Y(exu_n9176));
AND2X1 exu_U27296(.A(div_out64[60]), .B(exu_n16258), .Y(div_d_mux_n176));
INVX1 exu_U27297(.A(div_d_mux_n176), .Y(exu_n9177));
AND2X1 exu_U27298(.A(div_out64[5]), .B(exu_n16259), .Y(div_d_mux_n180));
INVX1 exu_U27299(.A(div_d_mux_n180), .Y(exu_n9178));
AND2X1 exu_U27300(.A(div_out64[59]), .B(exu_n16259), .Y(div_d_mux_n184));
INVX1 exu_U27301(.A(div_d_mux_n184), .Y(exu_n9179));
AND2X1 exu_U27302(.A(div_out64[58]), .B(exu_n16259), .Y(div_d_mux_n188));
INVX1 exu_U27303(.A(div_d_mux_n188), .Y(exu_n9180));
AND2X1 exu_U27304(.A(div_out64[57]), .B(exu_n16258), .Y(div_d_mux_n192));
INVX1 exu_U27305(.A(div_d_mux_n192), .Y(exu_n9181));
AND2X1 exu_U27306(.A(div_out64[56]), .B(exu_n16259), .Y(div_d_mux_n196));
INVX1 exu_U27307(.A(div_d_mux_n196), .Y(exu_n9182));
AND2X1 exu_U27308(.A(div_out64[55]), .B(exu_n16259), .Y(div_d_mux_n200));
INVX1 exu_U27309(.A(div_d_mux_n200), .Y(exu_n9183));
AND2X1 exu_U27310(.A(div_out64[54]), .B(exu_n16258), .Y(div_d_mux_n204));
INVX1 exu_U27311(.A(div_d_mux_n204), .Y(exu_n9184));
AND2X1 exu_U27312(.A(div_out64[53]), .B(exu_n16259), .Y(div_d_mux_n208));
INVX1 exu_U27313(.A(div_d_mux_n208), .Y(exu_n9185));
AND2X1 exu_U27314(.A(div_out64[52]), .B(exu_n16258), .Y(div_d_mux_n212));
INVX1 exu_U27315(.A(div_d_mux_n212), .Y(exu_n9186));
AND2X1 exu_U27316(.A(div_out64[51]), .B(exu_n16258), .Y(div_d_mux_n216));
INVX1 exu_U27317(.A(div_d_mux_n216), .Y(exu_n9187));
AND2X1 exu_U27318(.A(div_out64[50]), .B(exu_n16258), .Y(div_d_mux_n220));
INVX1 exu_U27319(.A(div_d_mux_n220), .Y(exu_n9188));
AND2X1 exu_U27320(.A(div_out64[4]), .B(exu_n16258), .Y(div_d_mux_n224));
INVX1 exu_U27321(.A(div_d_mux_n224), .Y(exu_n9189));
AND2X1 exu_U27322(.A(div_out64[49]), .B(exu_n16258), .Y(div_d_mux_n228));
INVX1 exu_U27323(.A(div_d_mux_n228), .Y(exu_n9190));
AND2X1 exu_U27324(.A(div_out64[48]), .B(exu_n16258), .Y(div_d_mux_n232));
INVX1 exu_U27325(.A(div_d_mux_n232), .Y(exu_n9191));
AND2X1 exu_U27326(.A(div_out64[47]), .B(exu_n16258), .Y(div_d_mux_n236));
INVX1 exu_U27327(.A(div_d_mux_n236), .Y(exu_n9192));
AND2X1 exu_U27328(.A(div_out64[46]), .B(exu_n16258), .Y(div_d_mux_n240));
INVX1 exu_U27329(.A(div_d_mux_n240), .Y(exu_n9193));
AND2X1 exu_U27330(.A(div_out64[45]), .B(exu_n16258), .Y(div_d_mux_n244));
INVX1 exu_U27331(.A(div_d_mux_n244), .Y(exu_n9194));
AND2X1 exu_U27332(.A(div_out64[44]), .B(exu_n16258), .Y(div_d_mux_n248));
INVX1 exu_U27333(.A(div_d_mux_n248), .Y(exu_n9195));
AND2X1 exu_U27334(.A(div_out64[43]), .B(exu_n16258), .Y(div_d_mux_n252));
INVX1 exu_U27335(.A(div_d_mux_n252), .Y(exu_n9196));
AND2X1 exu_U27336(.A(div_out64[42]), .B(exu_n16258), .Y(div_d_mux_n256));
INVX1 exu_U27337(.A(div_d_mux_n256), .Y(exu_n9197));
AND2X1 exu_U27338(.A(div_out64[41]), .B(exu_n16258), .Y(div_d_mux_n260));
INVX1 exu_U27339(.A(div_d_mux_n260), .Y(exu_n9198));
AND2X1 exu_U27340(.A(div_out64[40]), .B(exu_n16259), .Y(div_d_mux_n264));
INVX1 exu_U27341(.A(div_d_mux_n264), .Y(exu_n9199));
AND2X1 exu_U27342(.A(div_out64[3]), .B(exu_n16258), .Y(div_d_mux_n268));
INVX1 exu_U27343(.A(div_d_mux_n268), .Y(exu_n9200));
AND2X1 exu_U27344(.A(div_out64[39]), .B(exu_n16259), .Y(div_d_mux_n272));
INVX1 exu_U27345(.A(div_d_mux_n272), .Y(exu_n9201));
AND2X1 exu_U27346(.A(div_out64[38]), .B(exu_n16259), .Y(div_d_mux_n276));
INVX1 exu_U27347(.A(div_d_mux_n276), .Y(exu_n9202));
AND2X1 exu_U27348(.A(div_out64[37]), .B(exu_n16259), .Y(div_d_mux_n280));
INVX1 exu_U27349(.A(div_d_mux_n280), .Y(exu_n9203));
AND2X1 exu_U27350(.A(div_out64[36]), .B(exu_n16259), .Y(div_d_mux_n284));
INVX1 exu_U27351(.A(div_d_mux_n284), .Y(exu_n9204));
AND2X1 exu_U27352(.A(div_out64[35]), .B(exu_n16258), .Y(div_d_mux_n288));
INVX1 exu_U27353(.A(div_d_mux_n288), .Y(exu_n9205));
AND2X1 exu_U27354(.A(div_out64[34]), .B(exu_n16258), .Y(div_d_mux_n292));
INVX1 exu_U27355(.A(div_d_mux_n292), .Y(exu_n9206));
AND2X1 exu_U27356(.A(div_out64[33]), .B(exu_n16259), .Y(div_d_mux_n296));
INVX1 exu_U27357(.A(div_d_mux_n296), .Y(exu_n9207));
AND2X1 exu_U27358(.A(div_out64[32]), .B(exu_n16259), .Y(div_d_mux_n300));
INVX1 exu_U27359(.A(div_d_mux_n300), .Y(exu_n9208));
AND2X1 exu_U27360(.A(div_out64[31]), .B(exu_n16258), .Y(div_d_mux_n304));
INVX1 exu_U27361(.A(div_d_mux_n304), .Y(exu_n9209));
AND2X1 exu_U27362(.A(div_out64[30]), .B(exu_n16258), .Y(div_d_mux_n308));
INVX1 exu_U27363(.A(div_d_mux_n308), .Y(exu_n9210));
AND2X1 exu_U27364(.A(div_out64[2]), .B(exu_n16258), .Y(div_d_mux_n312));
INVX1 exu_U27365(.A(div_d_mux_n312), .Y(exu_n9211));
AND2X1 exu_U27366(.A(div_out64[29]), .B(exu_n16258), .Y(div_d_mux_n316));
INVX1 exu_U27367(.A(div_d_mux_n316), .Y(exu_n9212));
AND2X1 exu_U27368(.A(div_out64[28]), .B(exu_n16258), .Y(div_d_mux_n320));
INVX1 exu_U27369(.A(div_d_mux_n320), .Y(exu_n9213));
AND2X1 exu_U27370(.A(div_out64[27]), .B(exu_n16259), .Y(div_d_mux_n324));
INVX1 exu_U27371(.A(div_d_mux_n324), .Y(exu_n9214));
AND2X1 exu_U27372(.A(div_out64[26]), .B(exu_n16259), .Y(div_d_mux_n328));
INVX1 exu_U27373(.A(div_d_mux_n328), .Y(exu_n9215));
AND2X1 exu_U27374(.A(div_out64[25]), .B(exu_n16259), .Y(div_d_mux_n332));
INVX1 exu_U27375(.A(div_d_mux_n332), .Y(exu_n9216));
AND2X1 exu_U27376(.A(div_out64[24]), .B(exu_n16259), .Y(div_d_mux_n336));
INVX1 exu_U27377(.A(div_d_mux_n336), .Y(exu_n9217));
AND2X1 exu_U27378(.A(div_out64[23]), .B(exu_n16258), .Y(div_d_mux_n340));
INVX1 exu_U27379(.A(div_d_mux_n340), .Y(exu_n9218));
AND2X1 exu_U27380(.A(div_out64[22]), .B(exu_n16259), .Y(div_d_mux_n344));
INVX1 exu_U27381(.A(div_d_mux_n344), .Y(exu_n9219));
AND2X1 exu_U27382(.A(div_out64[21]), .B(exu_n16259), .Y(div_d_mux_n348));
INVX1 exu_U27383(.A(div_d_mux_n348), .Y(exu_n9220));
AND2X1 exu_U27384(.A(div_out64[20]), .B(exu_n16259), .Y(div_d_mux_n352));
INVX1 exu_U27385(.A(div_d_mux_n352), .Y(exu_n9221));
AND2X1 exu_U27386(.A(div_out64[1]), .B(exu_n16259), .Y(div_d_mux_n356));
INVX1 exu_U27387(.A(div_d_mux_n356), .Y(exu_n9222));
AND2X1 exu_U27388(.A(div_out64[19]), .B(exu_n16259), .Y(div_d_mux_n360));
INVX1 exu_U27389(.A(div_d_mux_n360), .Y(exu_n9223));
AND2X1 exu_U27390(.A(div_out64[18]), .B(exu_n16259), .Y(div_d_mux_n364));
INVX1 exu_U27391(.A(div_d_mux_n364), .Y(exu_n9224));
AND2X1 exu_U27392(.A(div_out64[17]), .B(exu_n16258), .Y(div_d_mux_n368));
INVX1 exu_U27393(.A(div_d_mux_n368), .Y(exu_n9225));
AND2X1 exu_U27394(.A(div_out64[16]), .B(exu_n16258), .Y(div_d_mux_n372));
INVX1 exu_U27395(.A(div_d_mux_n372), .Y(exu_n9226));
AND2X1 exu_U27396(.A(div_out64[15]), .B(exu_n16258), .Y(div_d_mux_n376));
INVX1 exu_U27397(.A(div_d_mux_n376), .Y(exu_n9227));
AND2X1 exu_U27398(.A(div_out64[14]), .B(exu_n16259), .Y(div_d_mux_n380));
INVX1 exu_U27399(.A(div_d_mux_n380), .Y(exu_n9228));
AND2X1 exu_U27400(.A(div_out64[13]), .B(exu_n16259), .Y(div_d_mux_n384));
INVX1 exu_U27401(.A(div_d_mux_n384), .Y(exu_n9229));
AND2X1 exu_U27402(.A(div_out64[12]), .B(exu_n16259), .Y(div_d_mux_n388));
INVX1 exu_U27403(.A(div_d_mux_n388), .Y(exu_n9230));
AND2X1 exu_U27404(.A(div_ecl_d_msb), .B(exu_n16258), .Y(div_d_mux_n392));
INVX1 exu_U27405(.A(div_d_mux_n392), .Y(exu_n9231));
AND2X1 exu_U27406(.A(div_curr_q[62]), .B(exu_n16259), .Y(div_d_mux_n396));
INVX1 exu_U27407(.A(div_d_mux_n396), .Y(exu_n9232));
AND2X1 exu_U27408(.A(div_curr_q[61]), .B(exu_n16258), .Y(div_d_mux_n400));
INVX1 exu_U27409(.A(div_d_mux_n400), .Y(exu_n9233));
AND2X1 exu_U27410(.A(div_curr_q[60]), .B(exu_n16258), .Y(div_d_mux_n404));
INVX1 exu_U27411(.A(div_d_mux_n404), .Y(exu_n9234));
AND2X1 exu_U27412(.A(div_curr_q[59]), .B(exu_n16258), .Y(div_d_mux_n408));
INVX1 exu_U27413(.A(div_d_mux_n408), .Y(exu_n9235));
AND2X1 exu_U27414(.A(div_curr_q[58]), .B(exu_n16259), .Y(div_d_mux_n412));
INVX1 exu_U27415(.A(div_d_mux_n412), .Y(exu_n9236));
AND2X1 exu_U27416(.A(div_curr_q[57]), .B(exu_n16259), .Y(div_d_mux_n416));
INVX1 exu_U27417(.A(div_d_mux_n416), .Y(exu_n9237));
AND2X1 exu_U27418(.A(div_curr_q[56]), .B(exu_n16259), .Y(div_d_mux_n420));
INVX1 exu_U27419(.A(div_d_mux_n420), .Y(exu_n9238));
AND2X1 exu_U27420(.A(div_out64[11]), .B(exu_n16259), .Y(div_d_mux_n424));
INVX1 exu_U27421(.A(div_d_mux_n424), .Y(exu_n9239));
AND2X1 exu_U27422(.A(div_curr_q[55]), .B(exu_n16259), .Y(div_d_mux_n428));
INVX1 exu_U27423(.A(div_d_mux_n428), .Y(exu_n9240));
AND2X1 exu_U27424(.A(div_curr_q[54]), .B(exu_n16258), .Y(div_d_mux_n432));
INVX1 exu_U27425(.A(div_d_mux_n432), .Y(exu_n9241));
AND2X1 exu_U27426(.A(div_curr_q[53]), .B(exu_n16259), .Y(div_d_mux_n436));
INVX1 exu_U27427(.A(div_d_mux_n436), .Y(exu_n9242));
AND2X1 exu_U27428(.A(div_curr_q[52]), .B(exu_n16259), .Y(div_d_mux_n440));
INVX1 exu_U27429(.A(div_d_mux_n440), .Y(exu_n9243));
AND2X1 exu_U27430(.A(div_curr_q[51]), .B(exu_n16259), .Y(div_d_mux_n444));
INVX1 exu_U27431(.A(div_d_mux_n444), .Y(exu_n9244));
AND2X1 exu_U27432(.A(div_curr_q[50]), .B(exu_n16258), .Y(div_d_mux_n448));
INVX1 exu_U27433(.A(div_d_mux_n448), .Y(exu_n9245));
AND2X1 exu_U27434(.A(div_curr_q[49]), .B(exu_n16258), .Y(div_d_mux_n452));
INVX1 exu_U27435(.A(div_d_mux_n452), .Y(exu_n9246));
AND2X1 exu_U27436(.A(div_curr_q[48]), .B(exu_n16258), .Y(div_d_mux_n456));
INVX1 exu_U27437(.A(div_d_mux_n456), .Y(exu_n9247));
AND2X1 exu_U27438(.A(div_curr_q[47]), .B(exu_n16258), .Y(div_d_mux_n460));
INVX1 exu_U27439(.A(div_d_mux_n460), .Y(exu_n9248));
AND2X1 exu_U27440(.A(div_curr_q[46]), .B(exu_n16259), .Y(div_d_mux_n464));
INVX1 exu_U27441(.A(div_d_mux_n464), .Y(exu_n9249));
AND2X1 exu_U27442(.A(div_out64[10]), .B(exu_n16259), .Y(div_d_mux_n468));
INVX1 exu_U27443(.A(div_d_mux_n468), .Y(exu_n9250));
AND2X1 exu_U27444(.A(div_curr_q[45]), .B(exu_n16258), .Y(div_d_mux_n472));
INVX1 exu_U27445(.A(div_d_mux_n472), .Y(exu_n9251));
AND2X1 exu_U27446(.A(div_curr_q[44]), .B(exu_n16259), .Y(div_d_mux_n476));
INVX1 exu_U27447(.A(div_d_mux_n476), .Y(exu_n9252));
AND2X1 exu_U27448(.A(div_curr_q[43]), .B(exu_n16259), .Y(div_d_mux_n480));
INVX1 exu_U27449(.A(div_d_mux_n480), .Y(exu_n9253));
AND2X1 exu_U27450(.A(div_curr_q[42]), .B(exu_n16258), .Y(div_d_mux_n484));
INVX1 exu_U27451(.A(div_d_mux_n484), .Y(exu_n9254));
AND2X1 exu_U27452(.A(div_curr_q[41]), .B(exu_n16259), .Y(div_d_mux_n488));
INVX1 exu_U27453(.A(div_d_mux_n488), .Y(exu_n9255));
AND2X1 exu_U27454(.A(div_curr_q[40]), .B(exu_n16259), .Y(div_d_mux_n492));
INVX1 exu_U27455(.A(div_d_mux_n492), .Y(exu_n9256));
AND2X1 exu_U27456(.A(div_curr_q[39]), .B(exu_n16258), .Y(div_d_mux_n496));
INVX1 exu_U27457(.A(div_d_mux_n496), .Y(exu_n9257));
AND2X1 exu_U27458(.A(div_curr_q[38]), .B(exu_n16258), .Y(div_d_mux_n500));
INVX1 exu_U27459(.A(div_d_mux_n500), .Y(exu_n9258));
AND2X1 exu_U27460(.A(div_curr_q[37]), .B(exu_n16259), .Y(div_d_mux_n504));
INVX1 exu_U27461(.A(div_d_mux_n504), .Y(exu_n9259));
AND2X1 exu_U27462(.A(div_curr_q[36]), .B(exu_n16258), .Y(div_d_mux_n508));
INVX1 exu_U27463(.A(div_d_mux_n508), .Y(exu_n9260));
AND2X1 exu_U27464(.A(div_out64[0]), .B(exu_n16258), .Y(div_d_mux_n512));
INVX1 exu_U27465(.A(div_d_mux_n512), .Y(exu_n9261));
OR2X1 exu_U27466(.A(exu_n12056), .B(exu_n14950), .Y(div_low32or_n4));
INVX1 exu_U27467(.A(div_low32or_n4), .Y(exu_n9262));
OR2X1 exu_U27468(.A(exu_n12001), .B(exu_n14889), .Y(div_low32or_n8));
INVX1 exu_U27469(.A(div_low32or_n8), .Y(exu_n9263));
OR2X1 exu_U27470(.A(exu_n11999), .B(exu_n14887), .Y(div_low32or_n10));
INVX1 exu_U27471(.A(div_low32or_n10), .Y(exu_n9264));
OR2X1 exu_U27472(.A(exu_n12005), .B(exu_n14893), .Y(div_low32or_n14));
INVX1 exu_U27473(.A(div_low32or_n14), .Y(exu_n9265));
OR2X1 exu_U27474(.A(exu_n12003), .B(exu_n14891), .Y(div_low32or_n16));
INVX1 exu_U27475(.A(div_low32or_n16), .Y(exu_n9266));
OR2X1 exu_U27476(.A(exu_n12058), .B(exu_n14952), .Y(div_low32or_n18));
INVX1 exu_U27477(.A(div_low32or_n18), .Y(exu_n9267));
OR2X1 exu_U27478(.A(exu_n11993), .B(exu_n14882), .Y(div_low32or_n22));
INVX1 exu_U27479(.A(div_low32or_n22), .Y(exu_n9268));
OR2X1 exu_U27480(.A(exu_n11991), .B(exu_n14880), .Y(div_low32or_n24));
INVX1 exu_U27481(.A(div_low32or_n24), .Y(exu_n9269));
OR2X1 exu_U27482(.A(exu_n11997), .B(exu_n14885), .Y(div_low32or_n28));
INVX1 exu_U27483(.A(div_low32or_n28), .Y(exu_n9270));
OR2X1 exu_U27484(.A(exu_n11995), .B(exu_n14883), .Y(div_low32or_n30));
INVX1 exu_U27485(.A(div_low32or_n30), .Y(exu_n9271));
AND2X1 exu_U27486(.A(alu_logic_rs1_data_bf1[41]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n3));
INVX1 exu_U27487(.A(shft_mux_rshift_extend_n3), .Y(exu_n9272));
AND2X1 exu_U27488(.A(alu_logic_rs1_data_bf1[40]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n5));
INVX1 exu_U27489(.A(shft_mux_rshift_extend_n5), .Y(exu_n9273));
AND2X1 exu_U27490(.A(alu_logic_rs1_data_bf1[39]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n7));
INVX1 exu_U27491(.A(shft_mux_rshift_extend_n7), .Y(exu_n9274));
AND2X1 exu_U27492(.A(alu_logic_rs1_data_bf1[38]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n9));
INVX1 exu_U27493(.A(shft_mux_rshift_extend_n9), .Y(exu_n9275));
AND2X1 exu_U27494(.A(alu_logic_rs1_data_bf1[37]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n11));
INVX1 exu_U27495(.A(shft_mux_rshift_extend_n11), .Y(exu_n9276));
AND2X1 exu_U27496(.A(alu_logic_rs1_data_bf1[36]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n13));
INVX1 exu_U27497(.A(shft_mux_rshift_extend_n13), .Y(exu_n9277));
AND2X1 exu_U27498(.A(alu_logic_rs1_data_bf1[35]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n15));
INVX1 exu_U27499(.A(shft_mux_rshift_extend_n15), .Y(exu_n9278));
AND2X1 exu_U27500(.A(alu_logic_rs1_data_bf1[63]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n17));
INVX1 exu_U27501(.A(shft_mux_rshift_extend_n17), .Y(exu_n9279));
AND2X1 exu_U27502(.A(alu_logic_rs1_data_bf1[62]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n19));
INVX1 exu_U27503(.A(shft_mux_rshift_extend_n19), .Y(exu_n9280));
AND2X1 exu_U27504(.A(alu_logic_rs1_data_bf1[34]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n21));
INVX1 exu_U27505(.A(shft_mux_rshift_extend_n21), .Y(exu_n9281));
AND2X1 exu_U27506(.A(alu_logic_rs1_data_bf1[61]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n23));
INVX1 exu_U27507(.A(shft_mux_rshift_extend_n23), .Y(exu_n9282));
AND2X1 exu_U27508(.A(alu_logic_rs1_data_bf1[60]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n25));
INVX1 exu_U27509(.A(shft_mux_rshift_extend_n25), .Y(exu_n9283));
AND2X1 exu_U27510(.A(alu_logic_rs1_data_bf1[59]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n27));
INVX1 exu_U27511(.A(shft_mux_rshift_extend_n27), .Y(exu_n9284));
AND2X1 exu_U27512(.A(alu_logic_rs1_data_bf1[58]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n29));
INVX1 exu_U27513(.A(shft_mux_rshift_extend_n29), .Y(exu_n9285));
AND2X1 exu_U27514(.A(alu_logic_rs1_data_bf1[57]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n31));
INVX1 exu_U27515(.A(shft_mux_rshift_extend_n31), .Y(exu_n9286));
AND2X1 exu_U27516(.A(alu_logic_rs1_data_bf1[56]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n33));
INVX1 exu_U27517(.A(shft_mux_rshift_extend_n33), .Y(exu_n9287));
AND2X1 exu_U27518(.A(alu_logic_rs1_data_bf1[55]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n35));
INVX1 exu_U27519(.A(shft_mux_rshift_extend_n35), .Y(exu_n9288));
AND2X1 exu_U27520(.A(alu_logic_rs1_data_bf1[54]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n37));
INVX1 exu_U27521(.A(shft_mux_rshift_extend_n37), .Y(exu_n9289));
AND2X1 exu_U27522(.A(alu_logic_rs1_data_bf1[53]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n39));
INVX1 exu_U27523(.A(shft_mux_rshift_extend_n39), .Y(exu_n9290));
AND2X1 exu_U27524(.A(alu_logic_rs1_data_bf1[52]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n41));
INVX1 exu_U27525(.A(shft_mux_rshift_extend_n41), .Y(exu_n9291));
AND2X1 exu_U27526(.A(alu_logic_rs1_data_bf1[33]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n43));
INVX1 exu_U27527(.A(shft_mux_rshift_extend_n43), .Y(exu_n9292));
AND2X1 exu_U27528(.A(alu_logic_rs1_data_bf1[51]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n45));
INVX1 exu_U27529(.A(shft_mux_rshift_extend_n45), .Y(exu_n9293));
AND2X1 exu_U27530(.A(alu_logic_rs1_data_bf1[50]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n47));
INVX1 exu_U27531(.A(shft_mux_rshift_extend_n47), .Y(exu_n9294));
AND2X1 exu_U27532(.A(alu_logic_rs1_data_bf1[49]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n49));
INVX1 exu_U27533(.A(shft_mux_rshift_extend_n49), .Y(exu_n9295));
AND2X1 exu_U27534(.A(alu_logic_rs1_data_bf1[48]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n51));
INVX1 exu_U27535(.A(shft_mux_rshift_extend_n51), .Y(exu_n9296));
AND2X1 exu_U27536(.A(alu_logic_rs1_data_bf1[47]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n53));
INVX1 exu_U27537(.A(shft_mux_rshift_extend_n53), .Y(exu_n9297));
AND2X1 exu_U27538(.A(alu_logic_rs1_data_bf1[46]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n55));
INVX1 exu_U27539(.A(shft_mux_rshift_extend_n55), .Y(exu_n9298));
AND2X1 exu_U27540(.A(alu_logic_rs1_data_bf1[45]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n57));
INVX1 exu_U27541(.A(shft_mux_rshift_extend_n57), .Y(exu_n9299));
AND2X1 exu_U27542(.A(alu_logic_rs1_data_bf1[44]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n59));
INVX1 exu_U27543(.A(shft_mux_rshift_extend_n59), .Y(exu_n9300));
AND2X1 exu_U27544(.A(alu_logic_rs1_data_bf1[43]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n61));
INVX1 exu_U27545(.A(shft_mux_rshift_extend_n61), .Y(exu_n9301));
AND2X1 exu_U27546(.A(alu_logic_rs1_data_bf1[42]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n63));
INVX1 exu_U27547(.A(shft_mux_rshift_extend_n63), .Y(exu_n9302));
AND2X1 exu_U27548(.A(alu_logic_rs1_data_bf1[32]), .B(ecl_shiftop_e[2]), .Y(shft_mux_rshift_extend_n65));
INVX1 exu_U27549(.A(shft_mux_rshift_extend_n65), .Y(exu_n9303));
OR2X1 exu_U27550(.A(exu_n12060), .B(exu_n14955), .Y(alu_chk_mem_addr_n4));
INVX1 exu_U27551(.A(alu_chk_mem_addr_n4), .Y(exu_n9304));
OR2X1 exu_U27552(.A(exu_n12063), .B(exu_n14957), .Y(alu_chk_mem_addr_n18));
INVX1 exu_U27553(.A(alu_chk_mem_addr_n18), .Y(exu_n9305));
AND2X1 exu_U27554(.A(exu_n11660), .B(ecl_mdqctl_n49), .Y(ecl_mdqctl_n47));
INVX1 exu_U27555(.A(ecl_mdqctl_n47), .Y(exu_n9306));
AND2X1 exu_U27556(.A(ecl_mdqctl_isdiv_w), .B(exu_n15395), .Y(ecl_mdqctl_n56));
INVX1 exu_U27557(.A(ecl_mdqctl_n56), .Y(exu_n9307));
AND2X1 exu_U27558(.A(exu_n16504), .B(ecl_divcntl_n26), .Y(ecl_divcntl_n25));
INVX1 exu_U27559(.A(ecl_divcntl_n25), .Y(exu_n9308));
AND2X1 exu_U27560(.A(exu_n16503), .B(exu_n10530), .Y(ecl_divcntl_n27));
INVX1 exu_U27561(.A(ecl_divcntl_n27), .Y(exu_n9309));
AND2X1 exu_U27562(.A(exu_n11664), .B(ecl_divcntl_n33), .Y(ecl_divcntl_n31));
INVX1 exu_U27563(.A(ecl_divcntl_n31), .Y(exu_n9310));
AND2X1 exu_U27564(.A(exu_n15398), .B(ecl_divcntl_div_state[5]), .Y(ecl_divcntl_n37));
INVX1 exu_U27565(.A(ecl_divcntl_n37), .Y(exu_n9311));
AND2X1 exu_U27566(.A(ecl_divcntl_subtract), .B(exu_n16257), .Y(ecl_divcntl_n64));
INVX1 exu_U27567(.A(ecl_divcntl_n64), .Y(exu_n9312));
AND2X1 exu_U27568(.A(ecl_divcntl_n66), .B(ecl_mdqctl_divcntl_muldone), .Y(ecl_divcntl_n65));
INVX1 exu_U27569(.A(ecl_divcntl_n65), .Y(exu_n9313));
AND2X1 exu_U27570(.A(ecl_divcntl_gencc_in_31_d1), .B(exu_n15684), .Y(ecl_divcntl_n71));
INVX1 exu_U27571(.A(ecl_divcntl_n71), .Y(exu_n9314));
AND2X1 exu_U27572(.A(ecl_divcntl_n76), .B(ecl_div_sel_neg32), .Y(ecl_divcntl_n75));
INVX1 exu_U27573(.A(ecl_divcntl_n75), .Y(exu_n9315));
AND2X1 exu_U27574(.A(exu_n15380), .B(ecl_byplog_rs2_n15), .Y(ecl_byplog_rs2_n13));
INVX1 exu_U27575(.A(ecl_byplog_rs2_n13), .Y(exu_n9316));
AND2X1 exu_U27576(.A(ecl_byplog_rs2_n29), .B(exu_n10536), .Y(ecl_byplog_rs2_n35));
INVX1 exu_U27577(.A(ecl_byplog_rs2_n35), .Y(exu_n9317));
AND2X1 exu_U27578(.A(exu_n15820), .B(exu_n15423), .Y(ecl_byplog_rs2_n38));
INVX1 exu_U27579(.A(ecl_byplog_rs2_n38), .Y(exu_n9318));
AND2X1 exu_U27580(.A(exu_n15464), .B(exu_n10537), .Y(ecl_byplog_rs2_n39));
INVX1 exu_U27581(.A(ecl_byplog_rs2_n39), .Y(exu_n9319));
AND2X1 exu_U27582(.A(exu_n11669), .B(exu_n10538), .Y(ecl_byplog_rs2_n48));
INVX1 exu_U27583(.A(ecl_byplog_rs2_n48), .Y(exu_n9320));
AND2X1 exu_U27584(.A(exu_n11670), .B(ecl_byplog_rs1_n20), .Y(ecl_byplog_rs1_n15));
INVX1 exu_U27585(.A(ecl_byplog_rs1_n15), .Y(exu_n9321));
OR2X1 exu_U27586(.A(ecl_ifu_exu_rs1_d[2]), .B(ecl_byplog_rs1_n41), .Y(ecl_byplog_rs1_n40));
INVX1 exu_U27587(.A(ecl_byplog_rs1_n40), .Y(exu_n9322));
AND2X1 exu_U27588(.A(exu_n15465), .B(exu_n10539), .Y(ecl_byplog_rs1_n43));
INVX1 exu_U27589(.A(ecl_byplog_rs1_n43), .Y(exu_n9323));
AND2X1 exu_U27590(.A(exu_n16592), .B(ecl_eccctl_n17), .Y(ecl_eccctl_n16));
INVX1 exu_U27591(.A(ecl_eccctl_n16), .Y(exu_n9324));
AND2X1 exu_U27592(.A(ecc_ecl_rs3_ce), .B(exu_n16394), .Y(ecl_eccctl_n22));
INVX1 exu_U27593(.A(ecl_eccctl_n22), .Y(exu_n9325));
AND2X1 exu_U27594(.A(ecl_eccctl_n35), .B(ecl_eccctl_rs1_ce_m), .Y(ecl_eccctl_n34));
INVX1 exu_U27595(.A(ecl_eccctl_n34), .Y(exu_n9326));
OR2X1 exu_U27596(.A(exu_n15356), .B(ecl_writeback_sraddr_w[1]), .Y(ecl_writeback_n43));
INVX1 exu_U27597(.A(ecl_writeback_n43), .Y(exu_n9327));
AND2X1 exu_U27598(.A(ecl_writeback_n130), .B(exu_n15482), .Y(ecl_writeback_n49));
INVX1 exu_U27599(.A(ecl_writeback_n49), .Y(exu_n9328));
OR2X1 exu_U27600(.A(ecl_writeback_sraddr_w[2]), .B(ecl_writeback_n57), .Y(ecl_writeback_n56));
INVX1 exu_U27601(.A(ecl_writeback_n56), .Y(exu_n9329));
INVX1 exu_U27602(.A(ecl_writeback_n182), .Y(exu_n9330));
OR2X1 exu_U27603(.A(ecl_writeback_n191), .B(exu_n16245), .Y(ecl_writeback_n182));
AND2X1 exu_U27604(.A(ecl_writeback_n101), .B(ecl_writeback_restore_tid[1]), .Y(ecl_writeback_n100));
INVX1 exu_U27605(.A(ecl_writeback_n100), .Y(exu_n9331));
AND2X1 exu_U27606(.A(exu_n11677), .B(ecl_writeback_restore_tid[1]), .Y(ecl_writeback_n108));
INVX1 exu_U27607(.A(ecl_writeback_n108), .Y(exu_n9332));
AND2X1 exu_U27608(.A(exu_n11678), .B(ecl_writeback_restore_tid[0]), .Y(ecl_writeback_n116));
INVX1 exu_U27609(.A(ecl_writeback_n116), .Y(exu_n9333));
AND2X1 exu_U27610(.A(ecl_mdqctl_wb_multhr_g[0]), .B(exu_n16199), .Y(ecl_writeback_n123));
INVX1 exu_U27611(.A(ecl_writeback_n123), .Y(exu_n9334));
AND2X1 exu_U27612(.A(ecl_mdqctl_wb_multhr_g[1]), .B(exu_n16199), .Y(ecl_writeback_n125));
INVX1 exu_U27613(.A(ecl_writeback_n125), .Y(exu_n9335));
AND2X1 exu_U27614(.A(exu_n11679), .B(ecl_writeback_n110), .Y(ecl_writeback_n127));
INVX1 exu_U27615(.A(ecl_writeback_n127), .Y(exu_n9336));
OR2X1 exu_U27616(.A(ecl_writeback_sraddr_e[6]), .B(ecl_writeback_sraddr_e[4]), .Y(ecl_writeback_n139));
INVX1 exu_U27617(.A(ecl_writeback_n139), .Y(exu_n9337));
AND2X1 exu_U27618(.A(exu_n16271), .B(ecl_writeback_n51), .Y(ecl_writeback_n154));
INVX1 exu_U27619(.A(ecl_writeback_n154), .Y(exu_n9338));
AND2X1 exu_U27620(.A(exu_n11682), .B(ecl_writeback_restore_w), .Y(ecl_writeback_n161));
INVX1 exu_U27621(.A(ecl_writeback_n161), .Y(exu_n9339));
AND2X1 exu_U27622(.A(ecl_writeback_restore_tid[1]), .B(exu_n15989), .Y(ecl_writeback_n169));
INVX1 exu_U27623(.A(ecl_writeback_n169), .Y(exu_n9340));
AND2X1 exu_U27624(.A(ecl_writeback_restore_tid[0]), .B(exu_n15989), .Y(ecl_writeback_n174));
INVX1 exu_U27625(.A(ecl_writeback_n174), .Y(exu_n9341));
OR2X1 exu_U27626(.A(exu_n16601), .B(exu_n14975), .Y(ecl_ccr_n22));
INVX1 exu_U27627(.A(ecl_ccr_n22), .Y(exu_n9342));
AND2X1 exu_U27628(.A(ecl_wb_ccr_wrccr_w), .B(exu_n16601), .Y(ecl_ccr_n37));
INVX1 exu_U27629(.A(ecl_ccr_n37), .Y(exu_n9343));
AND2X1 exu_U27630(.A(exu_n10761), .B(exu_n15029), .Y(ecl_ccr_n39));
INVX1 exu_U27631(.A(ecl_ccr_n39), .Y(exu_n9344));
AND2X1 exu_U27632(.A(exu_n10762), .B(exu_n15029), .Y(ecl_ccr_n42));
INVX1 exu_U27633(.A(ecl_ccr_n42), .Y(exu_n9345));
AND2X1 exu_U27634(.A(exu_n10763), .B(exu_n15029), .Y(ecl_ccr_n44));
INVX1 exu_U27635(.A(ecl_ccr_n44), .Y(exu_n9346));
AND2X1 exu_U27636(.A(exu_n10764), .B(exu_n15029), .Y(ecl_ccr_n46));
INVX1 exu_U27637(.A(ecl_ccr_n46), .Y(exu_n9347));
AND2X1 exu_U27638(.A(exu_n10765), .B(exu_n15029), .Y(ecl_ccr_n48));
INVX1 exu_U27639(.A(ecl_ccr_n48), .Y(exu_n9348));
AND2X1 exu_U27640(.A(exu_n10766), .B(exu_n15029), .Y(ecl_ccr_n50));
INVX1 exu_U27641(.A(ecl_ccr_n50), .Y(exu_n9349));
AND2X1 exu_U27642(.A(exu_n10767), .B(exu_n15029), .Y(ecl_ccr_n52));
INVX1 exu_U27643(.A(ecl_ccr_n52), .Y(exu_n9350));
AND2X1 exu_U27644(.A(exu_n10768), .B(exu_n15029), .Y(ecl_ccr_n54));
INVX1 exu_U27645(.A(ecl_ccr_n54), .Y(exu_n9351));
AND2X1 exu_U27646(.A(exu_n15030), .B(exu_n15930), .Y(ecl_ttype_mux_n12));
INVX1 exu_U27647(.A(ecl_ttype_mux_n12), .Y(exu_n9352));
AND2X1 exu_U27648(.A(exu_n11928), .B(exu_n15930), .Y(ecl_ttype_mux_n16));
INVX1 exu_U27649(.A(ecl_ttype_mux_n16), .Y(exu_n9353));
AND2X1 exu_U27650(.A(ecl_early1_ttype_e[4]), .B(exu_n15930), .Y(ecl_ttype_mux_n20));
INVX1 exu_U27651(.A(ecl_ttype_mux_n20), .Y(exu_n9354));
AND2X1 exu_U27652(.A(exu_n11930), .B(exu_n15930), .Y(ecl_ttype_mux_n24));
INVX1 exu_U27653(.A(ecl_ttype_mux_n24), .Y(exu_n9355));
AND2X1 exu_U27654(.A(exu_n11933), .B(exu_n15930), .Y(ecl_ttype_mux_n28));
INVX1 exu_U27655(.A(ecl_ttype_mux_n28), .Y(exu_n9356));
AND2X1 exu_U27656(.A(exu_n15337), .B(exu_n15930), .Y(ecl_ttype_mux_n36));
INVX1 exu_U27657(.A(ecl_ttype_mux_n36), .Y(exu_n9357));
AND2X1 exu_U27658(.A(exu_n15933), .B(div_yreg_div_ecl_yreg_0[2]), .Y(ecl_yreg0_mux_n4));
INVX1 exu_U27659(.A(ecl_yreg0_mux_n4), .Y(exu_n9358));
AND2X1 exu_U27660(.A(exu_n15935), .B(div_yreg_div_ecl_yreg_0[0]), .Y(ecl_yreg0_mux_n6));
INVX1 exu_U27661(.A(ecl_yreg0_mux_n6), .Y(exu_n9359));
AND2X1 exu_U27662(.A(ecl_ecc_sel_rs3_m_l), .B(ecc_rs3_err_m[6]), .Y(ecc_syn_mux_n2));
INVX1 exu_U27663(.A(ecc_syn_mux_n2), .Y(exu_n9360));
AND2X1 exu_U27664(.A(ecl_ecc_sel_rs1_m_l), .B(ecc_rs1_err_m[6]), .Y(ecc_syn_mux_n4));
INVX1 exu_U27665(.A(ecc_syn_mux_n4), .Y(exu_n9361));
AND2X1 exu_U27666(.A(ecc_rs3_err_m[5]), .B(ecl_ecc_sel_rs3_m_l), .Y(ecc_syn_mux_n6));
INVX1 exu_U27667(.A(ecc_syn_mux_n6), .Y(exu_n9362));
AND2X1 exu_U27668(.A(ecc_rs1_err_m[5]), .B(ecl_ecc_sel_rs1_m_l), .Y(ecc_syn_mux_n8));
INVX1 exu_U27669(.A(ecc_syn_mux_n8), .Y(exu_n9363));
AND2X1 exu_U27670(.A(ecc_rs3_err_m[4]), .B(ecl_ecc_sel_rs3_m_l), .Y(ecc_syn_mux_n10));
INVX1 exu_U27671(.A(ecc_syn_mux_n10), .Y(exu_n9364));
AND2X1 exu_U27672(.A(ecc_rs1_err_m[4]), .B(ecl_ecc_sel_rs1_m_l), .Y(ecc_syn_mux_n12));
INVX1 exu_U27673(.A(ecc_syn_mux_n12), .Y(exu_n9365));
AND2X1 exu_U27674(.A(ecc_rs3_err_m[3]), .B(ecl_ecc_sel_rs3_m_l), .Y(ecc_syn_mux_n14));
INVX1 exu_U27675(.A(ecc_syn_mux_n14), .Y(exu_n9366));
AND2X1 exu_U27676(.A(ecc_rs1_err_m[3]), .B(ecl_ecc_sel_rs1_m_l), .Y(ecc_syn_mux_n16));
INVX1 exu_U27677(.A(ecc_syn_mux_n16), .Y(exu_n9367));
AND2X1 exu_U27678(.A(ecc_rs3_err_m[2]), .B(ecl_ecc_sel_rs3_m_l), .Y(ecc_syn_mux_n18));
INVX1 exu_U27679(.A(ecc_syn_mux_n18), .Y(exu_n9368));
AND2X1 exu_U27680(.A(ecc_rs1_err_m[2]), .B(ecl_ecc_sel_rs1_m_l), .Y(ecc_syn_mux_n20));
INVX1 exu_U27681(.A(ecc_syn_mux_n20), .Y(exu_n9369));
AND2X1 exu_U27682(.A(ecc_rs3_err_m[1]), .B(ecl_ecc_sel_rs3_m_l), .Y(ecc_syn_mux_n22));
INVX1 exu_U27683(.A(ecc_syn_mux_n22), .Y(exu_n9370));
AND2X1 exu_U27684(.A(ecc_rs1_err_m[1]), .B(ecl_ecc_sel_rs1_m_l), .Y(ecc_syn_mux_n24));
INVX1 exu_U27685(.A(ecc_syn_mux_n24), .Y(exu_n9371));
AND2X1 exu_U27686(.A(ecc_rs3_err_m[0]), .B(ecl_ecc_sel_rs3_m_l), .Y(ecc_syn_mux_n26));
INVX1 exu_U27687(.A(ecc_syn_mux_n26), .Y(exu_n9372));
AND2X1 exu_U27688(.A(ecc_rs1_err_m[0]), .B(ecl_ecc_sel_rs1_m_l), .Y(ecc_syn_mux_n28));
INVX1 exu_U27689(.A(ecc_syn_mux_n28), .Y(exu_n9373));
OR2X1 exu_U27690(.A(ecc_rs1_err_e[6]), .B(ecc_rs1_err_e[5]), .Y(ecc_chk_rs1_n8));
INVX1 exu_U27691(.A(ecc_chk_rs1_n8), .Y(exu_n9374));
AND2X1 exu_U27692(.A(exu_n16286), .B(exu_tlu_wsr_data_m[9]), .Y(bypass_mux_rs3h_data_1_n6));
INVX1 exu_U27693(.A(bypass_mux_rs3h_data_1_n6), .Y(exu_n9375));
AND2X1 exu_U27694(.A(exu_tlu_wsr_data_m[8]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n12));
INVX1 exu_U27695(.A(bypass_mux_rs3h_data_1_n12), .Y(exu_n9376));
AND2X1 exu_U27696(.A(exu_tlu_wsr_data_m[7]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n18));
INVX1 exu_U27697(.A(bypass_mux_rs3h_data_1_n18), .Y(exu_n9377));
AND2X1 exu_U27698(.A(exu_tlu_wsr_data_m[6]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n24));
INVX1 exu_U27699(.A(bypass_mux_rs3h_data_1_n24), .Y(exu_n9378));
AND2X1 exu_U27700(.A(exu_tlu_wsr_data_m[5]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n30));
INVX1 exu_U27701(.A(bypass_mux_rs3h_data_1_n30), .Y(exu_n9379));
AND2X1 exu_U27702(.A(exu_tlu_wsr_data_m[4]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n36));
INVX1 exu_U27703(.A(bypass_mux_rs3h_data_1_n36), .Y(exu_n9380));
AND2X1 exu_U27704(.A(exu_tlu_wsr_data_m[3]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n42));
INVX1 exu_U27705(.A(bypass_mux_rs3h_data_1_n42), .Y(exu_n9381));
AND2X1 exu_U27706(.A(exu_tlu_wsr_data_m[31]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n48));
INVX1 exu_U27707(.A(bypass_mux_rs3h_data_1_n48), .Y(exu_n9382));
AND2X1 exu_U27708(.A(exu_tlu_wsr_data_m[30]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n54));
INVX1 exu_U27709(.A(bypass_mux_rs3h_data_1_n54), .Y(exu_n9383));
AND2X1 exu_U27710(.A(exu_tlu_wsr_data_m[2]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n60));
INVX1 exu_U27711(.A(bypass_mux_rs3h_data_1_n60), .Y(exu_n9384));
AND2X1 exu_U27712(.A(exu_tlu_wsr_data_m[29]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n66));
INVX1 exu_U27713(.A(bypass_mux_rs3h_data_1_n66), .Y(exu_n9385));
AND2X1 exu_U27714(.A(exu_tlu_wsr_data_m[28]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n72));
INVX1 exu_U27715(.A(bypass_mux_rs3h_data_1_n72), .Y(exu_n9386));
AND2X1 exu_U27716(.A(exu_tlu_wsr_data_m[27]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n78));
INVX1 exu_U27717(.A(bypass_mux_rs3h_data_1_n78), .Y(exu_n9387));
AND2X1 exu_U27718(.A(exu_tlu_wsr_data_m[26]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n84));
INVX1 exu_U27719(.A(bypass_mux_rs3h_data_1_n84), .Y(exu_n9388));
AND2X1 exu_U27720(.A(exu_tlu_wsr_data_m[25]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n90));
INVX1 exu_U27721(.A(bypass_mux_rs3h_data_1_n90), .Y(exu_n9389));
AND2X1 exu_U27722(.A(exu_tlu_wsr_data_m[24]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n96));
INVX1 exu_U27723(.A(bypass_mux_rs3h_data_1_n96), .Y(exu_n9390));
AND2X1 exu_U27724(.A(exu_tlu_wsr_data_m[23]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n102));
INVX1 exu_U27725(.A(bypass_mux_rs3h_data_1_n102), .Y(exu_n9391));
AND2X1 exu_U27726(.A(exu_tlu_wsr_data_m[22]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n108));
INVX1 exu_U27727(.A(bypass_mux_rs3h_data_1_n108), .Y(exu_n9392));
AND2X1 exu_U27728(.A(exu_tlu_wsr_data_m[21]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n114));
INVX1 exu_U27729(.A(bypass_mux_rs3h_data_1_n114), .Y(exu_n9393));
AND2X1 exu_U27730(.A(exu_tlu_wsr_data_m[20]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n120));
INVX1 exu_U27731(.A(bypass_mux_rs3h_data_1_n120), .Y(exu_n9394));
AND2X1 exu_U27732(.A(exu_tlu_wsr_data_m[1]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n126));
INVX1 exu_U27733(.A(bypass_mux_rs3h_data_1_n126), .Y(exu_n9395));
AND2X1 exu_U27734(.A(exu_tlu_wsr_data_m[19]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n132));
INVX1 exu_U27735(.A(bypass_mux_rs3h_data_1_n132), .Y(exu_n9396));
AND2X1 exu_U27736(.A(exu_tlu_wsr_data_m[18]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n138));
INVX1 exu_U27737(.A(bypass_mux_rs3h_data_1_n138), .Y(exu_n9397));
AND2X1 exu_U27738(.A(exu_tlu_wsr_data_m[17]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n144));
INVX1 exu_U27739(.A(bypass_mux_rs3h_data_1_n144), .Y(exu_n9398));
AND2X1 exu_U27740(.A(exu_tlu_wsr_data_m[16]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n150));
INVX1 exu_U27741(.A(bypass_mux_rs3h_data_1_n150), .Y(exu_n9399));
AND2X1 exu_U27742(.A(exu_tlu_wsr_data_m[15]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n156));
INVX1 exu_U27743(.A(bypass_mux_rs3h_data_1_n156), .Y(exu_n9400));
AND2X1 exu_U27744(.A(exu_tlu_wsr_data_m[14]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n162));
INVX1 exu_U27745(.A(bypass_mux_rs3h_data_1_n162), .Y(exu_n9401));
AND2X1 exu_U27746(.A(exu_tlu_wsr_data_m[13]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n168));
INVX1 exu_U27747(.A(bypass_mux_rs3h_data_1_n168), .Y(exu_n9402));
AND2X1 exu_U27748(.A(exu_tlu_wsr_data_m[12]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n174));
INVX1 exu_U27749(.A(bypass_mux_rs3h_data_1_n174), .Y(exu_n9403));
AND2X1 exu_U27750(.A(exu_tlu_wsr_data_m[11]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n180));
INVX1 exu_U27751(.A(bypass_mux_rs3h_data_1_n180), .Y(exu_n9404));
AND2X1 exu_U27752(.A(exu_tlu_wsr_data_m[10]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n186));
INVX1 exu_U27753(.A(bypass_mux_rs3h_data_1_n186), .Y(exu_n9405));
AND2X1 exu_U27754(.A(exu_tlu_wsr_data_m[0]), .B(exu_n16286), .Y(bypass_mux_rs3h_data_1_n192));
INVX1 exu_U27755(.A(bypass_mux_rs3h_data_1_n192), .Y(exu_n9406));
AND2X1 exu_U27756(.A(bypass_rs3h_w2_mux_n1), .B(exu_n10555), .Y(bypass_rs3h_data_w2[9]));
INVX1 exu_U27757(.A(bypass_rs3h_data_w2[9]), .Y(exu_n9407));
AND2X1 exu_U27758(.A(ecl_byp_rs3h_longmux_sel_w2), .B(byp_irf_rd_data_w2[9]), .Y(bypass_rs3h_w2_mux_n4));
INVX1 exu_U27759(.A(bypass_rs3h_w2_mux_n4), .Y(exu_n9408));
AND2X1 exu_U27760(.A(byp_irf_rd_data_w2[8]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n8));
INVX1 exu_U27761(.A(bypass_rs3h_w2_mux_n8), .Y(exu_n9409));
AND2X1 exu_U27762(.A(byp_irf_rd_data_w2[7]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n12));
INVX1 exu_U27763(.A(bypass_rs3h_w2_mux_n12), .Y(exu_n9410));
AND2X1 exu_U27764(.A(byp_irf_rd_data_w2[6]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n16));
INVX1 exu_U27765(.A(bypass_rs3h_w2_mux_n16), .Y(exu_n9411));
AND2X1 exu_U27766(.A(byp_irf_rd_data_w2[5]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n20));
INVX1 exu_U27767(.A(bypass_rs3h_w2_mux_n20), .Y(exu_n9412));
AND2X1 exu_U27768(.A(byp_irf_rd_data_w2[4]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n24));
INVX1 exu_U27769(.A(bypass_rs3h_w2_mux_n24), .Y(exu_n9413));
AND2X1 exu_U27770(.A(byp_irf_rd_data_w2[3]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n28));
INVX1 exu_U27771(.A(bypass_rs3h_w2_mux_n28), .Y(exu_n9414));
AND2X1 exu_U27772(.A(byp_irf_rd_data_w2[31]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n32));
INVX1 exu_U27773(.A(bypass_rs3h_w2_mux_n32), .Y(exu_n9415));
AND2X1 exu_U27774(.A(byp_irf_rd_data_w2[30]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n36));
INVX1 exu_U27775(.A(bypass_rs3h_w2_mux_n36), .Y(exu_n9416));
AND2X1 exu_U27776(.A(byp_irf_rd_data_w2[2]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n40));
INVX1 exu_U27777(.A(bypass_rs3h_w2_mux_n40), .Y(exu_n9417));
AND2X1 exu_U27778(.A(byp_irf_rd_data_w2[29]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n44));
INVX1 exu_U27779(.A(bypass_rs3h_w2_mux_n44), .Y(exu_n9418));
AND2X1 exu_U27780(.A(byp_irf_rd_data_w2[28]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n48));
INVX1 exu_U27781(.A(bypass_rs3h_w2_mux_n48), .Y(exu_n9419));
AND2X1 exu_U27782(.A(byp_irf_rd_data_w2[27]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n52));
INVX1 exu_U27783(.A(bypass_rs3h_w2_mux_n52), .Y(exu_n9420));
AND2X1 exu_U27784(.A(byp_irf_rd_data_w2[26]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n56));
INVX1 exu_U27785(.A(bypass_rs3h_w2_mux_n56), .Y(exu_n9421));
AND2X1 exu_U27786(.A(byp_irf_rd_data_w2[25]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n60));
INVX1 exu_U27787(.A(bypass_rs3h_w2_mux_n60), .Y(exu_n9422));
AND2X1 exu_U27788(.A(byp_irf_rd_data_w2[24]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n64));
INVX1 exu_U27789(.A(bypass_rs3h_w2_mux_n64), .Y(exu_n9423));
AND2X1 exu_U27790(.A(byp_irf_rd_data_w2[23]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n68));
INVX1 exu_U27791(.A(bypass_rs3h_w2_mux_n68), .Y(exu_n9424));
AND2X1 exu_U27792(.A(byp_irf_rd_data_w2[22]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n72));
INVX1 exu_U27793(.A(bypass_rs3h_w2_mux_n72), .Y(exu_n9425));
AND2X1 exu_U27794(.A(byp_irf_rd_data_w2[21]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n76));
INVX1 exu_U27795(.A(bypass_rs3h_w2_mux_n76), .Y(exu_n9426));
AND2X1 exu_U27796(.A(byp_irf_rd_data_w2[20]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n80));
INVX1 exu_U27797(.A(bypass_rs3h_w2_mux_n80), .Y(exu_n9427));
AND2X1 exu_U27798(.A(byp_irf_rd_data_w2[1]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n84));
INVX1 exu_U27799(.A(bypass_rs3h_w2_mux_n84), .Y(exu_n9428));
AND2X1 exu_U27800(.A(byp_irf_rd_data_w2[19]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n88));
INVX1 exu_U27801(.A(bypass_rs3h_w2_mux_n88), .Y(exu_n9429));
AND2X1 exu_U27802(.A(byp_irf_rd_data_w2[18]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n92));
INVX1 exu_U27803(.A(bypass_rs3h_w2_mux_n92), .Y(exu_n9430));
AND2X1 exu_U27804(.A(byp_irf_rd_data_w2[17]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n96));
INVX1 exu_U27805(.A(bypass_rs3h_w2_mux_n96), .Y(exu_n9431));
AND2X1 exu_U27806(.A(byp_irf_rd_data_w2[16]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n100));
INVX1 exu_U27807(.A(bypass_rs3h_w2_mux_n100), .Y(exu_n9432));
AND2X1 exu_U27808(.A(byp_irf_rd_data_w2[15]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n104));
INVX1 exu_U27809(.A(bypass_rs3h_w2_mux_n104), .Y(exu_n9433));
AND2X1 exu_U27810(.A(byp_irf_rd_data_w2[14]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n108));
INVX1 exu_U27811(.A(bypass_rs3h_w2_mux_n108), .Y(exu_n9434));
AND2X1 exu_U27812(.A(byp_irf_rd_data_w2[13]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n112));
INVX1 exu_U27813(.A(bypass_rs3h_w2_mux_n112), .Y(exu_n9435));
AND2X1 exu_U27814(.A(byp_irf_rd_data_w2[12]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n116));
INVX1 exu_U27815(.A(bypass_rs3h_w2_mux_n116), .Y(exu_n9436));
AND2X1 exu_U27816(.A(byp_irf_rd_data_w2[11]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n120));
INVX1 exu_U27817(.A(bypass_rs3h_w2_mux_n120), .Y(exu_n9437));
AND2X1 exu_U27818(.A(byp_irf_rd_data_w2[10]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n124));
INVX1 exu_U27819(.A(bypass_rs3h_w2_mux_n124), .Y(exu_n9438));
AND2X1 exu_U27820(.A(byp_irf_rd_data_w2[0]), .B(ecl_byp_rs3h_longmux_sel_w2), .Y(bypass_rs3h_w2_mux_n128));
INVX1 exu_U27821(.A(bypass_rs3h_w2_mux_n128), .Y(exu_n9439));
AND2X1 exu_U27822(.A(exu_n16264), .B(exu_tlu_wsr_data_m[9]), .Y(bypass_sr_out_mux_n4));
INVX1 exu_U27823(.A(bypass_sr_out_mux_n4), .Y(exu_n9440));
AND2X1 exu_U27824(.A(tlu_exu_rsr_data_m[8]), .B(exu_n16263), .Y(bypass_sr_out_mux_n6));
INVX1 exu_U27825(.A(bypass_sr_out_mux_n6), .Y(exu_n9441));
AND2X1 exu_U27826(.A(exu_tlu_wsr_data_m[8]), .B(exu_n16264), .Y(bypass_sr_out_mux_n8));
INVX1 exu_U27827(.A(bypass_sr_out_mux_n8), .Y(exu_n9442));
AND2X1 exu_U27828(.A(tlu_exu_rsr_data_m[7]), .B(exu_n16263), .Y(bypass_sr_out_mux_n10));
INVX1 exu_U27829(.A(bypass_sr_out_mux_n10), .Y(exu_n9443));
AND2X1 exu_U27830(.A(exu_tlu_wsr_data_m[7]), .B(exu_n16264), .Y(bypass_sr_out_mux_n12));
INVX1 exu_U27831(.A(bypass_sr_out_mux_n12), .Y(exu_n9444));
AND2X1 exu_U27832(.A(tlu_exu_rsr_data_m[6]), .B(exu_n16263), .Y(bypass_sr_out_mux_n14));
INVX1 exu_U27833(.A(bypass_sr_out_mux_n14), .Y(exu_n9445));
AND2X1 exu_U27834(.A(exu_tlu_wsr_data_m[6]), .B(exu_n16264), .Y(bypass_sr_out_mux_n16));
INVX1 exu_U27835(.A(bypass_sr_out_mux_n16), .Y(exu_n9446));
AND2X1 exu_U27836(.A(tlu_exu_rsr_data_m[63]), .B(exu_n16263), .Y(bypass_sr_out_mux_n18));
INVX1 exu_U27837(.A(bypass_sr_out_mux_n18), .Y(exu_n9447));
AND2X1 exu_U27838(.A(exu_tlu_wsr_data_m[63]), .B(exu_n16264), .Y(bypass_sr_out_mux_n20));
INVX1 exu_U27839(.A(bypass_sr_out_mux_n20), .Y(exu_n9448));
AND2X1 exu_U27840(.A(tlu_exu_rsr_data_m[62]), .B(exu_n16263), .Y(bypass_sr_out_mux_n22));
INVX1 exu_U27841(.A(bypass_sr_out_mux_n22), .Y(exu_n9449));
AND2X1 exu_U27842(.A(exu_tlu_wsr_data_m[62]), .B(exu_n16264), .Y(bypass_sr_out_mux_n24));
INVX1 exu_U27843(.A(bypass_sr_out_mux_n24), .Y(exu_n9450));
AND2X1 exu_U27844(.A(tlu_exu_rsr_data_m[61]), .B(exu_n16263), .Y(bypass_sr_out_mux_n26));
INVX1 exu_U27845(.A(bypass_sr_out_mux_n26), .Y(exu_n9451));
AND2X1 exu_U27846(.A(exu_tlu_wsr_data_m[61]), .B(exu_n16264), .Y(bypass_sr_out_mux_n28));
INVX1 exu_U27847(.A(bypass_sr_out_mux_n28), .Y(exu_n9452));
AND2X1 exu_U27848(.A(tlu_exu_rsr_data_m[60]), .B(exu_n16263), .Y(bypass_sr_out_mux_n30));
INVX1 exu_U27849(.A(bypass_sr_out_mux_n30), .Y(exu_n9453));
AND2X1 exu_U27850(.A(exu_tlu_wsr_data_m[60]), .B(exu_n16264), .Y(bypass_sr_out_mux_n32));
INVX1 exu_U27851(.A(bypass_sr_out_mux_n32), .Y(exu_n9454));
AND2X1 exu_U27852(.A(tlu_exu_rsr_data_m[5]), .B(exu_n16263), .Y(bypass_sr_out_mux_n34));
INVX1 exu_U27853(.A(bypass_sr_out_mux_n34), .Y(exu_n9455));
AND2X1 exu_U27854(.A(exu_tlu_wsr_data_m[5]), .B(exu_n16264), .Y(bypass_sr_out_mux_n36));
INVX1 exu_U27855(.A(bypass_sr_out_mux_n36), .Y(exu_n9456));
AND2X1 exu_U27856(.A(tlu_exu_rsr_data_m[59]), .B(exu_n16263), .Y(bypass_sr_out_mux_n38));
INVX1 exu_U27857(.A(bypass_sr_out_mux_n38), .Y(exu_n9457));
AND2X1 exu_U27858(.A(exu_tlu_wsr_data_m[59]), .B(exu_n16264), .Y(bypass_sr_out_mux_n40));
INVX1 exu_U27859(.A(bypass_sr_out_mux_n40), .Y(exu_n9458));
AND2X1 exu_U27860(.A(tlu_exu_rsr_data_m[58]), .B(exu_n16263), .Y(bypass_sr_out_mux_n42));
INVX1 exu_U27861(.A(bypass_sr_out_mux_n42), .Y(exu_n9459));
AND2X1 exu_U27862(.A(exu_tlu_wsr_data_m[58]), .B(exu_n16264), .Y(bypass_sr_out_mux_n44));
INVX1 exu_U27863(.A(bypass_sr_out_mux_n44), .Y(exu_n9460));
AND2X1 exu_U27864(.A(tlu_exu_rsr_data_m[57]), .B(exu_n16263), .Y(bypass_sr_out_mux_n46));
INVX1 exu_U27865(.A(bypass_sr_out_mux_n46), .Y(exu_n9461));
AND2X1 exu_U27866(.A(exu_tlu_wsr_data_m[57]), .B(exu_n16264), .Y(bypass_sr_out_mux_n48));
INVX1 exu_U27867(.A(bypass_sr_out_mux_n48), .Y(exu_n9462));
AND2X1 exu_U27868(.A(tlu_exu_rsr_data_m[56]), .B(exu_n16263), .Y(bypass_sr_out_mux_n50));
INVX1 exu_U27869(.A(bypass_sr_out_mux_n50), .Y(exu_n9463));
AND2X1 exu_U27870(.A(exu_tlu_wsr_data_m[56]), .B(exu_n16264), .Y(bypass_sr_out_mux_n52));
INVX1 exu_U27871(.A(bypass_sr_out_mux_n52), .Y(exu_n9464));
AND2X1 exu_U27872(.A(tlu_exu_rsr_data_m[55]), .B(exu_n16263), .Y(bypass_sr_out_mux_n54));
INVX1 exu_U27873(.A(bypass_sr_out_mux_n54), .Y(exu_n9465));
AND2X1 exu_U27874(.A(exu_tlu_wsr_data_m[55]), .B(exu_n16264), .Y(bypass_sr_out_mux_n56));
INVX1 exu_U27875(.A(bypass_sr_out_mux_n56), .Y(exu_n9466));
AND2X1 exu_U27876(.A(tlu_exu_rsr_data_m[54]), .B(exu_n16263), .Y(bypass_sr_out_mux_n58));
INVX1 exu_U27877(.A(bypass_sr_out_mux_n58), .Y(exu_n9467));
AND2X1 exu_U27878(.A(exu_tlu_wsr_data_m[54]), .B(exu_n16264), .Y(bypass_sr_out_mux_n60));
INVX1 exu_U27879(.A(bypass_sr_out_mux_n60), .Y(exu_n9468));
AND2X1 exu_U27880(.A(tlu_exu_rsr_data_m[53]), .B(exu_n16263), .Y(bypass_sr_out_mux_n62));
INVX1 exu_U27881(.A(bypass_sr_out_mux_n62), .Y(exu_n9469));
AND2X1 exu_U27882(.A(exu_tlu_wsr_data_m[53]), .B(exu_n16264), .Y(bypass_sr_out_mux_n64));
INVX1 exu_U27883(.A(bypass_sr_out_mux_n64), .Y(exu_n9470));
AND2X1 exu_U27884(.A(tlu_exu_rsr_data_m[52]), .B(exu_n16263), .Y(bypass_sr_out_mux_n66));
INVX1 exu_U27885(.A(bypass_sr_out_mux_n66), .Y(exu_n9471));
AND2X1 exu_U27886(.A(exu_tlu_wsr_data_m[52]), .B(exu_n16264), .Y(bypass_sr_out_mux_n68));
INVX1 exu_U27887(.A(bypass_sr_out_mux_n68), .Y(exu_n9472));
AND2X1 exu_U27888(.A(tlu_exu_rsr_data_m[51]), .B(exu_n16263), .Y(bypass_sr_out_mux_n70));
INVX1 exu_U27889(.A(bypass_sr_out_mux_n70), .Y(exu_n9473));
AND2X1 exu_U27890(.A(exu_tlu_wsr_data_m[51]), .B(exu_n16264), .Y(bypass_sr_out_mux_n72));
INVX1 exu_U27891(.A(bypass_sr_out_mux_n72), .Y(exu_n9474));
AND2X1 exu_U27892(.A(tlu_exu_rsr_data_m[50]), .B(exu_n16263), .Y(bypass_sr_out_mux_n74));
INVX1 exu_U27893(.A(bypass_sr_out_mux_n74), .Y(exu_n9475));
AND2X1 exu_U27894(.A(exu_tlu_wsr_data_m[50]), .B(exu_n16264), .Y(bypass_sr_out_mux_n76));
INVX1 exu_U27895(.A(bypass_sr_out_mux_n76), .Y(exu_n9476));
AND2X1 exu_U27896(.A(tlu_exu_rsr_data_m[4]), .B(exu_n16263), .Y(bypass_sr_out_mux_n78));
INVX1 exu_U27897(.A(bypass_sr_out_mux_n78), .Y(exu_n9477));
AND2X1 exu_U27898(.A(exu_tlu_wsr_data_m[4]), .B(exu_n16264), .Y(bypass_sr_out_mux_n80));
INVX1 exu_U27899(.A(bypass_sr_out_mux_n80), .Y(exu_n9478));
AND2X1 exu_U27900(.A(tlu_exu_rsr_data_m[49]), .B(exu_n16263), .Y(bypass_sr_out_mux_n82));
INVX1 exu_U27901(.A(bypass_sr_out_mux_n82), .Y(exu_n9479));
AND2X1 exu_U27902(.A(exu_tlu_wsr_data_m[49]), .B(exu_n16264), .Y(bypass_sr_out_mux_n84));
INVX1 exu_U27903(.A(bypass_sr_out_mux_n84), .Y(exu_n9480));
AND2X1 exu_U27904(.A(tlu_exu_rsr_data_m[48]), .B(exu_n16263), .Y(bypass_sr_out_mux_n86));
INVX1 exu_U27905(.A(bypass_sr_out_mux_n86), .Y(exu_n9481));
AND2X1 exu_U27906(.A(exu_tlu_wsr_data_m[48]), .B(exu_n16264), .Y(bypass_sr_out_mux_n88));
INVX1 exu_U27907(.A(bypass_sr_out_mux_n88), .Y(exu_n9482));
AND2X1 exu_U27908(.A(tlu_exu_rsr_data_m[47]), .B(exu_n16263), .Y(bypass_sr_out_mux_n90));
INVX1 exu_U27909(.A(bypass_sr_out_mux_n90), .Y(exu_n9483));
AND2X1 exu_U27910(.A(exu_tlu_wsr_data_m[47]), .B(exu_n16264), .Y(bypass_sr_out_mux_n92));
INVX1 exu_U27911(.A(bypass_sr_out_mux_n92), .Y(exu_n9484));
AND2X1 exu_U27912(.A(tlu_exu_rsr_data_m[46]), .B(exu_n16263), .Y(bypass_sr_out_mux_n94));
INVX1 exu_U27913(.A(bypass_sr_out_mux_n94), .Y(exu_n9485));
AND2X1 exu_U27914(.A(exu_tlu_wsr_data_m[46]), .B(exu_n16264), .Y(bypass_sr_out_mux_n96));
INVX1 exu_U27915(.A(bypass_sr_out_mux_n96), .Y(exu_n9486));
AND2X1 exu_U27916(.A(tlu_exu_rsr_data_m[45]), .B(exu_n16263), .Y(bypass_sr_out_mux_n98));
INVX1 exu_U27917(.A(bypass_sr_out_mux_n98), .Y(exu_n9487));
AND2X1 exu_U27918(.A(exu_tlu_wsr_data_m[45]), .B(exu_n16264), .Y(bypass_sr_out_mux_n100));
INVX1 exu_U27919(.A(bypass_sr_out_mux_n100), .Y(exu_n9488));
AND2X1 exu_U27920(.A(tlu_exu_rsr_data_m[44]), .B(exu_n16263), .Y(bypass_sr_out_mux_n102));
INVX1 exu_U27921(.A(bypass_sr_out_mux_n102), .Y(exu_n9489));
AND2X1 exu_U27922(.A(exu_tlu_wsr_data_m[44]), .B(exu_n16264), .Y(bypass_sr_out_mux_n104));
INVX1 exu_U27923(.A(bypass_sr_out_mux_n104), .Y(exu_n9490));
AND2X1 exu_U27924(.A(tlu_exu_rsr_data_m[43]), .B(exu_n16263), .Y(bypass_sr_out_mux_n106));
INVX1 exu_U27925(.A(bypass_sr_out_mux_n106), .Y(exu_n9491));
AND2X1 exu_U27926(.A(exu_tlu_wsr_data_m[43]), .B(exu_n16264), .Y(bypass_sr_out_mux_n108));
INVX1 exu_U27927(.A(bypass_sr_out_mux_n108), .Y(exu_n9492));
AND2X1 exu_U27928(.A(tlu_exu_rsr_data_m[42]), .B(exu_n16263), .Y(bypass_sr_out_mux_n110));
INVX1 exu_U27929(.A(bypass_sr_out_mux_n110), .Y(exu_n9493));
AND2X1 exu_U27930(.A(exu_tlu_wsr_data_m[42]), .B(exu_n16264), .Y(bypass_sr_out_mux_n112));
INVX1 exu_U27931(.A(bypass_sr_out_mux_n112), .Y(exu_n9494));
AND2X1 exu_U27932(.A(tlu_exu_rsr_data_m[41]), .B(exu_n16263), .Y(bypass_sr_out_mux_n114));
INVX1 exu_U27933(.A(bypass_sr_out_mux_n114), .Y(exu_n9495));
AND2X1 exu_U27934(.A(exu_tlu_wsr_data_m[41]), .B(exu_n16264), .Y(bypass_sr_out_mux_n116));
INVX1 exu_U27935(.A(bypass_sr_out_mux_n116), .Y(exu_n9496));
AND2X1 exu_U27936(.A(tlu_exu_rsr_data_m[40]), .B(exu_n16263), .Y(bypass_sr_out_mux_n118));
INVX1 exu_U27937(.A(bypass_sr_out_mux_n118), .Y(exu_n9497));
AND2X1 exu_U27938(.A(exu_tlu_wsr_data_m[40]), .B(exu_n16264), .Y(bypass_sr_out_mux_n120));
INVX1 exu_U27939(.A(bypass_sr_out_mux_n120), .Y(exu_n9498));
AND2X1 exu_U27940(.A(tlu_exu_rsr_data_m[3]), .B(exu_n16263), .Y(bypass_sr_out_mux_n122));
INVX1 exu_U27941(.A(bypass_sr_out_mux_n122), .Y(exu_n9499));
AND2X1 exu_U27942(.A(exu_tlu_wsr_data_m[3]), .B(exu_n16264), .Y(bypass_sr_out_mux_n124));
INVX1 exu_U27943(.A(bypass_sr_out_mux_n124), .Y(exu_n9500));
AND2X1 exu_U27944(.A(tlu_exu_rsr_data_m[39]), .B(exu_n16263), .Y(bypass_sr_out_mux_n126));
INVX1 exu_U27945(.A(bypass_sr_out_mux_n126), .Y(exu_n9501));
AND2X1 exu_U27946(.A(exu_tlu_wsr_data_m[39]), .B(exu_n16264), .Y(bypass_sr_out_mux_n128));
INVX1 exu_U27947(.A(bypass_sr_out_mux_n128), .Y(exu_n9502));
AND2X1 exu_U27948(.A(tlu_exu_rsr_data_m[38]), .B(exu_n16263), .Y(bypass_sr_out_mux_n130));
INVX1 exu_U27949(.A(bypass_sr_out_mux_n130), .Y(exu_n9503));
AND2X1 exu_U27950(.A(exu_tlu_wsr_data_m[38]), .B(exu_n16264), .Y(bypass_sr_out_mux_n132));
INVX1 exu_U27951(.A(bypass_sr_out_mux_n132), .Y(exu_n9504));
AND2X1 exu_U27952(.A(tlu_exu_rsr_data_m[37]), .B(exu_n16263), .Y(bypass_sr_out_mux_n134));
INVX1 exu_U27953(.A(bypass_sr_out_mux_n134), .Y(exu_n9505));
AND2X1 exu_U27954(.A(exu_tlu_wsr_data_m[37]), .B(exu_n16264), .Y(bypass_sr_out_mux_n136));
INVX1 exu_U27955(.A(bypass_sr_out_mux_n136), .Y(exu_n9506));
AND2X1 exu_U27956(.A(tlu_exu_rsr_data_m[36]), .B(exu_n16263), .Y(bypass_sr_out_mux_n138));
INVX1 exu_U27957(.A(bypass_sr_out_mux_n138), .Y(exu_n9507));
AND2X1 exu_U27958(.A(exu_tlu_wsr_data_m[36]), .B(exu_n16264), .Y(bypass_sr_out_mux_n140));
INVX1 exu_U27959(.A(bypass_sr_out_mux_n140), .Y(exu_n9508));
AND2X1 exu_U27960(.A(tlu_exu_rsr_data_m[35]), .B(exu_n16263), .Y(bypass_sr_out_mux_n142));
INVX1 exu_U27961(.A(bypass_sr_out_mux_n142), .Y(exu_n9509));
AND2X1 exu_U27962(.A(exu_tlu_wsr_data_m[35]), .B(exu_n16264), .Y(bypass_sr_out_mux_n144));
INVX1 exu_U27963(.A(bypass_sr_out_mux_n144), .Y(exu_n9510));
AND2X1 exu_U27964(.A(tlu_exu_rsr_data_m[34]), .B(exu_n16263), .Y(bypass_sr_out_mux_n146));
INVX1 exu_U27965(.A(bypass_sr_out_mux_n146), .Y(exu_n9511));
AND2X1 exu_U27966(.A(exu_tlu_wsr_data_m[34]), .B(exu_n16264), .Y(bypass_sr_out_mux_n148));
INVX1 exu_U27967(.A(bypass_sr_out_mux_n148), .Y(exu_n9512));
AND2X1 exu_U27968(.A(tlu_exu_rsr_data_m[33]), .B(exu_n16263), .Y(bypass_sr_out_mux_n150));
INVX1 exu_U27969(.A(bypass_sr_out_mux_n150), .Y(exu_n9513));
AND2X1 exu_U27970(.A(exu_tlu_wsr_data_m[33]), .B(exu_n16264), .Y(bypass_sr_out_mux_n152));
INVX1 exu_U27971(.A(bypass_sr_out_mux_n152), .Y(exu_n9514));
AND2X1 exu_U27972(.A(tlu_exu_rsr_data_m[32]), .B(exu_n16263), .Y(bypass_sr_out_mux_n154));
INVX1 exu_U27973(.A(bypass_sr_out_mux_n154), .Y(exu_n9515));
AND2X1 exu_U27974(.A(exu_tlu_wsr_data_m[32]), .B(exu_n16264), .Y(bypass_sr_out_mux_n156));
INVX1 exu_U27975(.A(bypass_sr_out_mux_n156), .Y(exu_n9516));
AND2X1 exu_U27976(.A(tlu_exu_rsr_data_m[31]), .B(exu_n16263), .Y(bypass_sr_out_mux_n158));
INVX1 exu_U27977(.A(bypass_sr_out_mux_n158), .Y(exu_n9517));
AND2X1 exu_U27978(.A(exu_tlu_wsr_data_m[31]), .B(exu_n16264), .Y(bypass_sr_out_mux_n160));
INVX1 exu_U27979(.A(bypass_sr_out_mux_n160), .Y(exu_n9518));
AND2X1 exu_U27980(.A(tlu_exu_rsr_data_m[30]), .B(exu_n16263), .Y(bypass_sr_out_mux_n162));
INVX1 exu_U27981(.A(bypass_sr_out_mux_n162), .Y(exu_n9519));
AND2X1 exu_U27982(.A(exu_tlu_wsr_data_m[30]), .B(exu_n16264), .Y(bypass_sr_out_mux_n164));
INVX1 exu_U27983(.A(bypass_sr_out_mux_n164), .Y(exu_n9520));
AND2X1 exu_U27984(.A(tlu_exu_rsr_data_m[2]), .B(exu_n16263), .Y(bypass_sr_out_mux_n166));
INVX1 exu_U27985(.A(bypass_sr_out_mux_n166), .Y(exu_n9521));
AND2X1 exu_U27986(.A(ecl_byp_3lsb_m[2]), .B(exu_n16264), .Y(bypass_sr_out_mux_n168));
INVX1 exu_U27987(.A(bypass_sr_out_mux_n168), .Y(exu_n9522));
AND2X1 exu_U27988(.A(tlu_exu_rsr_data_m[29]), .B(exu_n16263), .Y(bypass_sr_out_mux_n170));
INVX1 exu_U27989(.A(bypass_sr_out_mux_n170), .Y(exu_n9523));
AND2X1 exu_U27990(.A(exu_tlu_wsr_data_m[29]), .B(exu_n16264), .Y(bypass_sr_out_mux_n172));
INVX1 exu_U27991(.A(bypass_sr_out_mux_n172), .Y(exu_n9524));
AND2X1 exu_U27992(.A(tlu_exu_rsr_data_m[28]), .B(exu_n16263), .Y(bypass_sr_out_mux_n174));
INVX1 exu_U27993(.A(bypass_sr_out_mux_n174), .Y(exu_n9525));
AND2X1 exu_U27994(.A(exu_tlu_wsr_data_m[28]), .B(exu_n16264), .Y(bypass_sr_out_mux_n176));
INVX1 exu_U27995(.A(bypass_sr_out_mux_n176), .Y(exu_n9526));
AND2X1 exu_U27996(.A(tlu_exu_rsr_data_m[27]), .B(exu_n16263), .Y(bypass_sr_out_mux_n178));
INVX1 exu_U27997(.A(bypass_sr_out_mux_n178), .Y(exu_n9527));
AND2X1 exu_U27998(.A(exu_tlu_wsr_data_m[27]), .B(exu_n16264), .Y(bypass_sr_out_mux_n180));
INVX1 exu_U27999(.A(bypass_sr_out_mux_n180), .Y(exu_n9528));
AND2X1 exu_U28000(.A(tlu_exu_rsr_data_m[26]), .B(exu_n16263), .Y(bypass_sr_out_mux_n182));
INVX1 exu_U28001(.A(bypass_sr_out_mux_n182), .Y(exu_n9529));
AND2X1 exu_U28002(.A(exu_tlu_wsr_data_m[26]), .B(exu_n16264), .Y(bypass_sr_out_mux_n184));
INVX1 exu_U28003(.A(bypass_sr_out_mux_n184), .Y(exu_n9530));
AND2X1 exu_U28004(.A(tlu_exu_rsr_data_m[25]), .B(exu_n16263), .Y(bypass_sr_out_mux_n186));
INVX1 exu_U28005(.A(bypass_sr_out_mux_n186), .Y(exu_n9531));
AND2X1 exu_U28006(.A(exu_tlu_wsr_data_m[25]), .B(exu_n16264), .Y(bypass_sr_out_mux_n188));
INVX1 exu_U28007(.A(bypass_sr_out_mux_n188), .Y(exu_n9532));
AND2X1 exu_U28008(.A(tlu_exu_rsr_data_m[24]), .B(exu_n16263), .Y(bypass_sr_out_mux_n190));
INVX1 exu_U28009(.A(bypass_sr_out_mux_n190), .Y(exu_n9533));
AND2X1 exu_U28010(.A(exu_tlu_wsr_data_m[24]), .B(exu_n16264), .Y(bypass_sr_out_mux_n192));
INVX1 exu_U28011(.A(bypass_sr_out_mux_n192), .Y(exu_n9534));
AND2X1 exu_U28012(.A(tlu_exu_rsr_data_m[23]), .B(exu_n16263), .Y(bypass_sr_out_mux_n194));
INVX1 exu_U28013(.A(bypass_sr_out_mux_n194), .Y(exu_n9535));
AND2X1 exu_U28014(.A(exu_tlu_wsr_data_m[23]), .B(exu_n16264), .Y(bypass_sr_out_mux_n196));
INVX1 exu_U28015(.A(bypass_sr_out_mux_n196), .Y(exu_n9536));
AND2X1 exu_U28016(.A(tlu_exu_rsr_data_m[22]), .B(exu_n16263), .Y(bypass_sr_out_mux_n198));
INVX1 exu_U28017(.A(bypass_sr_out_mux_n198), .Y(exu_n9537));
AND2X1 exu_U28018(.A(exu_tlu_wsr_data_m[22]), .B(exu_n16264), .Y(bypass_sr_out_mux_n200));
INVX1 exu_U28019(.A(bypass_sr_out_mux_n200), .Y(exu_n9538));
AND2X1 exu_U28020(.A(tlu_exu_rsr_data_m[21]), .B(exu_n16263), .Y(bypass_sr_out_mux_n202));
INVX1 exu_U28021(.A(bypass_sr_out_mux_n202), .Y(exu_n9539));
AND2X1 exu_U28022(.A(exu_tlu_wsr_data_m[21]), .B(exu_n16264), .Y(bypass_sr_out_mux_n204));
INVX1 exu_U28023(.A(bypass_sr_out_mux_n204), .Y(exu_n9540));
AND2X1 exu_U28024(.A(tlu_exu_rsr_data_m[20]), .B(exu_n16263), .Y(bypass_sr_out_mux_n206));
INVX1 exu_U28025(.A(bypass_sr_out_mux_n206), .Y(exu_n9541));
AND2X1 exu_U28026(.A(exu_tlu_wsr_data_m[20]), .B(exu_n16264), .Y(bypass_sr_out_mux_n208));
INVX1 exu_U28027(.A(bypass_sr_out_mux_n208), .Y(exu_n9542));
AND2X1 exu_U28028(.A(tlu_exu_rsr_data_m[1]), .B(exu_n16263), .Y(bypass_sr_out_mux_n210));
INVX1 exu_U28029(.A(bypass_sr_out_mux_n210), .Y(exu_n9543));
AND2X1 exu_U28030(.A(ecl_byp_3lsb_m[1]), .B(exu_n16264), .Y(bypass_sr_out_mux_n212));
INVX1 exu_U28031(.A(bypass_sr_out_mux_n212), .Y(exu_n9544));
AND2X1 exu_U28032(.A(tlu_exu_rsr_data_m[19]), .B(exu_n16263), .Y(bypass_sr_out_mux_n214));
INVX1 exu_U28033(.A(bypass_sr_out_mux_n214), .Y(exu_n9545));
AND2X1 exu_U28034(.A(exu_tlu_wsr_data_m[19]), .B(exu_n16264), .Y(bypass_sr_out_mux_n216));
INVX1 exu_U28035(.A(bypass_sr_out_mux_n216), .Y(exu_n9546));
AND2X1 exu_U28036(.A(tlu_exu_rsr_data_m[18]), .B(exu_n16263), .Y(bypass_sr_out_mux_n218));
INVX1 exu_U28037(.A(bypass_sr_out_mux_n218), .Y(exu_n9547));
AND2X1 exu_U28038(.A(exu_tlu_wsr_data_m[18]), .B(exu_n16264), .Y(bypass_sr_out_mux_n220));
INVX1 exu_U28039(.A(bypass_sr_out_mux_n220), .Y(exu_n9548));
AND2X1 exu_U28040(.A(tlu_exu_rsr_data_m[17]), .B(exu_n16263), .Y(bypass_sr_out_mux_n222));
INVX1 exu_U28041(.A(bypass_sr_out_mux_n222), .Y(exu_n9549));
AND2X1 exu_U28042(.A(exu_tlu_wsr_data_m[17]), .B(exu_n16264), .Y(bypass_sr_out_mux_n224));
INVX1 exu_U28043(.A(bypass_sr_out_mux_n224), .Y(exu_n9550));
AND2X1 exu_U28044(.A(tlu_exu_rsr_data_m[16]), .B(exu_n16263), .Y(bypass_sr_out_mux_n226));
INVX1 exu_U28045(.A(bypass_sr_out_mux_n226), .Y(exu_n9551));
AND2X1 exu_U28046(.A(exu_tlu_wsr_data_m[16]), .B(exu_n16264), .Y(bypass_sr_out_mux_n228));
INVX1 exu_U28047(.A(bypass_sr_out_mux_n228), .Y(exu_n9552));
AND2X1 exu_U28048(.A(tlu_exu_rsr_data_m[15]), .B(exu_n16263), .Y(bypass_sr_out_mux_n230));
INVX1 exu_U28049(.A(bypass_sr_out_mux_n230), .Y(exu_n9553));
AND2X1 exu_U28050(.A(exu_tlu_wsr_data_m[15]), .B(exu_n16264), .Y(bypass_sr_out_mux_n232));
INVX1 exu_U28051(.A(bypass_sr_out_mux_n232), .Y(exu_n9554));
AND2X1 exu_U28052(.A(tlu_exu_rsr_data_m[14]), .B(exu_n16263), .Y(bypass_sr_out_mux_n234));
INVX1 exu_U28053(.A(bypass_sr_out_mux_n234), .Y(exu_n9555));
AND2X1 exu_U28054(.A(exu_tlu_wsr_data_m[14]), .B(exu_n16264), .Y(bypass_sr_out_mux_n236));
INVX1 exu_U28055(.A(bypass_sr_out_mux_n236), .Y(exu_n9556));
AND2X1 exu_U28056(.A(tlu_exu_rsr_data_m[13]), .B(exu_n16263), .Y(bypass_sr_out_mux_n238));
INVX1 exu_U28057(.A(bypass_sr_out_mux_n238), .Y(exu_n9557));
AND2X1 exu_U28058(.A(exu_tlu_wsr_data_m[13]), .B(exu_n16264), .Y(bypass_sr_out_mux_n240));
INVX1 exu_U28059(.A(bypass_sr_out_mux_n240), .Y(exu_n9558));
AND2X1 exu_U28060(.A(tlu_exu_rsr_data_m[12]), .B(exu_n16263), .Y(bypass_sr_out_mux_n242));
INVX1 exu_U28061(.A(bypass_sr_out_mux_n242), .Y(exu_n9559));
AND2X1 exu_U28062(.A(exu_tlu_wsr_data_m[12]), .B(exu_n16264), .Y(bypass_sr_out_mux_n244));
INVX1 exu_U28063(.A(bypass_sr_out_mux_n244), .Y(exu_n9560));
AND2X1 exu_U28064(.A(tlu_exu_rsr_data_m[11]), .B(exu_n16263), .Y(bypass_sr_out_mux_n246));
INVX1 exu_U28065(.A(bypass_sr_out_mux_n246), .Y(exu_n9561));
AND2X1 exu_U28066(.A(exu_tlu_wsr_data_m[11]), .B(exu_n16264), .Y(bypass_sr_out_mux_n248));
INVX1 exu_U28067(.A(bypass_sr_out_mux_n248), .Y(exu_n9562));
AND2X1 exu_U28068(.A(tlu_exu_rsr_data_m[10]), .B(exu_n16263), .Y(bypass_sr_out_mux_n250));
INVX1 exu_U28069(.A(bypass_sr_out_mux_n250), .Y(exu_n9563));
AND2X1 exu_U28070(.A(exu_tlu_wsr_data_m[10]), .B(exu_n16264), .Y(bypass_sr_out_mux_n252));
INVX1 exu_U28071(.A(bypass_sr_out_mux_n252), .Y(exu_n9564));
AND2X1 exu_U28072(.A(tlu_exu_rsr_data_m[0]), .B(exu_n16263), .Y(bypass_sr_out_mux_n254));
INVX1 exu_U28073(.A(bypass_sr_out_mux_n254), .Y(exu_n9565));
AND2X1 exu_U28074(.A(ecl_byp_3lsb_m[0]), .B(exu_n16264), .Y(bypass_sr_out_mux_n256));
INVX1 exu_U28075(.A(bypass_sr_out_mux_n256), .Y(exu_n9566));
AND2X1 exu_U28076(.A(exu_n16266), .B(ifu_exu_pcver_e[9]), .Y(bypass_ifu_exu_sr_mux_n4));
INVX1 exu_U28077(.A(bypass_ifu_exu_sr_mux_n4), .Y(exu_n9567));
AND2X1 exu_U28078(.A(ifu_exu_pcver_e[8]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n10));
INVX1 exu_U28079(.A(bypass_ifu_exu_sr_mux_n10), .Y(exu_n9568));
AND2X1 exu_U28080(.A(ifu_exu_pcver_e[7]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n16));
INVX1 exu_U28081(.A(bypass_ifu_exu_sr_mux_n16), .Y(exu_n9569));
AND2X1 exu_U28082(.A(div_byp_yreg_e[7]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n18));
INVX1 exu_U28083(.A(bypass_ifu_exu_sr_mux_n18), .Y(exu_n9570));
AND2X1 exu_U28084(.A(ifu_exu_pcver_e[6]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n22));
INVX1 exu_U28085(.A(bypass_ifu_exu_sr_mux_n22), .Y(exu_n9571));
AND2X1 exu_U28086(.A(div_byp_yreg_e[6]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n24));
INVX1 exu_U28087(.A(bypass_ifu_exu_sr_mux_n24), .Y(exu_n9572));
AND2X1 exu_U28088(.A(ifu_exu_pcver_e[5]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n52));
INVX1 exu_U28089(.A(bypass_ifu_exu_sr_mux_n52), .Y(exu_n9573));
AND2X1 exu_U28090(.A(div_byp_yreg_e[5]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n54));
INVX1 exu_U28091(.A(bypass_ifu_exu_sr_mux_n54), .Y(exu_n9574));
AND2X1 exu_U28092(.A(ifu_exu_pcver_e[4]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n118));
INVX1 exu_U28093(.A(bypass_ifu_exu_sr_mux_n118), .Y(exu_n9575));
AND2X1 exu_U28094(.A(div_byp_yreg_e[4]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n120));
INVX1 exu_U28095(.A(bypass_ifu_exu_sr_mux_n120), .Y(exu_n9576));
AND2X1 exu_U28096(.A(ifu_exu_pcver_e[3]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n184));
INVX1 exu_U28097(.A(bypass_ifu_exu_sr_mux_n184), .Y(exu_n9577));
AND2X1 exu_U28098(.A(div_byp_yreg_e[3]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n186));
INVX1 exu_U28099(.A(bypass_ifu_exu_sr_mux_n186), .Y(exu_n9578));
AND2X1 exu_U28100(.A(ifu_exu_pcver_e[31]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n238));
INVX1 exu_U28101(.A(bypass_ifu_exu_sr_mux_n238), .Y(exu_n9579));
AND2X1 exu_U28102(.A(ifu_exu_pcver_e[30]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n244));
INVX1 exu_U28103(.A(bypass_ifu_exu_sr_mux_n244), .Y(exu_n9580));
AND2X1 exu_U28104(.A(ifu_exu_pcver_e[2]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n250));
INVX1 exu_U28105(.A(bypass_ifu_exu_sr_mux_n250), .Y(exu_n9581));
AND2X1 exu_U28106(.A(div_byp_yreg_e[2]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n252));
INVX1 exu_U28107(.A(bypass_ifu_exu_sr_mux_n252), .Y(exu_n9582));
AND2X1 exu_U28108(.A(ifu_exu_pcver_e[29]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n256));
INVX1 exu_U28109(.A(bypass_ifu_exu_sr_mux_n256), .Y(exu_n9583));
AND2X1 exu_U28110(.A(ifu_exu_pcver_e[28]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n262));
INVX1 exu_U28111(.A(bypass_ifu_exu_sr_mux_n262), .Y(exu_n9584));
AND2X1 exu_U28112(.A(ifu_exu_pcver_e[27]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n268));
INVX1 exu_U28113(.A(bypass_ifu_exu_sr_mux_n268), .Y(exu_n9585));
AND2X1 exu_U28114(.A(ifu_exu_pcver_e[26]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n274));
INVX1 exu_U28115(.A(bypass_ifu_exu_sr_mux_n274), .Y(exu_n9586));
AND2X1 exu_U28116(.A(ifu_exu_pcver_e[25]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n280));
INVX1 exu_U28117(.A(bypass_ifu_exu_sr_mux_n280), .Y(exu_n9587));
AND2X1 exu_U28118(.A(ifu_exu_pcver_e[24]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n286));
INVX1 exu_U28119(.A(bypass_ifu_exu_sr_mux_n286), .Y(exu_n9588));
AND2X1 exu_U28120(.A(ifu_exu_pcver_e[23]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n292));
INVX1 exu_U28121(.A(bypass_ifu_exu_sr_mux_n292), .Y(exu_n9589));
AND2X1 exu_U28122(.A(ifu_exu_pcver_e[22]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n298));
INVX1 exu_U28123(.A(bypass_ifu_exu_sr_mux_n298), .Y(exu_n9590));
AND2X1 exu_U28124(.A(ifu_exu_pcver_e[21]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n304));
INVX1 exu_U28125(.A(bypass_ifu_exu_sr_mux_n304), .Y(exu_n9591));
AND2X1 exu_U28126(.A(ifu_exu_pcver_e[20]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n310));
INVX1 exu_U28127(.A(bypass_ifu_exu_sr_mux_n310), .Y(exu_n9592));
AND2X1 exu_U28128(.A(ifu_exu_pcver_e[1]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n316));
INVX1 exu_U28129(.A(bypass_ifu_exu_sr_mux_n316), .Y(exu_n9593));
AND2X1 exu_U28130(.A(div_byp_yreg_e[1]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n318));
INVX1 exu_U28131(.A(bypass_ifu_exu_sr_mux_n318), .Y(exu_n9594));
AND2X1 exu_U28132(.A(ifu_exu_pcver_e[19]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n322));
INVX1 exu_U28133(.A(bypass_ifu_exu_sr_mux_n322), .Y(exu_n9595));
AND2X1 exu_U28134(.A(ifu_exu_pcver_e[18]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n328));
INVX1 exu_U28135(.A(bypass_ifu_exu_sr_mux_n328), .Y(exu_n9596));
AND2X1 exu_U28136(.A(ifu_exu_pcver_e[17]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n334));
INVX1 exu_U28137(.A(bypass_ifu_exu_sr_mux_n334), .Y(exu_n9597));
AND2X1 exu_U28138(.A(ifu_exu_pcver_e[16]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n340));
INVX1 exu_U28139(.A(bypass_ifu_exu_sr_mux_n340), .Y(exu_n9598));
AND2X1 exu_U28140(.A(ifu_exu_pcver_e[15]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n346));
INVX1 exu_U28141(.A(bypass_ifu_exu_sr_mux_n346), .Y(exu_n9599));
AND2X1 exu_U28142(.A(ifu_exu_pcver_e[14]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n352));
INVX1 exu_U28143(.A(bypass_ifu_exu_sr_mux_n352), .Y(exu_n9600));
AND2X1 exu_U28144(.A(ifu_exu_pcver_e[13]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n358));
INVX1 exu_U28145(.A(bypass_ifu_exu_sr_mux_n358), .Y(exu_n9601));
AND2X1 exu_U28146(.A(ifu_exu_pcver_e[12]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n364));
INVX1 exu_U28147(.A(bypass_ifu_exu_sr_mux_n364), .Y(exu_n9602));
AND2X1 exu_U28148(.A(ifu_exu_pcver_e[11]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n370));
INVX1 exu_U28149(.A(bypass_ifu_exu_sr_mux_n370), .Y(exu_n9603));
AND2X1 exu_U28150(.A(ifu_exu_pcver_e[10]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n376));
INVX1 exu_U28151(.A(bypass_ifu_exu_sr_mux_n376), .Y(exu_n9604));
AND2X1 exu_U28152(.A(ifu_exu_pcver_e[0]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n382));
INVX1 exu_U28153(.A(bypass_ifu_exu_sr_mux_n382), .Y(exu_n9605));
AND2X1 exu_U28154(.A(div_byp_yreg_e[0]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n384));
INVX1 exu_U28155(.A(bypass_ifu_exu_sr_mux_n384), .Y(exu_n9606));
AND2X1 exu_U28156(.A(exu_n11850), .B(rml_rml_ecl_cwp_e[1]), .Y(rml_n39));
INVX1 exu_U28157(.A(rml_n39), .Y(exu_n9607));
AND2X1 exu_U28158(.A(rml_rml_ecl_cleanwin_e[1]), .B(rml_rml_ecl_cleanwin_e[0]), .Y(rml_n45));
INVX1 exu_U28159(.A(rml_n45), .Y(exu_n9608));
AND2X1 exu_U28160(.A(ifu_exu_flushw_e), .B(exu_n15685), .Y(rml_n61));
INVX1 exu_U28161(.A(rml_n61), .Y(exu_n9609));
AND2X1 exu_U28162(.A(rml_agp_thr2[1]), .B(exu_n15470), .Y(rml_n65));
INVX1 exu_U28163(.A(rml_n65), .Y(exu_n9610));
AND2X1 exu_U28164(.A(rml_agp_thr0[1]), .B(rml_n77), .Y(rml_n69));
INVX1 exu_U28165(.A(rml_n69), .Y(exu_n9611));
AND2X1 exu_U28166(.A(rml_agp_thr2[0]), .B(exu_n15470), .Y(rml_n74));
INVX1 exu_U28167(.A(rml_n74), .Y(exu_n9612));
AND2X1 exu_U28168(.A(rml_agp_thr0[0]), .B(rml_n77), .Y(rml_n76));
INVX1 exu_U28169(.A(rml_n76), .Y(exu_n9613));
AND2X1 exu_U28170(.A(exu_n16385), .B(exu_n16383), .Y(rml_n94));
INVX1 exu_U28171(.A(rml_n94), .Y(exu_n9614));
AND2X1 exu_U28172(.A(exu_n15383), .B(rml_exu_tlu_spill_e), .Y(rml_n98));
INVX1 exu_U28173(.A(rml_n98), .Y(exu_n9615));
AND2X1 exu_U28174(.A(rml_n101), .B(rml_rml_ecl_cleanwin_e[1]), .Y(rml_n100));
INVX1 exu_U28175(.A(rml_n100), .Y(exu_n9616));
AND2X1 exu_U28176(.A(exu_n11859), .B(rml_save_e), .Y(rml_n112));
INVX1 exu_U28177(.A(rml_n112), .Y(exu_n9617));
OR2X1 exu_U28178(.A(rml_n117), .B(exu_n14977), .Y(rml_n116));
INVX1 exu_U28179(.A(rml_n116), .Y(exu_n9618));
AND2X1 exu_U28180(.A(exu_n11860), .B(rml_rml_ecl_cansave_e[2]), .Y(rml_n119));
INVX1 exu_U28181(.A(rml_n119), .Y(exu_n9619));
OR2X1 exu_U28182(.A(exu_n12069), .B(exu_n14978), .Y(div_n40));
INVX1 exu_U28183(.A(div_n40), .Y(exu_n9620));
OR2X1 exu_U28184(.A(exu_n12033), .B(exu_n14921), .Y(div_n44));
INVX1 exu_U28185(.A(div_n44), .Y(exu_n9621));
OR2X1 exu_U28186(.A(exu_n12031), .B(exu_n14919), .Y(div_n46));
INVX1 exu_U28187(.A(div_n46), .Y(exu_n9622));
OR2X1 exu_U28188(.A(exu_n12037), .B(exu_n14925), .Y(div_n50));
INVX1 exu_U28189(.A(div_n50), .Y(exu_n9623));
OR2X1 exu_U28190(.A(exu_n12035), .B(exu_n14923), .Y(div_n52));
INVX1 exu_U28191(.A(div_n52), .Y(exu_n9624));
OR2X1 exu_U28192(.A(exu_n12071), .B(exu_n14980), .Y(div_n54));
INVX1 exu_U28193(.A(div_n54), .Y(exu_n9625));
OR2X1 exu_U28194(.A(exu_n12011), .B(exu_n14904), .Y(div_n58));
INVX1 exu_U28195(.A(div_n58), .Y(exu_n9626));
OR2X1 exu_U28196(.A(exu_n12007), .B(exu_n14895), .Y(div_n60));
INVX1 exu_U28197(.A(div_n60), .Y(exu_n9627));
OR2X1 exu_U28198(.A(exu_n12029), .B(exu_n14917), .Y(div_n64));
INVX1 exu_U28199(.A(div_n64), .Y(exu_n9628));
OR2X1 exu_U28200(.A(exu_n12027), .B(exu_n14915), .Y(div_n66));
INVX1 exu_U28201(.A(div_n66), .Y(exu_n9629));
OR2X1 exu_U28202(.A(exu_n12073), .B(exu_n14982), .Y(div_n70));
INVX1 exu_U28203(.A(div_n70), .Y(exu_n9630));
OR2X1 exu_U28204(.A(exu_n12020), .B(exu_n14908), .Y(div_n74));
INVX1 exu_U28205(.A(div_n74), .Y(exu_n9631));
OR2X1 exu_U28206(.A(exu_n12018), .B(exu_n14906), .Y(div_n76));
INVX1 exu_U28207(.A(div_n76), .Y(exu_n9632));
OR2X1 exu_U28208(.A(exu_n12025), .B(exu_n14912), .Y(div_n80));
INVX1 exu_U28209(.A(div_n80), .Y(exu_n9633));
OR2X1 exu_U28210(.A(exu_n12023), .B(exu_n14910), .Y(div_n82));
INVX1 exu_U28211(.A(div_n82), .Y(exu_n9634));
OR2X1 exu_U28212(.A(exu_n12075), .B(exu_n14984), .Y(div_n84));
INVX1 exu_U28213(.A(div_n84), .Y(exu_n9635));
OR2X1 exu_U28214(.A(exu_n12012), .B(exu_n14899), .Y(div_n88));
INVX1 exu_U28215(.A(div_n88), .Y(exu_n9636));
OR2X1 exu_U28216(.A(exu_n12009), .B(exu_n14897), .Y(div_n90));
INVX1 exu_U28217(.A(div_n90), .Y(exu_n9637));
OR2X1 exu_U28218(.A(exu_n12016), .B(exu_n14903), .Y(div_n94));
INVX1 exu_U28219(.A(div_n94), .Y(exu_n9638));
OR2X1 exu_U28220(.A(exu_n12014), .B(exu_n14901), .Y(div_n96));
INVX1 exu_U28221(.A(div_n96), .Y(exu_n9639));
OR2X1 exu_U28222(.A(exu_n12077), .B(exu_n14986), .Y(alu_n72));
INVX1 exu_U28223(.A(alu_n72), .Y(exu_n9640));
OR2X1 exu_U28224(.A(exu_n11985), .B(exu_n14874), .Y(alu_n76));
INVX1 exu_U28225(.A(alu_n76), .Y(exu_n9641));
OR2X1 exu_U28226(.A(exu_n11983), .B(exu_n14872), .Y(alu_n78));
INVX1 exu_U28227(.A(alu_n78), .Y(exu_n9642));
OR2X1 exu_U28228(.A(exu_n11989), .B(exu_n14878), .Y(alu_n82));
INVX1 exu_U28229(.A(alu_n82), .Y(exu_n9643));
OR2X1 exu_U28230(.A(exu_n11987), .B(exu_n14876), .Y(alu_n84));
INVX1 exu_U28231(.A(alu_n84), .Y(exu_n9644));
OR2X1 exu_U28232(.A(exu_n12079), .B(exu_n14988), .Y(alu_n86));
INVX1 exu_U28233(.A(alu_n86), .Y(exu_n9645));
OR2X1 exu_U28234(.A(exu_n11963), .B(exu_n14857), .Y(alu_n90));
INVX1 exu_U28235(.A(alu_n90), .Y(exu_n9646));
OR2X1 exu_U28236(.A(exu_n11959), .B(exu_n14848), .Y(alu_n92));
INVX1 exu_U28237(.A(alu_n92), .Y(exu_n9647));
OR2X1 exu_U28238(.A(exu_n11981), .B(exu_n14870), .Y(alu_n96));
INVX1 exu_U28239(.A(alu_n96), .Y(exu_n9648));
OR2X1 exu_U28240(.A(exu_n11979), .B(exu_n14868), .Y(alu_n98));
INVX1 exu_U28241(.A(alu_n98), .Y(exu_n9649));
OR2X1 exu_U28242(.A(exu_n12083), .B(exu_n14990), .Y(alu_ecl_zhigh_e));
INVX1 exu_U28243(.A(alu_ecl_zhigh_e), .Y(exu_n9650));
OR2X1 exu_U28244(.A(exu_n12081), .B(exu_n14991), .Y(alu_n102));
INVX1 exu_U28245(.A(alu_n102), .Y(exu_n9651));
OR2X1 exu_U28246(.A(exu_n11972), .B(exu_n14861), .Y(alu_n106));
INVX1 exu_U28247(.A(alu_n106), .Y(exu_n9652));
OR2X1 exu_U28248(.A(exu_n11970), .B(exu_n14859), .Y(alu_n108));
INVX1 exu_U28249(.A(alu_n108), .Y(exu_n9653));
OR2X1 exu_U28250(.A(exu_n11977), .B(exu_n14865), .Y(alu_n112));
INVX1 exu_U28251(.A(alu_n112), .Y(exu_n9654));
OR2X1 exu_U28252(.A(exu_n11975), .B(exu_n14863), .Y(alu_n114));
INVX1 exu_U28253(.A(alu_n114), .Y(exu_n9655));
OR2X1 exu_U28254(.A(exu_n12084), .B(exu_n14993), .Y(alu_n116));
INVX1 exu_U28255(.A(alu_n116), .Y(exu_n9656));
OR2X1 exu_U28256(.A(exu_n11964), .B(exu_n14852), .Y(alu_n120));
INVX1 exu_U28257(.A(alu_n120), .Y(exu_n9657));
OR2X1 exu_U28258(.A(exu_n11961), .B(exu_n14850), .Y(alu_n122));
INVX1 exu_U28259(.A(alu_n122), .Y(exu_n9658));
OR2X1 exu_U28260(.A(exu_n11968), .B(exu_n14856), .Y(alu_n126));
INVX1 exu_U28261(.A(alu_n126), .Y(exu_n9659));
OR2X1 exu_U28262(.A(exu_n11966), .B(exu_n14854), .Y(alu_n128));
INVX1 exu_U28263(.A(alu_n128), .Y(exu_n9660));
OR2X1 exu_U28264(.A(ifu_exu_enshift_d), .B(ifu_exu_aluop_d[2]), .Y(ecl_n78));
INVX1 exu_U28265(.A(ecl_n78), .Y(exu_n9661));
AND2X1 exu_U28266(.A(exu_n15921), .B(ecl_perr_store[3]), .Y(ecl_n85));
INVX1 exu_U28267(.A(ecl_n85), .Y(exu_n9662));
AND2X1 exu_U28268(.A(exu_n15923), .B(ecl_perr_store[1]), .Y(ecl_n87));
INVX1 exu_U28269(.A(ecl_n87), .Y(exu_n9663));
OR2X1 exu_U28270(.A(ifu_exu_ttype_vld_m), .B(exu_n14995), .Y(ecl_n89));
INVX1 exu_U28271(.A(ecl_n89), .Y(exu_n9664));
AND2X1 exu_U28272(.A(exu_n16372), .B(exu_n10706), .Y(ecl_n94));
INVX1 exu_U28273(.A(ecl_n94), .Y(exu_n9665));
AND2X1 exu_U28274(.A(ecl_n98), .B(tlu_exu_pic_onebelow_m), .Y(ecl_n100));
INVX1 exu_U28275(.A(ecl_n100), .Y(exu_n9666));
AND2X1 exu_U28276(.A(ecl_n104), .B(alu_logic_rs1_data_bf1[63]), .Y(ecl_n103));
INVX1 exu_U28277(.A(ecl_n103), .Y(exu_n9667));
AND2X1 exu_U28278(.A(exu_n16400), .B(exu_n16401), .Y(ecl_n108));
INVX1 exu_U28279(.A(ecl_n108), .Y(exu_n9668));
AND2X1 exu_U28280(.A(ecl_n116), .B(rml_ecl_fill_e), .Y(ecl_n115));
INVX1 exu_U28281(.A(ecl_n115), .Y(exu_n9669));
AND2X1 exu_U28282(.A(exu_n11931), .B(exu_n16213), .Y(ecl_n118));
INVX1 exu_U28283(.A(ecl_n118), .Y(exu_n9670));
AND2X1 exu_U28284(.A(rml_ecl_clean_window_e), .B(rml_ecl_fill_e), .Y(ecl_n122));
INVX1 exu_U28285(.A(ecl_n122), .Y(exu_n9671));
AND2X1 exu_U28286(.A(ifu_exu_dontmv_regz0_e), .B(exu_n31738), .Y(ecl_n125));
INVX1 exu_U28287(.A(ecl_n125), .Y(exu_n9672));
AND2X1 exu_U28288(.A(alu_ecl_add_n64_e), .B(exu_n16155), .Y(ecl_n127));
INVX1 exu_U28289(.A(ecl_n127), .Y(exu_n9673));
AND2X1 exu_U28290(.A(exu_ifu_brpc_e[31]), .B(exu_n16157), .Y(ecl_n129));
INVX1 exu_U28291(.A(ecl_n129), .Y(exu_n9674));
AND2X1 exu_U28292(.A(exu_n16627), .B(exu_n16560), .Y(exu_n16628));
INVX1 exu_U28293(.A(exu_n16628), .Y(exu_n9675));
AND2X1 exu_U28294(.A(ecl_wb_byplog_rd_g2[1]), .B(exu_n15222), .Y(exu_n16631));
INVX1 exu_U28295(.A(exu_n16631), .Y(exu_n9676));
AND2X1 exu_U28296(.A(exu_n16641), .B(exu_n16566), .Y(exu_n16642));
INVX1 exu_U28297(.A(exu_n16642), .Y(exu_n9677));
AND2X1 exu_U28298(.A(ecl_ld_rd_g[1]), .B(exu_n15223), .Y(exu_n16645));
INVX1 exu_U28299(.A(exu_n16645), .Y(exu_n9678));
AND2X1 exu_U28300(.A(exu_n16655), .B(exu_n16562), .Y(exu_n16656));
INVX1 exu_U28301(.A(exu_n16656), .Y(exu_n9679));
AND2X1 exu_U28302(.A(ecl_rd_m[1]), .B(exu_n15224), .Y(exu_n16659));
INVX1 exu_U28303(.A(exu_n16659), .Y(exu_n9680));
AND2X1 exu_U28304(.A(exu_n16669), .B(exu_n16564), .Y(exu_n16670));
INVX1 exu_U28305(.A(exu_n16670), .Y(exu_n9681));
AND2X1 exu_U28306(.A(ecl_rd_e[1]), .B(exu_n15225), .Y(exu_n16673));
INVX1 exu_U28307(.A(exu_n16673), .Y(exu_n9682));
AND2X1 exu_U28308(.A(exu_n16683), .B(exu_n16560), .Y(exu_n16684));
INVX1 exu_U28309(.A(exu_n16684), .Y(exu_n9683));
AND2X1 exu_U28310(.A(ecl_wb_byplog_rd_g2[1]), .B(exu_n15226), .Y(exu_n16687));
INVX1 exu_U28311(.A(exu_n16687), .Y(exu_n9684));
AND2X1 exu_U28312(.A(exu_n16697), .B(exu_n16566), .Y(exu_n16698));
INVX1 exu_U28313(.A(exu_n16698), .Y(exu_n9685));
AND2X1 exu_U28314(.A(ecl_ld_rd_g[1]), .B(exu_n15227), .Y(exu_n16701));
INVX1 exu_U28315(.A(exu_n16701), .Y(exu_n9686));
AND2X1 exu_U28316(.A(exu_n16711), .B(exu_n16562), .Y(exu_n16712));
INVX1 exu_U28317(.A(exu_n16712), .Y(exu_n9687));
AND2X1 exu_U28318(.A(ecl_rd_m[1]), .B(exu_n15228), .Y(exu_n16715));
INVX1 exu_U28319(.A(exu_n16715), .Y(exu_n9688));
AND2X1 exu_U28320(.A(exu_n16725), .B(exu_n16564), .Y(exu_n16726));
INVX1 exu_U28321(.A(exu_n16726), .Y(exu_n9689));
AND2X1 exu_U28322(.A(ecl_rd_e[1]), .B(exu_n15229), .Y(exu_n16729));
INVX1 exu_U28323(.A(exu_n16729), .Y(exu_n9690));
AND2X1 exu_U28324(.A(exu_n17403), .B(exu_n16560), .Y(exu_n17404));
INVX1 exu_U28325(.A(exu_n17404), .Y(exu_n9691));
AND2X1 exu_U28326(.A(ecl_wb_byplog_rd_g2[1]), .B(exu_n15230), .Y(exu_n17407));
INVX1 exu_U28327(.A(exu_n17407), .Y(exu_n9692));
AND2X1 exu_U28328(.A(exu_n17417), .B(exu_n16566), .Y(exu_n17418));
INVX1 exu_U28329(.A(exu_n17418), .Y(exu_n9693));
AND2X1 exu_U28330(.A(ecl_ld_rd_g[1]), .B(exu_n15231), .Y(exu_n17421));
INVX1 exu_U28331(.A(exu_n17421), .Y(exu_n9694));
AND2X1 exu_U28332(.A(exu_n17431), .B(exu_n16562), .Y(exu_n17432));
INVX1 exu_U28333(.A(exu_n17432), .Y(exu_n9695));
AND2X1 exu_U28334(.A(ecl_rd_m[1]), .B(exu_n15232), .Y(exu_n17435));
INVX1 exu_U28335(.A(exu_n17435), .Y(exu_n9696));
AND2X1 exu_U28336(.A(exu_n17445), .B(exu_n16564), .Y(exu_n17446));
INVX1 exu_U28337(.A(exu_n17446), .Y(exu_n9697));
AND2X1 exu_U28338(.A(ecl_rd_e[1]), .B(exu_n15233), .Y(exu_n17449));
INVX1 exu_U28339(.A(exu_n17449), .Y(exu_n9698));
AND2X1 exu_U28340(.A(rml_cwp_n43), .B(rml_cwp_swap_slot1_data[9]), .Y(exu_n17506));
INVX1 exu_U28341(.A(exu_n17506), .Y(exu_n9699));
AND2X1 exu_U28342(.A(rml_cwp_swap_slot1_data[8]), .B(rml_cwp_n43), .Y(exu_n17508));
INVX1 exu_U28343(.A(exu_n17508), .Y(exu_n9700));
AND2X1 exu_U28344(.A(rml_cwp_swap_slot1_data[7]), .B(rml_cwp_n43), .Y(exu_n17510));
INVX1 exu_U28345(.A(exu_n17510), .Y(exu_n9701));
AND2X1 exu_U28346(.A(rml_cwp_swap_slot1_data[6]), .B(rml_cwp_n43), .Y(exu_n17511));
INVX1 exu_U28347(.A(exu_n17511), .Y(exu_n9702));
AND2X1 exu_U28348(.A(rml_cwp_swap_slot1_data[5]), .B(rml_cwp_n43), .Y(exu_n17514));
INVX1 exu_U28349(.A(exu_n17514), .Y(exu_n9703));
AND2X1 exu_U28350(.A(rml_cwp_swap_slot1_data[4]), .B(rml_cwp_n43), .Y(exu_n17518));
INVX1 exu_U28351(.A(exu_n17518), .Y(exu_n9704));
AND2X1 exu_U28352(.A(rml_cwp_swap_slot1_data[3]), .B(rml_cwp_n43), .Y(exu_n17522));
INVX1 exu_U28353(.A(exu_n17522), .Y(exu_n9705));
AND2X1 exu_U28354(.A(rml_cwp_swap_slot1_data[2]), .B(rml_cwp_n43), .Y(exu_n17526));
INVX1 exu_U28355(.A(exu_n17526), .Y(exu_n9706));
AND2X1 exu_U28356(.A(rml_cwp_swap_slot1_data[1]), .B(rml_cwp_n43), .Y(exu_n17530));
INVX1 exu_U28357(.A(exu_n17530), .Y(exu_n9707));
AND2X1 exu_U28358(.A(rml_cwp_swap_slot1_data[12]), .B(rml_cwp_n43), .Y(exu_n17533));
INVX1 exu_U28359(.A(exu_n17533), .Y(exu_n9708));
AND2X1 exu_U28360(.A(rml_cwp_swap_slot1_data[11]), .B(rml_cwp_n43), .Y(exu_n17535));
INVX1 exu_U28361(.A(exu_n17535), .Y(exu_n9709));
AND2X1 exu_U28362(.A(rml_cwp_swap_slot1_data[10]), .B(rml_cwp_n43), .Y(exu_n17537));
INVX1 exu_U28363(.A(exu_n17537), .Y(exu_n9710));
AND2X1 exu_U28364(.A(rml_cwp_swap_slot1_data[0]), .B(rml_cwp_n43), .Y(exu_n17540));
INVX1 exu_U28365(.A(exu_n17540), .Y(exu_n9711));
AND2X1 exu_U28366(.A(rml_cwp_n41), .B(rml_cwp_swap_slot2_data[9]), .Y(exu_n17543));
INVX1 exu_U28367(.A(exu_n17543), .Y(exu_n9712));
AND2X1 exu_U28368(.A(rml_cwp_swap_slot2_data[8]), .B(rml_cwp_n41), .Y(exu_n17545));
INVX1 exu_U28369(.A(exu_n17545), .Y(exu_n9713));
AND2X1 exu_U28370(.A(rml_cwp_swap_slot2_data[7]), .B(rml_cwp_n41), .Y(exu_n17547));
INVX1 exu_U28371(.A(exu_n17547), .Y(exu_n9714));
AND2X1 exu_U28372(.A(rml_cwp_swap_slot2_data[6]), .B(rml_cwp_n41), .Y(exu_n17548));
INVX1 exu_U28373(.A(exu_n17548), .Y(exu_n9715));
AND2X1 exu_U28374(.A(rml_cwp_swap_slot2_data[5]), .B(rml_cwp_n41), .Y(exu_n17551));
INVX1 exu_U28375(.A(exu_n17551), .Y(exu_n9716));
AND2X1 exu_U28376(.A(rml_cwp_swap_slot2_data[4]), .B(rml_cwp_n41), .Y(exu_n17555));
INVX1 exu_U28377(.A(exu_n17555), .Y(exu_n9717));
AND2X1 exu_U28378(.A(rml_cwp_swap_slot2_data[3]), .B(rml_cwp_n41), .Y(exu_n17559));
INVX1 exu_U28379(.A(exu_n17559), .Y(exu_n9718));
AND2X1 exu_U28380(.A(rml_cwp_swap_slot2_data[2]), .B(rml_cwp_n41), .Y(exu_n17563));
INVX1 exu_U28381(.A(exu_n17563), .Y(exu_n9719));
AND2X1 exu_U28382(.A(rml_cwp_swap_slot2_data[1]), .B(rml_cwp_n41), .Y(exu_n17567));
INVX1 exu_U28383(.A(exu_n17567), .Y(exu_n9720));
AND2X1 exu_U28384(.A(rml_cwp_swap_slot2_data[12]), .B(rml_cwp_n41), .Y(exu_n17570));
INVX1 exu_U28385(.A(exu_n17570), .Y(exu_n9721));
AND2X1 exu_U28386(.A(rml_cwp_swap_slot2_data[11]), .B(rml_cwp_n41), .Y(exu_n17572));
INVX1 exu_U28387(.A(exu_n17572), .Y(exu_n9722));
AND2X1 exu_U28388(.A(rml_cwp_swap_slot2_data[10]), .B(rml_cwp_n41), .Y(exu_n17574));
INVX1 exu_U28389(.A(exu_n17574), .Y(exu_n9723));
AND2X1 exu_U28390(.A(rml_cwp_swap_slot2_data[0]), .B(rml_cwp_n41), .Y(exu_n17577));
INVX1 exu_U28391(.A(exu_n17577), .Y(exu_n9724));
AND2X1 exu_U28392(.A(rml_cwp_n39), .B(rml_cwp_swap_slot3_data[9]), .Y(exu_n17580));
INVX1 exu_U28393(.A(exu_n17580), .Y(exu_n9725));
AND2X1 exu_U28394(.A(rml_cwp_swap_slot3_data[8]), .B(rml_cwp_n39), .Y(exu_n17582));
INVX1 exu_U28395(.A(exu_n17582), .Y(exu_n9726));
AND2X1 exu_U28396(.A(rml_cwp_swap_slot3_data[7]), .B(rml_cwp_n39), .Y(exu_n17584));
INVX1 exu_U28397(.A(exu_n17584), .Y(exu_n9727));
AND2X1 exu_U28398(.A(rml_cwp_swap_slot3_data[6]), .B(rml_cwp_n39), .Y(exu_n17585));
INVX1 exu_U28399(.A(exu_n17585), .Y(exu_n9728));
AND2X1 exu_U28400(.A(rml_cwp_swap_slot3_data[5]), .B(rml_cwp_n39), .Y(exu_n17588));
INVX1 exu_U28401(.A(exu_n17588), .Y(exu_n9729));
AND2X1 exu_U28402(.A(rml_cwp_swap_slot3_data[4]), .B(rml_cwp_n39), .Y(exu_n17592));
INVX1 exu_U28403(.A(exu_n17592), .Y(exu_n9730));
AND2X1 exu_U28404(.A(rml_cwp_swap_slot3_data[3]), .B(rml_cwp_n39), .Y(exu_n17596));
INVX1 exu_U28405(.A(exu_n17596), .Y(exu_n9731));
AND2X1 exu_U28406(.A(rml_cwp_swap_slot3_data[2]), .B(rml_cwp_n39), .Y(exu_n17600));
INVX1 exu_U28407(.A(exu_n17600), .Y(exu_n9732));
AND2X1 exu_U28408(.A(rml_cwp_swap_slot3_data[1]), .B(rml_cwp_n39), .Y(exu_n17604));
INVX1 exu_U28409(.A(exu_n17604), .Y(exu_n9733));
AND2X1 exu_U28410(.A(rml_cwp_swap_slot3_data[12]), .B(rml_cwp_n39), .Y(exu_n17607));
INVX1 exu_U28411(.A(exu_n17607), .Y(exu_n9734));
AND2X1 exu_U28412(.A(rml_cwp_swap_slot3_data[11]), .B(rml_cwp_n39), .Y(exu_n17609));
INVX1 exu_U28413(.A(exu_n17609), .Y(exu_n9735));
AND2X1 exu_U28414(.A(rml_cwp_swap_slot3_data[10]), .B(rml_cwp_n39), .Y(exu_n17611));
INVX1 exu_U28415(.A(exu_n17611), .Y(exu_n9736));
AND2X1 exu_U28416(.A(rml_cwp_swap_slot3_data[0]), .B(rml_cwp_n39), .Y(exu_n17614));
INVX1 exu_U28417(.A(exu_n17614), .Y(exu_n9737));
AND2X1 exu_U28418(.A(exu_n10779), .B(div_ecl_cout64), .Y(exu_n17618));
INVX1 exu_U28419(.A(exu_n17618), .Y(exu_n9738));
AND2X1 exu_U28420(.A(ecl_ifu_exu_rs3_m[2]), .B(ecl_ecc_log_rs3_m), .Y(exu_n17717));
INVX1 exu_U28421(.A(exu_n17717), .Y(exu_n9739));
AND2X1 exu_U28422(.A(ecl_ifu_exu_rs3_m[1]), .B(ecl_ecc_log_rs3_m), .Y(exu_n17721));
INVX1 exu_U28423(.A(exu_n17721), .Y(exu_n9740));
AND2X1 exu_U28424(.A(ecl_ifu_exu_rs3_m[0]), .B(ecl_ecc_log_rs3_m), .Y(exu_n17725));
INVX1 exu_U28425(.A(exu_n17725), .Y(exu_n9741));
AND2X1 exu_U28426(.A(ecl_ccr_mux_ccrin1_sel2), .B(exu_tlu_ccr1_w[7]), .Y(exu_n18038));
INVX1 exu_U28427(.A(exu_n18038), .Y(exu_n9742));
AND2X1 exu_U28428(.A(exu_tlu_ccr1_w[6]), .B(ecl_ccr_mux_ccrin1_sel2), .Y(exu_n18042));
INVX1 exu_U28429(.A(exu_n18042), .Y(exu_n9743));
AND2X1 exu_U28430(.A(exu_tlu_ccr1_w[5]), .B(ecl_ccr_mux_ccrin1_sel2), .Y(exu_n18045));
INVX1 exu_U28431(.A(exu_n18045), .Y(exu_n9744));
AND2X1 exu_U28432(.A(exu_tlu_ccr1_w[4]), .B(ecl_ccr_mux_ccrin1_sel2), .Y(exu_n18047));
INVX1 exu_U28433(.A(exu_n18047), .Y(exu_n9745));
AND2X1 exu_U28434(.A(exu_tlu_ccr1_w[3]), .B(ecl_ccr_mux_ccrin1_sel2), .Y(exu_n18050));
INVX1 exu_U28435(.A(exu_n18050), .Y(exu_n9746));
AND2X1 exu_U28436(.A(exu_tlu_ccr1_w[2]), .B(ecl_ccr_mux_ccrin1_sel2), .Y(exu_n18054));
INVX1 exu_U28437(.A(exu_n18054), .Y(exu_n9747));
AND2X1 exu_U28438(.A(exu_tlu_ccr1_w[1]), .B(ecl_ccr_mux_ccrin1_sel2), .Y(exu_n18058));
INVX1 exu_U28439(.A(exu_n18058), .Y(exu_n9748));
AND2X1 exu_U28440(.A(exu_tlu_ccr1_w[0]), .B(ecl_ccr_mux_ccrin1_sel2), .Y(exu_n18062));
INVX1 exu_U28441(.A(exu_n18062), .Y(exu_n9749));
AND2X1 exu_U28442(.A(ecl_ccr_mux_ccrin2_sel2), .B(exu_tlu_ccr2_w[7]), .Y(exu_n18066));
INVX1 exu_U28443(.A(exu_n18066), .Y(exu_n9750));
AND2X1 exu_U28444(.A(exu_tlu_ccr2_w[6]), .B(ecl_ccr_mux_ccrin2_sel2), .Y(exu_n18070));
INVX1 exu_U28445(.A(exu_n18070), .Y(exu_n9751));
AND2X1 exu_U28446(.A(exu_tlu_ccr2_w[5]), .B(ecl_ccr_mux_ccrin2_sel2), .Y(exu_n18073));
INVX1 exu_U28447(.A(exu_n18073), .Y(exu_n9752));
AND2X1 exu_U28448(.A(exu_tlu_ccr2_w[4]), .B(ecl_ccr_mux_ccrin2_sel2), .Y(exu_n18075));
INVX1 exu_U28449(.A(exu_n18075), .Y(exu_n9753));
AND2X1 exu_U28450(.A(exu_tlu_ccr2_w[3]), .B(ecl_ccr_mux_ccrin2_sel2), .Y(exu_n18078));
INVX1 exu_U28451(.A(exu_n18078), .Y(exu_n9754));
AND2X1 exu_U28452(.A(exu_tlu_ccr2_w[2]), .B(ecl_ccr_mux_ccrin2_sel2), .Y(exu_n18082));
INVX1 exu_U28453(.A(exu_n18082), .Y(exu_n9755));
AND2X1 exu_U28454(.A(exu_tlu_ccr2_w[1]), .B(ecl_ccr_mux_ccrin2_sel2), .Y(exu_n18086));
INVX1 exu_U28455(.A(exu_n18086), .Y(exu_n9756));
AND2X1 exu_U28456(.A(exu_tlu_ccr2_w[0]), .B(ecl_ccr_mux_ccrin2_sel2), .Y(exu_n18090));
INVX1 exu_U28457(.A(exu_n18090), .Y(exu_n9757));
AND2X1 exu_U28458(.A(ecl_ccr_mux_ccrin3_sel2), .B(exu_tlu_ccr3_w[7]), .Y(exu_n18094));
INVX1 exu_U28459(.A(exu_n18094), .Y(exu_n9758));
AND2X1 exu_U28460(.A(exu_tlu_ccr3_w[6]), .B(ecl_ccr_mux_ccrin3_sel2), .Y(exu_n18098));
INVX1 exu_U28461(.A(exu_n18098), .Y(exu_n9759));
AND2X1 exu_U28462(.A(exu_tlu_ccr3_w[5]), .B(ecl_ccr_mux_ccrin3_sel2), .Y(exu_n18101));
INVX1 exu_U28463(.A(exu_n18101), .Y(exu_n9760));
AND2X1 exu_U28464(.A(exu_tlu_ccr3_w[4]), .B(ecl_ccr_mux_ccrin3_sel2), .Y(exu_n18103));
INVX1 exu_U28465(.A(exu_n18103), .Y(exu_n9761));
AND2X1 exu_U28466(.A(exu_tlu_ccr3_w[3]), .B(ecl_ccr_mux_ccrin3_sel2), .Y(exu_n18106));
INVX1 exu_U28467(.A(exu_n18106), .Y(exu_n9762));
AND2X1 exu_U28468(.A(exu_tlu_ccr3_w[2]), .B(ecl_ccr_mux_ccrin3_sel2), .Y(exu_n18110));
INVX1 exu_U28469(.A(exu_n18110), .Y(exu_n9763));
AND2X1 exu_U28470(.A(exu_tlu_ccr3_w[1]), .B(ecl_ccr_mux_ccrin3_sel2), .Y(exu_n18114));
INVX1 exu_U28471(.A(exu_n18114), .Y(exu_n9764));
AND2X1 exu_U28472(.A(exu_tlu_ccr3_w[0]), .B(ecl_ccr_mux_ccrin3_sel2), .Y(exu_n18118));
INVX1 exu_U28473(.A(exu_n18118), .Y(exu_n9765));
AND2X1 exu_U28474(.A(rml_agp_thr1[0]), .B(rml_agp_wen_thr1_w), .Y(exu_n18170));
INVX1 exu_U28475(.A(exu_n18170), .Y(exu_n9766));
AND2X1 exu_U28476(.A(rml_agp_thr1[1]), .B(rml_agp_wen_thr1_w), .Y(exu_n18172));
INVX1 exu_U28477(.A(exu_n18172), .Y(exu_n9767));
AND2X1 exu_U28478(.A(rml_agp_thr2[0]), .B(rml_agp_wen_thr2_w), .Y(exu_n18174));
INVX1 exu_U28479(.A(exu_n18174), .Y(exu_n9768));
AND2X1 exu_U28480(.A(rml_agp_thr2[1]), .B(rml_agp_wen_thr2_w), .Y(exu_n18176));
INVX1 exu_U28481(.A(exu_n18176), .Y(exu_n9769));
AND2X1 exu_U28482(.A(rml_agp_thr3[0]), .B(rml_agp_wen_thr3_w), .Y(exu_n18178));
INVX1 exu_U28483(.A(exu_n18178), .Y(exu_n9770));
AND2X1 exu_U28484(.A(rml_agp_thr3[1]), .B(rml_agp_wen_thr3_w), .Y(exu_n18180));
INVX1 exu_U28485(.A(exu_n18180), .Y(exu_n9771));
AND2X1 exu_U28486(.A(ecl_divcntl_subnext_mux_in1[0]), .B(exu_n16215), .Y(exu_n18181));
INVX1 exu_U28487(.A(exu_n18181), .Y(exu_n9772));
AND2X1 exu_U28488(.A(exu_n15334), .B(exu_n15979), .Y(exu_n18185));
INVX1 exu_U28489(.A(exu_n18185), .Y(exu_n9773));
AND2X1 exu_U28490(.A(rml_tid_e[0]), .B(exu_n15027), .Y(exu_n18188));
INVX1 exu_U28491(.A(exu_n18188), .Y(exu_n9774));
AND2X1 exu_U28492(.A(rml_tid_e[1]), .B(exu_n15027), .Y(exu_n18190));
INVX1 exu_U28493(.A(exu_n18190), .Y(exu_n9775));
AND2X1 exu_U28494(.A(rml_canrestore_reg_data_thr3[2]), .B(exu_n15745), .Y(exu_n18211));
INVX1 exu_U28495(.A(exu_n18211), .Y(exu_n9776));
AND2X1 exu_U28496(.A(rml_canrestore_reg_data_thr3[1]), .B(exu_n15745), .Y(exu_n18213));
INVX1 exu_U28497(.A(exu_n18213), .Y(exu_n9777));
AND2X1 exu_U28498(.A(rml_canrestore_reg_data_thr3[0]), .B(exu_n15745), .Y(exu_n18215));
INVX1 exu_U28499(.A(exu_n18215), .Y(exu_n9778));
AND2X1 exu_U28500(.A(rml_canrestore_reg_data_thr2[2]), .B(exu_n15746), .Y(exu_n18217));
INVX1 exu_U28501(.A(exu_n18217), .Y(exu_n9779));
AND2X1 exu_U28502(.A(rml_canrestore_reg_data_thr2[1]), .B(exu_n15746), .Y(exu_n18219));
INVX1 exu_U28503(.A(exu_n18219), .Y(exu_n9780));
AND2X1 exu_U28504(.A(rml_canrestore_reg_data_thr2[0]), .B(exu_n15746), .Y(exu_n18221));
INVX1 exu_U28505(.A(exu_n18221), .Y(exu_n9781));
AND2X1 exu_U28506(.A(rml_canrestore_reg_data_thr1[2]), .B(exu_n15747), .Y(exu_n18223));
INVX1 exu_U28507(.A(exu_n18223), .Y(exu_n9782));
AND2X1 exu_U28508(.A(rml_canrestore_reg_data_thr1[1]), .B(exu_n15747), .Y(exu_n18225));
INVX1 exu_U28509(.A(exu_n18225), .Y(exu_n9783));
AND2X1 exu_U28510(.A(rml_canrestore_reg_data_thr1[0]), .B(exu_n15747), .Y(exu_n18227));
INVX1 exu_U28511(.A(exu_n18227), .Y(exu_n9784));
AND2X1 exu_U28512(.A(rml_canrestore_reg_data_thr0[2]), .B(exu_n15748), .Y(exu_n18229));
INVX1 exu_U28513(.A(exu_n18229), .Y(exu_n9785));
AND2X1 exu_U28514(.A(rml_canrestore_reg_data_thr0[1]), .B(exu_n15748), .Y(exu_n18231));
INVX1 exu_U28515(.A(exu_n18231), .Y(exu_n9786));
AND2X1 exu_U28516(.A(rml_canrestore_reg_data_thr0[0]), .B(exu_n15748), .Y(exu_n18233));
INVX1 exu_U28517(.A(exu_n18233), .Y(exu_n9787));
AND2X1 exu_U28518(.A(rml_otherwin_reg_data_thr3[2]), .B(exu_n15749), .Y(exu_n18255));
INVX1 exu_U28519(.A(exu_n18255), .Y(exu_n9788));
AND2X1 exu_U28520(.A(rml_otherwin_reg_data_thr3[1]), .B(exu_n15749), .Y(exu_n18257));
INVX1 exu_U28521(.A(exu_n18257), .Y(exu_n9789));
AND2X1 exu_U28522(.A(rml_otherwin_reg_data_thr3[0]), .B(exu_n15749), .Y(exu_n18259));
INVX1 exu_U28523(.A(exu_n18259), .Y(exu_n9790));
AND2X1 exu_U28524(.A(rml_otherwin_reg_data_thr2[2]), .B(exu_n15750), .Y(exu_n18261));
INVX1 exu_U28525(.A(exu_n18261), .Y(exu_n9791));
AND2X1 exu_U28526(.A(rml_otherwin_reg_data_thr2[1]), .B(exu_n15750), .Y(exu_n18263));
INVX1 exu_U28527(.A(exu_n18263), .Y(exu_n9792));
AND2X1 exu_U28528(.A(rml_otherwin_reg_data_thr2[0]), .B(exu_n15750), .Y(exu_n18265));
INVX1 exu_U28529(.A(exu_n18265), .Y(exu_n9793));
AND2X1 exu_U28530(.A(rml_otherwin_reg_data_thr1[2]), .B(exu_n15751), .Y(exu_n18267));
INVX1 exu_U28531(.A(exu_n18267), .Y(exu_n9794));
AND2X1 exu_U28532(.A(rml_otherwin_reg_data_thr1[1]), .B(exu_n15751), .Y(exu_n18269));
INVX1 exu_U28533(.A(exu_n18269), .Y(exu_n9795));
AND2X1 exu_U28534(.A(rml_otherwin_reg_data_thr1[0]), .B(exu_n15751), .Y(exu_n18271));
INVX1 exu_U28535(.A(exu_n18271), .Y(exu_n9796));
AND2X1 exu_U28536(.A(rml_otherwin_reg_data_thr0[2]), .B(exu_n15752), .Y(exu_n18273));
INVX1 exu_U28537(.A(exu_n18273), .Y(exu_n9797));
AND2X1 exu_U28538(.A(rml_otherwin_reg_data_thr0[1]), .B(exu_n15752), .Y(exu_n18275));
INVX1 exu_U28539(.A(exu_n18275), .Y(exu_n9798));
AND2X1 exu_U28540(.A(rml_otherwin_reg_data_thr0[0]), .B(exu_n15752), .Y(exu_n18277));
INVX1 exu_U28541(.A(exu_n18277), .Y(exu_n9799));
AND2X1 exu_U28542(.A(rml_cleanwin_reg_data_thr3[2]), .B(exu_n15753), .Y(exu_n18299));
INVX1 exu_U28543(.A(exu_n18299), .Y(exu_n9800));
AND2X1 exu_U28544(.A(rml_cleanwin_reg_data_thr3[1]), .B(exu_n15753), .Y(exu_n18301));
INVX1 exu_U28545(.A(exu_n18301), .Y(exu_n9801));
AND2X1 exu_U28546(.A(rml_cleanwin_reg_data_thr3[0]), .B(exu_n15753), .Y(exu_n18303));
INVX1 exu_U28547(.A(exu_n18303), .Y(exu_n9802));
AND2X1 exu_U28548(.A(rml_cleanwin_reg_data_thr2[2]), .B(exu_n15754), .Y(exu_n18305));
INVX1 exu_U28549(.A(exu_n18305), .Y(exu_n9803));
AND2X1 exu_U28550(.A(rml_cleanwin_reg_data_thr2[1]), .B(exu_n15754), .Y(exu_n18307));
INVX1 exu_U28551(.A(exu_n18307), .Y(exu_n9804));
AND2X1 exu_U28552(.A(rml_cleanwin_reg_data_thr2[0]), .B(exu_n15754), .Y(exu_n18309));
INVX1 exu_U28553(.A(exu_n18309), .Y(exu_n9805));
AND2X1 exu_U28554(.A(rml_cleanwin_reg_data_thr1[2]), .B(exu_n15755), .Y(exu_n18311));
INVX1 exu_U28555(.A(exu_n18311), .Y(exu_n9806));
AND2X1 exu_U28556(.A(rml_cleanwin_reg_data_thr1[1]), .B(exu_n15755), .Y(exu_n18313));
INVX1 exu_U28557(.A(exu_n18313), .Y(exu_n9807));
AND2X1 exu_U28558(.A(rml_cleanwin_reg_data_thr1[0]), .B(exu_n15755), .Y(exu_n18315));
INVX1 exu_U28559(.A(exu_n18315), .Y(exu_n9808));
AND2X1 exu_U28560(.A(rml_cleanwin_reg_data_thr0[2]), .B(exu_n15756), .Y(exu_n18317));
INVX1 exu_U28561(.A(exu_n18317), .Y(exu_n9809));
AND2X1 exu_U28562(.A(rml_cleanwin_reg_data_thr0[1]), .B(exu_n15756), .Y(exu_n18319));
INVX1 exu_U28563(.A(exu_n18319), .Y(exu_n9810));
AND2X1 exu_U28564(.A(rml_cleanwin_reg_data_thr0[0]), .B(exu_n15756), .Y(exu_n18321));
INVX1 exu_U28565(.A(exu_n18321), .Y(exu_n9811));
INVX1 exu_U28566(.A(exu_n18343), .Y(exu_n9812));
INVX1 exu_U28567(.A(exu_n18345), .Y(exu_n9813));
AND2X1 exu_U28568(.A(rml_hi_wstate_reg_data_thr3[0]), .B(exu_n15194), .Y(exu_n18347));
INVX1 exu_U28569(.A(exu_n18347), .Y(exu_n9814));
INVX1 exu_U28570(.A(exu_n18349), .Y(exu_n9815));
INVX1 exu_U28571(.A(exu_n18351), .Y(exu_n9816));
AND2X1 exu_U28572(.A(rml_hi_wstate_reg_data_thr2[0]), .B(exu_n15195), .Y(exu_n18353));
INVX1 exu_U28573(.A(exu_n18353), .Y(exu_n9817));
INVX1 exu_U28574(.A(exu_n18355), .Y(exu_n9818));
INVX1 exu_U28575(.A(exu_n18357), .Y(exu_n9819));
AND2X1 exu_U28576(.A(rml_hi_wstate_reg_data_thr1[0]), .B(exu_n15196), .Y(exu_n18359));
INVX1 exu_U28577(.A(exu_n18359), .Y(exu_n9820));
INVX1 exu_U28578(.A(exu_n18361), .Y(exu_n9821));
INVX1 exu_U28579(.A(exu_n18363), .Y(exu_n9822));
AND2X1 exu_U28580(.A(rml_hi_wstate_reg_data_thr0[0]), .B(exu_n15197), .Y(exu_n18365));
INVX1 exu_U28581(.A(exu_n18365), .Y(exu_n9823));
AND2X1 exu_U28582(.A(rml_lo_wstate_reg_data_thr3[2]), .B(exu_n15194), .Y(exu_n18383));
INVX1 exu_U28583(.A(exu_n18383), .Y(exu_n9824));
AND2X1 exu_U28584(.A(rml_lo_wstate_reg_data_thr3[1]), .B(exu_n15194), .Y(exu_n18385));
INVX1 exu_U28585(.A(exu_n18385), .Y(exu_n9825));
AND2X1 exu_U28586(.A(rml_lo_wstate_reg_data_thr3[0]), .B(exu_n15194), .Y(exu_n18387));
INVX1 exu_U28587(.A(exu_n18387), .Y(exu_n9826));
AND2X1 exu_U28588(.A(rml_lo_wstate_reg_data_thr2[2]), .B(exu_n15195), .Y(exu_n18389));
INVX1 exu_U28589(.A(exu_n18389), .Y(exu_n9827));
AND2X1 exu_U28590(.A(rml_lo_wstate_reg_data_thr2[1]), .B(exu_n15195), .Y(exu_n18391));
INVX1 exu_U28591(.A(exu_n18391), .Y(exu_n9828));
AND2X1 exu_U28592(.A(rml_lo_wstate_reg_data_thr2[0]), .B(exu_n15195), .Y(exu_n18393));
INVX1 exu_U28593(.A(exu_n18393), .Y(exu_n9829));
AND2X1 exu_U28594(.A(rml_lo_wstate_reg_data_thr1[2]), .B(exu_n15196), .Y(exu_n18395));
INVX1 exu_U28595(.A(exu_n18395), .Y(exu_n9830));
AND2X1 exu_U28596(.A(rml_lo_wstate_reg_data_thr1[1]), .B(exu_n15196), .Y(exu_n18397));
INVX1 exu_U28597(.A(exu_n18397), .Y(exu_n9831));
AND2X1 exu_U28598(.A(rml_lo_wstate_reg_data_thr1[0]), .B(exu_n15196), .Y(exu_n18399));
INVX1 exu_U28599(.A(exu_n18399), .Y(exu_n9832));
AND2X1 exu_U28600(.A(rml_lo_wstate_reg_data_thr0[2]), .B(exu_n15197), .Y(exu_n18401));
INVX1 exu_U28601(.A(exu_n18401), .Y(exu_n9833));
AND2X1 exu_U28602(.A(rml_lo_wstate_reg_data_thr0[1]), .B(exu_n15197), .Y(exu_n18403));
INVX1 exu_U28603(.A(exu_n18403), .Y(exu_n9834));
AND2X1 exu_U28604(.A(rml_lo_wstate_reg_data_thr0[0]), .B(exu_n15197), .Y(exu_n18405));
INVX1 exu_U28605(.A(exu_n18405), .Y(exu_n9835));
AND2X1 exu_U28606(.A(ecl_rml_xor_data_e[0]), .B(exu_n16384), .Y(exu_n18433));
INVX1 exu_U28607(.A(exu_n18433), .Y(exu_n9836));
AND2X1 exu_U28608(.A(ecl_rml_xor_data_e[1]), .B(exu_n16384), .Y(exu_n18435));
INVX1 exu_U28609(.A(exu_n18435), .Y(exu_n9837));
AND2X1 exu_U28610(.A(ecl_rml_xor_data_e[2]), .B(exu_n16384), .Y(exu_n18437));
INVX1 exu_U28611(.A(exu_n18437), .Y(exu_n9838));
AND2X1 exu_U28612(.A(ecl_rml_xor_data_e[0]), .B(exu_n15762), .Y(exu_n18439));
INVX1 exu_U28613(.A(exu_n18439), .Y(exu_n9839));
AND2X1 exu_U28614(.A(ecl_rml_xor_data_e[1]), .B(exu_n15762), .Y(exu_n18441));
INVX1 exu_U28615(.A(exu_n18441), .Y(exu_n9840));
AND2X1 exu_U28616(.A(ecl_rml_xor_data_e[2]), .B(exu_n15762), .Y(exu_n18443));
INVX1 exu_U28617(.A(exu_n18443), .Y(exu_n9841));
AND2X1 exu_U28618(.A(ecl_rml_xor_data_e[0]), .B(exu_n15763), .Y(exu_n18445));
INVX1 exu_U28619(.A(exu_n18445), .Y(exu_n9842));
AND2X1 exu_U28620(.A(ecl_rml_xor_data_e[1]), .B(exu_n15763), .Y(exu_n18447));
INVX1 exu_U28621(.A(exu_n18447), .Y(exu_n9843));
AND2X1 exu_U28622(.A(ecl_rml_xor_data_e[2]), .B(exu_n15763), .Y(exu_n18449));
INVX1 exu_U28623(.A(exu_n18449), .Y(exu_n9844));
AND2X1 exu_U28624(.A(rml_cansave_reg_data_thr0[0]), .B(exu_n15760), .Y(exu_n18451));
INVX1 exu_U28625(.A(exu_n18451), .Y(exu_n9845));
AND2X1 exu_U28626(.A(rml_cansave_reg_data_thr0[1]), .B(exu_n15760), .Y(exu_n18453));
INVX1 exu_U28627(.A(exu_n18453), .Y(exu_n9846));
AND2X1 exu_U28628(.A(rml_cansave_reg_data_thr0[2]), .B(exu_n15760), .Y(exu_n18455));
INVX1 exu_U28629(.A(exu_n18455), .Y(exu_n9847));
AND2X1 exu_U28630(.A(rml_cansave_reg_data_thr1[0]), .B(exu_n15759), .Y(exu_n18457));
INVX1 exu_U28631(.A(exu_n18457), .Y(exu_n9848));
AND2X1 exu_U28632(.A(rml_cansave_reg_data_thr1[1]), .B(exu_n15759), .Y(exu_n18459));
INVX1 exu_U28633(.A(exu_n18459), .Y(exu_n9849));
AND2X1 exu_U28634(.A(rml_cansave_reg_data_thr1[2]), .B(exu_n15759), .Y(exu_n18461));
INVX1 exu_U28635(.A(exu_n18461), .Y(exu_n9850));
AND2X1 exu_U28636(.A(rml_cansave_reg_data_thr2[0]), .B(exu_n15758), .Y(exu_n18463));
INVX1 exu_U28637(.A(exu_n18463), .Y(exu_n9851));
AND2X1 exu_U28638(.A(rml_cansave_reg_data_thr2[1]), .B(exu_n15758), .Y(exu_n18465));
INVX1 exu_U28639(.A(exu_n18465), .Y(exu_n9852));
AND2X1 exu_U28640(.A(rml_cansave_reg_data_thr2[2]), .B(exu_n15758), .Y(exu_n18467));
INVX1 exu_U28641(.A(exu_n18467), .Y(exu_n9853));
AND2X1 exu_U28642(.A(rml_cansave_reg_data_thr3[0]), .B(exu_n15757), .Y(exu_n18469));
INVX1 exu_U28643(.A(exu_n18469), .Y(exu_n9854));
AND2X1 exu_U28644(.A(rml_cansave_reg_data_thr3[1]), .B(exu_n15757), .Y(exu_n18471));
INVX1 exu_U28645(.A(exu_n18471), .Y(exu_n9855));
AND2X1 exu_U28646(.A(rml_cansave_reg_data_thr3[2]), .B(exu_n15757), .Y(exu_n18473));
INVX1 exu_U28647(.A(exu_n18473), .Y(exu_n9856));
AND2X1 exu_U28648(.A(exu_n15986), .B(exu_mul_rs1_data[9]), .Y(exu_n18604));
INVX1 exu_U28649(.A(exu_n18604), .Y(exu_n9857));
AND2X1 exu_U28650(.A(exu_mul_rs2_data[35]), .B(exu_n15986), .Y(exu_n18608));
INVX1 exu_U28651(.A(exu_n18608), .Y(exu_n9858));
AND2X1 exu_U28652(.A(exu_mul_rs2_data[34]), .B(exu_n15986), .Y(exu_n18611));
INVX1 exu_U28653(.A(exu_n18611), .Y(exu_n9859));
AND2X1 exu_U28654(.A(exu_mul_rs2_data[33]), .B(exu_n15986), .Y(exu_n18614));
INVX1 exu_U28655(.A(exu_n18614), .Y(exu_n9860));
AND2X1 exu_U28656(.A(exu_mul_rs2_data[32]), .B(exu_n15985), .Y(exu_n18617));
INVX1 exu_U28657(.A(exu_n18617), .Y(exu_n9861));
AND2X1 exu_U28658(.A(exu_mul_rs2_data[31]), .B(exu_n15986), .Y(exu_n18620));
INVX1 exu_U28659(.A(exu_n18620), .Y(exu_n9862));
AND2X1 exu_U28660(.A(exu_mul_rs2_data[30]), .B(exu_n15986), .Y(exu_n18624));
INVX1 exu_U28661(.A(exu_n18624), .Y(exu_n9863));
AND2X1 exu_U28662(.A(exu_mul_rs2_data[29]), .B(exu_n15986), .Y(exu_n18628));
INVX1 exu_U28663(.A(exu_n18628), .Y(exu_n9864));
AND2X1 exu_U28664(.A(exu_mul_rs2_data[28]), .B(exu_n15985), .Y(exu_n18632));
INVX1 exu_U28665(.A(exu_n18632), .Y(exu_n9865));
AND2X1 exu_U28666(.A(exu_mul_rs2_data[27]), .B(exu_n15985), .Y(exu_n18636));
INVX1 exu_U28667(.A(exu_n18636), .Y(exu_n9866));
AND2X1 exu_U28668(.A(exu_mul_rs2_data[26]), .B(exu_n15986), .Y(exu_n18640));
INVX1 exu_U28669(.A(exu_n18640), .Y(exu_n9867));
AND2X1 exu_U28670(.A(exu_mul_rs1_data[8]), .B(exu_n15985), .Y(exu_n18644));
INVX1 exu_U28671(.A(exu_n18644), .Y(exu_n9868));
AND2X1 exu_U28672(.A(exu_mul_rs2_data[25]), .B(exu_n15986), .Y(exu_n18648));
INVX1 exu_U28673(.A(exu_n18648), .Y(exu_n9869));
AND2X1 exu_U28674(.A(exu_mul_rs2_data[24]), .B(exu_n15985), .Y(exu_n18652));
INVX1 exu_U28675(.A(exu_n18652), .Y(exu_n9870));
AND2X1 exu_U28676(.A(exu_mul_rs2_data[23]), .B(exu_n15986), .Y(exu_n18656));
INVX1 exu_U28677(.A(exu_n18656), .Y(exu_n9871));
AND2X1 exu_U28678(.A(exu_mul_rs2_data[22]), .B(exu_n15985), .Y(exu_n18660));
INVX1 exu_U28679(.A(exu_n18660), .Y(exu_n9872));
AND2X1 exu_U28680(.A(exu_mul_rs2_data[21]), .B(exu_n15985), .Y(exu_n18664));
INVX1 exu_U28681(.A(exu_n18664), .Y(exu_n9873));
AND2X1 exu_U28682(.A(exu_mul_rs2_data[20]), .B(exu_n15985), .Y(exu_n18668));
INVX1 exu_U28683(.A(exu_n18668), .Y(exu_n9874));
AND2X1 exu_U28684(.A(exu_mul_rs2_data[19]), .B(exu_n15985), .Y(exu_n18672));
INVX1 exu_U28685(.A(exu_n18672), .Y(exu_n9875));
AND2X1 exu_U28686(.A(exu_mul_rs2_data[18]), .B(exu_n15986), .Y(exu_n18676));
INVX1 exu_U28687(.A(exu_n18676), .Y(exu_n9876));
AND2X1 exu_U28688(.A(exu_mul_rs2_data[17]), .B(exu_n15985), .Y(exu_n18680));
INVX1 exu_U28689(.A(exu_n18680), .Y(exu_n9877));
AND2X1 exu_U28690(.A(exu_mul_rs2_data[16]), .B(exu_n15986), .Y(exu_n18684));
INVX1 exu_U28691(.A(exu_n18684), .Y(exu_n9878));
AND2X1 exu_U28692(.A(exu_mul_rs1_data[7]), .B(exu_n15985), .Y(exu_n18688));
INVX1 exu_U28693(.A(exu_n18688), .Y(exu_n9879));
AND2X1 exu_U28694(.A(exu_mul_rs2_data[15]), .B(exu_n15986), .Y(exu_n18692));
INVX1 exu_U28695(.A(exu_n18692), .Y(exu_n9880));
AND2X1 exu_U28696(.A(exu_mul_rs2_data[14]), .B(exu_n15985), .Y(exu_n18696));
INVX1 exu_U28697(.A(exu_n18696), .Y(exu_n9881));
AND2X1 exu_U28698(.A(exu_mul_rs2_data[13]), .B(exu_n15986), .Y(exu_n18700));
INVX1 exu_U28699(.A(exu_n18700), .Y(exu_n9882));
AND2X1 exu_U28700(.A(exu_mul_rs2_data[12]), .B(exu_n15985), .Y(exu_n18704));
INVX1 exu_U28701(.A(exu_n18704), .Y(exu_n9883));
AND2X1 exu_U28702(.A(exu_mul_rs2_data[11]), .B(exu_n15986), .Y(exu_n18708));
INVX1 exu_U28703(.A(exu_n18708), .Y(exu_n9884));
AND2X1 exu_U28704(.A(exu_mul_rs2_data[10]), .B(exu_n15985), .Y(exu_n18712));
INVX1 exu_U28705(.A(exu_n18712), .Y(exu_n9885));
AND2X1 exu_U28706(.A(exu_mul_rs2_data[9]), .B(exu_n15986), .Y(exu_n18716));
INVX1 exu_U28707(.A(exu_n18716), .Y(exu_n9886));
AND2X1 exu_U28708(.A(exu_mul_rs2_data[8]), .B(exu_n15985), .Y(exu_n18720));
INVX1 exu_U28709(.A(exu_n18720), .Y(exu_n9887));
AND2X1 exu_U28710(.A(exu_mul_rs2_data[7]), .B(exu_n15986), .Y(exu_n18724));
INVX1 exu_U28711(.A(exu_n18724), .Y(exu_n9888));
AND2X1 exu_U28712(.A(exu_mul_rs2_data[6]), .B(exu_n15985), .Y(exu_n18728));
INVX1 exu_U28713(.A(exu_n18728), .Y(exu_n9889));
AND2X1 exu_U28714(.A(exu_mul_rs1_data[6]), .B(exu_n15985), .Y(exu_n18732));
INVX1 exu_U28715(.A(exu_n18732), .Y(exu_n9890));
AND2X1 exu_U28716(.A(exu_mul_rs2_data[5]), .B(exu_n15986), .Y(exu_n18736));
INVX1 exu_U28717(.A(exu_n18736), .Y(exu_n9891));
AND2X1 exu_U28718(.A(exu_mul_rs2_data[4]), .B(exu_n15986), .Y(exu_n18740));
INVX1 exu_U28719(.A(exu_n18740), .Y(exu_n9892));
AND2X1 exu_U28720(.A(exu_mul_rs2_data[3]), .B(exu_n15985), .Y(exu_n18744));
INVX1 exu_U28721(.A(exu_n18744), .Y(exu_n9893));
AND2X1 exu_U28722(.A(exu_mul_rs2_data[2]), .B(exu_n15986), .Y(exu_n18748));
INVX1 exu_U28723(.A(exu_n18748), .Y(exu_n9894));
AND2X1 exu_U28724(.A(exu_mul_rs2_data[1]), .B(exu_n15986), .Y(exu_n18752));
INVX1 exu_U28725(.A(exu_n18752), .Y(exu_n9895));
AND2X1 exu_U28726(.A(exu_mul_rs2_data[0]), .B(exu_n15986), .Y(exu_n18756));
INVX1 exu_U28727(.A(exu_n18756), .Y(exu_n9896));
AND2X1 exu_U28728(.A(exu_mul_rs1_data[63]), .B(exu_n15986), .Y(exu_n18760));
INVX1 exu_U28729(.A(exu_n18760), .Y(exu_n9897));
AND2X1 exu_U28730(.A(exu_mul_rs1_data[62]), .B(exu_n15985), .Y(exu_n18763));
INVX1 exu_U28731(.A(exu_n18763), .Y(exu_n9898));
AND2X1 exu_U28732(.A(exu_mul_rs1_data[61]), .B(exu_n15985), .Y(exu_n18766));
INVX1 exu_U28733(.A(exu_n18766), .Y(exu_n9899));
AND2X1 exu_U28734(.A(exu_mul_rs1_data[60]), .B(exu_n15986), .Y(exu_n18769));
INVX1 exu_U28735(.A(exu_n18769), .Y(exu_n9900));
AND2X1 exu_U28736(.A(exu_mul_rs1_data[5]), .B(exu_n15986), .Y(exu_n18772));
INVX1 exu_U28737(.A(exu_n18772), .Y(exu_n9901));
AND2X1 exu_U28738(.A(exu_mul_rs1_data[59]), .B(exu_n15986), .Y(exu_n18776));
INVX1 exu_U28739(.A(exu_n18776), .Y(exu_n9902));
AND2X1 exu_U28740(.A(exu_mul_rs1_data[58]), .B(exu_n15985), .Y(exu_n18779));
INVX1 exu_U28741(.A(exu_n18779), .Y(exu_n9903));
AND2X1 exu_U28742(.A(exu_mul_rs1_data[57]), .B(exu_n15986), .Y(exu_n18782));
INVX1 exu_U28743(.A(exu_n18782), .Y(exu_n9904));
AND2X1 exu_U28744(.A(exu_mul_rs1_data[56]), .B(exu_n15985), .Y(exu_n18785));
INVX1 exu_U28745(.A(exu_n18785), .Y(exu_n9905));
AND2X1 exu_U28746(.A(exu_mul_rs1_data[55]), .B(exu_n15986), .Y(exu_n18788));
INVX1 exu_U28747(.A(exu_n18788), .Y(exu_n9906));
AND2X1 exu_U28748(.A(exu_mul_rs1_data[54]), .B(exu_n15986), .Y(exu_n18791));
INVX1 exu_U28749(.A(exu_n18791), .Y(exu_n9907));
AND2X1 exu_U28750(.A(exu_mul_rs1_data[53]), .B(exu_n15986), .Y(exu_n18794));
INVX1 exu_U28751(.A(exu_n18794), .Y(exu_n9908));
AND2X1 exu_U28752(.A(exu_mul_rs1_data[52]), .B(exu_n15985), .Y(exu_n18797));
INVX1 exu_U28753(.A(exu_n18797), .Y(exu_n9909));
AND2X1 exu_U28754(.A(exu_mul_rs1_data[51]), .B(exu_n15985), .Y(exu_n18800));
INVX1 exu_U28755(.A(exu_n18800), .Y(exu_n9910));
AND2X1 exu_U28756(.A(exu_mul_rs1_data[50]), .B(exu_n15986), .Y(exu_n18803));
INVX1 exu_U28757(.A(exu_n18803), .Y(exu_n9911));
AND2X1 exu_U28758(.A(exu_mul_rs1_data[4]), .B(exu_n15986), .Y(exu_n18806));
INVX1 exu_U28759(.A(exu_n18806), .Y(exu_n9912));
AND2X1 exu_U28760(.A(exu_mul_rs1_data[49]), .B(exu_n15986), .Y(exu_n18810));
INVX1 exu_U28761(.A(exu_n18810), .Y(exu_n9913));
AND2X1 exu_U28762(.A(exu_mul_rs1_data[48]), .B(exu_n15986), .Y(exu_n18813));
INVX1 exu_U28763(.A(exu_n18813), .Y(exu_n9914));
AND2X1 exu_U28764(.A(exu_mul_rs1_data[47]), .B(exu_n15985), .Y(exu_n18816));
INVX1 exu_U28765(.A(exu_n18816), .Y(exu_n9915));
AND2X1 exu_U28766(.A(exu_mul_rs1_data[46]), .B(exu_n15985), .Y(exu_n18819));
INVX1 exu_U28767(.A(exu_n18819), .Y(exu_n9916));
AND2X1 exu_U28768(.A(exu_mul_rs1_data[45]), .B(exu_n15985), .Y(exu_n18822));
INVX1 exu_U28769(.A(exu_n18822), .Y(exu_n9917));
AND2X1 exu_U28770(.A(exu_mul_rs1_data[44]), .B(exu_n15985), .Y(exu_n18825));
INVX1 exu_U28771(.A(exu_n18825), .Y(exu_n9918));
AND2X1 exu_U28772(.A(exu_mul_rs1_data[43]), .B(exu_n15986), .Y(exu_n18828));
INVX1 exu_U28773(.A(exu_n18828), .Y(exu_n9919));
AND2X1 exu_U28774(.A(exu_mul_rs1_data[42]), .B(exu_n15985), .Y(exu_n18831));
INVX1 exu_U28775(.A(exu_n18831), .Y(exu_n9920));
AND2X1 exu_U28776(.A(exu_mul_rs1_data[41]), .B(exu_n15986), .Y(exu_n18834));
INVX1 exu_U28777(.A(exu_n18834), .Y(exu_n9921));
AND2X1 exu_U28778(.A(exu_mul_rs1_data[40]), .B(exu_n15986), .Y(exu_n18837));
INVX1 exu_U28779(.A(exu_n18837), .Y(exu_n9922));
AND2X1 exu_U28780(.A(exu_mul_rs1_data[3]), .B(exu_n15986), .Y(exu_n18840));
INVX1 exu_U28781(.A(exu_n18840), .Y(exu_n9923));
AND2X1 exu_U28782(.A(exu_mul_rs1_data[39]), .B(exu_n15986), .Y(exu_n18844));
INVX1 exu_U28783(.A(exu_n18844), .Y(exu_n9924));
AND2X1 exu_U28784(.A(exu_mul_rs1_data[38]), .B(exu_n15986), .Y(exu_n18847));
INVX1 exu_U28785(.A(exu_n18847), .Y(exu_n9925));
AND2X1 exu_U28786(.A(exu_mul_rs1_data[37]), .B(exu_n15986), .Y(exu_n18850));
INVX1 exu_U28787(.A(exu_n18850), .Y(exu_n9926));
AND2X1 exu_U28788(.A(exu_mul_rs1_data[36]), .B(exu_n15986), .Y(exu_n18853));
INVX1 exu_U28789(.A(exu_n18853), .Y(exu_n9927));
AND2X1 exu_U28790(.A(exu_mul_rs1_data[35]), .B(exu_n15985), .Y(exu_n18856));
INVX1 exu_U28791(.A(exu_n18856), .Y(exu_n9928));
AND2X1 exu_U28792(.A(exu_mul_rs1_data[34]), .B(exu_n15985), .Y(exu_n18859));
INVX1 exu_U28793(.A(exu_n18859), .Y(exu_n9929));
AND2X1 exu_U28794(.A(exu_mul_rs1_data[33]), .B(exu_n15985), .Y(exu_n18862));
INVX1 exu_U28795(.A(exu_n18862), .Y(exu_n9930));
AND2X1 exu_U28796(.A(exu_mul_rs1_data[32]), .B(exu_n15985), .Y(exu_n18865));
INVX1 exu_U28797(.A(exu_n18865), .Y(exu_n9931));
AND2X1 exu_U28798(.A(exu_mul_rs1_data[31]), .B(exu_n15986), .Y(exu_n18869));
INVX1 exu_U28799(.A(exu_n18869), .Y(exu_n9932));
AND2X1 exu_U28800(.A(exu_mul_rs1_data[30]), .B(exu_n15986), .Y(exu_n18873));
INVX1 exu_U28801(.A(exu_n18873), .Y(exu_n9933));
AND2X1 exu_U28802(.A(exu_mul_rs1_data[2]), .B(exu_n15986), .Y(exu_n18877));
INVX1 exu_U28803(.A(exu_n18877), .Y(exu_n9934));
AND2X1 exu_U28804(.A(exu_mul_rs1_data[29]), .B(exu_n15986), .Y(exu_n18881));
INVX1 exu_U28805(.A(exu_n18881), .Y(exu_n9935));
AND2X1 exu_U28806(.A(exu_mul_rs1_data[28]), .B(exu_n15985), .Y(exu_n18885));
INVX1 exu_U28807(.A(exu_n18885), .Y(exu_n9936));
AND2X1 exu_U28808(.A(exu_mul_rs1_data[27]), .B(exu_n15985), .Y(exu_n18889));
INVX1 exu_U28809(.A(exu_n18889), .Y(exu_n9937));
AND2X1 exu_U28810(.A(exu_mul_rs1_data[26]), .B(exu_n15985), .Y(exu_n18893));
INVX1 exu_U28811(.A(exu_n18893), .Y(exu_n9938));
AND2X1 exu_U28812(.A(exu_mul_rs1_data[25]), .B(exu_n15986), .Y(exu_n18897));
INVX1 exu_U28813(.A(exu_n18897), .Y(exu_n9939));
AND2X1 exu_U28814(.A(exu_mul_rs1_data[24]), .B(exu_n15986), .Y(exu_n18901));
INVX1 exu_U28815(.A(exu_n18901), .Y(exu_n9940));
AND2X1 exu_U28816(.A(exu_mul_rs1_data[23]), .B(exu_n15986), .Y(exu_n18905));
INVX1 exu_U28817(.A(exu_n18905), .Y(exu_n9941));
AND2X1 exu_U28818(.A(exu_mul_rs1_data[22]), .B(exu_n15985), .Y(exu_n18909));
INVX1 exu_U28819(.A(exu_n18909), .Y(exu_n9942));
AND2X1 exu_U28820(.A(exu_mul_rs1_data[21]), .B(exu_n15985), .Y(exu_n18913));
INVX1 exu_U28821(.A(exu_n18913), .Y(exu_n9943));
AND2X1 exu_U28822(.A(exu_mul_rs1_data[20]), .B(exu_n15985), .Y(exu_n18917));
INVX1 exu_U28823(.A(exu_n18917), .Y(exu_n9944));
AND2X1 exu_U28824(.A(exu_mul_rs1_data[1]), .B(exu_n15985), .Y(exu_n18921));
INVX1 exu_U28825(.A(exu_n18921), .Y(exu_n9945));
AND2X1 exu_U28826(.A(exu_mul_rs1_data[19]), .B(exu_n15985), .Y(exu_n18925));
INVX1 exu_U28827(.A(exu_n18925), .Y(exu_n9946));
AND2X1 exu_U28828(.A(exu_mul_rs1_data[18]), .B(exu_n15985), .Y(exu_n18929));
INVX1 exu_U28829(.A(exu_n18929), .Y(exu_n9947));
AND2X1 exu_U28830(.A(exu_mul_rs1_data[17]), .B(exu_n15985), .Y(exu_n18933));
INVX1 exu_U28831(.A(exu_n18933), .Y(exu_n9948));
AND2X1 exu_U28832(.A(exu_mul_rs1_data[16]), .B(exu_n15985), .Y(exu_n18937));
INVX1 exu_U28833(.A(exu_n18937), .Y(exu_n9949));
AND2X1 exu_U28834(.A(exu_mul_rs1_data[15]), .B(exu_n15985), .Y(exu_n18941));
INVX1 exu_U28835(.A(exu_n18941), .Y(exu_n9950));
AND2X1 exu_U28836(.A(exu_mul_rs1_data[14]), .B(exu_n15985), .Y(exu_n18945));
INVX1 exu_U28837(.A(exu_n18945), .Y(exu_n9951));
AND2X1 exu_U28838(.A(exu_mul_rs1_data[13]), .B(exu_n15985), .Y(exu_n18949));
INVX1 exu_U28839(.A(exu_n18949), .Y(exu_n9952));
AND2X1 exu_U28840(.A(exu_mul_rs1_data[12]), .B(exu_n15985), .Y(exu_n18953));
INVX1 exu_U28841(.A(exu_n18953), .Y(exu_n9953));
AND2X1 exu_U28842(.A(exu_mul_rs2_data[63]), .B(exu_n15985), .Y(exu_n18957));
INVX1 exu_U28843(.A(exu_n18957), .Y(exu_n9954));
AND2X1 exu_U28844(.A(exu_mul_rs2_data[62]), .B(exu_n15985), .Y(exu_n18960));
INVX1 exu_U28845(.A(exu_n18960), .Y(exu_n9955));
AND2X1 exu_U28846(.A(exu_mul_rs2_data[61]), .B(exu_n15985), .Y(exu_n18963));
INVX1 exu_U28847(.A(exu_n18963), .Y(exu_n9956));
AND2X1 exu_U28848(.A(exu_mul_rs2_data[60]), .B(exu_n15985), .Y(exu_n18966));
INVX1 exu_U28849(.A(exu_n18966), .Y(exu_n9957));
AND2X1 exu_U28850(.A(exu_mul_rs2_data[59]), .B(exu_n15985), .Y(exu_n18969));
INVX1 exu_U28851(.A(exu_n18969), .Y(exu_n9958));
AND2X1 exu_U28852(.A(exu_mul_rs2_data[58]), .B(exu_n15986), .Y(exu_n18972));
INVX1 exu_U28853(.A(exu_n18972), .Y(exu_n9959));
AND2X1 exu_U28854(.A(exu_mul_rs2_data[57]), .B(exu_n15986), .Y(exu_n18975));
INVX1 exu_U28855(.A(exu_n18975), .Y(exu_n9960));
AND2X1 exu_U28856(.A(exu_mul_rs2_data[56]), .B(exu_n15986), .Y(exu_n18978));
INVX1 exu_U28857(.A(exu_n18978), .Y(exu_n9961));
AND2X1 exu_U28858(.A(exu_mul_rs1_data[11]), .B(exu_n15985), .Y(exu_n18981));
INVX1 exu_U28859(.A(exu_n18981), .Y(exu_n9962));
AND2X1 exu_U28860(.A(exu_mul_rs2_data[55]), .B(exu_n15986), .Y(exu_n18985));
INVX1 exu_U28861(.A(exu_n18985), .Y(exu_n9963));
AND2X1 exu_U28862(.A(exu_mul_rs2_data[54]), .B(exu_n15985), .Y(exu_n18988));
INVX1 exu_U28863(.A(exu_n18988), .Y(exu_n9964));
AND2X1 exu_U28864(.A(exu_mul_rs2_data[53]), .B(exu_n15985), .Y(exu_n18991));
INVX1 exu_U28865(.A(exu_n18991), .Y(exu_n9965));
AND2X1 exu_U28866(.A(exu_mul_rs2_data[52]), .B(exu_n15986), .Y(exu_n18994));
INVX1 exu_U28867(.A(exu_n18994), .Y(exu_n9966));
AND2X1 exu_U28868(.A(exu_mul_rs2_data[51]), .B(exu_n15986), .Y(exu_n18997));
INVX1 exu_U28869(.A(exu_n18997), .Y(exu_n9967));
AND2X1 exu_U28870(.A(exu_mul_rs2_data[50]), .B(exu_n15985), .Y(exu_n19000));
INVX1 exu_U28871(.A(exu_n19000), .Y(exu_n9968));
AND2X1 exu_U28872(.A(exu_mul_rs2_data[49]), .B(exu_n15986), .Y(exu_n19003));
INVX1 exu_U28873(.A(exu_n19003), .Y(exu_n9969));
AND2X1 exu_U28874(.A(exu_mul_rs2_data[48]), .B(exu_n15985), .Y(exu_n19006));
INVX1 exu_U28875(.A(exu_n19006), .Y(exu_n9970));
AND2X1 exu_U28876(.A(exu_mul_rs2_data[47]), .B(exu_n15986), .Y(exu_n19009));
INVX1 exu_U28877(.A(exu_n19009), .Y(exu_n9971));
AND2X1 exu_U28878(.A(exu_mul_rs2_data[46]), .B(exu_n15986), .Y(exu_n19012));
INVX1 exu_U28879(.A(exu_n19012), .Y(exu_n9972));
AND2X1 exu_U28880(.A(exu_mul_rs1_data[10]), .B(exu_n15986), .Y(exu_n19015));
INVX1 exu_U28881(.A(exu_n19015), .Y(exu_n9973));
AND2X1 exu_U28882(.A(exu_mul_rs2_data[45]), .B(exu_n15986), .Y(exu_n19019));
INVX1 exu_U28883(.A(exu_n19019), .Y(exu_n9974));
AND2X1 exu_U28884(.A(exu_mul_rs2_data[44]), .B(exu_n15985), .Y(exu_n19022));
INVX1 exu_U28885(.A(exu_n19022), .Y(exu_n9975));
AND2X1 exu_U28886(.A(exu_mul_rs2_data[43]), .B(exu_n15986), .Y(exu_n19025));
INVX1 exu_U28887(.A(exu_n19025), .Y(exu_n9976));
AND2X1 exu_U28888(.A(exu_mul_rs2_data[42]), .B(exu_n15985), .Y(exu_n19028));
INVX1 exu_U28889(.A(exu_n19028), .Y(exu_n9977));
AND2X1 exu_U28890(.A(exu_mul_rs2_data[41]), .B(exu_n15986), .Y(exu_n19031));
INVX1 exu_U28891(.A(exu_n19031), .Y(exu_n9978));
AND2X1 exu_U28892(.A(exu_mul_rs2_data[40]), .B(exu_n15986), .Y(exu_n19034));
INVX1 exu_U28893(.A(exu_n19034), .Y(exu_n9979));
AND2X1 exu_U28894(.A(exu_mul_rs2_data[39]), .B(exu_n15985), .Y(exu_n19037));
INVX1 exu_U28895(.A(exu_n19037), .Y(exu_n9980));
AND2X1 exu_U28896(.A(exu_mul_rs2_data[38]), .B(exu_n15985), .Y(exu_n19040));
INVX1 exu_U28897(.A(exu_n19040), .Y(exu_n9981));
AND2X1 exu_U28898(.A(exu_mul_rs2_data[37]), .B(exu_n15985), .Y(exu_n19043));
INVX1 exu_U28899(.A(exu_n19043), .Y(exu_n9982));
AND2X1 exu_U28900(.A(exu_mul_rs2_data[36]), .B(exu_n15985), .Y(exu_n19046));
INVX1 exu_U28901(.A(exu_n19046), .Y(exu_n9983));
AND2X1 exu_U28902(.A(exu_mul_rs1_data[0]), .B(exu_n15986), .Y(exu_n19050));
INVX1 exu_U28903(.A(exu_n19050), .Y(exu_n9984));
AND2X1 exu_U28904(.A(exu_n19199), .B(exu_n9986), .Y(exu_n19205));
INVX1 exu_U28905(.A(exu_n19205), .Y(exu_n9985));
AND2X1 exu_U28906(.A(exu_n19202), .B(exu_n15433), .Y(exu_n19206));
INVX1 exu_U28907(.A(exu_n19206), .Y(exu_n9986));
AND2X1 exu_U28908(.A(ecl_wb_byplog_wen_w2), .B(ecl_byplog_rs3_match_w2), .Y(exu_n19210));
INVX1 exu_U28909(.A(exu_n19210), .Y(exu_n9987));
OR2X1 exu_U28910(.A(ecl_ifu_exu_rs3_d[2]), .B(exu_n19219), .Y(exu_n19218));
INVX1 exu_U28911(.A(exu_n19218), .Y(exu_n9988));
AND2X1 exu_U28912(.A(exu_n19235), .B(exu_n9990), .Y(exu_n19241));
INVX1 exu_U28913(.A(exu_n19241), .Y(exu_n9989));
AND2X1 exu_U28914(.A(exu_n19238), .B(exu_n15434), .Y(exu_n19242));
INVX1 exu_U28915(.A(exu_n19242), .Y(exu_n9990));
AND2X1 exu_U28916(.A(ecl_wb_byplog_wen_w2), .B(ecl_byplog_rs3h_match_w2), .Y(exu_n19246));
INVX1 exu_U28917(.A(exu_n19246), .Y(exu_n9991));
AND2X1 exu_U28918(.A(ecl_ecc_log_rs3_m), .B(ecc_rs3_err_m[6]), .Y(exu_n19923));
INVX1 exu_U28919(.A(exu_n19923), .Y(exu_n9992));
AND2X1 exu_U28920(.A(ecc_rs3_err_m[5]), .B(ecl_ecc_log_rs3_m), .Y(exu_n19927));
INVX1 exu_U28921(.A(exu_n19927), .Y(exu_n9993));
AND2X1 exu_U28922(.A(ecc_rs3_err_m[4]), .B(ecl_ecc_log_rs3_m), .Y(exu_n19931));
INVX1 exu_U28923(.A(exu_n19931), .Y(exu_n9994));
AND2X1 exu_U28924(.A(ecc_rs3_err_m[3]), .B(ecl_ecc_log_rs3_m), .Y(exu_n19935));
INVX1 exu_U28925(.A(exu_n19935), .Y(exu_n9995));
AND2X1 exu_U28926(.A(ecc_rs3_err_m[2]), .B(ecl_ecc_log_rs3_m), .Y(exu_n19939));
INVX1 exu_U28927(.A(exu_n19939), .Y(exu_n9996));
AND2X1 exu_U28928(.A(ecc_rs3_err_m[1]), .B(ecl_ecc_log_rs3_m), .Y(exu_n19943));
INVX1 exu_U28929(.A(exu_n19943), .Y(exu_n9997));
AND2X1 exu_U28930(.A(ecc_rs3_err_m[0]), .B(ecl_ecc_log_rs3_m), .Y(exu_n19947));
INVX1 exu_U28931(.A(exu_n19947), .Y(exu_n9998));
AND2X1 exu_U28932(.A(exu_n22049), .B(exu_n10000), .Y(bypass_rs2_data_w2[9]));
INVX1 exu_U28933(.A(bypass_rs2_data_w2[9]), .Y(exu_n9999));
AND2X1 exu_U28934(.A(exu_n15966), .B(lsu_exu_ldxa_data_g[9]), .Y(exu_n22050));
INVX1 exu_U28935(.A(exu_n22050), .Y(exu_n10000));
AND2X1 exu_U28936(.A(exu_n15965), .B(lsu_exu_ldxa_data_g[9]), .Y(exu_n22306));
INVX1 exu_U28937(.A(exu_n22306), .Y(exu_n10001));
AND2X1 exu_U28938(.A(lsu_exu_ldxa_data_g[8]), .B(exu_n15965), .Y(exu_n22310));
INVX1 exu_U28939(.A(exu_n22310), .Y(exu_n10002));
AND2X1 exu_U28940(.A(lsu_exu_ldxa_data_g[7]), .B(exu_n15965), .Y(exu_n22314));
INVX1 exu_U28941(.A(exu_n22314), .Y(exu_n10003));
AND2X1 exu_U28942(.A(lsu_exu_ldxa_data_g[6]), .B(exu_n19191), .Y(exu_n22318));
INVX1 exu_U28943(.A(exu_n22318), .Y(exu_n10004));
AND2X1 exu_U28944(.A(lsu_exu_ldxa_data_g[63]), .B(exu_n19191), .Y(exu_n22322));
INVX1 exu_U28945(.A(exu_n22322), .Y(exu_n10005));
AND2X1 exu_U28946(.A(lsu_exu_ldxa_data_g[62]), .B(exu_n19191), .Y(exu_n22326));
INVX1 exu_U28947(.A(exu_n22326), .Y(exu_n10006));
AND2X1 exu_U28948(.A(lsu_exu_ldxa_data_g[61]), .B(exu_n15965), .Y(exu_n22330));
INVX1 exu_U28949(.A(exu_n22330), .Y(exu_n10007));
AND2X1 exu_U28950(.A(lsu_exu_ldxa_data_g[60]), .B(exu_n19191), .Y(exu_n22334));
INVX1 exu_U28951(.A(exu_n22334), .Y(exu_n10008));
AND2X1 exu_U28952(.A(lsu_exu_ldxa_data_g[5]), .B(exu_n19191), .Y(exu_n22338));
INVX1 exu_U28953(.A(exu_n22338), .Y(exu_n10009));
AND2X1 exu_U28954(.A(lsu_exu_ldxa_data_g[59]), .B(exu_n19191), .Y(exu_n22342));
INVX1 exu_U28955(.A(exu_n22342), .Y(exu_n10010));
AND2X1 exu_U28956(.A(lsu_exu_ldxa_data_g[58]), .B(exu_n15965), .Y(exu_n22346));
INVX1 exu_U28957(.A(exu_n22346), .Y(exu_n10011));
AND2X1 exu_U28958(.A(lsu_exu_ldxa_data_g[57]), .B(exu_n19191), .Y(exu_n22350));
INVX1 exu_U28959(.A(exu_n22350), .Y(exu_n10012));
AND2X1 exu_U28960(.A(lsu_exu_ldxa_data_g[56]), .B(exu_n15965), .Y(exu_n22354));
INVX1 exu_U28961(.A(exu_n22354), .Y(exu_n10013));
AND2X1 exu_U28962(.A(lsu_exu_ldxa_data_g[55]), .B(exu_n19191), .Y(exu_n22358));
INVX1 exu_U28963(.A(exu_n22358), .Y(exu_n10014));
AND2X1 exu_U28964(.A(lsu_exu_ldxa_data_g[54]), .B(exu_n15965), .Y(exu_n22362));
INVX1 exu_U28965(.A(exu_n22362), .Y(exu_n10015));
AND2X1 exu_U28966(.A(lsu_exu_ldxa_data_g[53]), .B(exu_n15965), .Y(exu_n22366));
INVX1 exu_U28967(.A(exu_n22366), .Y(exu_n10016));
AND2X1 exu_U28968(.A(lsu_exu_ldxa_data_g[52]), .B(exu_n19191), .Y(exu_n22370));
INVX1 exu_U28969(.A(exu_n22370), .Y(exu_n10017));
AND2X1 exu_U28970(.A(lsu_exu_ldxa_data_g[51]), .B(exu_n19191), .Y(exu_n22374));
INVX1 exu_U28971(.A(exu_n22374), .Y(exu_n10018));
AND2X1 exu_U28972(.A(lsu_exu_ldxa_data_g[50]), .B(exu_n15965), .Y(exu_n22378));
INVX1 exu_U28973(.A(exu_n22378), .Y(exu_n10019));
AND2X1 exu_U28974(.A(lsu_exu_ldxa_data_g[4]), .B(exu_n19191), .Y(exu_n22382));
INVX1 exu_U28975(.A(exu_n22382), .Y(exu_n10020));
AND2X1 exu_U28976(.A(lsu_exu_ldxa_data_g[49]), .B(exu_n15965), .Y(exu_n22386));
INVX1 exu_U28977(.A(exu_n22386), .Y(exu_n10021));
AND2X1 exu_U28978(.A(lsu_exu_ldxa_data_g[48]), .B(exu_n15965), .Y(exu_n22390));
INVX1 exu_U28979(.A(exu_n22390), .Y(exu_n10022));
AND2X1 exu_U28980(.A(lsu_exu_ldxa_data_g[47]), .B(exu_n19191), .Y(exu_n22394));
INVX1 exu_U28981(.A(exu_n22394), .Y(exu_n10023));
AND2X1 exu_U28982(.A(lsu_exu_ldxa_data_g[46]), .B(exu_n19191), .Y(exu_n22398));
INVX1 exu_U28983(.A(exu_n22398), .Y(exu_n10024));
AND2X1 exu_U28984(.A(lsu_exu_ldxa_data_g[45]), .B(exu_n15965), .Y(exu_n22402));
INVX1 exu_U28985(.A(exu_n22402), .Y(exu_n10025));
AND2X1 exu_U28986(.A(lsu_exu_ldxa_data_g[44]), .B(exu_n15965), .Y(exu_n22406));
INVX1 exu_U28987(.A(exu_n22406), .Y(exu_n10026));
AND2X1 exu_U28988(.A(lsu_exu_ldxa_data_g[43]), .B(exu_n19191), .Y(exu_n22410));
INVX1 exu_U28989(.A(exu_n22410), .Y(exu_n10027));
AND2X1 exu_U28990(.A(lsu_exu_ldxa_data_g[42]), .B(exu_n19191), .Y(exu_n22414));
INVX1 exu_U28991(.A(exu_n22414), .Y(exu_n10028));
AND2X1 exu_U28992(.A(lsu_exu_ldxa_data_g[41]), .B(exu_n19191), .Y(exu_n22418));
INVX1 exu_U28993(.A(exu_n22418), .Y(exu_n10029));
AND2X1 exu_U28994(.A(lsu_exu_ldxa_data_g[40]), .B(exu_n15965), .Y(exu_n22422));
INVX1 exu_U28995(.A(exu_n22422), .Y(exu_n10030));
AND2X1 exu_U28996(.A(lsu_exu_ldxa_data_g[3]), .B(exu_n19191), .Y(exu_n22426));
INVX1 exu_U28997(.A(exu_n22426), .Y(exu_n10031));
AND2X1 exu_U28998(.A(lsu_exu_ldxa_data_g[39]), .B(exu_n15965), .Y(exu_n22430));
INVX1 exu_U28999(.A(exu_n22430), .Y(exu_n10032));
AND2X1 exu_U29000(.A(lsu_exu_ldxa_data_g[38]), .B(exu_n19191), .Y(exu_n22434));
INVX1 exu_U29001(.A(exu_n22434), .Y(exu_n10033));
AND2X1 exu_U29002(.A(lsu_exu_ldxa_data_g[37]), .B(exu_n19191), .Y(exu_n22438));
INVX1 exu_U29003(.A(exu_n22438), .Y(exu_n10034));
AND2X1 exu_U29004(.A(lsu_exu_ldxa_data_g[36]), .B(exu_n15965), .Y(exu_n22442));
INVX1 exu_U29005(.A(exu_n22442), .Y(exu_n10035));
AND2X1 exu_U29006(.A(lsu_exu_ldxa_data_g[35]), .B(exu_n15965), .Y(exu_n22446));
INVX1 exu_U29007(.A(exu_n22446), .Y(exu_n10036));
AND2X1 exu_U29008(.A(lsu_exu_ldxa_data_g[34]), .B(exu_n19191), .Y(exu_n22450));
INVX1 exu_U29009(.A(exu_n22450), .Y(exu_n10037));
AND2X1 exu_U29010(.A(lsu_exu_ldxa_data_g[33]), .B(exu_n15965), .Y(exu_n22454));
INVX1 exu_U29011(.A(exu_n22454), .Y(exu_n10038));
AND2X1 exu_U29012(.A(lsu_exu_ldxa_data_g[32]), .B(exu_n19191), .Y(exu_n22458));
INVX1 exu_U29013(.A(exu_n22458), .Y(exu_n10039));
AND2X1 exu_U29014(.A(lsu_exu_ldxa_data_g[31]), .B(exu_n19191), .Y(exu_n22462));
INVX1 exu_U29015(.A(exu_n22462), .Y(exu_n10040));
AND2X1 exu_U29016(.A(lsu_exu_ldxa_data_g[30]), .B(exu_n19191), .Y(exu_n22466));
INVX1 exu_U29017(.A(exu_n22466), .Y(exu_n10041));
AND2X1 exu_U29018(.A(lsu_exu_ldxa_data_g[2]), .B(exu_n15965), .Y(exu_n22470));
INVX1 exu_U29019(.A(exu_n22470), .Y(exu_n10042));
AND2X1 exu_U29020(.A(lsu_exu_ldxa_data_g[29]), .B(exu_n19191), .Y(exu_n22474));
INVX1 exu_U29021(.A(exu_n22474), .Y(exu_n10043));
AND2X1 exu_U29022(.A(lsu_exu_ldxa_data_g[28]), .B(exu_n19191), .Y(exu_n22478));
INVX1 exu_U29023(.A(exu_n22478), .Y(exu_n10044));
AND2X1 exu_U29024(.A(lsu_exu_ldxa_data_g[27]), .B(exu_n19191), .Y(exu_n22482));
INVX1 exu_U29025(.A(exu_n22482), .Y(exu_n10045));
AND2X1 exu_U29026(.A(lsu_exu_ldxa_data_g[26]), .B(exu_n15965), .Y(exu_n22486));
INVX1 exu_U29027(.A(exu_n22486), .Y(exu_n10046));
AND2X1 exu_U29028(.A(lsu_exu_ldxa_data_g[25]), .B(exu_n19191), .Y(exu_n22490));
INVX1 exu_U29029(.A(exu_n22490), .Y(exu_n10047));
AND2X1 exu_U29030(.A(lsu_exu_ldxa_data_g[24]), .B(exu_n19191), .Y(exu_n22494));
INVX1 exu_U29031(.A(exu_n22494), .Y(exu_n10048));
AND2X1 exu_U29032(.A(lsu_exu_ldxa_data_g[23]), .B(exu_n19191), .Y(exu_n22498));
INVX1 exu_U29033(.A(exu_n22498), .Y(exu_n10049));
AND2X1 exu_U29034(.A(lsu_exu_ldxa_data_g[22]), .B(exu_n19191), .Y(exu_n22502));
INVX1 exu_U29035(.A(exu_n22502), .Y(exu_n10050));
AND2X1 exu_U29036(.A(lsu_exu_ldxa_data_g[21]), .B(exu_n15965), .Y(exu_n22506));
INVX1 exu_U29037(.A(exu_n22506), .Y(exu_n10051));
AND2X1 exu_U29038(.A(lsu_exu_ldxa_data_g[20]), .B(exu_n19191), .Y(exu_n22510));
INVX1 exu_U29039(.A(exu_n22510), .Y(exu_n10052));
AND2X1 exu_U29040(.A(lsu_exu_ldxa_data_g[1]), .B(exu_n19191), .Y(exu_n22514));
INVX1 exu_U29041(.A(exu_n22514), .Y(exu_n10053));
AND2X1 exu_U29042(.A(lsu_exu_ldxa_data_g[19]), .B(exu_n15965), .Y(exu_n22518));
INVX1 exu_U29043(.A(exu_n22518), .Y(exu_n10054));
AND2X1 exu_U29044(.A(lsu_exu_ldxa_data_g[18]), .B(exu_n15965), .Y(exu_n22522));
INVX1 exu_U29045(.A(exu_n22522), .Y(exu_n10055));
AND2X1 exu_U29046(.A(lsu_exu_ldxa_data_g[17]), .B(exu_n15965), .Y(exu_n22526));
INVX1 exu_U29047(.A(exu_n22526), .Y(exu_n10056));
AND2X1 exu_U29048(.A(lsu_exu_ldxa_data_g[16]), .B(exu_n15965), .Y(exu_n22530));
INVX1 exu_U29049(.A(exu_n22530), .Y(exu_n10057));
AND2X1 exu_U29050(.A(lsu_exu_ldxa_data_g[15]), .B(exu_n15965), .Y(exu_n22534));
INVX1 exu_U29051(.A(exu_n22534), .Y(exu_n10058));
AND2X1 exu_U29052(.A(lsu_exu_ldxa_data_g[14]), .B(exu_n15965), .Y(exu_n22538));
INVX1 exu_U29053(.A(exu_n22538), .Y(exu_n10059));
AND2X1 exu_U29054(.A(lsu_exu_ldxa_data_g[13]), .B(exu_n15965), .Y(exu_n22542));
INVX1 exu_U29055(.A(exu_n22542), .Y(exu_n10060));
AND2X1 exu_U29056(.A(lsu_exu_ldxa_data_g[12]), .B(exu_n15965), .Y(exu_n22546));
INVX1 exu_U29057(.A(exu_n22546), .Y(exu_n10061));
AND2X1 exu_U29058(.A(lsu_exu_ldxa_data_g[11]), .B(exu_n15965), .Y(exu_n22550));
INVX1 exu_U29059(.A(exu_n22550), .Y(exu_n10062));
AND2X1 exu_U29060(.A(lsu_exu_ldxa_data_g[10]), .B(exu_n15965), .Y(exu_n22554));
INVX1 exu_U29061(.A(exu_n22554), .Y(exu_n10063));
AND2X1 exu_U29062(.A(lsu_exu_ldxa_data_g[0]), .B(exu_n15965), .Y(exu_n22558));
INVX1 exu_U29063(.A(exu_n22558), .Y(exu_n10064));
AND2X1 exu_U29064(.A(bypass_restore_rd_data[9]), .B(exu_n16268), .Y(exu_n30146));
INVX1 exu_U29065(.A(exu_n30146), .Y(exu_n10065));
AND2X1 exu_U29066(.A(bypass_restore_rd_data[8]), .B(exu_n16268), .Y(exu_n30148));
INVX1 exu_U29067(.A(exu_n30148), .Y(exu_n10066));
AND2X1 exu_U29068(.A(bypass_restore_rd_data[7]), .B(exu_n16268), .Y(exu_n30150));
INVX1 exu_U29069(.A(exu_n30150), .Y(exu_n10067));
AND2X1 exu_U29070(.A(bypass_restore_rd_data[6]), .B(exu_n16268), .Y(exu_n30152));
INVX1 exu_U29071(.A(exu_n30152), .Y(exu_n10068));
AND2X1 exu_U29072(.A(bypass_restore_rd_data[63]), .B(exu_n16268), .Y(exu_n30154));
INVX1 exu_U29073(.A(exu_n30154), .Y(exu_n10069));
AND2X1 exu_U29074(.A(bypass_restore_rd_data[62]), .B(exu_n16268), .Y(exu_n30156));
INVX1 exu_U29075(.A(exu_n30156), .Y(exu_n10070));
AND2X1 exu_U29076(.A(bypass_restore_rd_data[61]), .B(exu_n16268), .Y(exu_n30158));
INVX1 exu_U29077(.A(exu_n30158), .Y(exu_n10071));
AND2X1 exu_U29078(.A(bypass_restore_rd_data[60]), .B(exu_n16268), .Y(exu_n30160));
INVX1 exu_U29079(.A(exu_n30160), .Y(exu_n10072));
AND2X1 exu_U29080(.A(bypass_restore_rd_data[5]), .B(exu_n16268), .Y(exu_n30162));
INVX1 exu_U29081(.A(exu_n30162), .Y(exu_n10073));
AND2X1 exu_U29082(.A(bypass_restore_rd_data[59]), .B(exu_n16268), .Y(exu_n30164));
INVX1 exu_U29083(.A(exu_n30164), .Y(exu_n10074));
AND2X1 exu_U29084(.A(bypass_restore_rd_data[58]), .B(exu_n16268), .Y(exu_n30166));
INVX1 exu_U29085(.A(exu_n30166), .Y(exu_n10075));
AND2X1 exu_U29086(.A(bypass_restore_rd_data[57]), .B(exu_n16268), .Y(exu_n30168));
INVX1 exu_U29087(.A(exu_n30168), .Y(exu_n10076));
AND2X1 exu_U29088(.A(bypass_restore_rd_data[56]), .B(exu_n16268), .Y(exu_n30170));
INVX1 exu_U29089(.A(exu_n30170), .Y(exu_n10077));
AND2X1 exu_U29090(.A(bypass_restore_rd_data[55]), .B(exu_n16268), .Y(exu_n30172));
INVX1 exu_U29091(.A(exu_n30172), .Y(exu_n10078));
AND2X1 exu_U29092(.A(bypass_restore_rd_data[54]), .B(exu_n16268), .Y(exu_n30174));
INVX1 exu_U29093(.A(exu_n30174), .Y(exu_n10079));
AND2X1 exu_U29094(.A(bypass_restore_rd_data[53]), .B(exu_n16268), .Y(exu_n30176));
INVX1 exu_U29095(.A(exu_n30176), .Y(exu_n10080));
AND2X1 exu_U29096(.A(bypass_restore_rd_data[52]), .B(exu_n16268), .Y(exu_n30178));
INVX1 exu_U29097(.A(exu_n30178), .Y(exu_n10081));
AND2X1 exu_U29098(.A(bypass_restore_rd_data[51]), .B(exu_n16268), .Y(exu_n30180));
INVX1 exu_U29099(.A(exu_n30180), .Y(exu_n10082));
AND2X1 exu_U29100(.A(bypass_restore_rd_data[50]), .B(exu_n16268), .Y(exu_n30182));
INVX1 exu_U29101(.A(exu_n30182), .Y(exu_n10083));
AND2X1 exu_U29102(.A(bypass_restore_rd_data[4]), .B(exu_n16268), .Y(exu_n30184));
INVX1 exu_U29103(.A(exu_n30184), .Y(exu_n10084));
AND2X1 exu_U29104(.A(bypass_restore_rd_data[49]), .B(exu_n16268), .Y(exu_n30186));
INVX1 exu_U29105(.A(exu_n30186), .Y(exu_n10085));
AND2X1 exu_U29106(.A(bypass_restore_rd_data[48]), .B(exu_n16268), .Y(exu_n30188));
INVX1 exu_U29107(.A(exu_n30188), .Y(exu_n10086));
AND2X1 exu_U29108(.A(bypass_restore_rd_data[47]), .B(exu_n16268), .Y(exu_n30190));
INVX1 exu_U29109(.A(exu_n30190), .Y(exu_n10087));
AND2X1 exu_U29110(.A(bypass_restore_rd_data[46]), .B(exu_n16268), .Y(exu_n30192));
INVX1 exu_U29111(.A(exu_n30192), .Y(exu_n10088));
AND2X1 exu_U29112(.A(bypass_restore_rd_data[45]), .B(exu_n16268), .Y(exu_n30194));
INVX1 exu_U29113(.A(exu_n30194), .Y(exu_n10089));
AND2X1 exu_U29114(.A(bypass_restore_rd_data[44]), .B(exu_n16268), .Y(exu_n30196));
INVX1 exu_U29115(.A(exu_n30196), .Y(exu_n10090));
AND2X1 exu_U29116(.A(bypass_restore_rd_data[43]), .B(exu_n16268), .Y(exu_n30198));
INVX1 exu_U29117(.A(exu_n30198), .Y(exu_n10091));
AND2X1 exu_U29118(.A(bypass_restore_rd_data[42]), .B(exu_n16268), .Y(exu_n30200));
INVX1 exu_U29119(.A(exu_n30200), .Y(exu_n10092));
AND2X1 exu_U29120(.A(bypass_restore_rd_data[41]), .B(exu_n16268), .Y(exu_n30202));
INVX1 exu_U29121(.A(exu_n30202), .Y(exu_n10093));
AND2X1 exu_U29122(.A(bypass_restore_rd_data[40]), .B(exu_n16268), .Y(exu_n30204));
INVX1 exu_U29123(.A(exu_n30204), .Y(exu_n10094));
AND2X1 exu_U29124(.A(bypass_restore_rd_data[3]), .B(exu_n16268), .Y(exu_n30206));
INVX1 exu_U29125(.A(exu_n30206), .Y(exu_n10095));
AND2X1 exu_U29126(.A(bypass_restore_rd_data[39]), .B(exu_n16268), .Y(exu_n30208));
INVX1 exu_U29127(.A(exu_n30208), .Y(exu_n10096));
AND2X1 exu_U29128(.A(bypass_restore_rd_data[38]), .B(exu_n16268), .Y(exu_n30210));
INVX1 exu_U29129(.A(exu_n30210), .Y(exu_n10097));
AND2X1 exu_U29130(.A(bypass_restore_rd_data[37]), .B(exu_n16268), .Y(exu_n30212));
INVX1 exu_U29131(.A(exu_n30212), .Y(exu_n10098));
AND2X1 exu_U29132(.A(bypass_restore_rd_data[36]), .B(exu_n16268), .Y(exu_n30214));
INVX1 exu_U29133(.A(exu_n30214), .Y(exu_n10099));
AND2X1 exu_U29134(.A(bypass_restore_rd_data[35]), .B(exu_n16268), .Y(exu_n30216));
INVX1 exu_U29135(.A(exu_n30216), .Y(exu_n10100));
AND2X1 exu_U29136(.A(bypass_restore_rd_data[34]), .B(exu_n16268), .Y(exu_n30218));
INVX1 exu_U29137(.A(exu_n30218), .Y(exu_n10101));
AND2X1 exu_U29138(.A(bypass_restore_rd_data[33]), .B(exu_n16268), .Y(exu_n30220));
INVX1 exu_U29139(.A(exu_n30220), .Y(exu_n10102));
AND2X1 exu_U29140(.A(bypass_restore_rd_data[32]), .B(exu_n16268), .Y(exu_n30222));
INVX1 exu_U29141(.A(exu_n30222), .Y(exu_n10103));
AND2X1 exu_U29142(.A(bypass_restore_rd_data[31]), .B(exu_n16268), .Y(exu_n30224));
INVX1 exu_U29143(.A(exu_n30224), .Y(exu_n10104));
AND2X1 exu_U29144(.A(bypass_restore_rd_data[30]), .B(exu_n16268), .Y(exu_n30226));
INVX1 exu_U29145(.A(exu_n30226), .Y(exu_n10105));
AND2X1 exu_U29146(.A(bypass_restore_rd_data[2]), .B(exu_n16268), .Y(exu_n30228));
INVX1 exu_U29147(.A(exu_n30228), .Y(exu_n10106));
AND2X1 exu_U29148(.A(bypass_restore_rd_data[29]), .B(exu_n16268), .Y(exu_n30230));
INVX1 exu_U29149(.A(exu_n30230), .Y(exu_n10107));
AND2X1 exu_U29150(.A(bypass_restore_rd_data[28]), .B(exu_n16268), .Y(exu_n30232));
INVX1 exu_U29151(.A(exu_n30232), .Y(exu_n10108));
AND2X1 exu_U29152(.A(bypass_restore_rd_data[27]), .B(exu_n16268), .Y(exu_n30234));
INVX1 exu_U29153(.A(exu_n30234), .Y(exu_n10109));
AND2X1 exu_U29154(.A(bypass_restore_rd_data[26]), .B(exu_n16268), .Y(exu_n30236));
INVX1 exu_U29155(.A(exu_n30236), .Y(exu_n10110));
AND2X1 exu_U29156(.A(bypass_restore_rd_data[25]), .B(exu_n16268), .Y(exu_n30238));
INVX1 exu_U29157(.A(exu_n30238), .Y(exu_n10111));
AND2X1 exu_U29158(.A(bypass_restore_rd_data[24]), .B(exu_n16268), .Y(exu_n30240));
INVX1 exu_U29159(.A(exu_n30240), .Y(exu_n10112));
AND2X1 exu_U29160(.A(bypass_restore_rd_data[23]), .B(exu_n16268), .Y(exu_n30242));
INVX1 exu_U29161(.A(exu_n30242), .Y(exu_n10113));
AND2X1 exu_U29162(.A(bypass_restore_rd_data[22]), .B(exu_n16268), .Y(exu_n30244));
INVX1 exu_U29163(.A(exu_n30244), .Y(exu_n10114));
AND2X1 exu_U29164(.A(bypass_restore_rd_data[21]), .B(exu_n16268), .Y(exu_n30246));
INVX1 exu_U29165(.A(exu_n30246), .Y(exu_n10115));
AND2X1 exu_U29166(.A(bypass_restore_rd_data[20]), .B(exu_n16268), .Y(exu_n30248));
INVX1 exu_U29167(.A(exu_n30248), .Y(exu_n10116));
AND2X1 exu_U29168(.A(bypass_restore_rd_data[1]), .B(exu_n16268), .Y(exu_n30250));
INVX1 exu_U29169(.A(exu_n30250), .Y(exu_n10117));
AND2X1 exu_U29170(.A(bypass_restore_rd_data[19]), .B(exu_n16268), .Y(exu_n30252));
INVX1 exu_U29171(.A(exu_n30252), .Y(exu_n10118));
AND2X1 exu_U29172(.A(bypass_restore_rd_data[18]), .B(exu_n16268), .Y(exu_n30254));
INVX1 exu_U29173(.A(exu_n30254), .Y(exu_n10119));
AND2X1 exu_U29174(.A(bypass_restore_rd_data[17]), .B(exu_n16268), .Y(exu_n30256));
INVX1 exu_U29175(.A(exu_n30256), .Y(exu_n10120));
AND2X1 exu_U29176(.A(bypass_restore_rd_data[16]), .B(exu_n16268), .Y(exu_n30258));
INVX1 exu_U29177(.A(exu_n30258), .Y(exu_n10121));
AND2X1 exu_U29178(.A(bypass_restore_rd_data[15]), .B(exu_n16268), .Y(exu_n30260));
INVX1 exu_U29179(.A(exu_n30260), .Y(exu_n10122));
AND2X1 exu_U29180(.A(bypass_restore_rd_data[14]), .B(exu_n16268), .Y(exu_n30262));
INVX1 exu_U29181(.A(exu_n30262), .Y(exu_n10123));
AND2X1 exu_U29182(.A(bypass_restore_rd_data[13]), .B(exu_n16268), .Y(exu_n30264));
INVX1 exu_U29183(.A(exu_n30264), .Y(exu_n10124));
AND2X1 exu_U29184(.A(bypass_restore_rd_data[12]), .B(exu_n16268), .Y(exu_n30266));
INVX1 exu_U29185(.A(exu_n30266), .Y(exu_n10125));
AND2X1 exu_U29186(.A(bypass_restore_rd_data[11]), .B(exu_n16268), .Y(exu_n30268));
INVX1 exu_U29187(.A(exu_n30268), .Y(exu_n10126));
AND2X1 exu_U29188(.A(bypass_restore_rd_data[10]), .B(exu_n16268), .Y(exu_n30270));
INVX1 exu_U29189(.A(exu_n30270), .Y(exu_n10127));
AND2X1 exu_U29190(.A(bypass_restore_rd_data[0]), .B(exu_n16268), .Y(exu_n30272));
INVX1 exu_U29191(.A(exu_n30272), .Y(exu_n10128));
AND2X1 exu_U29192(.A(div_input_data_e[73]), .B(exu_n16168), .Y(exu_n30274));
INVX1 exu_U29193(.A(exu_n30274), .Y(exu_n10129));
AND2X1 exu_U29194(.A(div_input_data_e[72]), .B(exu_n16168), .Y(exu_n30276));
INVX1 exu_U29195(.A(exu_n30276), .Y(exu_n10130));
AND2X1 exu_U29196(.A(div_input_data_e[71]), .B(exu_n16169), .Y(exu_n30278));
INVX1 exu_U29197(.A(exu_n30278), .Y(exu_n10131));
AND2X1 exu_U29198(.A(div_input_data_e[70]), .B(exu_n16168), .Y(exu_n30280));
INVX1 exu_U29199(.A(exu_n30280), .Y(exu_n10132));
AND2X1 exu_U29200(.A(div_input_data_e[127]), .B(exu_n16167), .Y(exu_n30282));
INVX1 exu_U29201(.A(exu_n30282), .Y(exu_n10133));
AND2X1 exu_U29202(.A(div_input_data_e[126]), .B(exu_n16169), .Y(exu_n30284));
INVX1 exu_U29203(.A(exu_n30284), .Y(exu_n10134));
AND2X1 exu_U29204(.A(div_input_data_e[125]), .B(exu_n16170), .Y(exu_n30286));
INVX1 exu_U29205(.A(exu_n30286), .Y(exu_n10135));
AND2X1 exu_U29206(.A(div_input_data_e[124]), .B(exu_n16168), .Y(exu_n30288));
INVX1 exu_U29207(.A(exu_n30288), .Y(exu_n10136));
AND2X1 exu_U29208(.A(div_input_data_e[69]), .B(exu_n16167), .Y(exu_n30290));
INVX1 exu_U29209(.A(exu_n30290), .Y(exu_n10137));
AND2X1 exu_U29210(.A(div_input_data_e[123]), .B(exu_n16169), .Y(exu_n30292));
INVX1 exu_U29211(.A(exu_n30292), .Y(exu_n10138));
AND2X1 exu_U29212(.A(div_input_data_e[122]), .B(exu_n16167), .Y(exu_n30294));
INVX1 exu_U29213(.A(exu_n30294), .Y(exu_n10139));
AND2X1 exu_U29214(.A(div_input_data_e[121]), .B(exu_n16169), .Y(exu_n30296));
INVX1 exu_U29215(.A(exu_n30296), .Y(exu_n10140));
AND2X1 exu_U29216(.A(div_input_data_e[120]), .B(exu_n16170), .Y(exu_n30298));
INVX1 exu_U29217(.A(exu_n30298), .Y(exu_n10141));
AND2X1 exu_U29218(.A(div_input_data_e[119]), .B(exu_n16167), .Y(exu_n30300));
INVX1 exu_U29219(.A(exu_n30300), .Y(exu_n10142));
AND2X1 exu_U29220(.A(div_input_data_e[118]), .B(exu_n16168), .Y(exu_n30302));
INVX1 exu_U29221(.A(exu_n30302), .Y(exu_n10143));
AND2X1 exu_U29222(.A(div_input_data_e[117]), .B(exu_n16170), .Y(exu_n30304));
INVX1 exu_U29223(.A(exu_n30304), .Y(exu_n10144));
AND2X1 exu_U29224(.A(div_input_data_e[116]), .B(exu_n16169), .Y(exu_n30306));
INVX1 exu_U29225(.A(exu_n30306), .Y(exu_n10145));
AND2X1 exu_U29226(.A(div_input_data_e[115]), .B(exu_n16167), .Y(exu_n30308));
INVX1 exu_U29227(.A(exu_n30308), .Y(exu_n10146));
AND2X1 exu_U29228(.A(div_input_data_e[114]), .B(exu_n16168), .Y(exu_n30310));
INVX1 exu_U29229(.A(exu_n30310), .Y(exu_n10147));
AND2X1 exu_U29230(.A(div_input_data_e[68]), .B(exu_n16170), .Y(exu_n30312));
INVX1 exu_U29231(.A(exu_n30312), .Y(exu_n10148));
AND2X1 exu_U29232(.A(div_input_data_e[113]), .B(exu_n16169), .Y(exu_n30314));
INVX1 exu_U29233(.A(exu_n30314), .Y(exu_n10149));
AND2X1 exu_U29234(.A(div_input_data_e[112]), .B(exu_n16167), .Y(exu_n30316));
INVX1 exu_U29235(.A(exu_n30316), .Y(exu_n10150));
AND2X1 exu_U29236(.A(div_input_data_e[111]), .B(exu_n16168), .Y(exu_n30318));
INVX1 exu_U29237(.A(exu_n30318), .Y(exu_n10151));
AND2X1 exu_U29238(.A(div_input_data_e[110]), .B(exu_n16170), .Y(exu_n30320));
INVX1 exu_U29239(.A(exu_n30320), .Y(exu_n10152));
AND2X1 exu_U29240(.A(div_input_data_e[109]), .B(exu_n16169), .Y(exu_n30322));
INVX1 exu_U29241(.A(exu_n30322), .Y(exu_n10153));
AND2X1 exu_U29242(.A(div_input_data_e[108]), .B(exu_n16167), .Y(exu_n30324));
INVX1 exu_U29243(.A(exu_n30324), .Y(exu_n10154));
AND2X1 exu_U29244(.A(div_input_data_e[107]), .B(exu_n16168), .Y(exu_n30326));
INVX1 exu_U29245(.A(exu_n30326), .Y(exu_n10155));
AND2X1 exu_U29246(.A(div_input_data_e[106]), .B(exu_n16169), .Y(exu_n30328));
INVX1 exu_U29247(.A(exu_n30328), .Y(exu_n10156));
AND2X1 exu_U29248(.A(div_input_data_e[105]), .B(exu_n16169), .Y(exu_n30330));
INVX1 exu_U29249(.A(exu_n30330), .Y(exu_n10157));
AND2X1 exu_U29250(.A(div_input_data_e[104]), .B(exu_n16169), .Y(exu_n30332));
INVX1 exu_U29251(.A(exu_n30332), .Y(exu_n10158));
AND2X1 exu_U29252(.A(div_input_data_e[67]), .B(exu_n16169), .Y(exu_n30334));
INVX1 exu_U29253(.A(exu_n30334), .Y(exu_n10159));
AND2X1 exu_U29254(.A(div_input_data_e[103]), .B(exu_n16169), .Y(exu_n30336));
INVX1 exu_U29255(.A(exu_n30336), .Y(exu_n10160));
AND2X1 exu_U29256(.A(div_input_data_e[102]), .B(exu_n16169), .Y(exu_n30338));
INVX1 exu_U29257(.A(exu_n30338), .Y(exu_n10161));
AND2X1 exu_U29258(.A(div_input_data_e[101]), .B(exu_n16169), .Y(exu_n30340));
INVX1 exu_U29259(.A(exu_n30340), .Y(exu_n10162));
AND2X1 exu_U29260(.A(div_input_data_e[100]), .B(exu_n16169), .Y(exu_n30342));
INVX1 exu_U29261(.A(exu_n30342), .Y(exu_n10163));
AND2X1 exu_U29262(.A(div_input_data_e[99]), .B(exu_n16169), .Y(exu_n30344));
INVX1 exu_U29263(.A(exu_n30344), .Y(exu_n10164));
AND2X1 exu_U29264(.A(div_input_data_e[98]), .B(exu_n16169), .Y(exu_n30346));
INVX1 exu_U29265(.A(exu_n30346), .Y(exu_n10165));
AND2X1 exu_U29266(.A(div_input_data_e[97]), .B(exu_n16169), .Y(exu_n30348));
INVX1 exu_U29267(.A(exu_n30348), .Y(exu_n10166));
AND2X1 exu_U29268(.A(div_input_data_e[96]), .B(exu_n16169), .Y(exu_n30350));
INVX1 exu_U29269(.A(exu_n30350), .Y(exu_n10167));
AND2X1 exu_U29270(.A(div_input_data_e[95]), .B(exu_n16169), .Y(exu_n30352));
INVX1 exu_U29271(.A(exu_n30352), .Y(exu_n10168));
AND2X1 exu_U29272(.A(div_input_data_e[94]), .B(exu_n16170), .Y(exu_n30354));
INVX1 exu_U29273(.A(exu_n30354), .Y(exu_n10169));
AND2X1 exu_U29274(.A(div_input_data_e[66]), .B(exu_n16170), .Y(exu_n30356));
INVX1 exu_U29275(.A(exu_n30356), .Y(exu_n10170));
AND2X1 exu_U29276(.A(div_input_data_e[93]), .B(exu_n16170), .Y(exu_n30358));
INVX1 exu_U29277(.A(exu_n30358), .Y(exu_n10171));
AND2X1 exu_U29278(.A(div_input_data_e[92]), .B(exu_n16170), .Y(exu_n30360));
INVX1 exu_U29279(.A(exu_n30360), .Y(exu_n10172));
AND2X1 exu_U29280(.A(div_input_data_e[91]), .B(exu_n16170), .Y(exu_n30362));
INVX1 exu_U29281(.A(exu_n30362), .Y(exu_n10173));
AND2X1 exu_U29282(.A(div_input_data_e[90]), .B(exu_n16170), .Y(exu_n30364));
INVX1 exu_U29283(.A(exu_n30364), .Y(exu_n10174));
AND2X1 exu_U29284(.A(div_input_data_e[89]), .B(exu_n16170), .Y(exu_n30366));
INVX1 exu_U29285(.A(exu_n30366), .Y(exu_n10175));
AND2X1 exu_U29286(.A(div_input_data_e[88]), .B(exu_n16170), .Y(exu_n30368));
INVX1 exu_U29287(.A(exu_n30368), .Y(exu_n10176));
AND2X1 exu_U29288(.A(div_input_data_e[87]), .B(exu_n16170), .Y(exu_n30370));
INVX1 exu_U29289(.A(exu_n30370), .Y(exu_n10177));
AND2X1 exu_U29290(.A(div_input_data_e[86]), .B(exu_n16170), .Y(exu_n30372));
INVX1 exu_U29291(.A(exu_n30372), .Y(exu_n10178));
AND2X1 exu_U29292(.A(div_input_data_e[85]), .B(exu_n16170), .Y(exu_n30374));
INVX1 exu_U29293(.A(exu_n30374), .Y(exu_n10179));
AND2X1 exu_U29294(.A(div_input_data_e[84]), .B(exu_n16170), .Y(exu_n30376));
INVX1 exu_U29295(.A(exu_n30376), .Y(exu_n10180));
AND2X1 exu_U29296(.A(div_input_data_e[65]), .B(exu_n16170), .Y(exu_n30378));
INVX1 exu_U29297(.A(exu_n30378), .Y(exu_n10181));
AND2X1 exu_U29298(.A(div_input_data_e[83]), .B(exu_n16167), .Y(exu_n30380));
INVX1 exu_U29299(.A(exu_n30380), .Y(exu_n10182));
AND2X1 exu_U29300(.A(div_input_data_e[82]), .B(exu_n16167), .Y(exu_n30382));
INVX1 exu_U29301(.A(exu_n30382), .Y(exu_n10183));
AND2X1 exu_U29302(.A(div_input_data_e[81]), .B(exu_n16167), .Y(exu_n30384));
INVX1 exu_U29303(.A(exu_n30384), .Y(exu_n10184));
AND2X1 exu_U29304(.A(div_input_data_e[80]), .B(exu_n16167), .Y(exu_n30386));
INVX1 exu_U29305(.A(exu_n30386), .Y(exu_n10185));
AND2X1 exu_U29306(.A(div_input_data_e[79]), .B(exu_n16167), .Y(exu_n30388));
INVX1 exu_U29307(.A(exu_n30388), .Y(exu_n10186));
AND2X1 exu_U29308(.A(div_input_data_e[78]), .B(exu_n16167), .Y(exu_n30390));
INVX1 exu_U29309(.A(exu_n30390), .Y(exu_n10187));
AND2X1 exu_U29310(.A(div_input_data_e[77]), .B(exu_n16167), .Y(exu_n30392));
INVX1 exu_U29311(.A(exu_n30392), .Y(exu_n10188));
AND2X1 exu_U29312(.A(div_input_data_e[76]), .B(exu_n16167), .Y(exu_n30394));
INVX1 exu_U29313(.A(exu_n30394), .Y(exu_n10189));
AND2X1 exu_U29314(.A(div_input_data_e[75]), .B(exu_n16167), .Y(exu_n30396));
INVX1 exu_U29315(.A(exu_n30396), .Y(exu_n10190));
AND2X1 exu_U29316(.A(div_input_data_e[74]), .B(exu_n16167), .Y(exu_n30398));
INVX1 exu_U29317(.A(exu_n30398), .Y(exu_n10191));
AND2X1 exu_U29318(.A(div_input_data_e[64]), .B(exu_n16167), .Y(exu_n30400));
INVX1 exu_U29319(.A(exu_n30400), .Y(exu_n10192));
AND2X1 exu_U29320(.A(exu_ifu_brpc_e[9]), .B(exu_n16262), .Y(exu_n30498));
INVX1 exu_U29321(.A(exu_n30498), .Y(exu_n10193));
AND2X1 exu_U29322(.A(exu_ifu_brpc_e[8]), .B(exu_n16262), .Y(exu_n30500));
INVX1 exu_U29323(.A(exu_n30500), .Y(exu_n10194));
AND2X1 exu_U29324(.A(exu_ifu_brpc_e[7]), .B(exu_n16262), .Y(exu_n30502));
INVX1 exu_U29325(.A(exu_n30502), .Y(exu_n10195));
AND2X1 exu_U29326(.A(exu_ifu_brpc_e[6]), .B(exu_n16262), .Y(exu_n30504));
INVX1 exu_U29327(.A(exu_n30504), .Y(exu_n10196));
AND2X1 exu_U29328(.A(exu_ifu_brpc_e[5]), .B(exu_n16262), .Y(exu_n30514));
INVX1 exu_U29329(.A(exu_n30514), .Y(exu_n10197));
AND2X1 exu_U29330(.A(exu_ifu_brpc_e[4]), .B(exu_n16262), .Y(exu_n30536));
INVX1 exu_U29331(.A(exu_n30536), .Y(exu_n10198));
AND2X1 exu_U29332(.A(exu_ifu_brpc_e[46]), .B(exu_n16262), .Y(exu_n30544));
INVX1 exu_U29333(.A(exu_n30544), .Y(exu_n10199));
AND2X1 exu_U29334(.A(exu_ifu_brpc_e[45]), .B(exu_n16262), .Y(exu_n30546));
INVX1 exu_U29335(.A(exu_n30546), .Y(exu_n10200));
AND2X1 exu_U29336(.A(exu_ifu_brpc_e[44]), .B(exu_n16262), .Y(exu_n30548));
INVX1 exu_U29337(.A(exu_n30548), .Y(exu_n10201));
AND2X1 exu_U29338(.A(exu_ifu_brpc_e[43]), .B(exu_n16262), .Y(exu_n30550));
INVX1 exu_U29339(.A(exu_n30550), .Y(exu_n10202));
AND2X1 exu_U29340(.A(exu_ifu_brpc_e[42]), .B(exu_n16262), .Y(exu_n30552));
INVX1 exu_U29341(.A(exu_n30552), .Y(exu_n10203));
AND2X1 exu_U29342(.A(exu_ifu_brpc_e[41]), .B(exu_n16262), .Y(exu_n30554));
INVX1 exu_U29343(.A(exu_n30554), .Y(exu_n10204));
AND2X1 exu_U29344(.A(exu_ifu_brpc_e[40]), .B(exu_n16262), .Y(exu_n30556));
INVX1 exu_U29345(.A(exu_n30556), .Y(exu_n10205));
AND2X1 exu_U29346(.A(exu_ifu_brpc_e[3]), .B(exu_n16262), .Y(exu_n30558));
INVX1 exu_U29347(.A(exu_n30558), .Y(exu_n10206));
AND2X1 exu_U29348(.A(exu_ifu_brpc_e[39]), .B(exu_n16262), .Y(exu_n30560));
INVX1 exu_U29349(.A(exu_n30560), .Y(exu_n10207));
AND2X1 exu_U29350(.A(exu_ifu_brpc_e[38]), .B(exu_n16262), .Y(exu_n30562));
INVX1 exu_U29351(.A(exu_n30562), .Y(exu_n10208));
AND2X1 exu_U29352(.A(exu_ifu_brpc_e[37]), .B(exu_n16262), .Y(exu_n30564));
INVX1 exu_U29353(.A(exu_n30564), .Y(exu_n10209));
AND2X1 exu_U29354(.A(exu_ifu_brpc_e[36]), .B(exu_n16262), .Y(exu_n30566));
INVX1 exu_U29355(.A(exu_n30566), .Y(exu_n10210));
AND2X1 exu_U29356(.A(exu_ifu_brpc_e[35]), .B(exu_n16262), .Y(exu_n30568));
INVX1 exu_U29357(.A(exu_n30568), .Y(exu_n10211));
AND2X1 exu_U29358(.A(exu_ifu_brpc_e[34]), .B(exu_n16262), .Y(exu_n30570));
INVX1 exu_U29359(.A(exu_n30570), .Y(exu_n10212));
AND2X1 exu_U29360(.A(exu_ifu_brpc_e[33]), .B(exu_n16262), .Y(exu_n30572));
INVX1 exu_U29361(.A(exu_n30572), .Y(exu_n10213));
AND2X1 exu_U29362(.A(exu_ifu_brpc_e[32]), .B(exu_n16262), .Y(exu_n30574));
INVX1 exu_U29363(.A(exu_n30574), .Y(exu_n10214));
AND2X1 exu_U29364(.A(exu_ifu_brpc_e[31]), .B(exu_n16262), .Y(exu_n30576));
INVX1 exu_U29365(.A(exu_n30576), .Y(exu_n10215));
AND2X1 exu_U29366(.A(exu_ifu_brpc_e[30]), .B(exu_n16262), .Y(exu_n30578));
INVX1 exu_U29367(.A(exu_n30578), .Y(exu_n10216));
AND2X1 exu_U29368(.A(exu_ifu_brpc_e[2]), .B(exu_n16262), .Y(exu_n30580));
INVX1 exu_U29369(.A(exu_n30580), .Y(exu_n10217));
AND2X1 exu_U29370(.A(exu_ifu_brpc_e[29]), .B(exu_n16262), .Y(exu_n30582));
INVX1 exu_U29371(.A(exu_n30582), .Y(exu_n10218));
AND2X1 exu_U29372(.A(exu_ifu_brpc_e[28]), .B(exu_n16262), .Y(exu_n30584));
INVX1 exu_U29373(.A(exu_n30584), .Y(exu_n10219));
AND2X1 exu_U29374(.A(exu_ifu_brpc_e[27]), .B(exu_n16262), .Y(exu_n30586));
INVX1 exu_U29375(.A(exu_n30586), .Y(exu_n10220));
AND2X1 exu_U29376(.A(exu_ifu_brpc_e[26]), .B(exu_n16262), .Y(exu_n30588));
INVX1 exu_U29377(.A(exu_n30588), .Y(exu_n10221));
AND2X1 exu_U29378(.A(exu_ifu_brpc_e[25]), .B(exu_n16262), .Y(exu_n30590));
INVX1 exu_U29379(.A(exu_n30590), .Y(exu_n10222));
AND2X1 exu_U29380(.A(exu_ifu_brpc_e[24]), .B(exu_n16262), .Y(exu_n30592));
INVX1 exu_U29381(.A(exu_n30592), .Y(exu_n10223));
AND2X1 exu_U29382(.A(exu_ifu_brpc_e[23]), .B(exu_n16262), .Y(exu_n30594));
INVX1 exu_U29383(.A(exu_n30594), .Y(exu_n10224));
AND2X1 exu_U29384(.A(exu_ifu_brpc_e[22]), .B(exu_n16262), .Y(exu_n30596));
INVX1 exu_U29385(.A(exu_n30596), .Y(exu_n10225));
AND2X1 exu_U29386(.A(exu_ifu_brpc_e[21]), .B(exu_n16262), .Y(exu_n30598));
INVX1 exu_U29387(.A(exu_n30598), .Y(exu_n10226));
AND2X1 exu_U29388(.A(exu_ifu_brpc_e[20]), .B(exu_n16262), .Y(exu_n30600));
INVX1 exu_U29389(.A(exu_n30600), .Y(exu_n10227));
AND2X1 exu_U29390(.A(exu_ifu_brpc_e[1]), .B(exu_n16262), .Y(exu_n30602));
INVX1 exu_U29391(.A(exu_n30602), .Y(exu_n10228));
AND2X1 exu_U29392(.A(exu_ifu_brpc_e[19]), .B(exu_n16262), .Y(exu_n30604));
INVX1 exu_U29393(.A(exu_n30604), .Y(exu_n10229));
AND2X1 exu_U29394(.A(exu_ifu_brpc_e[18]), .B(exu_n16262), .Y(exu_n30606));
INVX1 exu_U29395(.A(exu_n30606), .Y(exu_n10230));
AND2X1 exu_U29396(.A(exu_ifu_brpc_e[17]), .B(exu_n16262), .Y(exu_n30608));
INVX1 exu_U29397(.A(exu_n30608), .Y(exu_n10231));
AND2X1 exu_U29398(.A(exu_ifu_brpc_e[16]), .B(exu_n16262), .Y(exu_n30610));
INVX1 exu_U29399(.A(exu_n30610), .Y(exu_n10232));
AND2X1 exu_U29400(.A(exu_ifu_brpc_e[15]), .B(exu_n16262), .Y(exu_n30612));
INVX1 exu_U29401(.A(exu_n30612), .Y(exu_n10233));
AND2X1 exu_U29402(.A(exu_ifu_brpc_e[14]), .B(exu_n16262), .Y(exu_n30614));
INVX1 exu_U29403(.A(exu_n30614), .Y(exu_n10234));
AND2X1 exu_U29404(.A(exu_ifu_brpc_e[13]), .B(exu_n16262), .Y(exu_n30616));
INVX1 exu_U29405(.A(exu_n30616), .Y(exu_n10235));
AND2X1 exu_U29406(.A(exu_ifu_brpc_e[12]), .B(exu_n16262), .Y(exu_n30618));
INVX1 exu_U29407(.A(exu_n30618), .Y(exu_n10236));
AND2X1 exu_U29408(.A(exu_ifu_brpc_e[11]), .B(exu_n16262), .Y(exu_n30620));
INVX1 exu_U29409(.A(exu_n30620), .Y(exu_n10237));
AND2X1 exu_U29410(.A(exu_ifu_brpc_e[10]), .B(exu_n16262), .Y(exu_n30622));
INVX1 exu_U29411(.A(exu_n30622), .Y(exu_n10238));
AND2X1 exu_U29412(.A(exu_ifu_brpc_e[0]), .B(exu_n16262), .Y(exu_n30624));
INVX1 exu_U29413(.A(exu_n30624), .Y(exu_n10239));
AND2X1 exu_U29414(.A(exu_n11234), .B(exu_n10241), .Y(shft_alu_shift_out_e[9]));
INVX1 exu_U29415(.A(shft_alu_shift_out_e[9]), .Y(exu_n10240));
AND2X1 exu_U29416(.A(shft_lshift1[9]), .B(exu_n16236), .Y(exu_n30754));
INVX1 exu_U29417(.A(exu_n30754), .Y(exu_n10241));
AND2X1 exu_U29418(.A(exu_n11361), .B(exu_n10243), .Y(div_byp_muldivout_g[9]));
INVX1 exu_U29419(.A(div_byp_muldivout_g[9]), .Y(exu_n10242));
AND2X1 exu_U29420(.A(div_mul_result[9]), .B(exu_n16199), .Y(exu_n30882));
INVX1 exu_U29421(.A(exu_n30882), .Y(exu_n10243));
AND2X1 exu_U29422(.A(div_mul_result[9]), .B(exu_n16186), .Y(exu_n31330));
INVX1 exu_U29423(.A(exu_n31330), .Y(exu_n10244));
AND2X1 exu_U29424(.A(div_mul_result[8]), .B(exu_n16186), .Y(exu_n31332));
INVX1 exu_U29425(.A(exu_n31332), .Y(exu_n10245));
AND2X1 exu_U29426(.A(div_mul_result[7]), .B(exu_n16186), .Y(exu_n31334));
INVX1 exu_U29427(.A(exu_n31334), .Y(exu_n10246));
AND2X1 exu_U29428(.A(div_mul_result[6]), .B(exu_n16186), .Y(exu_n31336));
INVX1 exu_U29429(.A(exu_n31336), .Y(exu_n10247));
AND2X1 exu_U29430(.A(div_mul_result[63]), .B(exu_n16186), .Y(exu_n31338));
INVX1 exu_U29431(.A(exu_n31338), .Y(exu_n10248));
AND2X1 exu_U29432(.A(div_mul_result[62]), .B(exu_n16186), .Y(exu_n31340));
INVX1 exu_U29433(.A(exu_n31340), .Y(exu_n10249));
AND2X1 exu_U29434(.A(div_mul_result[61]), .B(exu_n16186), .Y(exu_n31342));
INVX1 exu_U29435(.A(exu_n31342), .Y(exu_n10250));
AND2X1 exu_U29436(.A(div_mul_result[60]), .B(exu_n16186), .Y(exu_n31344));
INVX1 exu_U29437(.A(exu_n31344), .Y(exu_n10251));
AND2X1 exu_U29438(.A(div_mul_result[5]), .B(exu_n16186), .Y(exu_n31346));
INVX1 exu_U29439(.A(exu_n31346), .Y(exu_n10252));
AND2X1 exu_U29440(.A(div_mul_result[59]), .B(exu_n16186), .Y(exu_n31348));
INVX1 exu_U29441(.A(exu_n31348), .Y(exu_n10253));
AND2X1 exu_U29442(.A(div_mul_result[58]), .B(exu_n16186), .Y(exu_n31350));
INVX1 exu_U29443(.A(exu_n31350), .Y(exu_n10254));
AND2X1 exu_U29444(.A(div_mul_result[57]), .B(exu_n16186), .Y(exu_n31352));
INVX1 exu_U29445(.A(exu_n31352), .Y(exu_n10255));
AND2X1 exu_U29446(.A(div_mul_result[56]), .B(exu_n16186), .Y(exu_n31354));
INVX1 exu_U29447(.A(exu_n31354), .Y(exu_n10256));
AND2X1 exu_U29448(.A(div_mul_result[55]), .B(exu_n16186), .Y(exu_n31356));
INVX1 exu_U29449(.A(exu_n31356), .Y(exu_n10257));
AND2X1 exu_U29450(.A(div_mul_result[54]), .B(exu_n16186), .Y(exu_n31358));
INVX1 exu_U29451(.A(exu_n31358), .Y(exu_n10258));
AND2X1 exu_U29452(.A(div_mul_result[53]), .B(exu_n16186), .Y(exu_n31360));
INVX1 exu_U29453(.A(exu_n31360), .Y(exu_n10259));
AND2X1 exu_U29454(.A(div_mul_result[52]), .B(exu_n16186), .Y(exu_n31362));
INVX1 exu_U29455(.A(exu_n31362), .Y(exu_n10260));
AND2X1 exu_U29456(.A(div_mul_result[51]), .B(exu_n16186), .Y(exu_n31364));
INVX1 exu_U29457(.A(exu_n31364), .Y(exu_n10261));
AND2X1 exu_U29458(.A(div_mul_result[50]), .B(exu_n16186), .Y(exu_n31366));
INVX1 exu_U29459(.A(exu_n31366), .Y(exu_n10262));
AND2X1 exu_U29460(.A(div_mul_result[4]), .B(exu_n16186), .Y(exu_n31368));
INVX1 exu_U29461(.A(exu_n31368), .Y(exu_n10263));
AND2X1 exu_U29462(.A(div_mul_result[49]), .B(exu_n16186), .Y(exu_n31370));
INVX1 exu_U29463(.A(exu_n31370), .Y(exu_n10264));
AND2X1 exu_U29464(.A(div_mul_result[48]), .B(exu_n16186), .Y(exu_n31372));
INVX1 exu_U29465(.A(exu_n31372), .Y(exu_n10265));
AND2X1 exu_U29466(.A(div_mul_result[47]), .B(exu_n16186), .Y(exu_n31374));
INVX1 exu_U29467(.A(exu_n31374), .Y(exu_n10266));
AND2X1 exu_U29468(.A(div_mul_result[46]), .B(exu_n16186), .Y(exu_n31376));
INVX1 exu_U29469(.A(exu_n31376), .Y(exu_n10267));
AND2X1 exu_U29470(.A(div_mul_result[45]), .B(exu_n16186), .Y(exu_n31378));
INVX1 exu_U29471(.A(exu_n31378), .Y(exu_n10268));
AND2X1 exu_U29472(.A(div_mul_result[44]), .B(exu_n16186), .Y(exu_n31380));
INVX1 exu_U29473(.A(exu_n31380), .Y(exu_n10269));
AND2X1 exu_U29474(.A(div_mul_result[43]), .B(exu_n16186), .Y(exu_n31382));
INVX1 exu_U29475(.A(exu_n31382), .Y(exu_n10270));
AND2X1 exu_U29476(.A(div_mul_result[42]), .B(exu_n16186), .Y(exu_n31384));
INVX1 exu_U29477(.A(exu_n31384), .Y(exu_n10271));
AND2X1 exu_U29478(.A(div_mul_result[41]), .B(exu_n16186), .Y(exu_n31386));
INVX1 exu_U29479(.A(exu_n31386), .Y(exu_n10272));
AND2X1 exu_U29480(.A(div_mul_result[40]), .B(exu_n16186), .Y(exu_n31388));
INVX1 exu_U29481(.A(exu_n31388), .Y(exu_n10273));
AND2X1 exu_U29482(.A(div_mul_result[3]), .B(exu_n16186), .Y(exu_n31390));
INVX1 exu_U29483(.A(exu_n31390), .Y(exu_n10274));
AND2X1 exu_U29484(.A(div_mul_result[39]), .B(exu_n16186), .Y(exu_n31392));
INVX1 exu_U29485(.A(exu_n31392), .Y(exu_n10275));
AND2X1 exu_U29486(.A(div_mul_result[38]), .B(exu_n16186), .Y(exu_n31394));
INVX1 exu_U29487(.A(exu_n31394), .Y(exu_n10276));
AND2X1 exu_U29488(.A(div_mul_result[37]), .B(exu_n16186), .Y(exu_n31396));
INVX1 exu_U29489(.A(exu_n31396), .Y(exu_n10277));
AND2X1 exu_U29490(.A(div_mul_result[36]), .B(exu_n16186), .Y(exu_n31398));
INVX1 exu_U29491(.A(exu_n31398), .Y(exu_n10278));
AND2X1 exu_U29492(.A(div_mul_result[35]), .B(exu_n16186), .Y(exu_n31400));
INVX1 exu_U29493(.A(exu_n31400), .Y(exu_n10279));
AND2X1 exu_U29494(.A(div_mul_result[34]), .B(exu_n16186), .Y(exu_n31402));
INVX1 exu_U29495(.A(exu_n31402), .Y(exu_n10280));
AND2X1 exu_U29496(.A(div_mul_result[33]), .B(exu_n16186), .Y(exu_n31404));
INVX1 exu_U29497(.A(exu_n31404), .Y(exu_n10281));
AND2X1 exu_U29498(.A(div_mul_result[32]), .B(exu_n16186), .Y(exu_n31406));
INVX1 exu_U29499(.A(exu_n31406), .Y(exu_n10282));
AND2X1 exu_U29500(.A(div_mul_result[31]), .B(exu_n16186), .Y(exu_n31408));
INVX1 exu_U29501(.A(exu_n31408), .Y(exu_n10283));
AND2X1 exu_U29502(.A(div_mul_result[30]), .B(exu_n16186), .Y(exu_n31410));
INVX1 exu_U29503(.A(exu_n31410), .Y(exu_n10284));
AND2X1 exu_U29504(.A(div_mul_result[2]), .B(exu_n16186), .Y(exu_n31412));
INVX1 exu_U29505(.A(exu_n31412), .Y(exu_n10285));
AND2X1 exu_U29506(.A(div_mul_result[29]), .B(exu_n16186), .Y(exu_n31414));
INVX1 exu_U29507(.A(exu_n31414), .Y(exu_n10286));
AND2X1 exu_U29508(.A(div_mul_result[28]), .B(exu_n16186), .Y(exu_n31416));
INVX1 exu_U29509(.A(exu_n31416), .Y(exu_n10287));
AND2X1 exu_U29510(.A(div_mul_result[27]), .B(exu_n16186), .Y(exu_n31418));
INVX1 exu_U29511(.A(exu_n31418), .Y(exu_n10288));
AND2X1 exu_U29512(.A(div_mul_result[26]), .B(exu_n16186), .Y(exu_n31420));
INVX1 exu_U29513(.A(exu_n31420), .Y(exu_n10289));
AND2X1 exu_U29514(.A(div_mul_result[25]), .B(exu_n16186), .Y(exu_n31422));
INVX1 exu_U29515(.A(exu_n31422), .Y(exu_n10290));
AND2X1 exu_U29516(.A(div_mul_result[24]), .B(exu_n16186), .Y(exu_n31424));
INVX1 exu_U29517(.A(exu_n31424), .Y(exu_n10291));
AND2X1 exu_U29518(.A(div_mul_result[23]), .B(exu_n16186), .Y(exu_n31426));
INVX1 exu_U29519(.A(exu_n31426), .Y(exu_n10292));
AND2X1 exu_U29520(.A(div_mul_result[22]), .B(exu_n16186), .Y(exu_n31428));
INVX1 exu_U29521(.A(exu_n31428), .Y(exu_n10293));
AND2X1 exu_U29522(.A(div_mul_result[21]), .B(exu_n16186), .Y(exu_n31430));
INVX1 exu_U29523(.A(exu_n31430), .Y(exu_n10294));
AND2X1 exu_U29524(.A(div_mul_result[20]), .B(exu_n16186), .Y(exu_n31432));
INVX1 exu_U29525(.A(exu_n31432), .Y(exu_n10295));
AND2X1 exu_U29526(.A(div_mul_result[1]), .B(exu_n16186), .Y(exu_n31434));
INVX1 exu_U29527(.A(exu_n31434), .Y(exu_n10296));
AND2X1 exu_U29528(.A(div_mul_result[19]), .B(exu_n16186), .Y(exu_n31436));
INVX1 exu_U29529(.A(exu_n31436), .Y(exu_n10297));
AND2X1 exu_U29530(.A(div_mul_result[18]), .B(exu_n16186), .Y(exu_n31438));
INVX1 exu_U29531(.A(exu_n31438), .Y(exu_n10298));
AND2X1 exu_U29532(.A(div_mul_result[17]), .B(exu_n16186), .Y(exu_n31440));
INVX1 exu_U29533(.A(exu_n31440), .Y(exu_n10299));
AND2X1 exu_U29534(.A(div_mul_result[16]), .B(exu_n16186), .Y(exu_n31442));
INVX1 exu_U29535(.A(exu_n31442), .Y(exu_n10300));
AND2X1 exu_U29536(.A(div_mul_result[15]), .B(exu_n16186), .Y(exu_n31444));
INVX1 exu_U29537(.A(exu_n31444), .Y(exu_n10301));
AND2X1 exu_U29538(.A(div_mul_result[14]), .B(exu_n16186), .Y(exu_n31446));
INVX1 exu_U29539(.A(exu_n31446), .Y(exu_n10302));
AND2X1 exu_U29540(.A(div_mul_result[13]), .B(exu_n16186), .Y(exu_n31448));
INVX1 exu_U29541(.A(exu_n31448), .Y(exu_n10303));
AND2X1 exu_U29542(.A(div_mul_result[12]), .B(exu_n16186), .Y(exu_n31450));
INVX1 exu_U29543(.A(exu_n31450), .Y(exu_n10304));
AND2X1 exu_U29544(.A(div_mul_result[11]), .B(exu_n16186), .Y(exu_n31452));
INVX1 exu_U29545(.A(exu_n31452), .Y(exu_n10305));
AND2X1 exu_U29546(.A(div_mul_result[10]), .B(exu_n16186), .Y(exu_n31454));
INVX1 exu_U29547(.A(exu_n31454), .Y(exu_n10306));
AND2X1 exu_U29548(.A(div_mul_result[0]), .B(exu_n16186), .Y(exu_n31456));
INVX1 exu_U29549(.A(exu_n31456), .Y(exu_n10307));
AND2X1 exu_U29550(.A(rml_cwp_N99), .B(rml_cwp_next_swap_thr[3]), .Y(rml_cwp_cwp_output_queue_n11));
INVX1 exu_U29551(.A(rml_cwp_cwp_output_queue_n11), .Y(exu_n10308));
AND2X1 exu_U29552(.A(rml_cwp_next_swap_thr[2]), .B(rml_cwp_N99), .Y(rml_cwp_cwp_output_queue_n13));
INVX1 exu_U29553(.A(rml_cwp_cwp_output_queue_n13), .Y(exu_n10309));
AND2X1 exu_U29554(.A(rml_cwp_next_swap_thr[1]), .B(rml_cwp_N99), .Y(rml_cwp_cwp_output_queue_n15));
INVX1 exu_U29555(.A(rml_cwp_cwp_output_queue_n15), .Y(exu_n10310));
AND2X1 exu_U29556(.A(rml_cwp_N99), .B(exu_n15234), .Y(rml_cwp_cwp_output_queue_n17));
INVX1 exu_U29557(.A(rml_cwp_cwp_output_queue_n17), .Y(exu_n10311));
AND2X1 exu_U29558(.A(rml_cwp_cwp_output_queue_n20), .B(exu_n10313), .Y(rml_cwp_cwp_output_queue_n19));
INVX1 exu_U29559(.A(rml_cwp_cwp_output_queue_n19), .Y(exu_n10312));
AND2X1 exu_U29560(.A(rml_cwp_swap_req_vec[0]), .B(exu_n16616), .Y(rml_cwp_cwp_output_queue_n21));
INVX1 exu_U29561(.A(rml_cwp_cwp_output_queue_n21), .Y(exu_n10313));
AND2X1 exu_U29562(.A(exu_n11556), .B(exu_n16626), .Y(rml_cwp_cwp_output_queue_n24));
INVX1 exu_U29563(.A(rml_cwp_cwp_output_queue_n24), .Y(exu_n10314));
AND2X1 exu_U29564(.A(rml_cwp_cwp_output_queue_n30), .B(exu_n10316), .Y(rml_cwp_cwp_output_queue_n29));
INVX1 exu_U29565(.A(rml_cwp_cwp_output_queue_n29), .Y(exu_n10315));
AND2X1 exu_U29566(.A(rml_cwp_swap_req_vec[2]), .B(exu_n16618), .Y(rml_cwp_cwp_output_queue_n31));
INVX1 exu_U29567(.A(rml_cwp_cwp_output_queue_n31), .Y(exu_n10316));
AND2X1 exu_U29568(.A(exu_n15026), .B(rml_cwp_swap_slot0_data[9]), .Y(rml_cwp_slot0_data_mux_n2));
INVX1 exu_U29569(.A(rml_cwp_slot0_data_mux_n2), .Y(exu_n10317));
AND2X1 exu_U29570(.A(rml_cwp_swap_slot0_data[8]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n6));
INVX1 exu_U29571(.A(rml_cwp_slot0_data_mux_n6), .Y(exu_n10318));
AND2X1 exu_U29572(.A(rml_cwp_swap_slot0_data[7]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n10));
INVX1 exu_U29573(.A(rml_cwp_slot0_data_mux_n10), .Y(exu_n10319));
AND2X1 exu_U29574(.A(rml_cwp_swap_slot0_data[6]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n14));
INVX1 exu_U29575(.A(rml_cwp_slot0_data_mux_n14), .Y(exu_n10320));
AND2X1 exu_U29576(.A(rml_cwp_swap_slot0_data[5]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n18));
INVX1 exu_U29577(.A(rml_cwp_slot0_data_mux_n18), .Y(exu_n10321));
AND2X1 exu_U29578(.A(rml_cwp_swap_slot0_data[4]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n22));
INVX1 exu_U29579(.A(rml_cwp_slot0_data_mux_n22), .Y(exu_n10322));
AND2X1 exu_U29580(.A(rml_cwp_swap_slot0_data[3]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n26));
INVX1 exu_U29581(.A(rml_cwp_slot0_data_mux_n26), .Y(exu_n10323));
AND2X1 exu_U29582(.A(rml_cwp_swap_slot0_data[2]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n30));
INVX1 exu_U29583(.A(rml_cwp_slot0_data_mux_n30), .Y(exu_n10324));
AND2X1 exu_U29584(.A(rml_cwp_swap_slot0_data[1]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n34));
INVX1 exu_U29585(.A(rml_cwp_slot0_data_mux_n34), .Y(exu_n10325));
AND2X1 exu_U29586(.A(rml_cwp_swap_slot0_data[12]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n38));
INVX1 exu_U29587(.A(rml_cwp_slot0_data_mux_n38), .Y(exu_n10326));
AND2X1 exu_U29588(.A(rml_cwp_swap_slot0_data[11]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n42));
INVX1 exu_U29589(.A(rml_cwp_slot0_data_mux_n42), .Y(exu_n10327));
AND2X1 exu_U29590(.A(rml_cwp_swap_slot0_data[10]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n46));
INVX1 exu_U29591(.A(rml_cwp_slot0_data_mux_n46), .Y(exu_n10328));
AND2X1 exu_U29592(.A(rml_cwp_swap_slot0_data[0]), .B(exu_n15026), .Y(rml_cwp_slot0_data_mux_n50));
INVX1 exu_U29593(.A(rml_cwp_slot0_data_mux_n50), .Y(exu_n10329));
AND2X1 exu_U29594(.A(ecl_mdqctl_wb_divthr_g[0]), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n3));
INVX1 exu_U29595(.A(ecl_mdqctl_div_data_mux_n3), .Y(exu_n10330));
AND2X1 exu_U29596(.A(ecl_mdqctl_wb_divthr_g[1]), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n5));
INVX1 exu_U29597(.A(ecl_mdqctl_div_data_mux_n5), .Y(exu_n10331));
AND2X1 exu_U29598(.A(ecl_mdqctl_wb_divrd_g[0]), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n7));
INVX1 exu_U29599(.A(ecl_mdqctl_div_data_mux_n7), .Y(exu_n10332));
AND2X1 exu_U29600(.A(ecl_mdqctl_wb_divrd_g[1]), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n9));
INVX1 exu_U29601(.A(ecl_mdqctl_div_data_mux_n9), .Y(exu_n10333));
AND2X1 exu_U29602(.A(ecl_mdqctl_wb_divrd_g[2]), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n11));
INVX1 exu_U29603(.A(ecl_mdqctl_div_data_mux_n11), .Y(exu_n10334));
AND2X1 exu_U29604(.A(ecl_mdqctl_wb_divrd_g[3]), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n13));
INVX1 exu_U29605(.A(ecl_mdqctl_div_data_mux_n13), .Y(exu_n10335));
AND2X1 exu_U29606(.A(ecl_mdqctl_wb_divrd_g[4]), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n15));
INVX1 exu_U29607(.A(ecl_mdqctl_div_data_mux_n15), .Y(exu_n10336));
AND2X1 exu_U29608(.A(ecl_mdqctl_div_data_7), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n17));
INVX1 exu_U29609(.A(ecl_mdqctl_div_data_mux_n17), .Y(exu_n10337));
AND2X1 exu_U29610(.A(ecl_ecl_div_signed_div), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n19));
INVX1 exu_U29611(.A(ecl_mdqctl_div_data_mux_n19), .Y(exu_n10338));
AND2X1 exu_U29612(.A(ecl_div_div64), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n21));
INVX1 exu_U29613(.A(ecl_mdqctl_div_data_mux_n21), .Y(exu_n10339));
AND2X1 exu_U29614(.A(ecl_div_muls), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n23));
INVX1 exu_U29615(.A(ecl_mdqctl_div_data_mux_n23), .Y(exu_n10340));
AND2X1 exu_U29616(.A(exu_n11661), .B(exu_n16387), .Y(ecl_mdqctl_div_data_mux_n25));
INVX1 exu_U29617(.A(ecl_mdqctl_div_data_mux_n25), .Y(exu_n10341));
AND2X1 exu_U29618(.A(ecl_divcntl_inputs_neg_dff_n8), .B(ecl_divcntl_inputs_neg_dff_n6), .Y(ecl_divcntl_inputs_neg_dff_n4));
INVX1 exu_U29619(.A(ecl_divcntl_inputs_neg_dff_n4), .Y(exu_n10342));
AND2X1 exu_U29620(.A(exu_n10775), .B(div_ecl_cout64), .Y(ecl_divcntl_qnext_cout_mux_n3));
INVX1 exu_U29621(.A(ecl_divcntl_qnext_cout_mux_n3), .Y(exu_n10343));
AND2X1 exu_U29622(.A(exu_n16623), .B(ecl_divcntl_div_state_1), .Y(ecl_divcntl_cnt6_n19));
INVX1 exu_U29623(.A(ecl_divcntl_cnt6_n19), .Y(exu_n10344));
AND2X1 exu_U29624(.A(ecl_divcntl_cnt6_n23), .B(exu_n16622), .Y(ecl_divcntl_cnt6_n28));
INVX1 exu_U29625(.A(ecl_divcntl_cnt6_n28), .Y(exu_n10345));
AND2X1 exu_U29626(.A(ecl_ecc_log_rs3_m), .B(exu_n16592), .Y(ecl_eccctl_ecc_synd7_mux_n2));
INVX1 exu_U29627(.A(ecl_eccctl_ecc_synd7_mux_n2), .Y(exu_n10346));
AND2X1 exu_U29628(.A(ecl_eccctl_ecc_rd_mux_n1), .B(exu_n10348), .Y(ecl_eccctl_wb_rd_m[4]));
INVX1 exu_U29629(.A(ecl_eccctl_wb_rd_m[4]), .Y(exu_n10347));
AND2X1 exu_U29630(.A(exu_n15973), .B(ecl_ifu_exu_rs3_m[4]), .Y(ecl_eccctl_ecc_rd_mux_n2));
INVX1 exu_U29631(.A(ecl_eccctl_ecc_rd_mux_n2), .Y(exu_n10348));
AND2X1 exu_U29632(.A(ecl_writeback_restore_rd[0]), .B(exu_n15839), .Y(ecl_writeback_restore_rd_dff_n2));
INVX1 exu_U29633(.A(ecl_writeback_restore_rd_dff_n2), .Y(exu_n10349));
AND2X1 exu_U29634(.A(ecl_writeback_restore_rd[1]), .B(exu_n15839), .Y(ecl_writeback_restore_rd_dff_n8));
INVX1 exu_U29635(.A(ecl_writeback_restore_rd_dff_n8), .Y(exu_n10350));
AND2X1 exu_U29636(.A(ecl_writeback_restore_rd[2]), .B(exu_n15839), .Y(ecl_writeback_restore_rd_dff_n12));
INVX1 exu_U29637(.A(ecl_writeback_restore_rd_dff_n12), .Y(exu_n10351));
AND2X1 exu_U29638(.A(ecl_writeback_restore_rd[3]), .B(exu_n15839), .Y(ecl_writeback_restore_rd_dff_n16));
INVX1 exu_U29639(.A(ecl_writeback_restore_rd_dff_n16), .Y(exu_n10352));
AND2X1 exu_U29640(.A(ecl_writeback_restore_rd[4]), .B(exu_n15839), .Y(ecl_writeback_restore_rd_dff_n20));
INVX1 exu_U29641(.A(ecl_writeback_restore_rd_dff_n20), .Y(exu_n10353));
AND2X1 U29642 ( .A(ecl_writeback_restore_tid_dff_n8 ), .B(ecl_writeback_restore_tid_dff_n6 ), .Y(
        ecl_writeback_restore_tid_dff_n4 ) );
INVX1 exu_U29643(.A(ecl_writeback_restore_tid_dff_n4), .Y(exu_n10354));
AND2X1 U29644 ( .A(ecl_writeback_restore_tid_dff_n13 ), .B(ecl_writeback_restore_tid_dff_n6 ), .Y(
        ecl_writeback_restore_tid_dff_n10 ) );
INVX1 exu_U29645(.A(ecl_writeback_restore_tid_dff_n10), .Y(exu_n10355));
AND2X1 exu_U29646(.A(ecl_mdqctl_wb_mulsetcc_g), .B(exu_n16199), .Y(ecl_writeback_setcc_g_mux_n3));
INVX1 exu_U29647(.A(ecl_writeback_setcc_g_mux_n3), .Y(exu_n10356));
AND2X1 exu_U29648(.A(ecl_ccr_mux_ccrin0_sel2), .B(exu_tlu_ccr0_w[7]), .Y(ecl_ccr_mux_ccrin0_n2));
INVX1 exu_U29649(.A(ecl_ccr_mux_ccrin0_n2), .Y(exu_n10357));
AND2X1 exu_U29650(.A(exu_tlu_ccr0_w[6]), .B(ecl_ccr_mux_ccrin0_sel2), .Y(ecl_ccr_mux_ccrin0_n6));
INVX1 exu_U29651(.A(ecl_ccr_mux_ccrin0_n6), .Y(exu_n10358));
AND2X1 exu_U29652(.A(exu_tlu_ccr0_w[5]), .B(ecl_ccr_mux_ccrin0_sel2), .Y(ecl_ccr_mux_ccrin0_n10));
INVX1 exu_U29653(.A(ecl_ccr_mux_ccrin0_n10), .Y(exu_n10359));
AND2X1 exu_U29654(.A(exu_tlu_ccr0_w[4]), .B(ecl_ccr_mux_ccrin0_sel2), .Y(ecl_ccr_mux_ccrin0_n14));
INVX1 exu_U29655(.A(ecl_ccr_mux_ccrin0_n14), .Y(exu_n10360));
AND2X1 exu_U29656(.A(exu_tlu_ccr0_w[3]), .B(ecl_ccr_mux_ccrin0_sel2), .Y(ecl_ccr_mux_ccrin0_n18));
INVX1 exu_U29657(.A(ecl_ccr_mux_ccrin0_n18), .Y(exu_n10361));
AND2X1 exu_U29658(.A(exu_tlu_ccr0_w[2]), .B(ecl_ccr_mux_ccrin0_sel2), .Y(ecl_ccr_mux_ccrin0_n22));
INVX1 exu_U29659(.A(ecl_ccr_mux_ccrin0_n22), .Y(exu_n10362));
AND2X1 exu_U29660(.A(exu_tlu_ccr0_w[1]), .B(ecl_ccr_mux_ccrin0_sel2), .Y(ecl_ccr_mux_ccrin0_n26));
INVX1 exu_U29661(.A(ecl_ccr_mux_ccrin0_n26), .Y(exu_n10363));
AND2X1 exu_U29662(.A(exu_tlu_ccr0_w[0]), .B(ecl_ccr_mux_ccrin0_sel2), .Y(ecl_ccr_mux_ccrin0_n30));
INVX1 exu_U29663(.A(ecl_ccr_mux_ccrin0_n30), .Y(exu_n10364));
AND2X1 exu_U29664(.A(ecl_ccr_alu_cc_m[0]), .B(exu_n16319), .Y(ecl_ccr_mux_ccr_m_n3));
INVX1 exu_U29665(.A(ecl_ccr_mux_ccr_m_n3), .Y(exu_n10365));
AND2X1 exu_U29666(.A(ecl_ccr_alu_cc_m[1]), .B(exu_n16319), .Y(ecl_ccr_mux_ccr_m_n5));
INVX1 exu_U29667(.A(ecl_ccr_mux_ccr_m_n5), .Y(exu_n10366));
AND2X1 exu_U29668(.A(ecl_ccr_alu_cc_m[2]), .B(exu_n16319), .Y(ecl_ccr_mux_ccr_m_n7));
INVX1 exu_U29669(.A(ecl_ccr_mux_ccr_m_n7), .Y(exu_n10367));
AND2X1 exu_U29670(.A(ecl_ccr_alu_cc_m[3]), .B(exu_n16319), .Y(ecl_ccr_mux_ccr_m_n9));
INVX1 exu_U29671(.A(ecl_ccr_mux_ccr_m_n9), .Y(exu_n10368));
AND2X1 exu_U29672(.A(ecl_ccr_alu_cc_m[4]), .B(exu_n16319), .Y(ecl_ccr_mux_ccr_m_n11));
INVX1 exu_U29673(.A(ecl_ccr_mux_ccr_m_n11), .Y(exu_n10369));
AND2X1 exu_U29674(.A(ecl_ccr_alu_cc_m[5]), .B(exu_n16319), .Y(ecl_ccr_mux_ccr_m_n13));
INVX1 exu_U29675(.A(ecl_ccr_mux_ccr_m_n13), .Y(exu_n10370));
AND2X1 exu_U29676(.A(ecl_ccr_alu_cc_m[6]), .B(exu_n16319), .Y(ecl_ccr_mux_ccr_m_n15));
INVX1 exu_U29677(.A(ecl_ccr_mux_ccr_m_n15), .Y(exu_n10371));
AND2X1 exu_U29678(.A(ecl_ccr_alu_cc_m[7]), .B(exu_n16319), .Y(ecl_ccr_mux_ccr_m_n17));
INVX1 exu_U29679(.A(ecl_ccr_mux_ccr_m_n17), .Y(exu_n10372));
AND2X1 exu_U29680(.A(rml_agp_thr0[0]), .B(rml_agp_wen_thr0_w), .Y(rml_agp_next0_mux_n3));
INVX1 exu_U29681(.A(rml_agp_next0_mux_n3), .Y(exu_n10373));
AND2X1 exu_U29682(.A(rml_agp_thr0[1]), .B(rml_agp_wen_thr0_w), .Y(rml_agp_next0_mux_n5));
INVX1 exu_U29683(.A(rml_agp_next0_mux_n5), .Y(exu_n10374));
AND2X1 exu_U29684(.A(ecl_rml_xor_data_e[0]), .B(exu_n16382), .Y(rml_next_cansave_mux_n3));
INVX1 exu_U29685(.A(rml_next_cansave_mux_n3), .Y(exu_n10375));
AND2X1 exu_U29686(.A(ecl_rml_xor_data_e[1]), .B(exu_n16382), .Y(rml_next_cansave_mux_n5));
INVX1 exu_U29687(.A(rml_next_cansave_mux_n5), .Y(exu_n10376));
AND2X1 exu_U29688(.A(ecl_rml_xor_data_e[2]), .B(exu_n16382), .Y(rml_next_cansave_mux_n7));
INVX1 exu_U29689(.A(rml_next_cansave_mux_n7), .Y(exu_n10377));
OR2X1 exu_U29690(.A(rml_cwp_full_swap_m), .B(exu_n15925), .Y(rml_cwp_n26));
INVX1 exu_U29691(.A(rml_cwp_n26), .Y(exu_n10378));
AND2X1 exu_U29692(.A(rml_cwp_old_swap_cwp[2]), .B(rml_cwp_N99), .Y(rml_cwp_n54));
INVX1 exu_U29693(.A(rml_cwp_n54), .Y(exu_n10379));
AND2X1 exu_U29694(.A(rml_cwp_old_swap_cwp[1]), .B(rml_cwp_N99), .Y(rml_cwp_n56));
INVX1 exu_U29695(.A(rml_cwp_n56), .Y(exu_n10380));
AND2X1 exu_U29696(.A(rml_cwp_old_swap_cwp[0]), .B(rml_cwp_N99), .Y(rml_cwp_n58));
INVX1 exu_U29697(.A(rml_cwp_n58), .Y(exu_n10381));
AND2X1 exu_U29698(.A(rml_cwp_new_swap_cwp[2]), .B(rml_cwp_N99), .Y(rml_cwp_n60));
INVX1 exu_U29699(.A(rml_cwp_n60), .Y(exu_n10382));
AND2X1 exu_U29700(.A(rml_cwp_new_swap_cwp[1]), .B(rml_cwp_N99), .Y(rml_cwp_n62));
INVX1 exu_U29701(.A(rml_cwp_n62), .Y(exu_n10383));
AND2X1 exu_U29702(.A(rml_cwp_new_swap_cwp[0]), .B(rml_cwp_N99), .Y(rml_cwp_n64));
INVX1 exu_U29703(.A(rml_cwp_n64), .Y(exu_n10384));
AND2X1 exu_U29704(.A(exu_n16213), .B(alu_logic_rs1_data_bf1[9]), .Y(div_d_mux_n2));
INVX1 exu_U29705(.A(div_d_mux_n2), .Y(exu_n10385));
INVX1 exu_U29706(.A(exu_n10389), .Y(exu_n10386));
INVX1 exu_U29707(.A(exu_n10386), .Y(exu_n10387));
INVX1 exu_U29708(.A(exu_n10391), .Y(exu_n10388));
INVX1 exu_U29709(.A(exu_n10388), .Y(exu_n10389));
INVX1 exu_U29710(.A(exu_n10484), .Y(exu_n10390));
INVX1 exu_U29711(.A(exu_n10390), .Y(exu_n10391));
AND2X1 exu_U29712(.A(exu_n10941), .B(exu_n16213), .Y(div_d_mux_n26));
INVX1 exu_U29713(.A(div_d_mux_n26), .Y(exu_n10392));
AND2X1 exu_U29714(.A(exu_n10943), .B(exu_n16212), .Y(div_d_mux_n30));
INVX1 exu_U29715(.A(div_d_mux_n30), .Y(exu_n10393));
AND2X1 exu_U29716(.A(exu_n10947), .B(exu_n16212), .Y(div_d_mux_n34));
INVX1 exu_U29717(.A(div_d_mux_n34), .Y(exu_n10394));
AND2X1 exu_U29718(.A(exu_n10949), .B(exu_n16212), .Y(div_d_mux_n38));
INVX1 exu_U29719(.A(div_d_mux_n38), .Y(exu_n10395));
AND2X1 exu_U29720(.A(exu_n10951), .B(exu_n16212), .Y(div_d_mux_n42));
INVX1 exu_U29721(.A(div_d_mux_n42), .Y(exu_n10396));
AND2X1 exu_U29722(.A(alu_logic_rs1_data_bf1[8]), .B(exu_n16212), .Y(div_d_mux_n46));
INVX1 exu_U29723(.A(div_d_mux_n46), .Y(exu_n10397));
AND2X1 exu_U29724(.A(exu_n10953), .B(exu_n16212), .Y(div_d_mux_n50));
INVX1 exu_U29725(.A(div_d_mux_n50), .Y(exu_n10398));
AND2X1 exu_U29726(.A(exu_n10955), .B(exu_n16212), .Y(div_d_mux_n54));
INVX1 exu_U29727(.A(div_d_mux_n54), .Y(exu_n10399));
AND2X1 exu_U29728(.A(exu_n10957), .B(exu_n16212), .Y(div_d_mux_n58));
INVX1 exu_U29729(.A(div_d_mux_n58), .Y(exu_n10400));
AND2X1 exu_U29730(.A(exu_n10959), .B(exu_n16212), .Y(div_d_mux_n62));
INVX1 exu_U29731(.A(div_d_mux_n62), .Y(exu_n10401));
AND2X1 exu_U29732(.A(exu_n10961), .B(exu_n16212), .Y(div_d_mux_n66));
INVX1 exu_U29733(.A(div_d_mux_n66), .Y(exu_n10402));
AND2X1 exu_U29734(.A(exu_n10963), .B(exu_n16212), .Y(div_d_mux_n70));
INVX1 exu_U29735(.A(div_d_mux_n70), .Y(exu_n10403));
AND2X1 exu_U29736(.A(exu_n10965), .B(exu_n16212), .Y(div_d_mux_n74));
INVX1 exu_U29737(.A(div_d_mux_n74), .Y(exu_n10404));
AND2X1 exu_U29738(.A(exu_n10969), .B(exu_n16212), .Y(div_d_mux_n78));
INVX1 exu_U29739(.A(div_d_mux_n78), .Y(exu_n10405));
AND2X1 exu_U29740(.A(exu_n10971), .B(exu_n16212), .Y(div_d_mux_n82));
INVX1 exu_U29741(.A(div_d_mux_n82), .Y(exu_n10406));
AND2X1 exu_U29742(.A(exu_n10973), .B(exu_n16211), .Y(div_d_mux_n86));
INVX1 exu_U29743(.A(div_d_mux_n86), .Y(exu_n10407));
AND2X1 exu_U29744(.A(alu_logic_rs1_data_bf1[7]), .B(exu_n16211), .Y(div_d_mux_n90));
INVX1 exu_U29745(.A(div_d_mux_n90), .Y(exu_n10408));
AND2X1 exu_U29746(.A(exu_n10975), .B(exu_n16211), .Y(div_d_mux_n94));
INVX1 exu_U29747(.A(div_d_mux_n94), .Y(exu_n10409));
AND2X1 exu_U29748(.A(exu_n10977), .B(exu_n16211), .Y(div_d_mux_n98));
INVX1 exu_U29749(.A(div_d_mux_n98), .Y(exu_n10410));
AND2X1 exu_U29750(.A(exu_n10979), .B(exu_n16211), .Y(div_d_mux_n102));
INVX1 exu_U29751(.A(div_d_mux_n102), .Y(exu_n10411));
AND2X1 exu_U29752(.A(exu_n10981), .B(exu_n16211), .Y(div_d_mux_n106));
INVX1 exu_U29753(.A(div_d_mux_n106), .Y(exu_n10412));
AND2X1 exu_U29754(.A(exu_n10983), .B(exu_n16211), .Y(div_d_mux_n110));
INVX1 exu_U29755(.A(div_d_mux_n110), .Y(exu_n10413));
AND2X1 exu_U29756(.A(exu_n10985), .B(exu_n16211), .Y(div_d_mux_n114));
INVX1 exu_U29757(.A(div_d_mux_n114), .Y(exu_n10414));
AND2X1 exu_U29758(.A(exu_n10987), .B(exu_n16211), .Y(div_d_mux_n118));
INVX1 exu_U29759(.A(div_d_mux_n118), .Y(exu_n10415));
AND2X1 exu_U29760(.A(exu_n10927), .B(exu_n16211), .Y(div_d_mux_n122));
INVX1 exu_U29761(.A(div_d_mux_n122), .Y(exu_n10416));
AND2X1 exu_U29762(.A(exu_n10929), .B(exu_n16211), .Y(div_d_mux_n126));
INVX1 exu_U29763(.A(div_d_mux_n126), .Y(exu_n10417));
AND2X1 exu_U29764(.A(exu_n10931), .B(exu_n16211), .Y(div_d_mux_n130));
INVX1 exu_U29765(.A(div_d_mux_n130), .Y(exu_n10418));
AND2X1 exu_U29766(.A(alu_logic_rs1_data_bf1[6]), .B(exu_n16211), .Y(div_d_mux_n134));
INVX1 exu_U29767(.A(div_d_mux_n134), .Y(exu_n10419));
AND2X1 exu_U29768(.A(exu_n10933), .B(exu_n16211), .Y(div_d_mux_n138));
INVX1 exu_U29769(.A(div_d_mux_n138), .Y(exu_n10420));
AND2X1 exu_U29770(.A(exu_n10935), .B(exu_n16210), .Y(div_d_mux_n142));
INVX1 exu_U29771(.A(div_d_mux_n142), .Y(exu_n10421));
AND2X1 exu_U29772(.A(exu_n10937), .B(exu_n16210), .Y(div_d_mux_n146));
INVX1 exu_U29773(.A(div_d_mux_n146), .Y(exu_n10422));
AND2X1 exu_U29774(.A(exu_n10939), .B(exu_n16210), .Y(div_d_mux_n150));
INVX1 exu_U29775(.A(div_d_mux_n150), .Y(exu_n10423));
AND2X1 exu_U29776(.A(exu_n10945), .B(exu_n16210), .Y(div_d_mux_n154));
INVX1 exu_U29777(.A(div_d_mux_n154), .Y(exu_n10424));
AND2X1 exu_U29778(.A(exu_n10967), .B(exu_n16210), .Y(div_d_mux_n158));
INVX1 exu_U29779(.A(div_d_mux_n158), .Y(exu_n10425));
AND2X1 exu_U29780(.A(exu_n10989), .B(exu_n16210), .Y(div_d_mux_n162));
INVX1 exu_U29781(.A(div_d_mux_n162), .Y(exu_n10426));
AND2X1 exu_U29782(.A(exu_n10879), .B(exu_n16210), .Y(div_d_mux_n166));
INVX1 exu_U29783(.A(div_d_mux_n166), .Y(exu_n10427));
AND2X1 exu_U29784(.A(exu_n10883), .B(exu_n16210), .Y(div_d_mux_n170));
INVX1 exu_U29785(.A(div_d_mux_n170), .Y(exu_n10428));
AND2X1 exu_U29786(.A(exu_n10885), .B(exu_n16210), .Y(div_d_mux_n174));
INVX1 exu_U29787(.A(div_d_mux_n174), .Y(exu_n10429));
AND2X1 exu_U29788(.A(alu_logic_rs1_data_bf1[5]), .B(exu_n16210), .Y(div_d_mux_n178));
INVX1 exu_U29789(.A(div_d_mux_n178), .Y(exu_n10430));
AND2X1 exu_U29790(.A(exu_n10887), .B(exu_n16210), .Y(div_d_mux_n182));
INVX1 exu_U29791(.A(div_d_mux_n182), .Y(exu_n10431));
AND2X1 exu_U29792(.A(exu_n10889), .B(exu_n16210), .Y(div_d_mux_n186));
INVX1 exu_U29793(.A(div_d_mux_n186), .Y(exu_n10432));
AND2X1 exu_U29794(.A(exu_n10891), .B(exu_n16210), .Y(div_d_mux_n190));
INVX1 exu_U29795(.A(div_d_mux_n190), .Y(exu_n10433));
AND2X1 exu_U29796(.A(exu_n10893), .B(exu_n16210), .Y(div_d_mux_n194));
INVX1 exu_U29797(.A(div_d_mux_n194), .Y(exu_n10434));
AND2X1 exu_U29798(.A(exu_n10895), .B(exu_n16209), .Y(div_d_mux_n198));
INVX1 exu_U29799(.A(div_d_mux_n198), .Y(exu_n10435));
AND2X1 exu_U29800(.A(exu_n10897), .B(exu_n16209), .Y(div_d_mux_n202));
INVX1 exu_U29801(.A(div_d_mux_n202), .Y(exu_n10436));
AND2X1 exu_U29802(.A(exu_n10899), .B(exu_n16209), .Y(div_d_mux_n206));
INVX1 exu_U29803(.A(div_d_mux_n206), .Y(exu_n10437));
AND2X1 exu_U29804(.A(exu_n10901), .B(exu_n16209), .Y(div_d_mux_n210));
INVX1 exu_U29805(.A(div_d_mux_n210), .Y(exu_n10438));
AND2X1 exu_U29806(.A(exu_n10905), .B(exu_n16209), .Y(div_d_mux_n214));
INVX1 exu_U29807(.A(div_d_mux_n214), .Y(exu_n10439));
AND2X1 exu_U29808(.A(exu_n10907), .B(exu_n16209), .Y(div_d_mux_n218));
INVX1 exu_U29809(.A(div_d_mux_n218), .Y(exu_n10440));
AND2X1 exu_U29810(.A(alu_logic_rs1_data_bf1[4]), .B(exu_n16209), .Y(div_d_mux_n222));
INVX1 exu_U29811(.A(div_d_mux_n222), .Y(exu_n10441));
AND2X1 exu_U29812(.A(exu_n10909), .B(exu_n16209), .Y(div_d_mux_n226));
INVX1 exu_U29813(.A(div_d_mux_n226), .Y(exu_n10442));
AND2X1 exu_U29814(.A(exu_n10911), .B(exu_n16209), .Y(div_d_mux_n230));
INVX1 exu_U29815(.A(div_d_mux_n230), .Y(exu_n10443));
AND2X1 exu_U29816(.A(exu_n10913), .B(exu_n16209), .Y(div_d_mux_n234));
INVX1 exu_U29817(.A(div_d_mux_n234), .Y(exu_n10444));
AND2X1 exu_U29818(.A(exu_n10915), .B(exu_n16209), .Y(div_d_mux_n238));
INVX1 exu_U29819(.A(div_d_mux_n238), .Y(exu_n10445));
AND2X1 exu_U29820(.A(exu_n10917), .B(exu_n16209), .Y(div_d_mux_n242));
INVX1 exu_U29821(.A(div_d_mux_n242), .Y(exu_n10446));
AND2X1 exu_U29822(.A(exu_n10919), .B(exu_n16209), .Y(div_d_mux_n246));
INVX1 exu_U29823(.A(div_d_mux_n246), .Y(exu_n10447));
AND2X1 exu_U29824(.A(exu_n10921), .B(exu_n16209), .Y(div_d_mux_n250));
INVX1 exu_U29825(.A(div_d_mux_n250), .Y(exu_n10448));
AND2X1 exu_U29826(.A(exu_n10923), .B(exu_n16203), .Y(div_d_mux_n254));
INVX1 exu_U29827(.A(div_d_mux_n254), .Y(exu_n10449));
AND2X1 exu_U29828(.A(exu_n10865), .B(exu_n16203), .Y(div_d_mux_n258));
INVX1 exu_U29829(.A(div_d_mux_n258), .Y(exu_n10450));
AND2X1 exu_U29830(.A(exu_n10867), .B(exu_n16203), .Y(div_d_mux_n262));
INVX1 exu_U29831(.A(div_d_mux_n262), .Y(exu_n10451));
AND2X1 exu_U29832(.A(alu_logic_rs1_data_bf1[3]), .B(exu_n16203), .Y(div_d_mux_n266));
INVX1 exu_U29833(.A(div_d_mux_n266), .Y(exu_n10452));
AND2X1 exu_U29834(.A(exu_n10869), .B(exu_n16204), .Y(div_d_mux_n270));
INVX1 exu_U29835(.A(div_d_mux_n270), .Y(exu_n10453));
AND2X1 exu_U29836(.A(exu_n10871), .B(exu_n16207), .Y(div_d_mux_n274));
INVX1 exu_U29837(.A(div_d_mux_n274), .Y(exu_n10454));
AND2X1 exu_U29838(.A(exu_n10873), .B(ecl_div_ld_inputs), .Y(div_d_mux_n278));
INVX1 exu_U29839(.A(div_d_mux_n278), .Y(exu_n10455));
AND2X1 exu_U29840(.A(exu_n10875), .B(exu_n16204), .Y(div_d_mux_n282));
INVX1 exu_U29841(.A(div_d_mux_n282), .Y(exu_n10456));
AND2X1 exu_U29842(.A(exu_n10877), .B(exu_n16203), .Y(div_d_mux_n286));
INVX1 exu_U29843(.A(div_d_mux_n286), .Y(exu_n10457));
AND2X1 exu_U29844(.A(exu_n10881), .B(exu_n16213), .Y(div_d_mux_n290));
INVX1 exu_U29845(.A(div_d_mux_n290), .Y(exu_n10458));
AND2X1 exu_U29846(.A(exu_n10903), .B(exu_n16204), .Y(div_d_mux_n294));
INVX1 exu_U29847(.A(div_d_mux_n294), .Y(exu_n10459));
AND2X1 exu_U29848(.A(exu_n10925), .B(exu_n16207), .Y(div_d_mux_n298));
INVX1 exu_U29849(.A(div_d_mux_n298), .Y(exu_n10460));
AND2X1 exu_U29850(.A(alu_logic_rs1_data_bf1[31]), .B(ecl_div_ld_inputs), .Y(div_d_mux_n302));
INVX1 exu_U29851(.A(div_d_mux_n302), .Y(exu_n10461));
AND2X1 exu_U29852(.A(alu_logic_rs1_data_bf1[30]), .B(exu_n16208), .Y(div_d_mux_n306));
INVX1 exu_U29853(.A(div_d_mux_n306), .Y(exu_n10462));
AND2X1 exu_U29854(.A(alu_logic_rs1_data_bf1[2]), .B(exu_n16208), .Y(div_d_mux_n310));
INVX1 exu_U29855(.A(div_d_mux_n310), .Y(exu_n10463));
AND2X1 exu_U29856(.A(alu_logic_rs1_data_bf1[29]), .B(exu_n16208), .Y(div_d_mux_n314));
INVX1 exu_U29857(.A(div_d_mux_n314), .Y(exu_n10464));
AND2X1 exu_U29858(.A(alu_logic_rs1_data_bf1[28]), .B(exu_n16208), .Y(div_d_mux_n318));
INVX1 exu_U29859(.A(div_d_mux_n318), .Y(exu_n10465));
AND2X1 exu_U29860(.A(alu_logic_rs1_data_bf1[27]), .B(exu_n16208), .Y(div_d_mux_n322));
INVX1 exu_U29861(.A(div_d_mux_n322), .Y(exu_n10466));
AND2X1 exu_U29862(.A(alu_logic_rs1_data_bf1[26]), .B(exu_n16208), .Y(div_d_mux_n326));
INVX1 exu_U29863(.A(div_d_mux_n326), .Y(exu_n10467));
AND2X1 exu_U29864(.A(alu_logic_rs1_data_bf1[25]), .B(exu_n16208), .Y(div_d_mux_n330));
INVX1 exu_U29865(.A(div_d_mux_n330), .Y(exu_n10468));
AND2X1 exu_U29866(.A(alu_logic_rs1_data_bf1[24]), .B(exu_n16208), .Y(div_d_mux_n334));
INVX1 exu_U29867(.A(div_d_mux_n334), .Y(exu_n10469));
AND2X1 exu_U29868(.A(alu_logic_rs1_data_bf1[23]), .B(exu_n16208), .Y(div_d_mux_n338));
INVX1 exu_U29869(.A(div_d_mux_n338), .Y(exu_n10470));
AND2X1 exu_U29870(.A(alu_logic_rs1_data_bf1[22]), .B(exu_n16208), .Y(div_d_mux_n342));
INVX1 exu_U29871(.A(div_d_mux_n342), .Y(exu_n10471));
AND2X1 exu_U29872(.A(alu_logic_rs1_data_bf1[21]), .B(exu_n16208), .Y(div_d_mux_n346));
INVX1 exu_U29873(.A(div_d_mux_n346), .Y(exu_n10472));
AND2X1 exu_U29874(.A(alu_logic_rs1_data_bf1[20]), .B(exu_n16208), .Y(div_d_mux_n350));
INVX1 exu_U29875(.A(div_d_mux_n350), .Y(exu_n10473));
AND2X1 exu_U29876(.A(alu_logic_rs1_data_bf1[1]), .B(exu_n16208), .Y(div_d_mux_n354));
INVX1 exu_U29877(.A(div_d_mux_n354), .Y(exu_n10474));
AND2X1 exu_U29878(.A(alu_logic_rs1_data_bf1[19]), .B(exu_n16208), .Y(div_d_mux_n358));
INVX1 exu_U29879(.A(div_d_mux_n358), .Y(exu_n10475));
AND2X1 exu_U29880(.A(alu_logic_rs1_data_bf1[18]), .B(exu_n16207), .Y(div_d_mux_n362));
INVX1 exu_U29881(.A(div_d_mux_n362), .Y(exu_n10476));
AND2X1 exu_U29882(.A(alu_logic_rs1_data_bf1[17]), .B(exu_n16207), .Y(div_d_mux_n366));
INVX1 exu_U29883(.A(div_d_mux_n366), .Y(exu_n10477));
AND2X1 exu_U29884(.A(alu_logic_rs1_data_bf1[16]), .B(exu_n16207), .Y(div_d_mux_n370));
INVX1 exu_U29885(.A(div_d_mux_n370), .Y(exu_n10478));
AND2X1 exu_U29886(.A(alu_logic_rs1_data_bf1[15]), .B(exu_n16207), .Y(div_d_mux_n374));
INVX1 exu_U29887(.A(div_d_mux_n374), .Y(exu_n10479));
AND2X1 exu_U29888(.A(alu_logic_rs1_data_bf1[14]), .B(exu_n16207), .Y(div_d_mux_n378));
INVX1 exu_U29889(.A(div_d_mux_n378), .Y(exu_n10480));
AND2X1 exu_U29890(.A(alu_logic_rs1_data_bf1[13]), .B(exu_n16207), .Y(div_d_mux_n382));
INVX1 exu_U29891(.A(div_d_mux_n382), .Y(exu_n10481));
AND2X1 exu_U29892(.A(alu_logic_rs1_data_bf1[12]), .B(exu_n16207), .Y(div_d_mux_n386));
INVX1 exu_U29893(.A(div_d_mux_n386), .Y(exu_n10482));
INVX1 exu_U29894(.A(exu_n10486), .Y(exu_n10483));
INVX1 exu_U29895(.A(exu_n10483), .Y(exu_n10484));
INVX1 exu_U29896(.A(exu_n10488), .Y(exu_n10485));
INVX1 exu_U29897(.A(exu_n10485), .Y(exu_n10486));
INVX1 exu_U29898(.A(exu_n10490), .Y(exu_n10487));
INVX1 exu_U29899(.A(exu_n10487), .Y(exu_n10488));
INVX1 exu_U29900(.A(exu_n10492), .Y(exu_n10489));
INVX1 exu_U29901(.A(exu_n10489), .Y(exu_n10490));
INVX1 exu_U29902(.A(exu_n10494), .Y(exu_n10491));
INVX1 exu_U29903(.A(exu_n10491), .Y(exu_n10492));
INVX1 exu_U29904(.A(exu_n10496), .Y(exu_n10493));
INVX1 exu_U29905(.A(exu_n10493), .Y(exu_n10494));
INVX1 exu_U29906(.A(exu_n10498), .Y(exu_n10495));
INVX1 exu_U29907(.A(exu_n10495), .Y(exu_n10496));
INVX1 exu_U29908(.A(exu_n10501), .Y(exu_n10497));
INVX1 exu_U29909(.A(exu_n10497), .Y(exu_n10498));
AND2X1 exu_U29910(.A(alu_logic_rs1_data_bf1[11]), .B(exu_n16213), .Y(div_d_mux_n422));
INVX1 exu_U29911(.A(div_d_mux_n422), .Y(exu_n10499));
INVX1 exu_U29912(.A(exu_n10503), .Y(exu_n10500));
INVX1 exu_U29913(.A(exu_n10500), .Y(exu_n10501));
INVX1 exu_U29914(.A(exu_n10505), .Y(exu_n10502));
INVX1 exu_U29915(.A(exu_n10502), .Y(exu_n10503));
INVX1 exu_U29916(.A(exu_n10507), .Y(exu_n10504));
INVX1 exu_U29917(.A(exu_n10504), .Y(exu_n10505));
INVX1 exu_U29918(.A(exu_n10509), .Y(exu_n10506));
INVX1 exu_U29919(.A(exu_n10506), .Y(exu_n10507));
INVX1 exu_U29920(.A(exu_n10511), .Y(exu_n10508));
INVX1 exu_U29921(.A(exu_n10508), .Y(exu_n10509));
INVX1 exu_U29922(.A(exu_n10513), .Y(exu_n10510));
INVX1 exu_U29923(.A(exu_n10510), .Y(exu_n10511));
INVX1 exu_U29924(.A(exu_n10515), .Y(exu_n10512));
INVX1 exu_U29925(.A(exu_n10512), .Y(exu_n10513));
INVX1 exu_U29926(.A(exu_n10778), .Y(exu_n10514));
INVX1 exu_U29927(.A(exu_n10514), .Y(exu_n10515));
AND2X1 exu_U29928(.A(alu_logic_rs1_data_bf1[10]), .B(exu_n16213), .Y(div_d_mux_n466));
INVX1 exu_U29929(.A(div_d_mux_n466), .Y(exu_n10516));
AND2X1 exu_U29930(.A(alu_logic_rs1_data_bf1[0]), .B(exu_n16203), .Y(div_d_mux_n510));
INVX1 exu_U29931(.A(div_d_mux_n510), .Y(exu_n10517));
AND2X1 exu_U29932(.A(ecl_mdqctl_divcntl_muldone), .B(exu_n10519), .Y(ecl_mdqctl_n14));
INVX1 exu_U29933(.A(ecl_mdqctl_n14), .Y(exu_n10518));
AND2X1 exu_U29934(.A(exu_n15398), .B(exu_n16199), .Y(ecl_mdqctl_n15));
INVX1 exu_U29935(.A(ecl_mdqctl_n15), .Y(exu_n10519));
AND2X1 exu_U29936(.A(ifu_exu_muldivop_d[4]), .B(ifu_exu_muldivop_d[2]), .Y(ecl_mdqctl_n27));
INVX1 exu_U29937(.A(ecl_mdqctl_n27), .Y(exu_n10520));
AND2X1 exu_U29938(.A(ifu_exu_muldivop_d[1]), .B(ifu_exu_muldivop_d[4]), .Y(ecl_mdqctl_n29));
INVX1 exu_U29939(.A(ecl_mdqctl_n29), .Y(exu_n10521));
AND2X1 exu_U29940(.A(ifu_exu_muldivop_d[0]), .B(ifu_exu_muldivop_d[4]), .Y(ecl_mdqctl_n31));
INVX1 exu_U29941(.A(ecl_mdqctl_n31), .Y(exu_n10522));
AND2X1 exu_U29942(.A(ecl_mdqctl_wb_mulrd_g[4]), .B(exu_n16388), .Y(ecl_mdqctl_n33));
INVX1 exu_U29943(.A(ecl_mdqctl_n33), .Y(exu_n10523));
AND2X1 exu_U29944(.A(ecl_mdqctl_wb_mulrd_g[3]), .B(exu_n16388), .Y(ecl_mdqctl_n35));
INVX1 exu_U29945(.A(ecl_mdqctl_n35), .Y(exu_n10524));
AND2X1 exu_U29946(.A(ecl_mdqctl_wb_mulrd_g[2]), .B(exu_n16388), .Y(ecl_mdqctl_n37));
INVX1 exu_U29947(.A(ecl_mdqctl_n37), .Y(exu_n10525));
AND2X1 exu_U29948(.A(ecl_mdqctl_wb_mulrd_g[1]), .B(exu_n16388), .Y(ecl_mdqctl_n39));
INVX1 exu_U29949(.A(ecl_mdqctl_n39), .Y(exu_n10526));
AND2X1 exu_U29950(.A(ecl_mdqctl_wb_mulrd_g[0]), .B(exu_n16388), .Y(ecl_mdqctl_n41));
INVX1 exu_U29951(.A(ecl_mdqctl_n41), .Y(exu_n10527));
AND2X1 exu_U29952(.A(ecl_mdqctl_wb_multhr_g[1]), .B(exu_n16388), .Y(ecl_mdqctl_n43));
INVX1 exu_U29953(.A(ecl_mdqctl_n43), .Y(exu_n10528));
AND2X1 exu_U29954(.A(ecl_mdqctl_wb_multhr_g[0]), .B(exu_n16388), .Y(ecl_mdqctl_n45));
INVX1 exu_U29955(.A(ecl_mdqctl_n45), .Y(exu_n10529));
AND2X1 exu_U29956(.A(ecl_div_muls), .B(ecl_divcntl_div_state_1), .Y(ecl_divcntl_n28));
INVX1 exu_U29957(.A(ecl_divcntl_n28), .Y(exu_n10530));
AND2X1 exu_U29958(.A(ecl_divcntl_div_state[4]), .B(exu_n10532), .Y(ecl_divcntl_n39));
INVX1 exu_U29959(.A(ecl_divcntl_n39), .Y(exu_n10531));
AND2X1 exu_U29960(.A(exu_n11665), .B(exu_n10533), .Y(ecl_divcntl_n40));
INVX1 exu_U29961(.A(ecl_divcntl_n40), .Y(exu_n10532));
AND2X1 exu_U29962(.A(ecl_divcntl_n43), .B(ecl_divcntl_rs2_data_31_w), .Y(ecl_divcntl_n42));
INVX1 exu_U29963(.A(ecl_divcntl_n42), .Y(exu_n10533));
AND2X1 exu_U29964(.A(exu_n15558), .B(ecl_divcntl_div_state_1), .Y(ecl_divcntl_n46));
INVX1 exu_U29965(.A(ecl_divcntl_n46), .Y(exu_n10534));
AND2X1 exu_U29966(.A(ecl_byplog_rs2_n18), .B(ecl_byplog_rs2_n19), .Y(ecl_byplog_rs2_n17));
INVX1 exu_U29967(.A(ecl_byplog_rs2_n17), .Y(exu_n10535));
AND2X1 exu_U29968(.A(ecl_byplog_rs2_n32), .B(exu_n15435), .Y(ecl_byplog_rs2_n36));
INVX1 exu_U29969(.A(ecl_byplog_rs2_n36), .Y(exu_n10536));
AND2X1 exu_U29970(.A(ecl_wb_byplog_wen_w2), .B(ecl_byplog_rs2_match_w2), .Y(ecl_byplog_rs2_n40));
INVX1 exu_U29971(.A(ecl_byplog_rs2_n40), .Y(exu_n10537));
OR2X1 exu_U29972(.A(ecl_ifu_exu_rs2_d[2]), .B(ecl_byplog_rs2_n51), .Y(ecl_byplog_rs2_n50));
INVX1 exu_U29973(.A(ecl_byplog_rs2_n50), .Y(exu_n10538));
AND2X1 exu_U29974(.A(ecl_wb_byplog_wen_w2), .B(ecl_byplog_rs1_match_w2), .Y(ecl_byplog_rs1_n44));
INVX1 exu_U29975(.A(ecl_byplog_rs1_n44), .Y(exu_n10539));
OR2X1 exu_U29976(.A(ecc_ecl_rs2_ue), .B(ecc_ecl_rs1_ue), .Y(ecl_eccctl_n19));
INVX1 exu_U29977(.A(ecl_eccctl_n19), .Y(exu_n10540));
AND2X1 exu_U29978(.A(ecl_eccctl_cwp_m[1]), .B(ecl_eccctl_n25), .Y(ecl_eccctl_n24));
INVX1 exu_U29979(.A(ecl_eccctl_n24), .Y(exu_n10541));
AND2X1 exu_U29980(.A(ecl_eccctl_cwp_m[0]), .B(ecl_eccctl_n25), .Y(ecl_eccctl_n27));
INVX1 exu_U29981(.A(ecl_eccctl_n27), .Y(exu_n10542));
AND2X1 exu_U29982(.A(exu_n11673), .B(ecl_eccctl_rs2_ce_m), .Y(ecl_eccctl_n32));
INVX1 exu_U29983(.A(ecl_eccctl_n32), .Y(exu_n10543));
AND2X1 exu_U29984(.A(exu_n11674), .B(ecl_writeback_n19), .Y(ecl_writeback_n46));
INVX1 exu_U29985(.A(ecl_writeback_n46), .Y(exu_n10544));
AND2X1 exu_U29986(.A(ifu_tlu_sraddr_d[2]), .B(exu_n16375), .Y(ecl_writeback_n90));
INVX1 exu_U29987(.A(ecl_writeback_n90), .Y(exu_n10545));
OR2X1 exu_U29988(.A(rml_ecl_swap_done[3]), .B(exu_n14964), .Y(ecl_writeback_n93));
INVX1 exu_U29989(.A(ecl_writeback_n93), .Y(exu_n10546));
OR2X1 exu_U29990(.A(rml_ecl_swap_done[2]), .B(exu_n14966), .Y(ecl_writeback_n104));
INVX1 exu_U29991(.A(ecl_writeback_n104), .Y(exu_n10547));
OR2X1 exu_U29992(.A(rml_ecl_swap_done[1]), .B(exu_n14968), .Y(ecl_writeback_n112));
INVX1 exu_U29993(.A(ecl_writeback_n112), .Y(exu_n10548));
OR2X1 exu_U29994(.A(rml_ecl_swap_done[0]), .B(exu_n14970), .Y(ecl_writeback_n119));
INVX1 exu_U29995(.A(ecl_writeback_n119), .Y(exu_n10549));
AND2X1 exu_U29996(.A(ecl_writeback_inst_vld_noflush_wen_w), .B(ifu_exu_inst_vld_w), .Y(ecl_writeback_n147));
INVX1 exu_U29997(.A(ecl_writeback_n147), .Y(exu_n10550));
AND2X1 exu_U29998(.A(exu_n11681), .B(ecl_writeback_n19), .Y(ecl_writeback_n151));
INVX1 exu_U29999(.A(ecl_writeback_n151), .Y(exu_n10551));
AND2X1 exu_U30000(.A(exu_n11684), .B(exu_n15765), .Y(ecl_writeback_n165));
INVX1 exu_U30001(.A(ecl_writeback_n165), .Y(exu_n10552));
AND2X1 exu_U30002(.A(exu_n11687), .B(exu_n15765), .Y(ecl_writeback_n171));
INVX1 exu_U30003(.A(ecl_writeback_n171), .Y(exu_n10553));
AND2X1 exu_U30004(.A(exu_n15477), .B(exu_n16600), .Y(ecl_writeback_n197));
INVX1 exu_U30005(.A(ecl_writeback_n197), .Y(exu_n10554));
AND2X1 exu_U30006(.A(exu_n19227), .B(lsu_exu_ldxa_data_g[9]), .Y(bypass_rs3h_w2_mux_n2));
INVX1 exu_U30007(.A(bypass_rs3h_w2_mux_n2), .Y(exu_n10555));
AND2X1 exu_U30008(.A(lsu_exu_ldxa_data_g[8]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n6));
INVX1 exu_U30009(.A(bypass_rs3h_w2_mux_n6), .Y(exu_n10556));
AND2X1 exu_U30010(.A(lsu_exu_ldxa_data_g[7]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n10));
INVX1 exu_U30011(.A(bypass_rs3h_w2_mux_n10), .Y(exu_n10557));
AND2X1 exu_U30012(.A(lsu_exu_ldxa_data_g[6]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n14));
INVX1 exu_U30013(.A(bypass_rs3h_w2_mux_n14), .Y(exu_n10558));
AND2X1 exu_U30014(.A(lsu_exu_ldxa_data_g[5]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n18));
INVX1 exu_U30015(.A(bypass_rs3h_w2_mux_n18), .Y(exu_n10559));
AND2X1 exu_U30016(.A(lsu_exu_ldxa_data_g[4]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n22));
INVX1 exu_U30017(.A(bypass_rs3h_w2_mux_n22), .Y(exu_n10560));
AND2X1 exu_U30018(.A(lsu_exu_ldxa_data_g[3]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n26));
INVX1 exu_U30019(.A(bypass_rs3h_w2_mux_n26), .Y(exu_n10561));
AND2X1 exu_U30020(.A(lsu_exu_ldxa_data_g[31]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n30));
INVX1 exu_U30021(.A(bypass_rs3h_w2_mux_n30), .Y(exu_n10562));
AND2X1 exu_U30022(.A(lsu_exu_ldxa_data_g[30]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n34));
INVX1 exu_U30023(.A(bypass_rs3h_w2_mux_n34), .Y(exu_n10563));
AND2X1 exu_U30024(.A(lsu_exu_ldxa_data_g[2]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n38));
INVX1 exu_U30025(.A(bypass_rs3h_w2_mux_n38), .Y(exu_n10564));
AND2X1 exu_U30026(.A(lsu_exu_ldxa_data_g[29]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n42));
INVX1 exu_U30027(.A(bypass_rs3h_w2_mux_n42), .Y(exu_n10565));
AND2X1 exu_U30028(.A(lsu_exu_ldxa_data_g[28]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n46));
INVX1 exu_U30029(.A(bypass_rs3h_w2_mux_n46), .Y(exu_n10566));
AND2X1 exu_U30030(.A(lsu_exu_ldxa_data_g[27]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n50));
INVX1 exu_U30031(.A(bypass_rs3h_w2_mux_n50), .Y(exu_n10567));
AND2X1 exu_U30032(.A(lsu_exu_ldxa_data_g[26]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n54));
INVX1 exu_U30033(.A(bypass_rs3h_w2_mux_n54), .Y(exu_n10568));
AND2X1 exu_U30034(.A(lsu_exu_ldxa_data_g[25]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n58));
INVX1 exu_U30035(.A(bypass_rs3h_w2_mux_n58), .Y(exu_n10569));
AND2X1 exu_U30036(.A(lsu_exu_ldxa_data_g[24]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n62));
INVX1 exu_U30037(.A(bypass_rs3h_w2_mux_n62), .Y(exu_n10570));
AND2X1 exu_U30038(.A(lsu_exu_ldxa_data_g[23]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n66));
INVX1 exu_U30039(.A(bypass_rs3h_w2_mux_n66), .Y(exu_n10571));
AND2X1 exu_U30040(.A(lsu_exu_ldxa_data_g[22]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n70));
INVX1 exu_U30041(.A(bypass_rs3h_w2_mux_n70), .Y(exu_n10572));
AND2X1 exu_U30042(.A(lsu_exu_ldxa_data_g[21]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n74));
INVX1 exu_U30043(.A(bypass_rs3h_w2_mux_n74), .Y(exu_n10573));
AND2X1 exu_U30044(.A(lsu_exu_ldxa_data_g[20]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n78));
INVX1 exu_U30045(.A(bypass_rs3h_w2_mux_n78), .Y(exu_n10574));
AND2X1 exu_U30046(.A(lsu_exu_ldxa_data_g[1]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n82));
INVX1 exu_U30047(.A(bypass_rs3h_w2_mux_n82), .Y(exu_n10575));
AND2X1 exu_U30048(.A(lsu_exu_ldxa_data_g[19]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n86));
INVX1 exu_U30049(.A(bypass_rs3h_w2_mux_n86), .Y(exu_n10576));
AND2X1 exu_U30050(.A(lsu_exu_ldxa_data_g[18]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n90));
INVX1 exu_U30051(.A(bypass_rs3h_w2_mux_n90), .Y(exu_n10577));
AND2X1 exu_U30052(.A(lsu_exu_ldxa_data_g[17]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n94));
INVX1 exu_U30053(.A(bypass_rs3h_w2_mux_n94), .Y(exu_n10578));
AND2X1 exu_U30054(.A(lsu_exu_ldxa_data_g[16]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n98));
INVX1 exu_U30055(.A(bypass_rs3h_w2_mux_n98), .Y(exu_n10579));
AND2X1 exu_U30056(.A(lsu_exu_ldxa_data_g[15]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n102));
INVX1 exu_U30057(.A(bypass_rs3h_w2_mux_n102), .Y(exu_n10580));
AND2X1 exu_U30058(.A(lsu_exu_ldxa_data_g[14]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n106));
INVX1 exu_U30059(.A(bypass_rs3h_w2_mux_n106), .Y(exu_n10581));
AND2X1 exu_U30060(.A(lsu_exu_ldxa_data_g[13]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n110));
INVX1 exu_U30061(.A(bypass_rs3h_w2_mux_n110), .Y(exu_n10582));
AND2X1 exu_U30062(.A(lsu_exu_ldxa_data_g[12]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n114));
INVX1 exu_U30063(.A(bypass_rs3h_w2_mux_n114), .Y(exu_n10583));
AND2X1 exu_U30064(.A(lsu_exu_ldxa_data_g[11]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n118));
INVX1 exu_U30065(.A(bypass_rs3h_w2_mux_n118), .Y(exu_n10584));
AND2X1 exu_U30066(.A(lsu_exu_ldxa_data_g[10]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n122));
INVX1 exu_U30067(.A(bypass_rs3h_w2_mux_n122), .Y(exu_n10585));
AND2X1 exu_U30068(.A(lsu_exu_ldxa_data_g[0]), .B(exu_n19227), .Y(bypass_rs3h_w2_mux_n126));
INVX1 exu_U30069(.A(bypass_rs3h_w2_mux_n126), .Y(exu_n10586));
AND2X1 exu_U30070(.A(bypass_sr_out_mux_n1), .B(exu_n10588), .Y(bypass_full_rd_data_m[9]));
INVX1 exu_U30071(.A(bypass_full_rd_data_m[9]), .Y(exu_n10587));
AND2X1 exu_U30072(.A(exu_n16263), .B(tlu_exu_rsr_data_m[9]), .Y(bypass_sr_out_mux_n2));
INVX1 exu_U30073(.A(bypass_sr_out_mux_n2), .Y(exu_n10588));
AND2X1 exu_U30074(.A(ifu_exu_pcver_e[63]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n28));
INVX1 exu_U30075(.A(bypass_ifu_exu_sr_mux_n28), .Y(exu_n10589));
AND2X1 exu_U30076(.A(ifu_exu_pcver_e[62]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n34));
INVX1 exu_U30077(.A(bypass_ifu_exu_sr_mux_n34), .Y(exu_n10590));
AND2X1 exu_U30078(.A(ifu_exu_pcver_e[61]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n40));
INVX1 exu_U30079(.A(bypass_ifu_exu_sr_mux_n40), .Y(exu_n10591));
AND2X1 exu_U30080(.A(ifu_exu_pcver_e[60]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n46));
INVX1 exu_U30081(.A(bypass_ifu_exu_sr_mux_n46), .Y(exu_n10592));
AND2X1 exu_U30082(.A(ifu_exu_pcver_e[59]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n58));
INVX1 exu_U30083(.A(bypass_ifu_exu_sr_mux_n58), .Y(exu_n10593));
AND2X1 exu_U30084(.A(ifu_exu_pcver_e[58]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n64));
INVX1 exu_U30085(.A(bypass_ifu_exu_sr_mux_n64), .Y(exu_n10594));
AND2X1 exu_U30086(.A(ifu_exu_pcver_e[57]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n70));
INVX1 exu_U30087(.A(bypass_ifu_exu_sr_mux_n70), .Y(exu_n10595));
AND2X1 exu_U30088(.A(ifu_exu_pcver_e[56]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n76));
INVX1 exu_U30089(.A(bypass_ifu_exu_sr_mux_n76), .Y(exu_n10596));
AND2X1 exu_U30090(.A(ifu_exu_pcver_e[55]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n82));
INVX1 exu_U30091(.A(bypass_ifu_exu_sr_mux_n82), .Y(exu_n10597));
AND2X1 exu_U30092(.A(ifu_exu_pcver_e[54]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n88));
INVX1 exu_U30093(.A(bypass_ifu_exu_sr_mux_n88), .Y(exu_n10598));
AND2X1 exu_U30094(.A(ifu_exu_pcver_e[53]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n94));
INVX1 exu_U30095(.A(bypass_ifu_exu_sr_mux_n94), .Y(exu_n10599));
AND2X1 exu_U30096(.A(ifu_exu_pcver_e[52]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n100));
INVX1 exu_U30097(.A(bypass_ifu_exu_sr_mux_n100), .Y(exu_n10600));
AND2X1 exu_U30098(.A(ifu_exu_pcver_e[51]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n106));
INVX1 exu_U30099(.A(bypass_ifu_exu_sr_mux_n106), .Y(exu_n10601));
AND2X1 exu_U30100(.A(ifu_exu_pcver_e[50]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n112));
INVX1 exu_U30101(.A(bypass_ifu_exu_sr_mux_n112), .Y(exu_n10602));
AND2X1 exu_U30102(.A(ifu_exu_pcver_e[49]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n124));
INVX1 exu_U30103(.A(bypass_ifu_exu_sr_mux_n124), .Y(exu_n10603));
AND2X1 exu_U30104(.A(ifu_exu_pcver_e[48]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n130));
INVX1 exu_U30105(.A(bypass_ifu_exu_sr_mux_n130), .Y(exu_n10604));
AND2X1 exu_U30106(.A(ifu_exu_pcver_e[47]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n136));
INVX1 exu_U30107(.A(bypass_ifu_exu_sr_mux_n136), .Y(exu_n10605));
AND2X1 exu_U30108(.A(ifu_exu_pcver_e[46]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n142));
INVX1 exu_U30109(.A(bypass_ifu_exu_sr_mux_n142), .Y(exu_n10606));
AND2X1 exu_U30110(.A(ifu_exu_pcver_e[45]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n148));
INVX1 exu_U30111(.A(bypass_ifu_exu_sr_mux_n148), .Y(exu_n10607));
AND2X1 exu_U30112(.A(ifu_exu_pcver_e[44]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n154));
INVX1 exu_U30113(.A(bypass_ifu_exu_sr_mux_n154), .Y(exu_n10608));
AND2X1 exu_U30114(.A(ifu_exu_pcver_e[43]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n160));
INVX1 exu_U30115(.A(bypass_ifu_exu_sr_mux_n160), .Y(exu_n10609));
AND2X1 exu_U30116(.A(ifu_exu_pcver_e[42]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n166));
INVX1 exu_U30117(.A(bypass_ifu_exu_sr_mux_n166), .Y(exu_n10610));
AND2X1 exu_U30118(.A(ifu_exu_pcver_e[41]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n172));
INVX1 exu_U30119(.A(bypass_ifu_exu_sr_mux_n172), .Y(exu_n10611));
AND2X1 exu_U30120(.A(ifu_exu_pcver_e[40]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n178));
INVX1 exu_U30121(.A(bypass_ifu_exu_sr_mux_n178), .Y(exu_n10612));
AND2X1 exu_U30122(.A(ifu_exu_pcver_e[39]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n190));
INVX1 exu_U30123(.A(bypass_ifu_exu_sr_mux_n190), .Y(exu_n10613));
AND2X1 exu_U30124(.A(ifu_exu_pcver_e[38]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n196));
INVX1 exu_U30125(.A(bypass_ifu_exu_sr_mux_n196), .Y(exu_n10614));
AND2X1 exu_U30126(.A(ifu_exu_pcver_e[37]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n202));
INVX1 exu_U30127(.A(bypass_ifu_exu_sr_mux_n202), .Y(exu_n10615));
AND2X1 exu_U30128(.A(ifu_exu_pcver_e[36]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n208));
INVX1 exu_U30129(.A(bypass_ifu_exu_sr_mux_n208), .Y(exu_n10616));
AND2X1 exu_U30130(.A(ifu_exu_pcver_e[35]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n214));
INVX1 exu_U30131(.A(bypass_ifu_exu_sr_mux_n214), .Y(exu_n10617));
AND2X1 exu_U30132(.A(ifu_exu_pcver_e[34]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n220));
INVX1 exu_U30133(.A(bypass_ifu_exu_sr_mux_n220), .Y(exu_n10618));
AND2X1 exu_U30134(.A(ifu_exu_pcver_e[33]), .B(exu_n16266), .Y(bypass_ifu_exu_sr_mux_n226));
INVX1 exu_U30135(.A(bypass_ifu_exu_sr_mux_n226), .Y(exu_n10619));
AND2X1 exu_U30136(.A(ifu_exu_pcver_e[32]), .B(ecl_byp_sel_ifusr_e), .Y(bypass_ifu_exu_sr_mux_n232));
INVX1 exu_U30137(.A(bypass_ifu_exu_sr_mux_n232), .Y(exu_n10620));
AND2X1 exu_U30138(.A(lsu_exu_dfill_data_g[9]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n3));
INVX1 exu_U30139(.A(bypass_dfill_data_mux_n3), .Y(exu_n10621));
AND2X1 exu_U30140(.A(lsu_exu_dfill_data_g[8]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n5));
INVX1 exu_U30141(.A(bypass_dfill_data_mux_n5), .Y(exu_n10622));
AND2X1 exu_U30142(.A(lsu_exu_dfill_data_g[7]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n7));
INVX1 exu_U30143(.A(bypass_dfill_data_mux_n7), .Y(exu_n10623));
AND2X1 exu_U30144(.A(lsu_exu_dfill_data_g[6]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n9));
INVX1 exu_U30145(.A(bypass_dfill_data_mux_n9), .Y(exu_n10624));
AND2X1 exu_U30146(.A(lsu_exu_dfill_data_g[63]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n11));
INVX1 exu_U30147(.A(bypass_dfill_data_mux_n11), .Y(exu_n10625));
AND2X1 exu_U30148(.A(lsu_exu_dfill_data_g[62]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n13));
INVX1 exu_U30149(.A(bypass_dfill_data_mux_n13), .Y(exu_n10626));
AND2X1 exu_U30150(.A(lsu_exu_dfill_data_g[61]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n15));
INVX1 exu_U30151(.A(bypass_dfill_data_mux_n15), .Y(exu_n10627));
AND2X1 exu_U30152(.A(lsu_exu_dfill_data_g[60]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n17));
INVX1 exu_U30153(.A(bypass_dfill_data_mux_n17), .Y(exu_n10628));
AND2X1 exu_U30154(.A(lsu_exu_dfill_data_g[5]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n19));
INVX1 exu_U30155(.A(bypass_dfill_data_mux_n19), .Y(exu_n10629));
AND2X1 exu_U30156(.A(lsu_exu_dfill_data_g[59]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n21));
INVX1 exu_U30157(.A(bypass_dfill_data_mux_n21), .Y(exu_n10630));
AND2X1 exu_U30158(.A(lsu_exu_dfill_data_g[58]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n23));
INVX1 exu_U30159(.A(bypass_dfill_data_mux_n23), .Y(exu_n10631));
AND2X1 exu_U30160(.A(lsu_exu_dfill_data_g[57]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n25));
INVX1 exu_U30161(.A(bypass_dfill_data_mux_n25), .Y(exu_n10632));
AND2X1 exu_U30162(.A(lsu_exu_dfill_data_g[56]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n27));
INVX1 exu_U30163(.A(bypass_dfill_data_mux_n27), .Y(exu_n10633));
AND2X1 exu_U30164(.A(lsu_exu_dfill_data_g[55]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n29));
INVX1 exu_U30165(.A(bypass_dfill_data_mux_n29), .Y(exu_n10634));
AND2X1 exu_U30166(.A(lsu_exu_dfill_data_g[54]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n31));
INVX1 exu_U30167(.A(bypass_dfill_data_mux_n31), .Y(exu_n10635));
AND2X1 exu_U30168(.A(lsu_exu_dfill_data_g[53]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n33));
INVX1 exu_U30169(.A(bypass_dfill_data_mux_n33), .Y(exu_n10636));
AND2X1 exu_U30170(.A(lsu_exu_dfill_data_g[52]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n35));
INVX1 exu_U30171(.A(bypass_dfill_data_mux_n35), .Y(exu_n10637));
AND2X1 exu_U30172(.A(lsu_exu_dfill_data_g[51]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n37));
INVX1 exu_U30173(.A(bypass_dfill_data_mux_n37), .Y(exu_n10638));
AND2X1 exu_U30174(.A(lsu_exu_dfill_data_g[50]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n39));
INVX1 exu_U30175(.A(bypass_dfill_data_mux_n39), .Y(exu_n10639));
AND2X1 exu_U30176(.A(lsu_exu_dfill_data_g[4]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n41));
INVX1 exu_U30177(.A(bypass_dfill_data_mux_n41), .Y(exu_n10640));
AND2X1 exu_U30178(.A(lsu_exu_dfill_data_g[49]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n43));
INVX1 exu_U30179(.A(bypass_dfill_data_mux_n43), .Y(exu_n10641));
AND2X1 exu_U30180(.A(lsu_exu_dfill_data_g[48]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n45));
INVX1 exu_U30181(.A(bypass_dfill_data_mux_n45), .Y(exu_n10642));
AND2X1 exu_U30182(.A(lsu_exu_dfill_data_g[47]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n47));
INVX1 exu_U30183(.A(bypass_dfill_data_mux_n47), .Y(exu_n10643));
AND2X1 exu_U30184(.A(lsu_exu_dfill_data_g[46]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n49));
INVX1 exu_U30185(.A(bypass_dfill_data_mux_n49), .Y(exu_n10644));
AND2X1 exu_U30186(.A(lsu_exu_dfill_data_g[45]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n51));
INVX1 exu_U30187(.A(bypass_dfill_data_mux_n51), .Y(exu_n10645));
AND2X1 exu_U30188(.A(lsu_exu_dfill_data_g[44]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n53));
INVX1 exu_U30189(.A(bypass_dfill_data_mux_n53), .Y(exu_n10646));
AND2X1 exu_U30190(.A(lsu_exu_dfill_data_g[43]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n55));
INVX1 exu_U30191(.A(bypass_dfill_data_mux_n55), .Y(exu_n10647));
AND2X1 exu_U30192(.A(lsu_exu_dfill_data_g[42]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n57));
INVX1 exu_U30193(.A(bypass_dfill_data_mux_n57), .Y(exu_n10648));
AND2X1 exu_U30194(.A(lsu_exu_dfill_data_g[41]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n59));
INVX1 exu_U30195(.A(bypass_dfill_data_mux_n59), .Y(exu_n10649));
AND2X1 exu_U30196(.A(lsu_exu_dfill_data_g[40]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n61));
INVX1 exu_U30197(.A(bypass_dfill_data_mux_n61), .Y(exu_n10650));
AND2X1 exu_U30198(.A(lsu_exu_dfill_data_g[3]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n63));
INVX1 exu_U30199(.A(bypass_dfill_data_mux_n63), .Y(exu_n10651));
AND2X1 exu_U30200(.A(lsu_exu_dfill_data_g[39]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n65));
INVX1 exu_U30201(.A(bypass_dfill_data_mux_n65), .Y(exu_n10652));
AND2X1 exu_U30202(.A(lsu_exu_dfill_data_g[38]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n67));
INVX1 exu_U30203(.A(bypass_dfill_data_mux_n67), .Y(exu_n10653));
AND2X1 exu_U30204(.A(lsu_exu_dfill_data_g[37]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n69));
INVX1 exu_U30205(.A(bypass_dfill_data_mux_n69), .Y(exu_n10654));
AND2X1 exu_U30206(.A(lsu_exu_dfill_data_g[36]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n71));
INVX1 exu_U30207(.A(bypass_dfill_data_mux_n71), .Y(exu_n10655));
AND2X1 exu_U30208(.A(lsu_exu_dfill_data_g[35]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n73));
INVX1 exu_U30209(.A(bypass_dfill_data_mux_n73), .Y(exu_n10656));
AND2X1 exu_U30210(.A(lsu_exu_dfill_data_g[34]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n75));
INVX1 exu_U30211(.A(bypass_dfill_data_mux_n75), .Y(exu_n10657));
AND2X1 exu_U30212(.A(lsu_exu_dfill_data_g[33]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n77));
INVX1 exu_U30213(.A(bypass_dfill_data_mux_n77), .Y(exu_n10658));
AND2X1 exu_U30214(.A(lsu_exu_dfill_data_g[32]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n79));
INVX1 exu_U30215(.A(bypass_dfill_data_mux_n79), .Y(exu_n10659));
AND2X1 exu_U30216(.A(lsu_exu_dfill_data_g[31]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n81));
INVX1 exu_U30217(.A(bypass_dfill_data_mux_n81), .Y(exu_n10660));
AND2X1 exu_U30218(.A(lsu_exu_dfill_data_g[30]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n83));
INVX1 exu_U30219(.A(bypass_dfill_data_mux_n83), .Y(exu_n10661));
AND2X1 exu_U30220(.A(lsu_exu_dfill_data_g[2]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n85));
INVX1 exu_U30221(.A(bypass_dfill_data_mux_n85), .Y(exu_n10662));
AND2X1 exu_U30222(.A(lsu_exu_dfill_data_g[29]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n87));
INVX1 exu_U30223(.A(bypass_dfill_data_mux_n87), .Y(exu_n10663));
AND2X1 exu_U30224(.A(lsu_exu_dfill_data_g[28]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n89));
INVX1 exu_U30225(.A(bypass_dfill_data_mux_n89), .Y(exu_n10664));
AND2X1 exu_U30226(.A(lsu_exu_dfill_data_g[27]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n91));
INVX1 exu_U30227(.A(bypass_dfill_data_mux_n91), .Y(exu_n10665));
AND2X1 exu_U30228(.A(lsu_exu_dfill_data_g[26]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n93));
INVX1 exu_U30229(.A(bypass_dfill_data_mux_n93), .Y(exu_n10666));
AND2X1 exu_U30230(.A(lsu_exu_dfill_data_g[25]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n95));
INVX1 exu_U30231(.A(bypass_dfill_data_mux_n95), .Y(exu_n10667));
AND2X1 exu_U30232(.A(lsu_exu_dfill_data_g[24]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n97));
INVX1 exu_U30233(.A(bypass_dfill_data_mux_n97), .Y(exu_n10668));
AND2X1 exu_U30234(.A(lsu_exu_dfill_data_g[23]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n99));
INVX1 exu_U30235(.A(bypass_dfill_data_mux_n99), .Y(exu_n10669));
AND2X1 exu_U30236(.A(lsu_exu_dfill_data_g[22]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n101));
INVX1 exu_U30237(.A(bypass_dfill_data_mux_n101), .Y(exu_n10670));
AND2X1 exu_U30238(.A(lsu_exu_dfill_data_g[21]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n103));
INVX1 exu_U30239(.A(bypass_dfill_data_mux_n103), .Y(exu_n10671));
AND2X1 exu_U30240(.A(lsu_exu_dfill_data_g[20]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n105));
INVX1 exu_U30241(.A(bypass_dfill_data_mux_n105), .Y(exu_n10672));
AND2X1 exu_U30242(.A(lsu_exu_dfill_data_g[1]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n107));
INVX1 exu_U30243(.A(bypass_dfill_data_mux_n107), .Y(exu_n10673));
AND2X1 exu_U30244(.A(lsu_exu_dfill_data_g[19]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n109));
INVX1 exu_U30245(.A(bypass_dfill_data_mux_n109), .Y(exu_n10674));
AND2X1 exu_U30246(.A(lsu_exu_dfill_data_g[18]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n111));
INVX1 exu_U30247(.A(bypass_dfill_data_mux_n111), .Y(exu_n10675));
AND2X1 exu_U30248(.A(lsu_exu_dfill_data_g[17]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n113));
INVX1 exu_U30249(.A(bypass_dfill_data_mux_n113), .Y(exu_n10676));
AND2X1 exu_U30250(.A(lsu_exu_dfill_data_g[16]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n115));
INVX1 exu_U30251(.A(bypass_dfill_data_mux_n115), .Y(exu_n10677));
AND2X1 exu_U30252(.A(lsu_exu_dfill_data_g[15]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n117));
INVX1 exu_U30253(.A(bypass_dfill_data_mux_n117), .Y(exu_n10678));
AND2X1 exu_U30254(.A(lsu_exu_dfill_data_g[14]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n119));
INVX1 exu_U30255(.A(bypass_dfill_data_mux_n119), .Y(exu_n10679));
AND2X1 exu_U30256(.A(lsu_exu_dfill_data_g[13]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n121));
INVX1 exu_U30257(.A(bypass_dfill_data_mux_n121), .Y(exu_n10680));
AND2X1 exu_U30258(.A(lsu_exu_dfill_data_g[12]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n123));
INVX1 exu_U30259(.A(bypass_dfill_data_mux_n123), .Y(exu_n10681));
AND2X1 exu_U30260(.A(lsu_exu_dfill_data_g[11]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n125));
INVX1 exu_U30261(.A(bypass_dfill_data_mux_n125), .Y(exu_n10682));
AND2X1 exu_U30262(.A(lsu_exu_dfill_data_g[10]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n127));
INVX1 exu_U30263(.A(bypass_dfill_data_mux_n127), .Y(exu_n10683));
AND2X1 exu_U30264(.A(lsu_exu_dfill_data_g[0]), .B(exu_n16270), .Y(bypass_dfill_data_mux_n129));
INVX1 exu_U30265(.A(bypass_dfill_data_mux_n129), .Y(exu_n10684));
AND2X1 exu_U30266(.A(rml_n48), .B(exu_n15856), .Y(rml_n47));
INVX1 exu_U30267(.A(rml_n47), .Y(exu_n10685));
AND2X1 exu_U30268(.A(exu_n15857), .B(rml_n48), .Y(rml_n54));
INVX1 exu_U30269(.A(rml_n54), .Y(exu_n10686));
AND2X1 exu_U30270(.A(rml_oddwin_w[3]), .B(exu_n10688), .Y(rml_n82));
INVX1 exu_U30271(.A(rml_n82), .Y(exu_n10687));
AND2X1 exu_U30272(.A(rml_rml_cwp_wen_m), .B(exu_n15921), .Y(rml_n83));
INVX1 exu_U30273(.A(rml_n83), .Y(exu_n10688));
AND2X1 exu_U30274(.A(rml_oddwin_w[2]), .B(exu_n10690), .Y(rml_n86));
INVX1 exu_U30275(.A(rml_n86), .Y(exu_n10689));
AND2X1 exu_U30276(.A(exu_n15922), .B(rml_rml_cwp_wen_m), .Y(rml_n87));
INVX1 exu_U30277(.A(rml_n87), .Y(exu_n10690));
AND2X1 exu_U30278(.A(rml_oddwin_w[1]), .B(exu_n10692), .Y(rml_n89));
INVX1 exu_U30279(.A(rml_n89), .Y(exu_n10691));
AND2X1 exu_U30280(.A(exu_n15923), .B(rml_rml_cwp_wen_m), .Y(rml_n90));
INVX1 exu_U30281(.A(rml_n90), .Y(exu_n10692));
AND2X1 exu_U30282(.A(rml_oddwin_w[0]), .B(exu_n10694), .Y(rml_n92));
INVX1 exu_U30283(.A(rml_n92), .Y(exu_n10693));
AND2X1 exu_U30284(.A(exu_n15924), .B(rml_rml_cwp_wen_m), .Y(rml_n93));
INVX1 exu_U30285(.A(rml_n93), .Y(exu_n10694));
AND2X1 exu_U30286(.A(ecl_divcntl_n70), .B(exu_n16413), .Y(div_u32[9]));
INVX1 exu_U30287(.A(div_u32[9]), .Y(exu_n10695));
AND2X1 exu_U30288(.A(exu_n16246), .B(exu_n16413), .Y(div_pos32[9]));
INVX1 exu_U30289(.A(div_pos32[9]), .Y(exu_n10696));
AND2X1 exu_U30290(.A(ecl_perr_store[3]), .B(exu_n10698), .Y(ecl_n50));
INVX1 exu_U30291(.A(ecl_n50), .Y(exu_n10697));
AND2X1 exu_U30292(.A(ecl_rml_thr_w[3]), .B(exu_n15817), .Y(ecl_n51));
INVX1 exu_U30293(.A(ecl_n51), .Y(exu_n10698));
AND2X1 exu_U30294(.A(ecl_perr_store[2]), .B(exu_n10700), .Y(ecl_n53));
INVX1 exu_U30295(.A(ecl_n53), .Y(exu_n10699));
AND2X1 exu_U30296(.A(ecl_rml_thr_w[2]), .B(exu_n15817), .Y(ecl_n54));
INVX1 exu_U30297(.A(ecl_n54), .Y(exu_n10700));
AND2X1 exu_U30298(.A(ecl_perr_store[1]), .B(exu_n10702), .Y(ecl_n56));
INVX1 exu_U30299(.A(ecl_n56), .Y(exu_n10701));
AND2X1 exu_U30300(.A(exu_n15958), .B(exu_n15817), .Y(ecl_n57));
INVX1 exu_U30301(.A(ecl_n57), .Y(exu_n10702));
AND2X1 exu_U30302(.A(ecl_perr_store[0]), .B(exu_n10704), .Y(ecl_n59));
INVX1 exu_U30303(.A(ecl_n59), .Y(exu_n10703));
AND2X1 exu_U30304(.A(exu_n15960), .B(exu_n15817), .Y(ecl_n60));
INVX1 exu_U30305(.A(ecl_n60), .Y(exu_n10704));
AND2X1 exu_U30306(.A(ecl_muls_e), .B(alu_logic_rs1_data_bf1[0]), .Y(ecl_n64));
INVX1 exu_U30307(.A(ecl_n64), .Y(exu_n10705));
AND2X1 exu_U30308(.A(ifu_exu_inst_vld_w), .B(exu_n10707), .Y(ecl_n95));
INVX1 exu_U30309(.A(ecl_n95), .Y(exu_n10706));
AND2X1 exu_U30310(.A(exu_n16318), .B(exu_n10708), .Y(ecl_n96));
INVX1 exu_U30311(.A(ecl_n96), .Y(exu_n10707));
AND2X1 exu_U30312(.A(ecl_n98), .B(tlu_exu_pic_twobelow_m), .Y(ecl_n97));
INVX1 exu_U30313(.A(ecl_n97), .Y(exu_n10708));
AND2X1 exu_U30314(.A(exu_n11935), .B(alu_ecl_adderin2_63_e), .Y(ecl_n132));
INVX1 exu_U30315(.A(ecl_n132), .Y(exu_n10709));
AND2X1 exu_U30316(.A(ecl_ifu_exu_tagop_e), .B(exu_n10711), .Y(ecl_n138));
INVX1 exu_U30317(.A(ecl_n138), .Y(exu_n10710));
AND2X1 exu_U30318(.A(exu_n11938), .B(exu_n16224), .Y(ecl_n139));
INVX1 exu_U30319(.A(ecl_n139), .Y(exu_n10711));
AND2X1 exu_U30320(.A(ecl_ifu_exu_rs1_d[1]), .B(exu_n16627), .Y(exu_n16629));
INVX1 exu_U30321(.A(exu_n16629), .Y(exu_n10712));
AND2X1 exu_U30322(.A(exu_n15222), .B(exu_n16399), .Y(exu_n16632));
INVX1 exu_U30323(.A(exu_n16632), .Y(exu_n10713));
AND2X1 exu_U30324(.A(ecl_ifu_exu_rs1_d[1]), .B(exu_n16641), .Y(exu_n16643));
INVX1 exu_U30325(.A(exu_n16643), .Y(exu_n10714));
AND2X1 exu_U30326(.A(exu_n15223), .B(exu_n16399), .Y(exu_n16646));
INVX1 exu_U30327(.A(exu_n16646), .Y(exu_n10715));
AND2X1 exu_U30328(.A(ecl_ifu_exu_rs1_d[1]), .B(exu_n16655), .Y(exu_n16657));
INVX1 exu_U30329(.A(exu_n16657), .Y(exu_n10716));
AND2X1 exu_U30330(.A(exu_n15224), .B(exu_n16399), .Y(exu_n16660));
INVX1 exu_U30331(.A(exu_n16660), .Y(exu_n10717));
AND2X1 exu_U30332(.A(ecl_ifu_exu_rs1_d[1]), .B(exu_n16669), .Y(exu_n16671));
INVX1 exu_U30333(.A(exu_n16671), .Y(exu_n10718));
AND2X1 exu_U30334(.A(exu_n15225), .B(exu_n16399), .Y(exu_n16674));
INVX1 exu_U30335(.A(exu_n16674), .Y(exu_n10719));
AND2X1 exu_U30336(.A(ecl_ifu_exu_rs2_d[1]), .B(exu_n16683), .Y(exu_n16685));
INVX1 exu_U30337(.A(exu_n16685), .Y(exu_n10720));
AND2X1 exu_U30338(.A(exu_n15226), .B(exu_n16568), .Y(exu_n16688));
INVX1 exu_U30339(.A(exu_n16688), .Y(exu_n10721));
AND2X1 exu_U30340(.A(ecl_ifu_exu_rs2_d[1]), .B(exu_n16697), .Y(exu_n16699));
INVX1 exu_U30341(.A(exu_n16699), .Y(exu_n10722));
AND2X1 exu_U30342(.A(exu_n15227), .B(exu_n16568), .Y(exu_n16702));
INVX1 exu_U30343(.A(exu_n16702), .Y(exu_n10723));
AND2X1 exu_U30344(.A(ecl_ifu_exu_rs2_d[1]), .B(exu_n16711), .Y(exu_n16713));
INVX1 exu_U30345(.A(exu_n16713), .Y(exu_n10724));
AND2X1 exu_U30346(.A(exu_n15228), .B(exu_n16568), .Y(exu_n16716));
INVX1 exu_U30347(.A(exu_n16716), .Y(exu_n10725));
AND2X1 exu_U30348(.A(ecl_ifu_exu_rs2_d[1]), .B(exu_n16725), .Y(exu_n16727));
INVX1 exu_U30349(.A(exu_n16727), .Y(exu_n10726));
AND2X1 exu_U30350(.A(exu_n15229), .B(exu_n16568), .Y(exu_n16730));
INVX1 exu_U30351(.A(exu_n16730), .Y(exu_n10727));
AND2X1 exu_U30352(.A(ecl_ifu_exu_rs3_d[1]), .B(exu_n17403), .Y(exu_n17405));
INVX1 exu_U30353(.A(exu_n17405), .Y(exu_n10728));
AND2X1 exu_U30354(.A(exu_n15230), .B(exu_n16567), .Y(exu_n17408));
INVX1 exu_U30355(.A(exu_n17408), .Y(exu_n10729));
AND2X1 exu_U30356(.A(ecl_ifu_exu_rs3_d[1]), .B(exu_n17417), .Y(exu_n17419));
INVX1 exu_U30357(.A(exu_n17419), .Y(exu_n10730));
AND2X1 exu_U30358(.A(exu_n15231), .B(exu_n16567), .Y(exu_n17422));
INVX1 exu_U30359(.A(exu_n17422), .Y(exu_n10731));
AND2X1 exu_U30360(.A(ecl_ifu_exu_rs3_d[1]), .B(exu_n17431), .Y(exu_n17433));
INVX1 exu_U30361(.A(exu_n17433), .Y(exu_n10732));
AND2X1 exu_U30362(.A(exu_n15232), .B(exu_n16567), .Y(exu_n17436));
INVX1 exu_U30363(.A(exu_n17436), .Y(exu_n10733));
AND2X1 exu_U30364(.A(ecl_ifu_exu_rs3_d[1]), .B(exu_n17445), .Y(exu_n17447));
INVX1 exu_U30365(.A(exu_n17447), .Y(exu_n10734));
AND2X1 exu_U30366(.A(exu_n15233), .B(exu_n16567), .Y(exu_n17450));
INVX1 exu_U30367(.A(exu_n17450), .Y(exu_n10735));
AND2X1 exu_U30368(.A(rml_cwp_n37), .B(rml_ecl_wtype_e[0]), .Y(exu_n17507));
INVX1 exu_U30369(.A(exu_n17507), .Y(exu_n10736));
AND2X1 exu_U30370(.A(rml_ecl_other_e), .B(rml_cwp_n37), .Y(exu_n17509));
INVX1 exu_U30371(.A(exu_n17509), .Y(exu_n10737));
AND2X1 exu_U30372(.A(exu_n15940), .B(rml_cwp_n37), .Y(exu_n17512));
INVX1 exu_U30373(.A(exu_n17512), .Y(exu_n10738));
AND2X1 exu_U30374(.A(rml_cwp_tlu_swap_data[12]), .B(rml_cwp_n34), .Y(exu_n17534));
INVX1 exu_U30375(.A(exu_n17534), .Y(exu_n10739));
AND2X1 exu_U30376(.A(rml_ecl_wtype_e[2]), .B(rml_cwp_n37), .Y(exu_n17536));
INVX1 exu_U30377(.A(exu_n17536), .Y(exu_n10740));
AND2X1 exu_U30378(.A(rml_ecl_wtype_e[1]), .B(rml_cwp_n37), .Y(exu_n17538));
INVX1 exu_U30379(.A(exu_n17538), .Y(exu_n10741));
AND2X1 exu_U30380(.A(rml_cwp_n36), .B(rml_ecl_wtype_e[0]), .Y(exu_n17544));
INVX1 exu_U30381(.A(exu_n17544), .Y(exu_n10742));
AND2X1 exu_U30382(.A(rml_ecl_other_e), .B(rml_cwp_n36), .Y(exu_n17546));
INVX1 exu_U30383(.A(exu_n17546), .Y(exu_n10743));
AND2X1 exu_U30384(.A(exu_n15940), .B(rml_cwp_n36), .Y(exu_n17549));
INVX1 exu_U30385(.A(exu_n17549), .Y(exu_n10744));
AND2X1 exu_U30386(.A(rml_cwp_tlu_swap_data[12]), .B(rml_cwp_n33), .Y(exu_n17571));
INVX1 exu_U30387(.A(exu_n17571), .Y(exu_n10745));
AND2X1 exu_U30388(.A(rml_ecl_wtype_e[2]), .B(rml_cwp_n36), .Y(exu_n17573));
INVX1 exu_U30389(.A(exu_n17573), .Y(exu_n10746));
AND2X1 exu_U30390(.A(rml_ecl_wtype_e[1]), .B(rml_cwp_n36), .Y(exu_n17575));
INVX1 exu_U30391(.A(exu_n17575), .Y(exu_n10747));
AND2X1 exu_U30392(.A(rml_cwp_n35), .B(rml_ecl_wtype_e[0]), .Y(exu_n17581));
INVX1 exu_U30393(.A(exu_n17581), .Y(exu_n10748));
AND2X1 exu_U30394(.A(rml_ecl_other_e), .B(rml_cwp_n35), .Y(exu_n17583));
INVX1 exu_U30395(.A(exu_n17583), .Y(exu_n10749));
AND2X1 exu_U30396(.A(exu_n15940), .B(rml_cwp_n35), .Y(exu_n17586));
INVX1 exu_U30397(.A(exu_n17586), .Y(exu_n10750));
AND2X1 exu_U30398(.A(rml_cwp_tlu_swap_data[12]), .B(rml_cwp_n32), .Y(exu_n17608));
INVX1 exu_U30399(.A(exu_n17608), .Y(exu_n10751));
AND2X1 exu_U30400(.A(rml_ecl_wtype_e[2]), .B(rml_cwp_n35), .Y(exu_n17610));
INVX1 exu_U30401(.A(exu_n17610), .Y(exu_n10752));
AND2X1 exu_U30402(.A(rml_ecl_wtype_e[1]), .B(rml_cwp_n35), .Y(exu_n17612));
INVX1 exu_U30403(.A(exu_n17612), .Y(exu_n10753));
INVX1 exu_U30404(.A(exu_n17617), .Y(exu_n10754));
AND2X1 exu_U30405(.A(exu_n15701), .B(ecl_ccr_wen_thr1_w), .Y(exu_n18046));
INVX1 exu_U30406(.A(exu_n18046), .Y(exu_n10755));
AND2X1 exu_U30407(.A(exu_n15700), .B(ecl_ccr_wen_thr1_w), .Y(exu_n18048));
INVX1 exu_U30408(.A(exu_n18048), .Y(exu_n10756));
AND2X1 exu_U30409(.A(exu_n15701), .B(ecl_ccr_wen_thr2_w), .Y(exu_n18074));
INVX1 exu_U30410(.A(exu_n18074), .Y(exu_n10757));
AND2X1 exu_U30411(.A(exu_n15700), .B(ecl_ccr_wen_thr2_w), .Y(exu_n18076));
INVX1 exu_U30412(.A(exu_n18076), .Y(exu_n10758));
AND2X1 exu_U30413(.A(exu_n15701), .B(ecl_ccr_wen_thr3_w), .Y(exu_n18102));
INVX1 exu_U30414(.A(exu_n18102), .Y(exu_n10759));
AND2X1 exu_U30415(.A(exu_n15700), .B(ecl_ccr_wen_thr3_w), .Y(exu_n18104));
INVX1 exu_U30416(.A(exu_n18104), .Y(exu_n10760));
INVX1 exu_U30417(.A(ecl_ccr_partial_cc_d[7]), .Y(exu_n10761));
INVX1 exu_U30418(.A(ecl_ccr_partial_cc_d[6]), .Y(exu_n10762));
INVX1 exu_U30419(.A(ecl_ccr_partial_cc_d[5]), .Y(exu_n10763));
INVX1 exu_U30420(.A(ecl_ccr_partial_cc_d[4]), .Y(exu_n10764));
INVX1 exu_U30421(.A(ecl_ccr_partial_cc_d[3]), .Y(exu_n10765));
INVX1 exu_U30422(.A(ecl_ccr_partial_cc_d[2]), .Y(exu_n10766));
INVX1 exu_U30423(.A(ecl_ccr_partial_cc_d[1]), .Y(exu_n10767));
INVX1 exu_U30424(.A(ecl_ccr_partial_cc_d[0]), .Y(exu_n10768));
AND2X1 exu_U30425(.A(rml_new_agp[0]), .B(exu_n15485), .Y(exu_n18169));
INVX1 exu_U30426(.A(exu_n18169), .Y(exu_n10769));
AND2X1 exu_U30427(.A(rml_new_agp[1]), .B(exu_n15485), .Y(exu_n18171));
INVX1 exu_U30428(.A(exu_n18171), .Y(exu_n10770));
AND2X1 exu_U30429(.A(rml_new_agp[0]), .B(exu_n15484), .Y(exu_n18173));
INVX1 exu_U30430(.A(exu_n18173), .Y(exu_n10771));
AND2X1 exu_U30431(.A(rml_new_agp[1]), .B(exu_n15484), .Y(exu_n18175));
INVX1 exu_U30432(.A(exu_n18175), .Y(exu_n10772));
AND2X1 exu_U30433(.A(rml_new_agp[0]), .B(exu_n15483), .Y(exu_n18177));
INVX1 exu_U30434(.A(exu_n18177), .Y(exu_n10773));
AND2X1 exu_U30435(.A(rml_new_agp[1]), .B(exu_n15483), .Y(exu_n18179));
INVX1 exu_U30436(.A(exu_n18179), .Y(exu_n10774));
INVX1 exu_U30437(.A(ecl_divcntl_q_next_nocout[1]), .Y(exu_n10775));
INVX1 exu_U30438(.A(exu_n10778), .Y(exu_n10776));
INVX1 exu_U30439(.A(exu_n10776), .Y(exu_n10777));
AND2X1 exu_U30440(.A(exu_n16260), .B(exu_n16214), .Y(exu_n18182));
INVX1 exu_U30441(.A(exu_n18182), .Y(exu_n10778));
INVX1 exu_U30442(.A(ecl_divcntl_sub_next_nocout[1]), .Y(exu_n10779));
AND2X1 exu_U30443(.A(ecl_divcntl_subnext_mux_in1[0]), .B(ecl_divcntl_N56), .Y(exu_n18184));
INVX1 exu_U30444(.A(exu_n18184), .Y(exu_n10780));
AND2X1 exu_U30445(.A(exu_n16437), .B(ecl_divcntl_N56), .Y(exu_n18186));
INVX1 exu_U30446(.A(exu_n18186), .Y(exu_n10781));
AND2X1 exu_U30447(.A(rml_cwp_swap_tid[0]), .B(rml_cwp_N99), .Y(exu_n18187));
INVX1 exu_U30448(.A(exu_n18187), .Y(exu_n10782));
AND2X1 exu_U30449(.A(rml_cwp_swap_tid[1]), .B(rml_cwp_N99), .Y(exu_n18189));
INVX1 exu_U30450(.A(exu_n18189), .Y(exu_n10783));
AND2X1 exu_U30451(.A(rml_next_canrestore_w[2]), .B(exu_n18191), .Y(exu_n18212));
INVX1 exu_U30452(.A(exu_n18212), .Y(exu_n10784));
AND2X1 exu_U30453(.A(rml_next_canrestore_w[1]), .B(exu_n18191), .Y(exu_n18214));
INVX1 exu_U30454(.A(exu_n18214), .Y(exu_n10785));
AND2X1 exu_U30455(.A(rml_next_canrestore_w[0]), .B(exu_n18191), .Y(exu_n18216));
INVX1 exu_U30456(.A(exu_n18216), .Y(exu_n10786));
AND2X1 exu_U30457(.A(rml_next_canrestore_w[2]), .B(exu_n18192), .Y(exu_n18218));
INVX1 exu_U30458(.A(exu_n18218), .Y(exu_n10787));
AND2X1 exu_U30459(.A(rml_next_canrestore_w[1]), .B(exu_n18192), .Y(exu_n18220));
INVX1 exu_U30460(.A(exu_n18220), .Y(exu_n10788));
AND2X1 exu_U30461(.A(rml_next_canrestore_w[0]), .B(exu_n18192), .Y(exu_n18222));
INVX1 exu_U30462(.A(exu_n18222), .Y(exu_n10789));
AND2X1 exu_U30463(.A(rml_next_canrestore_w[2]), .B(exu_n18193), .Y(exu_n18224));
INVX1 exu_U30464(.A(exu_n18224), .Y(exu_n10790));
AND2X1 exu_U30465(.A(rml_next_canrestore_w[1]), .B(exu_n18193), .Y(exu_n18226));
INVX1 exu_U30466(.A(exu_n18226), .Y(exu_n10791));
AND2X1 exu_U30467(.A(rml_next_canrestore_w[0]), .B(exu_n18193), .Y(exu_n18228));
INVX1 exu_U30468(.A(exu_n18228), .Y(exu_n10792));
AND2X1 exu_U30469(.A(rml_next_canrestore_w[2]), .B(exu_n18194), .Y(exu_n18230));
INVX1 exu_U30470(.A(exu_n18230), .Y(exu_n10793));
AND2X1 exu_U30471(.A(rml_next_canrestore_w[1]), .B(exu_n18194), .Y(exu_n18232));
INVX1 exu_U30472(.A(exu_n18232), .Y(exu_n10794));
AND2X1 exu_U30473(.A(rml_next_canrestore_w[0]), .B(exu_n18194), .Y(exu_n18234));
INVX1 exu_U30474(.A(exu_n18234), .Y(exu_n10795));
AND2X1 exu_U30475(.A(rml_next_otherwin_w[2]), .B(exu_n18235), .Y(exu_n18256));
INVX1 exu_U30476(.A(exu_n18256), .Y(exu_n10796));
AND2X1 exu_U30477(.A(rml_next_otherwin_w[1]), .B(exu_n18235), .Y(exu_n18258));
INVX1 exu_U30478(.A(exu_n18258), .Y(exu_n10797));
AND2X1 exu_U30479(.A(rml_next_otherwin_w[0]), .B(exu_n18235), .Y(exu_n18260));
INVX1 exu_U30480(.A(exu_n18260), .Y(exu_n10798));
AND2X1 exu_U30481(.A(rml_next_otherwin_w[2]), .B(exu_n18236), .Y(exu_n18262));
INVX1 exu_U30482(.A(exu_n18262), .Y(exu_n10799));
AND2X1 exu_U30483(.A(rml_next_otherwin_w[1]), .B(exu_n18236), .Y(exu_n18264));
INVX1 exu_U30484(.A(exu_n18264), .Y(exu_n10800));
AND2X1 exu_U30485(.A(rml_next_otherwin_w[0]), .B(exu_n18236), .Y(exu_n18266));
INVX1 exu_U30486(.A(exu_n18266), .Y(exu_n10801));
AND2X1 exu_U30487(.A(rml_next_otherwin_w[2]), .B(exu_n18237), .Y(exu_n18268));
INVX1 exu_U30488(.A(exu_n18268), .Y(exu_n10802));
AND2X1 exu_U30489(.A(rml_next_otherwin_w[1]), .B(exu_n18237), .Y(exu_n18270));
INVX1 exu_U30490(.A(exu_n18270), .Y(exu_n10803));
AND2X1 exu_U30491(.A(rml_next_otherwin_w[0]), .B(exu_n18237), .Y(exu_n18272));
INVX1 exu_U30492(.A(exu_n18272), .Y(exu_n10804));
AND2X1 exu_U30493(.A(rml_next_otherwin_w[2]), .B(exu_n18238), .Y(exu_n18274));
INVX1 exu_U30494(.A(exu_n18274), .Y(exu_n10805));
AND2X1 exu_U30495(.A(rml_next_otherwin_w[1]), .B(exu_n18238), .Y(exu_n18276));
INVX1 exu_U30496(.A(exu_n18276), .Y(exu_n10806));
AND2X1 exu_U30497(.A(rml_next_otherwin_w[0]), .B(exu_n18238), .Y(exu_n18278));
INVX1 exu_U30498(.A(exu_n18278), .Y(exu_n10807));
AND2X1 exu_U30499(.A(rml_next_cleanwin_w[2]), .B(exu_n18279), .Y(exu_n18300));
INVX1 exu_U30500(.A(exu_n18300), .Y(exu_n10808));
AND2X1 exu_U30501(.A(rml_next_cleanwin_w[1]), .B(exu_n18279), .Y(exu_n18302));
INVX1 exu_U30502(.A(exu_n18302), .Y(exu_n10809));
AND2X1 exu_U30503(.A(rml_next_cleanwin_w[0]), .B(exu_n18279), .Y(exu_n18304));
INVX1 exu_U30504(.A(exu_n18304), .Y(exu_n10810));
AND2X1 exu_U30505(.A(rml_next_cleanwin_w[2]), .B(exu_n18280), .Y(exu_n18306));
INVX1 exu_U30506(.A(exu_n18306), .Y(exu_n10811));
AND2X1 exu_U30507(.A(rml_next_cleanwin_w[1]), .B(exu_n18280), .Y(exu_n18308));
INVX1 exu_U30508(.A(exu_n18308), .Y(exu_n10812));
AND2X1 exu_U30509(.A(rml_next_cleanwin_w[0]), .B(exu_n18280), .Y(exu_n18310));
INVX1 exu_U30510(.A(exu_n18310), .Y(exu_n10813));
AND2X1 exu_U30511(.A(rml_next_cleanwin_w[2]), .B(exu_n18281), .Y(exu_n18312));
INVX1 exu_U30512(.A(exu_n18312), .Y(exu_n10814));
AND2X1 exu_U30513(.A(rml_next_cleanwin_w[1]), .B(exu_n18281), .Y(exu_n18314));
INVX1 exu_U30514(.A(exu_n18314), .Y(exu_n10815));
AND2X1 exu_U30515(.A(rml_next_cleanwin_w[0]), .B(exu_n18281), .Y(exu_n18316));
INVX1 exu_U30516(.A(exu_n18316), .Y(exu_n10816));
AND2X1 exu_U30517(.A(rml_next_cleanwin_w[2]), .B(exu_n18282), .Y(exu_n18318));
INVX1 exu_U30518(.A(exu_n18318), .Y(exu_n10817));
AND2X1 exu_U30519(.A(rml_next_cleanwin_w[1]), .B(exu_n18282), .Y(exu_n18320));
INVX1 exu_U30520(.A(exu_n18320), .Y(exu_n10818));
AND2X1 exu_U30521(.A(rml_next_cleanwin_w[0]), .B(exu_n18282), .Y(exu_n18322));
INVX1 exu_U30522(.A(exu_n18322), .Y(exu_n10819));
AND2X1 exu_U30523(.A(byp_irf_rd_data_w[5]), .B(exu_n18323), .Y(exu_n18344));
INVX1 exu_U30524(.A(exu_n18344), .Y(exu_n10820));
AND2X1 exu_U30525(.A(byp_irf_rd_data_w[4]), .B(exu_n18323), .Y(exu_n18346));
INVX1 exu_U30526(.A(exu_n18346), .Y(exu_n10821));
AND2X1 exu_U30527(.A(byp_irf_rd_data_w[3]), .B(exu_n18323), .Y(exu_n18348));
INVX1 exu_U30528(.A(exu_n18348), .Y(exu_n10822));
AND2X1 exu_U30529(.A(byp_irf_rd_data_w[5]), .B(exu_n18324), .Y(exu_n18350));
INVX1 exu_U30530(.A(exu_n18350), .Y(exu_n10823));
AND2X1 exu_U30531(.A(byp_irf_rd_data_w[4]), .B(exu_n18324), .Y(exu_n18352));
INVX1 exu_U30532(.A(exu_n18352), .Y(exu_n10824));
AND2X1 exu_U30533(.A(byp_irf_rd_data_w[3]), .B(exu_n18324), .Y(exu_n18354));
INVX1 exu_U30534(.A(exu_n18354), .Y(exu_n10825));
AND2X1 exu_U30535(.A(byp_irf_rd_data_w[5]), .B(exu_n18325), .Y(exu_n18356));
INVX1 exu_U30536(.A(exu_n18356), .Y(exu_n10826));
AND2X1 exu_U30537(.A(byp_irf_rd_data_w[4]), .B(exu_n18325), .Y(exu_n18358));
INVX1 exu_U30538(.A(exu_n18358), .Y(exu_n10827));
AND2X1 exu_U30539(.A(byp_irf_rd_data_w[3]), .B(exu_n18325), .Y(exu_n18360));
INVX1 exu_U30540(.A(exu_n18360), .Y(exu_n10828));
AND2X1 exu_U30541(.A(byp_irf_rd_data_w[5]), .B(exu_n18326), .Y(exu_n18362));
INVX1 exu_U30542(.A(exu_n18362), .Y(exu_n10829));
AND2X1 exu_U30543(.A(byp_irf_rd_data_w[4]), .B(exu_n18326), .Y(exu_n18364));
INVX1 exu_U30544(.A(exu_n18364), .Y(exu_n10830));
AND2X1 exu_U30545(.A(byp_irf_rd_data_w[3]), .B(exu_n18326), .Y(exu_n18366));
INVX1 exu_U30546(.A(exu_n18366), .Y(exu_n10831));
AND2X1 exu_U30547(.A(byp_irf_rd_data_w[2]), .B(exu_n18323), .Y(exu_n18384));
INVX1 exu_U30548(.A(exu_n18384), .Y(exu_n10832));
AND2X1 exu_U30549(.A(byp_irf_rd_data_w[1]), .B(exu_n18323), .Y(exu_n18386));
INVX1 exu_U30550(.A(exu_n18386), .Y(exu_n10833));
AND2X1 exu_U30551(.A(byp_irf_rd_data_w[0]), .B(exu_n18323), .Y(exu_n18388));
INVX1 exu_U30552(.A(exu_n18388), .Y(exu_n10834));
AND2X1 exu_U30553(.A(byp_irf_rd_data_w[2]), .B(exu_n18324), .Y(exu_n18390));
INVX1 exu_U30554(.A(exu_n18390), .Y(exu_n10835));
AND2X1 exu_U30555(.A(byp_irf_rd_data_w[1]), .B(exu_n18324), .Y(exu_n18392));
INVX1 exu_U30556(.A(exu_n18392), .Y(exu_n10836));
AND2X1 exu_U30557(.A(byp_irf_rd_data_w[0]), .B(exu_n18324), .Y(exu_n18394));
INVX1 exu_U30558(.A(exu_n18394), .Y(exu_n10837));
AND2X1 exu_U30559(.A(byp_irf_rd_data_w[2]), .B(exu_n18325), .Y(exu_n18396));
INVX1 exu_U30560(.A(exu_n18396), .Y(exu_n10838));
AND2X1 exu_U30561(.A(byp_irf_rd_data_w[1]), .B(exu_n18325), .Y(exu_n18398));
INVX1 exu_U30562(.A(exu_n18398), .Y(exu_n10839));
AND2X1 exu_U30563(.A(byp_irf_rd_data_w[0]), .B(exu_n18325), .Y(exu_n18400));
INVX1 exu_U30564(.A(exu_n18400), .Y(exu_n10840));
AND2X1 exu_U30565(.A(byp_irf_rd_data_w[2]), .B(exu_n18326), .Y(exu_n18402));
INVX1 exu_U30566(.A(exu_n18402), .Y(exu_n10841));
AND2X1 exu_U30567(.A(byp_irf_rd_data_w[1]), .B(exu_n18326), .Y(exu_n18404));
INVX1 exu_U30568(.A(exu_n18404), .Y(exu_n10842));
AND2X1 exu_U30569(.A(byp_irf_rd_data_w[0]), .B(exu_n18326), .Y(exu_n18406));
INVX1 exu_U30570(.A(exu_n18406), .Y(exu_n10843));
AND2X1 exu_U30571(.A(exu_n16588), .B(rml_canrestore_wen_e), .Y(exu_n18432));
INVX1 exu_U30572(.A(exu_n18432), .Y(exu_n10844));
AND2X1 exu_U30573(.A(rml_rml_next_canrestore_e[1]), .B(rml_canrestore_wen_e), .Y(exu_n18434));
INVX1 exu_U30574(.A(exu_n18434), .Y(exu_n10845));
AND2X1 exu_U30575(.A(rml_rml_next_canrestore_e[2]), .B(rml_canrestore_wen_e), .Y(exu_n18436));
INVX1 exu_U30576(.A(exu_n18436), .Y(exu_n10846));
AND2X1 exu_U30577(.A(exu_n16587), .B(rml_n130), .Y(exu_n18438));
INVX1 exu_U30578(.A(exu_n18438), .Y(exu_n10847));
AND2X1 exu_U30579(.A(rml_rml_next_otherwin_e[1]), .B(rml_n130), .Y(exu_n18440));
INVX1 exu_U30580(.A(exu_n18440), .Y(exu_n10848));
AND2X1 exu_U30581(.A(rml_rml_next_otherwin_e[2]), .B(rml_n130), .Y(exu_n18442));
INVX1 exu_U30582(.A(exu_n18442), .Y(exu_n10849));
AND2X1 exu_U30583(.A(exu_n16585), .B(rml_n131), .Y(exu_n18444));
INVX1 exu_U30584(.A(exu_n18444), .Y(exu_n10850));
AND2X1 exu_U30585(.A(rml_rml_next_cleanwin_e[1]), .B(rml_n131), .Y(exu_n18446));
INVX1 exu_U30586(.A(exu_n18446), .Y(exu_n10851));
AND2X1 exu_U30587(.A(exu_n11852), .B(rml_n131), .Y(exu_n18448));
INVX1 exu_U30588(.A(exu_n18448), .Y(exu_n10852));
AND2X1 exu_U30589(.A(rml_next_cansave_w[0]), .B(rml_cansave_reg_n8), .Y(exu_n18450));
INVX1 exu_U30590(.A(exu_n18450), .Y(exu_n10853));
AND2X1 exu_U30591(.A(rml_next_cansave_w[1]), .B(rml_cansave_reg_n8), .Y(exu_n18452));
INVX1 exu_U30592(.A(exu_n18452), .Y(exu_n10854));
AND2X1 exu_U30593(.A(rml_next_cansave_w[2]), .B(rml_cansave_reg_n8), .Y(exu_n18454));
INVX1 exu_U30594(.A(exu_n18454), .Y(exu_n10855));
AND2X1 exu_U30595(.A(rml_next_cansave_w[0]), .B(rml_cansave_reg_n7), .Y(exu_n18456));
INVX1 exu_U30596(.A(exu_n18456), .Y(exu_n10856));
AND2X1 exu_U30597(.A(rml_next_cansave_w[1]), .B(rml_cansave_reg_n7), .Y(exu_n18458));
INVX1 exu_U30598(.A(exu_n18458), .Y(exu_n10857));
AND2X1 exu_U30599(.A(rml_next_cansave_w[2]), .B(rml_cansave_reg_n7), .Y(exu_n18460));
INVX1 exu_U30600(.A(exu_n18460), .Y(exu_n10858));
AND2X1 exu_U30601(.A(rml_next_cansave_w[0]), .B(rml_cansave_reg_n6), .Y(exu_n18462));
INVX1 exu_U30602(.A(exu_n18462), .Y(exu_n10859));
AND2X1 exu_U30603(.A(rml_next_cansave_w[1]), .B(rml_cansave_reg_n6), .Y(exu_n18464));
INVX1 exu_U30604(.A(exu_n18464), .Y(exu_n10860));
AND2X1 exu_U30605(.A(rml_next_cansave_w[2]), .B(rml_cansave_reg_n6), .Y(exu_n18466));
INVX1 exu_U30606(.A(exu_n18466), .Y(exu_n10861));
AND2X1 exu_U30607(.A(rml_next_cansave_w[0]), .B(rml_cansave_reg_n5), .Y(exu_n18468));
INVX1 exu_U30608(.A(exu_n18468), .Y(exu_n10862));
AND2X1 exu_U30609(.A(rml_next_cansave_w[1]), .B(rml_cansave_reg_n5), .Y(exu_n18470));
INVX1 exu_U30610(.A(exu_n18470), .Y(exu_n10863));
AND2X1 exu_U30611(.A(rml_next_cansave_w[2]), .B(rml_cansave_reg_n5), .Y(exu_n18472));
INVX1 exu_U30612(.A(exu_n18472), .Y(exu_n10864));
INVX1 exu_U30613(.A(div_dividend[41]), .Y(exu_n10865));
AND2X1 exu_U30614(.A(ecl_div_div64), .B(alu_logic_rs1_data_bf1[41]), .Y(exu_n19053));
INVX1 exu_U30615(.A(exu_n19053), .Y(exu_n10866));
INVX1 exu_U30616(.A(div_dividend[40]), .Y(exu_n10867));
AND2X1 exu_U30617(.A(alu_logic_rs1_data_bf1[40]), .B(ecl_div_div64), .Y(exu_n19055));
INVX1 exu_U30618(.A(exu_n19055), .Y(exu_n10868));
INVX1 exu_U30619(.A(div_dividend[39]), .Y(exu_n10869));
AND2X1 exu_U30620(.A(alu_logic_rs1_data_bf1[39]), .B(ecl_div_div64), .Y(exu_n19057));
INVX1 exu_U30621(.A(exu_n19057), .Y(exu_n10870));
INVX1 exu_U30622(.A(div_dividend[38]), .Y(exu_n10871));
AND2X1 exu_U30623(.A(alu_logic_rs1_data_bf1[38]), .B(ecl_div_div64), .Y(exu_n19059));
INVX1 exu_U30624(.A(exu_n19059), .Y(exu_n10872));
INVX1 exu_U30625(.A(div_dividend[37]), .Y(exu_n10873));
AND2X1 exu_U30626(.A(alu_logic_rs1_data_bf1[37]), .B(ecl_div_div64), .Y(exu_n19061));
INVX1 exu_U30627(.A(exu_n19061), .Y(exu_n10874));
INVX1 exu_U30628(.A(div_dividend[36]), .Y(exu_n10875));
AND2X1 exu_U30629(.A(alu_logic_rs1_data_bf1[36]), .B(ecl_div_div64), .Y(exu_n19063));
INVX1 exu_U30630(.A(exu_n19063), .Y(exu_n10876));
INVX1 exu_U30631(.A(div_dividend[35]), .Y(exu_n10877));
AND2X1 exu_U30632(.A(alu_logic_rs1_data_bf1[35]), .B(ecl_div_div64), .Y(exu_n19065));
INVX1 exu_U30633(.A(exu_n19065), .Y(exu_n10878));
INVX1 exu_U30634(.A(div_dividend[62]), .Y(exu_n10879));
AND2X1 exu_U30635(.A(alu_logic_rs1_data_bf1[62]), .B(ecl_div_div64), .Y(exu_n19069));
INVX1 exu_U30636(.A(exu_n19069), .Y(exu_n10880));
INVX1 exu_U30637(.A(div_dividend[34]), .Y(exu_n10881));
AND2X1 exu_U30638(.A(alu_logic_rs1_data_bf1[34]), .B(ecl_div_div64), .Y(exu_n19071));
INVX1 exu_U30639(.A(exu_n19071), .Y(exu_n10882));
INVX1 exu_U30640(.A(div_dividend[61]), .Y(exu_n10883));
AND2X1 exu_U30641(.A(alu_logic_rs1_data_bf1[61]), .B(ecl_div_div64), .Y(exu_n19073));
INVX1 exu_U30642(.A(exu_n19073), .Y(exu_n10884));
INVX1 exu_U30643(.A(div_dividend[60]), .Y(exu_n10885));
AND2X1 exu_U30644(.A(alu_logic_rs1_data_bf1[60]), .B(ecl_div_div64), .Y(exu_n19075));
INVX1 exu_U30645(.A(exu_n19075), .Y(exu_n10886));
INVX1 exu_U30646(.A(div_dividend[59]), .Y(exu_n10887));
AND2X1 exu_U30647(.A(alu_logic_rs1_data_bf1[59]), .B(ecl_div_div64), .Y(exu_n19077));
INVX1 exu_U30648(.A(exu_n19077), .Y(exu_n10888));
INVX1 exu_U30649(.A(div_dividend[58]), .Y(exu_n10889));
AND2X1 exu_U30650(.A(alu_logic_rs1_data_bf1[58]), .B(ecl_div_div64), .Y(exu_n19079));
INVX1 exu_U30651(.A(exu_n19079), .Y(exu_n10890));
INVX1 exu_U30652(.A(div_dividend[57]), .Y(exu_n10891));
AND2X1 exu_U30653(.A(alu_logic_rs1_data_bf1[57]), .B(ecl_div_div64), .Y(exu_n19081));
INVX1 exu_U30654(.A(exu_n19081), .Y(exu_n10892));
INVX1 exu_U30655(.A(div_dividend[56]), .Y(exu_n10893));
AND2X1 exu_U30656(.A(alu_logic_rs1_data_bf1[56]), .B(ecl_div_div64), .Y(exu_n19083));
INVX1 exu_U30657(.A(exu_n19083), .Y(exu_n10894));
INVX1 exu_U30658(.A(div_dividend[55]), .Y(exu_n10895));
AND2X1 exu_U30659(.A(alu_logic_rs1_data_bf1[55]), .B(ecl_div_div64), .Y(exu_n19085));
INVX1 exu_U30660(.A(exu_n19085), .Y(exu_n10896));
INVX1 exu_U30661(.A(div_dividend[54]), .Y(exu_n10897));
AND2X1 exu_U30662(.A(alu_logic_rs1_data_bf1[54]), .B(ecl_div_div64), .Y(exu_n19087));
INVX1 exu_U30663(.A(exu_n19087), .Y(exu_n10898));
INVX1 exu_U30664(.A(div_dividend[53]), .Y(exu_n10899));
AND2X1 exu_U30665(.A(alu_logic_rs1_data_bf1[53]), .B(ecl_div_div64), .Y(exu_n19089));
INVX1 exu_U30666(.A(exu_n19089), .Y(exu_n10900));
INVX1 exu_U30667(.A(div_dividend[52]), .Y(exu_n10901));
AND2X1 exu_U30668(.A(alu_logic_rs1_data_bf1[52]), .B(ecl_div_div64), .Y(exu_n19091));
INVX1 exu_U30669(.A(exu_n19091), .Y(exu_n10902));
INVX1 exu_U30670(.A(div_dividend[33]), .Y(exu_n10903));
AND2X1 exu_U30671(.A(alu_logic_rs1_data_bf1[33]), .B(ecl_div_div64), .Y(exu_n19093));
INVX1 exu_U30672(.A(exu_n19093), .Y(exu_n10904));
INVX1 exu_U30673(.A(div_dividend[51]), .Y(exu_n10905));
AND2X1 exu_U30674(.A(alu_logic_rs1_data_bf1[51]), .B(ecl_div_div64), .Y(exu_n19095));
INVX1 exu_U30675(.A(exu_n19095), .Y(exu_n10906));
INVX1 exu_U30676(.A(div_dividend[50]), .Y(exu_n10907));
AND2X1 exu_U30677(.A(alu_logic_rs1_data_bf1[50]), .B(ecl_div_div64), .Y(exu_n19097));
INVX1 exu_U30678(.A(exu_n19097), .Y(exu_n10908));
INVX1 exu_U30679(.A(div_dividend[49]), .Y(exu_n10909));
AND2X1 exu_U30680(.A(alu_logic_rs1_data_bf1[49]), .B(ecl_div_div64), .Y(exu_n19099));
INVX1 exu_U30681(.A(exu_n19099), .Y(exu_n10910));
INVX1 exu_U30682(.A(div_dividend[48]), .Y(exu_n10911));
AND2X1 exu_U30683(.A(alu_logic_rs1_data_bf1[48]), .B(ecl_div_div64), .Y(exu_n19101));
INVX1 exu_U30684(.A(exu_n19101), .Y(exu_n10912));
INVX1 exu_U30685(.A(div_dividend[47]), .Y(exu_n10913));
AND2X1 exu_U30686(.A(alu_logic_rs1_data_bf1[47]), .B(ecl_div_div64), .Y(exu_n19103));
INVX1 exu_U30687(.A(exu_n19103), .Y(exu_n10914));
INVX1 exu_U30688(.A(div_dividend[46]), .Y(exu_n10915));
AND2X1 exu_U30689(.A(alu_logic_rs1_data_bf1[46]), .B(ecl_div_div64), .Y(exu_n19105));
INVX1 exu_U30690(.A(exu_n19105), .Y(exu_n10916));
INVX1 exu_U30691(.A(div_dividend[45]), .Y(exu_n10917));
AND2X1 exu_U30692(.A(alu_logic_rs1_data_bf1[45]), .B(ecl_div_div64), .Y(exu_n19107));
INVX1 exu_U30693(.A(exu_n19107), .Y(exu_n10918));
INVX1 exu_U30694(.A(div_dividend[44]), .Y(exu_n10919));
AND2X1 exu_U30695(.A(alu_logic_rs1_data_bf1[44]), .B(ecl_div_div64), .Y(exu_n19109));
INVX1 exu_U30696(.A(exu_n19109), .Y(exu_n10920));
INVX1 exu_U30697(.A(div_dividend[43]), .Y(exu_n10921));
AND2X1 exu_U30698(.A(alu_logic_rs1_data_bf1[43]), .B(ecl_div_div64), .Y(exu_n19111));
INVX1 exu_U30699(.A(exu_n19111), .Y(exu_n10922));
INVX1 exu_U30700(.A(div_dividend[42]), .Y(exu_n10923));
AND2X1 exu_U30701(.A(alu_logic_rs1_data_bf1[42]), .B(ecl_div_div64), .Y(exu_n19113));
INVX1 exu_U30702(.A(exu_n19113), .Y(exu_n10924));
INVX1 exu_U30703(.A(div_dividend[32]), .Y(exu_n10925));
AND2X1 exu_U30704(.A(alu_logic_rs1_data_bf1[32]), .B(ecl_div_div64), .Y(exu_n19115));
INVX1 exu_U30705(.A(exu_n19115), .Y(exu_n10926));
INVX1 exu_U30706(.A(div_din[72]), .Y(exu_n10927));
AND2X1 exu_U30707(.A(ecl_div_muls), .B(alu_logic_rs1_data_bf1[10]), .Y(exu_n19117));
INVX1 exu_U30708(.A(exu_n19117), .Y(exu_n10928));
INVX1 exu_U30709(.A(div_din[71]), .Y(exu_n10929));
AND2X1 exu_U30710(.A(alu_logic_rs1_data_bf1[9]), .B(ecl_div_muls), .Y(exu_n19118));
INVX1 exu_U30711(.A(exu_n19118), .Y(exu_n10930));
INVX1 exu_U30712(.A(div_din[70]), .Y(exu_n10931));
AND2X1 exu_U30713(.A(alu_logic_rs1_data_bf1[8]), .B(ecl_div_muls), .Y(exu_n19119));
INVX1 exu_U30714(.A(exu_n19119), .Y(exu_n10932));
INVX1 exu_U30715(.A(div_din[69]), .Y(exu_n10933));
AND2X1 exu_U30716(.A(alu_logic_rs1_data_bf1[7]), .B(ecl_div_muls), .Y(exu_n19120));
INVX1 exu_U30717(.A(exu_n19120), .Y(exu_n10934));
INVX1 exu_U30718(.A(div_din[68]), .Y(exu_n10935));
AND2X1 exu_U30719(.A(alu_logic_rs1_data_bf1[6]), .B(ecl_div_muls), .Y(exu_n19121));
INVX1 exu_U30720(.A(exu_n19121), .Y(exu_n10936));
INVX1 exu_U30721(.A(div_din[67]), .Y(exu_n10937));
AND2X1 exu_U30722(.A(alu_logic_rs1_data_bf1[5]), .B(ecl_div_muls), .Y(exu_n19122));
INVX1 exu_U30723(.A(exu_n19122), .Y(exu_n10938));
INVX1 exu_U30724(.A(div_din[66]), .Y(exu_n10939));
AND2X1 exu_U30725(.A(alu_logic_rs1_data_bf1[4]), .B(ecl_div_muls), .Y(exu_n19123));
INVX1 exu_U30726(.A(exu_n19123), .Y(exu_n10940));
INVX1 exu_U30727(.A(div_din[94]), .Y(exu_n10941));
AND2X1 exu_U30728(.A(exu_n16581), .B(ecl_div_muls), .Y(exu_n19124));
INVX1 exu_U30729(.A(exu_n19124), .Y(exu_n10942));
INVX1 exu_U30730(.A(div_din[93]), .Y(exu_n10943));
AND2X1 exu_U30731(.A(alu_logic_rs1_data_bf1[31]), .B(ecl_div_muls), .Y(exu_n19125));
INVX1 exu_U30732(.A(exu_n19125), .Y(exu_n10944));
INVX1 exu_U30733(.A(div_din[65]), .Y(exu_n10945));
AND2X1 exu_U30734(.A(alu_logic_rs1_data_bf1[3]), .B(ecl_div_muls), .Y(exu_n19126));
INVX1 exu_U30735(.A(exu_n19126), .Y(exu_n10946));
INVX1 exu_U30736(.A(div_din[92]), .Y(exu_n10947));
AND2X1 exu_U30737(.A(alu_logic_rs1_data_bf1[30]), .B(ecl_div_muls), .Y(exu_n19127));
INVX1 exu_U30738(.A(exu_n19127), .Y(exu_n10948));
INVX1 exu_U30739(.A(div_din[91]), .Y(exu_n10949));
AND2X1 exu_U30740(.A(alu_logic_rs1_data_bf1[29]), .B(ecl_div_muls), .Y(exu_n19128));
INVX1 exu_U30741(.A(exu_n19128), .Y(exu_n10950));
INVX1 exu_U30742(.A(div_din[90]), .Y(exu_n10951));
AND2X1 exu_U30743(.A(alu_logic_rs1_data_bf1[28]), .B(ecl_div_muls), .Y(exu_n19129));
INVX1 exu_U30744(.A(exu_n19129), .Y(exu_n10952));
INVX1 exu_U30745(.A(div_din[89]), .Y(exu_n10953));
AND2X1 exu_U30746(.A(alu_logic_rs1_data_bf1[27]), .B(ecl_div_muls), .Y(exu_n19130));
INVX1 exu_U30747(.A(exu_n19130), .Y(exu_n10954));
INVX1 exu_U30748(.A(div_din[88]), .Y(exu_n10955));
AND2X1 exu_U30749(.A(alu_logic_rs1_data_bf1[26]), .B(ecl_div_muls), .Y(exu_n19131));
INVX1 exu_U30750(.A(exu_n19131), .Y(exu_n10956));
INVX1 exu_U30751(.A(div_din[87]), .Y(exu_n10957));
AND2X1 exu_U30752(.A(alu_logic_rs1_data_bf1[25]), .B(ecl_div_muls), .Y(exu_n19132));
INVX1 exu_U30753(.A(exu_n19132), .Y(exu_n10958));
INVX1 exu_U30754(.A(div_din[86]), .Y(exu_n10959));
AND2X1 exu_U30755(.A(alu_logic_rs1_data_bf1[24]), .B(ecl_div_muls), .Y(exu_n19133));
INVX1 exu_U30756(.A(exu_n19133), .Y(exu_n10960));
INVX1 exu_U30757(.A(div_din[85]), .Y(exu_n10961));
AND2X1 exu_U30758(.A(alu_logic_rs1_data_bf1[23]), .B(ecl_div_muls), .Y(exu_n19134));
INVX1 exu_U30759(.A(exu_n19134), .Y(exu_n10962));
INVX1 exu_U30760(.A(div_din[84]), .Y(exu_n10963));
AND2X1 exu_U30761(.A(alu_logic_rs1_data_bf1[22]), .B(ecl_div_muls), .Y(exu_n19135));
INVX1 exu_U30762(.A(exu_n19135), .Y(exu_n10964));
INVX1 exu_U30763(.A(div_din[83]), .Y(exu_n10965));
AND2X1 exu_U30764(.A(alu_logic_rs1_data_bf1[21]), .B(ecl_div_muls), .Y(exu_n19136));
INVX1 exu_U30765(.A(exu_n19136), .Y(exu_n10966));
INVX1 exu_U30766(.A(div_din[64]), .Y(exu_n10967));
AND2X1 exu_U30767(.A(alu_logic_rs1_data_bf1[2]), .B(ecl_div_muls), .Y(exu_n19137));
INVX1 exu_U30768(.A(exu_n19137), .Y(exu_n10968));
INVX1 exu_U30769(.A(div_din[82]), .Y(exu_n10969));
AND2X1 exu_U30770(.A(alu_logic_rs1_data_bf1[20]), .B(ecl_div_muls), .Y(exu_n19138));
INVX1 exu_U30771(.A(exu_n19138), .Y(exu_n10970));
INVX1 exu_U30772(.A(div_din[81]), .Y(exu_n10971));
AND2X1 exu_U30773(.A(alu_logic_rs1_data_bf1[19]), .B(ecl_div_muls), .Y(exu_n19139));
INVX1 exu_U30774(.A(exu_n19139), .Y(exu_n10972));
INVX1 exu_U30775(.A(div_din[80]), .Y(exu_n10973));
AND2X1 exu_U30776(.A(alu_logic_rs1_data_bf1[18]), .B(ecl_div_muls), .Y(exu_n19140));
INVX1 exu_U30777(.A(exu_n19140), .Y(exu_n10974));
INVX1 exu_U30778(.A(div_din[79]), .Y(exu_n10975));
AND2X1 exu_U30779(.A(alu_logic_rs1_data_bf1[17]), .B(ecl_div_muls), .Y(exu_n19141));
INVX1 exu_U30780(.A(exu_n19141), .Y(exu_n10976));
INVX1 exu_U30781(.A(div_din[78]), .Y(exu_n10977));
AND2X1 exu_U30782(.A(alu_logic_rs1_data_bf1[16]), .B(ecl_div_muls), .Y(exu_n19142));
INVX1 exu_U30783(.A(exu_n19142), .Y(exu_n10978));
INVX1 exu_U30784(.A(div_din[77]), .Y(exu_n10979));
AND2X1 exu_U30785(.A(alu_logic_rs1_data_bf1[15]), .B(ecl_div_muls), .Y(exu_n19143));
INVX1 exu_U30786(.A(exu_n19143), .Y(exu_n10980));
INVX1 exu_U30787(.A(div_din[76]), .Y(exu_n10981));
AND2X1 exu_U30788(.A(alu_logic_rs1_data_bf1[14]), .B(ecl_div_muls), .Y(exu_n19144));
INVX1 exu_U30789(.A(exu_n19144), .Y(exu_n10982));
INVX1 exu_U30790(.A(div_din[75]), .Y(exu_n10983));
AND2X1 exu_U30791(.A(alu_logic_rs1_data_bf1[13]), .B(ecl_div_muls), .Y(exu_n19145));
INVX1 exu_U30792(.A(exu_n19145), .Y(exu_n10984));
INVX1 exu_U30793(.A(div_din[74]), .Y(exu_n10985));
AND2X1 exu_U30794(.A(alu_logic_rs1_data_bf1[12]), .B(ecl_div_muls), .Y(exu_n19146));
INVX1 exu_U30795(.A(exu_n19146), .Y(exu_n10986));
INVX1 exu_U30796(.A(div_din[73]), .Y(exu_n10987));
AND2X1 exu_U30797(.A(alu_logic_rs1_data_bf1[11]), .B(ecl_div_muls), .Y(exu_n19147));
INVX1 exu_U30798(.A(exu_n19147), .Y(exu_n10988));
INVX1 exu_U30799(.A(div_din[63]), .Y(exu_n10989));
AND2X1 exu_U30800(.A(alu_logic_rs1_data_bf1[1]), .B(ecl_div_muls), .Y(exu_n19149));
INVX1 exu_U30801(.A(exu_n19149), .Y(exu_n10990));
OR2X1 exu_U30802(.A(ecl_ifu_exu_rs3_d[1]), .B(ecl_ifu_exu_rs3_d[0]), .Y(exu_n19217));
INVX1 exu_U30803(.A(exu_n19217), .Y(exu_n10991));
OR2X1 exu_U30804(.A(ecc_rs2_err_e[0]), .B(exu_n20002), .Y(exu_n19998));
INVX1 exu_U30805(.A(exu_n19998), .Y(exu_n10992));
OR2X1 exu_U30806(.A(ecc_rs3_err_e[0]), .B(exu_n20138), .Y(exu_n20134));
INVX1 exu_U30807(.A(exu_n20134), .Y(exu_n10993));
INVX1 exu_U30808(.A(bypass_rs2_data_w2[8]), .Y(exu_n10994));
INVX1 exu_U30809(.A(bypass_rs2_data_w2[7]), .Y(exu_n10995));
INVX1 exu_U30810(.A(bypass_rs2_data_w2[6]), .Y(exu_n10996));
INVX1 exu_U30811(.A(bypass_rs2_data_w2[63]), .Y(exu_n10997));
INVX1 exu_U30812(.A(bypass_rs2_data_w2[62]), .Y(exu_n10998));
INVX1 exu_U30813(.A(bypass_rs2_data_w2[61]), .Y(exu_n10999));
INVX1 exu_U30814(.A(bypass_rs2_data_w2[60]), .Y(exu_n11000));
INVX1 exu_U30815(.A(bypass_rs2_data_w2[5]), .Y(exu_n11001));
INVX1 exu_U30816(.A(bypass_rs2_data_w2[59]), .Y(exu_n11002));
INVX1 exu_U30817(.A(bypass_rs2_data_w2[58]), .Y(exu_n11003));
INVX1 exu_U30818(.A(bypass_rs2_data_w2[57]), .Y(exu_n11004));
INVX1 exu_U30819(.A(bypass_rs2_data_w2[56]), .Y(exu_n11005));
INVX1 exu_U30820(.A(bypass_rs2_data_w2[55]), .Y(exu_n11006));
INVX1 exu_U30821(.A(bypass_rs2_data_w2[54]), .Y(exu_n11007));
INVX1 exu_U30822(.A(bypass_rs2_data_w2[53]), .Y(exu_n11008));
INVX1 exu_U30823(.A(bypass_rs2_data_w2[52]), .Y(exu_n11009));
INVX1 exu_U30824(.A(bypass_rs2_data_w2[51]), .Y(exu_n11010));
INVX1 exu_U30825(.A(bypass_rs2_data_w2[50]), .Y(exu_n11011));
INVX1 exu_U30826(.A(bypass_rs2_data_w2[4]), .Y(exu_n11012));
INVX1 exu_U30827(.A(bypass_rs2_data_w2[49]), .Y(exu_n11013));
INVX1 exu_U30828(.A(bypass_rs2_data_w2[48]), .Y(exu_n11014));
INVX1 exu_U30829(.A(bypass_rs2_data_w2[47]), .Y(exu_n11015));
INVX1 exu_U30830(.A(bypass_rs2_data_w2[46]), .Y(exu_n11016));
INVX1 exu_U30831(.A(bypass_rs2_data_w2[45]), .Y(exu_n11017));
INVX1 exu_U30832(.A(bypass_rs2_data_w2[44]), .Y(exu_n11018));
INVX1 exu_U30833(.A(bypass_rs2_data_w2[43]), .Y(exu_n11019));
INVX1 exu_U30834(.A(bypass_rs2_data_w2[42]), .Y(exu_n11020));
INVX1 exu_U30835(.A(bypass_rs2_data_w2[41]), .Y(exu_n11021));
INVX1 exu_U30836(.A(bypass_rs2_data_w2[40]), .Y(exu_n11022));
INVX1 exu_U30837(.A(bypass_rs2_data_w2[3]), .Y(exu_n11023));
INVX1 exu_U30838(.A(bypass_rs2_data_w2[39]), .Y(exu_n11024));
INVX1 exu_U30839(.A(bypass_rs2_data_w2[38]), .Y(exu_n11025));
INVX1 exu_U30840(.A(bypass_rs2_data_w2[37]), .Y(exu_n11026));
INVX1 exu_U30841(.A(bypass_rs2_data_w2[36]), .Y(exu_n11027));
INVX1 exu_U30842(.A(bypass_rs2_data_w2[35]), .Y(exu_n11028));
INVX1 exu_U30843(.A(bypass_rs2_data_w2[34]), .Y(exu_n11029));
INVX1 exu_U30844(.A(bypass_rs2_data_w2[33]), .Y(exu_n11030));
INVX1 exu_U30845(.A(bypass_rs2_data_w2[32]), .Y(exu_n11031));
INVX1 exu_U30846(.A(bypass_rs2_data_w2[31]), .Y(exu_n11032));
INVX1 exu_U30847(.A(bypass_rs2_data_w2[30]), .Y(exu_n11033));
INVX1 exu_U30848(.A(bypass_rs2_data_w2[2]), .Y(exu_n11034));
INVX1 exu_U30849(.A(bypass_rs2_data_w2[29]), .Y(exu_n11035));
INVX1 exu_U30850(.A(bypass_rs2_data_w2[28]), .Y(exu_n11036));
INVX1 exu_U30851(.A(bypass_rs2_data_w2[27]), .Y(exu_n11037));
INVX1 exu_U30852(.A(bypass_rs2_data_w2[26]), .Y(exu_n11038));
INVX1 exu_U30853(.A(bypass_rs2_data_w2[25]), .Y(exu_n11039));
INVX1 exu_U30854(.A(bypass_rs2_data_w2[24]), .Y(exu_n11040));
INVX1 exu_U30855(.A(bypass_rs2_data_w2[23]), .Y(exu_n11041));
INVX1 exu_U30856(.A(bypass_rs2_data_w2[22]), .Y(exu_n11042));
INVX1 exu_U30857(.A(bypass_rs2_data_w2[21]), .Y(exu_n11043));
INVX1 exu_U30858(.A(bypass_rs2_data_w2[20]), .Y(exu_n11044));
INVX1 exu_U30859(.A(bypass_rs2_data_w2[1]), .Y(exu_n11045));
INVX1 exu_U30860(.A(bypass_rs2_data_w2[19]), .Y(exu_n11046));
INVX1 exu_U30861(.A(bypass_rs2_data_w2[18]), .Y(exu_n11047));
INVX1 exu_U30862(.A(bypass_rs2_data_w2[17]), .Y(exu_n11048));
INVX1 exu_U30863(.A(bypass_rs2_data_w2[16]), .Y(exu_n11049));
INVX1 exu_U30864(.A(bypass_rs2_data_w2[15]), .Y(exu_n11050));
INVX1 exu_U30865(.A(bypass_rs2_data_w2[14]), .Y(exu_n11051));
INVX1 exu_U30866(.A(bypass_rs2_data_w2[13]), .Y(exu_n11052));
INVX1 exu_U30867(.A(bypass_rs2_data_w2[12]), .Y(exu_n11053));
INVX1 exu_U30868(.A(bypass_rs2_data_w2[11]), .Y(exu_n11054));
INVX1 exu_U30869(.A(bypass_rs2_data_w2[10]), .Y(exu_n11055));
INVX1 exu_U30870(.A(bypass_rs2_data_w2[0]), .Y(exu_n11056));
INVX1 exu_U30871(.A(exu_n28632), .Y(exu_n11057));
AND2X1 exu_U30872(.A(exu_n28264), .B(exu_n16223), .Y(exu_n28633));
INVX1 exu_U30873(.A(exu_n28633), .Y(exu_n11058));
AND2X1 exu_U30874(.A(ecl_byp_restore_m), .B(exu_tlu_wsr_data_m[9]), .Y(exu_n30145));
INVX1 exu_U30875(.A(exu_n30145), .Y(exu_n11059));
AND2X1 exu_U30876(.A(exu_tlu_wsr_data_m[8]), .B(ecl_byp_restore_m), .Y(exu_n30147));
INVX1 exu_U30877(.A(exu_n30147), .Y(exu_n11060));
AND2X1 exu_U30878(.A(exu_tlu_wsr_data_m[7]), .B(ecl_byp_restore_m), .Y(exu_n30149));
INVX1 exu_U30879(.A(exu_n30149), .Y(exu_n11061));
AND2X1 exu_U30880(.A(exu_tlu_wsr_data_m[6]), .B(ecl_byp_restore_m), .Y(exu_n30151));
INVX1 exu_U30881(.A(exu_n30151), .Y(exu_n11062));
AND2X1 exu_U30882(.A(exu_tlu_wsr_data_m[63]), .B(ecl_byp_restore_m), .Y(exu_n30153));
INVX1 exu_U30883(.A(exu_n30153), .Y(exu_n11063));
AND2X1 exu_U30884(.A(exu_tlu_wsr_data_m[62]), .B(ecl_byp_restore_m), .Y(exu_n30155));
INVX1 exu_U30885(.A(exu_n30155), .Y(exu_n11064));
AND2X1 exu_U30886(.A(exu_tlu_wsr_data_m[61]), .B(ecl_byp_restore_m), .Y(exu_n30157));
INVX1 exu_U30887(.A(exu_n30157), .Y(exu_n11065));
AND2X1 exu_U30888(.A(exu_tlu_wsr_data_m[60]), .B(ecl_byp_restore_m), .Y(exu_n30159));
INVX1 exu_U30889(.A(exu_n30159), .Y(exu_n11066));
AND2X1 exu_U30890(.A(exu_tlu_wsr_data_m[5]), .B(ecl_byp_restore_m), .Y(exu_n30161));
INVX1 exu_U30891(.A(exu_n30161), .Y(exu_n11067));
AND2X1 exu_U30892(.A(exu_tlu_wsr_data_m[59]), .B(ecl_byp_restore_m), .Y(exu_n30163));
INVX1 exu_U30893(.A(exu_n30163), .Y(exu_n11068));
AND2X1 exu_U30894(.A(exu_tlu_wsr_data_m[58]), .B(ecl_byp_restore_m), .Y(exu_n30165));
INVX1 exu_U30895(.A(exu_n30165), .Y(exu_n11069));
AND2X1 exu_U30896(.A(exu_tlu_wsr_data_m[57]), .B(ecl_byp_restore_m), .Y(exu_n30167));
INVX1 exu_U30897(.A(exu_n30167), .Y(exu_n11070));
AND2X1 exu_U30898(.A(exu_tlu_wsr_data_m[56]), .B(ecl_byp_restore_m), .Y(exu_n30169));
INVX1 exu_U30899(.A(exu_n30169), .Y(exu_n11071));
AND2X1 exu_U30900(.A(exu_tlu_wsr_data_m[55]), .B(ecl_byp_restore_m), .Y(exu_n30171));
INVX1 exu_U30901(.A(exu_n30171), .Y(exu_n11072));
AND2X1 exu_U30902(.A(exu_tlu_wsr_data_m[54]), .B(ecl_byp_restore_m), .Y(exu_n30173));
INVX1 exu_U30903(.A(exu_n30173), .Y(exu_n11073));
AND2X1 exu_U30904(.A(exu_tlu_wsr_data_m[53]), .B(ecl_byp_restore_m), .Y(exu_n30175));
INVX1 exu_U30905(.A(exu_n30175), .Y(exu_n11074));
AND2X1 exu_U30906(.A(exu_tlu_wsr_data_m[52]), .B(ecl_byp_restore_m), .Y(exu_n30177));
INVX1 exu_U30907(.A(exu_n30177), .Y(exu_n11075));
AND2X1 exu_U30908(.A(exu_tlu_wsr_data_m[51]), .B(ecl_byp_restore_m), .Y(exu_n30179));
INVX1 exu_U30909(.A(exu_n30179), .Y(exu_n11076));
AND2X1 exu_U30910(.A(exu_tlu_wsr_data_m[50]), .B(ecl_byp_restore_m), .Y(exu_n30181));
INVX1 exu_U30911(.A(exu_n30181), .Y(exu_n11077));
AND2X1 exu_U30912(.A(exu_tlu_wsr_data_m[4]), .B(ecl_byp_restore_m), .Y(exu_n30183));
INVX1 exu_U30913(.A(exu_n30183), .Y(exu_n11078));
AND2X1 exu_U30914(.A(exu_tlu_wsr_data_m[49]), .B(ecl_byp_restore_m), .Y(exu_n30185));
INVX1 exu_U30915(.A(exu_n30185), .Y(exu_n11079));
AND2X1 exu_U30916(.A(exu_tlu_wsr_data_m[48]), .B(ecl_byp_restore_m), .Y(exu_n30187));
INVX1 exu_U30917(.A(exu_n30187), .Y(exu_n11080));
AND2X1 exu_U30918(.A(exu_tlu_wsr_data_m[47]), .B(ecl_byp_restore_m), .Y(exu_n30189));
INVX1 exu_U30919(.A(exu_n30189), .Y(exu_n11081));
AND2X1 exu_U30920(.A(exu_tlu_wsr_data_m[46]), .B(ecl_byp_restore_m), .Y(exu_n30191));
INVX1 exu_U30921(.A(exu_n30191), .Y(exu_n11082));
AND2X1 exu_U30922(.A(exu_tlu_wsr_data_m[45]), .B(ecl_byp_restore_m), .Y(exu_n30193));
INVX1 exu_U30923(.A(exu_n30193), .Y(exu_n11083));
AND2X1 exu_U30924(.A(exu_tlu_wsr_data_m[44]), .B(ecl_byp_restore_m), .Y(exu_n30195));
INVX1 exu_U30925(.A(exu_n30195), .Y(exu_n11084));
AND2X1 exu_U30926(.A(exu_tlu_wsr_data_m[43]), .B(ecl_byp_restore_m), .Y(exu_n30197));
INVX1 exu_U30927(.A(exu_n30197), .Y(exu_n11085));
AND2X1 exu_U30928(.A(exu_tlu_wsr_data_m[42]), .B(ecl_byp_restore_m), .Y(exu_n30199));
INVX1 exu_U30929(.A(exu_n30199), .Y(exu_n11086));
AND2X1 exu_U30930(.A(exu_tlu_wsr_data_m[41]), .B(ecl_byp_restore_m), .Y(exu_n30201));
INVX1 exu_U30931(.A(exu_n30201), .Y(exu_n11087));
AND2X1 exu_U30932(.A(exu_tlu_wsr_data_m[40]), .B(ecl_byp_restore_m), .Y(exu_n30203));
INVX1 exu_U30933(.A(exu_n30203), .Y(exu_n11088));
AND2X1 exu_U30934(.A(exu_tlu_wsr_data_m[3]), .B(ecl_byp_restore_m), .Y(exu_n30205));
INVX1 exu_U30935(.A(exu_n30205), .Y(exu_n11089));
AND2X1 exu_U30936(.A(exu_tlu_wsr_data_m[39]), .B(ecl_byp_restore_m), .Y(exu_n30207));
INVX1 exu_U30937(.A(exu_n30207), .Y(exu_n11090));
AND2X1 exu_U30938(.A(exu_tlu_wsr_data_m[38]), .B(ecl_byp_restore_m), .Y(exu_n30209));
INVX1 exu_U30939(.A(exu_n30209), .Y(exu_n11091));
AND2X1 exu_U30940(.A(exu_tlu_wsr_data_m[37]), .B(ecl_byp_restore_m), .Y(exu_n30211));
INVX1 exu_U30941(.A(exu_n30211), .Y(exu_n11092));
AND2X1 exu_U30942(.A(exu_tlu_wsr_data_m[36]), .B(ecl_byp_restore_m), .Y(exu_n30213));
INVX1 exu_U30943(.A(exu_n30213), .Y(exu_n11093));
AND2X1 exu_U30944(.A(exu_tlu_wsr_data_m[35]), .B(ecl_byp_restore_m), .Y(exu_n30215));
INVX1 exu_U30945(.A(exu_n30215), .Y(exu_n11094));
AND2X1 exu_U30946(.A(exu_tlu_wsr_data_m[34]), .B(ecl_byp_restore_m), .Y(exu_n30217));
INVX1 exu_U30947(.A(exu_n30217), .Y(exu_n11095));
AND2X1 exu_U30948(.A(exu_tlu_wsr_data_m[33]), .B(ecl_byp_restore_m), .Y(exu_n30219));
INVX1 exu_U30949(.A(exu_n30219), .Y(exu_n11096));
AND2X1 exu_U30950(.A(exu_tlu_wsr_data_m[32]), .B(ecl_byp_restore_m), .Y(exu_n30221));
INVX1 exu_U30951(.A(exu_n30221), .Y(exu_n11097));
AND2X1 exu_U30952(.A(exu_tlu_wsr_data_m[31]), .B(ecl_byp_restore_m), .Y(exu_n30223));
INVX1 exu_U30953(.A(exu_n30223), .Y(exu_n11098));
AND2X1 exu_U30954(.A(exu_tlu_wsr_data_m[30]), .B(ecl_byp_restore_m), .Y(exu_n30225));
INVX1 exu_U30955(.A(exu_n30225), .Y(exu_n11099));
AND2X1 exu_U30956(.A(exu_tlu_wsr_data_m[2]), .B(ecl_byp_restore_m), .Y(exu_n30227));
INVX1 exu_U30957(.A(exu_n30227), .Y(exu_n11100));
AND2X1 exu_U30958(.A(exu_tlu_wsr_data_m[29]), .B(ecl_byp_restore_m), .Y(exu_n30229));
INVX1 exu_U30959(.A(exu_n30229), .Y(exu_n11101));
AND2X1 exu_U30960(.A(exu_tlu_wsr_data_m[28]), .B(ecl_byp_restore_m), .Y(exu_n30231));
INVX1 exu_U30961(.A(exu_n30231), .Y(exu_n11102));
AND2X1 exu_U30962(.A(exu_tlu_wsr_data_m[27]), .B(ecl_byp_restore_m), .Y(exu_n30233));
INVX1 exu_U30963(.A(exu_n30233), .Y(exu_n11103));
AND2X1 exu_U30964(.A(exu_tlu_wsr_data_m[26]), .B(ecl_byp_restore_m), .Y(exu_n30235));
INVX1 exu_U30965(.A(exu_n30235), .Y(exu_n11104));
AND2X1 exu_U30966(.A(exu_tlu_wsr_data_m[25]), .B(ecl_byp_restore_m), .Y(exu_n30237));
INVX1 exu_U30967(.A(exu_n30237), .Y(exu_n11105));
AND2X1 exu_U30968(.A(exu_tlu_wsr_data_m[24]), .B(ecl_byp_restore_m), .Y(exu_n30239));
INVX1 exu_U30969(.A(exu_n30239), .Y(exu_n11106));
AND2X1 exu_U30970(.A(exu_tlu_wsr_data_m[23]), .B(ecl_byp_restore_m), .Y(exu_n30241));
INVX1 exu_U30971(.A(exu_n30241), .Y(exu_n11107));
AND2X1 exu_U30972(.A(exu_tlu_wsr_data_m[22]), .B(ecl_byp_restore_m), .Y(exu_n30243));
INVX1 exu_U30973(.A(exu_n30243), .Y(exu_n11108));
AND2X1 exu_U30974(.A(exu_tlu_wsr_data_m[21]), .B(ecl_byp_restore_m), .Y(exu_n30245));
INVX1 exu_U30975(.A(exu_n30245), .Y(exu_n11109));
AND2X1 exu_U30976(.A(exu_tlu_wsr_data_m[20]), .B(ecl_byp_restore_m), .Y(exu_n30247));
INVX1 exu_U30977(.A(exu_n30247), .Y(exu_n11110));
AND2X1 exu_U30978(.A(exu_tlu_wsr_data_m[1]), .B(ecl_byp_restore_m), .Y(exu_n30249));
INVX1 exu_U30979(.A(exu_n30249), .Y(exu_n11111));
AND2X1 exu_U30980(.A(exu_tlu_wsr_data_m[19]), .B(ecl_byp_restore_m), .Y(exu_n30251));
INVX1 exu_U30981(.A(exu_n30251), .Y(exu_n11112));
AND2X1 exu_U30982(.A(exu_tlu_wsr_data_m[18]), .B(ecl_byp_restore_m), .Y(exu_n30253));
INVX1 exu_U30983(.A(exu_n30253), .Y(exu_n11113));
AND2X1 exu_U30984(.A(exu_tlu_wsr_data_m[17]), .B(ecl_byp_restore_m), .Y(exu_n30255));
INVX1 exu_U30985(.A(exu_n30255), .Y(exu_n11114));
AND2X1 exu_U30986(.A(exu_tlu_wsr_data_m[16]), .B(ecl_byp_restore_m), .Y(exu_n30257));
INVX1 exu_U30987(.A(exu_n30257), .Y(exu_n11115));
AND2X1 exu_U30988(.A(exu_tlu_wsr_data_m[15]), .B(ecl_byp_restore_m), .Y(exu_n30259));
INVX1 exu_U30989(.A(exu_n30259), .Y(exu_n11116));
AND2X1 exu_U30990(.A(exu_tlu_wsr_data_m[14]), .B(ecl_byp_restore_m), .Y(exu_n30261));
INVX1 exu_U30991(.A(exu_n30261), .Y(exu_n11117));
AND2X1 exu_U30992(.A(exu_tlu_wsr_data_m[13]), .B(ecl_byp_restore_m), .Y(exu_n30263));
INVX1 exu_U30993(.A(exu_n30263), .Y(exu_n11118));
AND2X1 exu_U30994(.A(exu_tlu_wsr_data_m[12]), .B(ecl_byp_restore_m), .Y(exu_n30265));
INVX1 exu_U30995(.A(exu_n30265), .Y(exu_n11119));
AND2X1 exu_U30996(.A(exu_tlu_wsr_data_m[11]), .B(ecl_byp_restore_m), .Y(exu_n30267));
INVX1 exu_U30997(.A(exu_n30267), .Y(exu_n11120));
AND2X1 exu_U30998(.A(exu_tlu_wsr_data_m[10]), .B(ecl_byp_restore_m), .Y(exu_n30269));
INVX1 exu_U30999(.A(exu_n30269), .Y(exu_n11121));
AND2X1 exu_U31000(.A(exu_tlu_wsr_data_m[0]), .B(ecl_byp_restore_m), .Y(exu_n30271));
INVX1 exu_U31001(.A(exu_n30271), .Y(exu_n11122));
AND2X1 exu_U31002(.A(exu_n16164), .B(exu_spu_rs3_data_e[9]), .Y(exu_n30273));
INVX1 exu_U31003(.A(exu_n30273), .Y(exu_n11123));
AND2X1 exu_U31004(.A(exu_spu_rs3_data_e[8]), .B(exu_n16165), .Y(exu_n30275));
INVX1 exu_U31005(.A(exu_n30275), .Y(exu_n11124));
AND2X1 exu_U31006(.A(exu_spu_rs3_data_e[7]), .B(exu_n16165), .Y(exu_n30277));
INVX1 exu_U31007(.A(exu_n30277), .Y(exu_n11125));
AND2X1 exu_U31008(.A(exu_spu_rs3_data_e[6]), .B(exu_n16165), .Y(exu_n30279));
INVX1 exu_U31009(.A(exu_n30279), .Y(exu_n11126));
AND2X1 exu_U31010(.A(exu_spu_rs3_data_e[63]), .B(exu_n16165), .Y(exu_n30281));
INVX1 exu_U31011(.A(exu_n30281), .Y(exu_n11127));
AND2X1 exu_U31012(.A(exu_spu_rs3_data_e[62]), .B(exu_n16165), .Y(exu_n30283));
INVX1 exu_U31013(.A(exu_n30283), .Y(exu_n11128));
AND2X1 exu_U31014(.A(exu_spu_rs3_data_e[61]), .B(exu_n16165), .Y(exu_n30285));
INVX1 exu_U31015(.A(exu_n30285), .Y(exu_n11129));
AND2X1 exu_U31016(.A(exu_spu_rs3_data_e[60]), .B(exu_n16165), .Y(exu_n30287));
INVX1 exu_U31017(.A(exu_n30287), .Y(exu_n11130));
AND2X1 exu_U31018(.A(exu_spu_rs3_data_e[5]), .B(exu_n16165), .Y(exu_n30289));
INVX1 exu_U31019(.A(exu_n30289), .Y(exu_n11131));
AND2X1 exu_U31020(.A(exu_spu_rs3_data_e[59]), .B(exu_n16165), .Y(exu_n30291));
INVX1 exu_U31021(.A(exu_n30291), .Y(exu_n11132));
AND2X1 exu_U31022(.A(exu_spu_rs3_data_e[58]), .B(exu_n16165), .Y(exu_n30293));
INVX1 exu_U31023(.A(exu_n30293), .Y(exu_n11133));
AND2X1 exu_U31024(.A(exu_spu_rs3_data_e[57]), .B(ecl_std_e), .Y(exu_n30295));
INVX1 exu_U31025(.A(exu_n30295), .Y(exu_n11134));
AND2X1 exu_U31026(.A(exu_spu_rs3_data_e[56]), .B(ecl_std_e), .Y(exu_n30297));
INVX1 exu_U31027(.A(exu_n30297), .Y(exu_n11135));
AND2X1 exu_U31028(.A(exu_spu_rs3_data_e[55]), .B(ecl_std_e), .Y(exu_n30299));
INVX1 exu_U31029(.A(exu_n30299), .Y(exu_n11136));
AND2X1 exu_U31030(.A(exu_spu_rs3_data_e[54]), .B(ecl_std_e), .Y(exu_n30301));
INVX1 exu_U31031(.A(exu_n30301), .Y(exu_n11137));
AND2X1 exu_U31032(.A(exu_spu_rs3_data_e[53]), .B(exu_n16163), .Y(exu_n30303));
INVX1 exu_U31033(.A(exu_n30303), .Y(exu_n11138));
AND2X1 exu_U31034(.A(exu_spu_rs3_data_e[52]), .B(ecl_std_e), .Y(exu_n30305));
INVX1 exu_U31035(.A(exu_n30305), .Y(exu_n11139));
AND2X1 exu_U31036(.A(exu_spu_rs3_data_e[51]), .B(exu_n16163), .Y(exu_n30307));
INVX1 exu_U31037(.A(exu_n30307), .Y(exu_n11140));
AND2X1 exu_U31038(.A(exu_spu_rs3_data_e[50]), .B(ecl_std_e), .Y(exu_n30309));
INVX1 exu_U31039(.A(exu_n30309), .Y(exu_n11141));
AND2X1 exu_U31040(.A(exu_spu_rs3_data_e[4]), .B(exu_n16163), .Y(exu_n30311));
INVX1 exu_U31041(.A(exu_n30311), .Y(exu_n11142));
AND2X1 exu_U31042(.A(exu_spu_rs3_data_e[49]), .B(ecl_std_e), .Y(exu_n30313));
INVX1 exu_U31043(.A(exu_n30313), .Y(exu_n11143));
AND2X1 exu_U31044(.A(exu_spu_rs3_data_e[48]), .B(exu_n16163), .Y(exu_n30315));
INVX1 exu_U31045(.A(exu_n30315), .Y(exu_n11144));
AND2X1 exu_U31046(.A(exu_spu_rs3_data_e[47]), .B(ecl_std_e), .Y(exu_n30317));
INVX1 exu_U31047(.A(exu_n30317), .Y(exu_n11145));
AND2X1 exu_U31048(.A(exu_spu_rs3_data_e[46]), .B(exu_n16163), .Y(exu_n30319));
INVX1 exu_U31049(.A(exu_n30319), .Y(exu_n11146));
AND2X1 exu_U31050(.A(exu_spu_rs3_data_e[45]), .B(exu_n16166), .Y(exu_n30321));
INVX1 exu_U31051(.A(exu_n30321), .Y(exu_n11147));
AND2X1 exu_U31052(.A(exu_spu_rs3_data_e[44]), .B(exu_n16166), .Y(exu_n30323));
INVX1 exu_U31053(.A(exu_n30323), .Y(exu_n11148));
AND2X1 exu_U31054(.A(exu_spu_rs3_data_e[43]), .B(exu_n16166), .Y(exu_n30325));
INVX1 exu_U31055(.A(exu_n30325), .Y(exu_n11149));
AND2X1 exu_U31056(.A(exu_spu_rs3_data_e[42]), .B(exu_n16166), .Y(exu_n30327));
INVX1 exu_U31057(.A(exu_n30327), .Y(exu_n11150));
AND2X1 exu_U31058(.A(exu_spu_rs3_data_e[41]), .B(exu_n16166), .Y(exu_n30329));
INVX1 exu_U31059(.A(exu_n30329), .Y(exu_n11151));
AND2X1 exu_U31060(.A(exu_spu_rs3_data_e[40]), .B(exu_n16166), .Y(exu_n30331));
INVX1 exu_U31061(.A(exu_n30331), .Y(exu_n11152));
AND2X1 exu_U31062(.A(exu_spu_rs3_data_e[3]), .B(exu_n16166), .Y(exu_n30333));
INVX1 exu_U31063(.A(exu_n30333), .Y(exu_n11153));
AND2X1 exu_U31064(.A(exu_spu_rs3_data_e[39]), .B(exu_n16166), .Y(exu_n30335));
INVX1 exu_U31065(.A(exu_n30335), .Y(exu_n11154));
AND2X1 exu_U31066(.A(exu_spu_rs3_data_e[38]), .B(exu_n16166), .Y(exu_n30337));
INVX1 exu_U31067(.A(exu_n30337), .Y(exu_n11155));
AND2X1 exu_U31068(.A(exu_spu_rs3_data_e[37]), .B(exu_n16166), .Y(exu_n30339));
INVX1 exu_U31069(.A(exu_n30339), .Y(exu_n11156));
AND2X1 exu_U31070(.A(exu_spu_rs3_data_e[36]), .B(exu_n16166), .Y(exu_n30341));
INVX1 exu_U31071(.A(exu_n30341), .Y(exu_n11157));
AND2X1 exu_U31072(.A(exu_spu_rs3_data_e[35]), .B(exu_n16166), .Y(exu_n30343));
INVX1 exu_U31073(.A(exu_n30343), .Y(exu_n11158));
AND2X1 exu_U31074(.A(exu_spu_rs3_data_e[34]), .B(exu_n16166), .Y(exu_n30345));
INVX1 exu_U31075(.A(exu_n30345), .Y(exu_n11159));
AND2X1 exu_U31076(.A(exu_spu_rs3_data_e[33]), .B(exu_n16166), .Y(exu_n30347));
INVX1 exu_U31077(.A(exu_n30347), .Y(exu_n11160));
AND2X1 exu_U31078(.A(exu_spu_rs3_data_e[32]), .B(exu_n16166), .Y(exu_n30349));
INVX1 exu_U31079(.A(exu_n30349), .Y(exu_n11161));
AND2X1 exu_U31080(.A(exu_spu_rs3_data_e[31]), .B(exu_n16166), .Y(exu_n30351));
INVX1 exu_U31081(.A(exu_n30351), .Y(exu_n11162));
AND2X1 exu_U31082(.A(exu_spu_rs3_data_e[30]), .B(ecl_std_e), .Y(exu_n30353));
INVX1 exu_U31083(.A(exu_n30353), .Y(exu_n11163));
AND2X1 exu_U31084(.A(exu_spu_rs3_data_e[2]), .B(ecl_std_e), .Y(exu_n30355));
INVX1 exu_U31085(.A(exu_n30355), .Y(exu_n11164));
AND2X1 exu_U31086(.A(exu_spu_rs3_data_e[29]), .B(ecl_std_e), .Y(exu_n30357));
INVX1 exu_U31087(.A(exu_n30357), .Y(exu_n11165));
AND2X1 exu_U31088(.A(exu_spu_rs3_data_e[28]), .B(ecl_std_e), .Y(exu_n30359));
INVX1 exu_U31089(.A(exu_n30359), .Y(exu_n11166));
AND2X1 exu_U31090(.A(exu_spu_rs3_data_e[27]), .B(exu_n16165), .Y(exu_n30361));
INVX1 exu_U31091(.A(exu_n30361), .Y(exu_n11167));
AND2X1 exu_U31092(.A(exu_spu_rs3_data_e[26]), .B(ecl_std_e), .Y(exu_n30363));
INVX1 exu_U31093(.A(exu_n30363), .Y(exu_n11168));
AND2X1 exu_U31094(.A(exu_spu_rs3_data_e[25]), .B(exu_n16162), .Y(exu_n30365));
INVX1 exu_U31095(.A(exu_n30365), .Y(exu_n11169));
AND2X1 exu_U31096(.A(exu_spu_rs3_data_e[24]), .B(ecl_std_e), .Y(exu_n30367));
INVX1 exu_U31097(.A(exu_n30367), .Y(exu_n11170));
AND2X1 exu_U31098(.A(exu_spu_rs3_data_e[23]), .B(exu_n16163), .Y(exu_n30369));
INVX1 exu_U31099(.A(exu_n30369), .Y(exu_n11171));
AND2X1 exu_U31100(.A(exu_spu_rs3_data_e[22]), .B(exu_n16164), .Y(exu_n30371));
INVX1 exu_U31101(.A(exu_n30371), .Y(exu_n11172));
AND2X1 exu_U31102(.A(exu_spu_rs3_data_e[21]), .B(exu_n16165), .Y(exu_n30373));
INVX1 exu_U31103(.A(exu_n30373), .Y(exu_n11173));
AND2X1 exu_U31104(.A(exu_spu_rs3_data_e[20]), .B(exu_n16163), .Y(exu_n30375));
INVX1 exu_U31105(.A(exu_n30375), .Y(exu_n11174));
AND2X1 exu_U31106(.A(exu_spu_rs3_data_e[1]), .B(exu_n16166), .Y(exu_n30377));
INVX1 exu_U31107(.A(exu_n30377), .Y(exu_n11175));
AND2X1 exu_U31108(.A(exu_spu_rs3_data_e[19]), .B(ecl_std_e), .Y(exu_n30379));
INVX1 exu_U31109(.A(exu_n30379), .Y(exu_n11176));
AND2X1 exu_U31110(.A(exu_spu_rs3_data_e[18]), .B(exu_n16162), .Y(exu_n30381));
INVX1 exu_U31111(.A(exu_n30381), .Y(exu_n11177));
AND2X1 exu_U31112(.A(exu_spu_rs3_data_e[17]), .B(ecl_std_e), .Y(exu_n30383));
INVX1 exu_U31113(.A(exu_n30383), .Y(exu_n11178));
AND2X1 exu_U31114(.A(exu_spu_rs3_data_e[16]), .B(exu_n16162), .Y(exu_n30385));
INVX1 exu_U31115(.A(exu_n30385), .Y(exu_n11179));
AND2X1 exu_U31116(.A(exu_spu_rs3_data_e[15]), .B(ecl_std_e), .Y(exu_n30387));
INVX1 exu_U31117(.A(exu_n30387), .Y(exu_n11180));
AND2X1 exu_U31118(.A(exu_spu_rs3_data_e[14]), .B(exu_n16163), .Y(exu_n30389));
INVX1 exu_U31119(.A(exu_n30389), .Y(exu_n11181));
AND2X1 exu_U31120(.A(exu_spu_rs3_data_e[13]), .B(exu_n16166), .Y(exu_n30391));
INVX1 exu_U31121(.A(exu_n30391), .Y(exu_n11182));
AND2X1 exu_U31122(.A(exu_spu_rs3_data_e[12]), .B(exu_n16162), .Y(exu_n30393));
INVX1 exu_U31123(.A(exu_n30393), .Y(exu_n11183));
AND2X1 exu_U31124(.A(exu_spu_rs3_data_e[11]), .B(exu_n16162), .Y(exu_n30395));
INVX1 exu_U31125(.A(exu_n30395), .Y(exu_n11184));
AND2X1 exu_U31126(.A(exu_spu_rs3_data_e[10]), .B(exu_n16164), .Y(exu_n30397));
INVX1 exu_U31127(.A(exu_n30397), .Y(exu_n11185));
AND2X1 exu_U31128(.A(exu_spu_rs3_data_e[0]), .B(exu_n16163), .Y(exu_n30399));
INVX1 exu_U31129(.A(exu_n30399), .Y(exu_n11186));
AND2X1 exu_U31130(.A(ecl_alu_casa_e), .B(alu_logic_rs1_data_bf1[9]), .Y(exu_n30497));
INVX1 exu_U31131(.A(exu_n30497), .Y(exu_n11187));
AND2X1 exu_U31132(.A(alu_logic_rs1_data_bf1[8]), .B(ecl_alu_casa_e), .Y(exu_n30499));
INVX1 exu_U31133(.A(exu_n30499), .Y(exu_n11188));
AND2X1 exu_U31134(.A(alu_logic_rs1_data_bf1[7]), .B(ecl_alu_casa_e), .Y(exu_n30501));
INVX1 exu_U31135(.A(exu_n30501), .Y(exu_n11189));
AND2X1 exu_U31136(.A(alu_logic_rs1_data_bf1[6]), .B(ecl_alu_casa_e), .Y(exu_n30503));
INVX1 exu_U31137(.A(exu_n30503), .Y(exu_n11190));
AND2X1 exu_U31138(.A(alu_logic_rs1_data_bf1[5]), .B(ecl_alu_casa_e), .Y(exu_n30513));
INVX1 exu_U31139(.A(exu_n30513), .Y(exu_n11191));
AND2X1 exu_U31140(.A(alu_logic_rs1_data_bf1[4]), .B(ecl_alu_casa_e), .Y(exu_n30535));
INVX1 exu_U31141(.A(exu_n30535), .Y(exu_n11192));
AND2X1 exu_U31142(.A(alu_logic_rs1_data_bf1[46]), .B(ecl_alu_casa_e), .Y(exu_n30543));
INVX1 exu_U31143(.A(exu_n30543), .Y(exu_n11193));
AND2X1 exu_U31144(.A(alu_logic_rs1_data_bf1[45]), .B(ecl_alu_casa_e), .Y(exu_n30545));
INVX1 exu_U31145(.A(exu_n30545), .Y(exu_n11194));
AND2X1 exu_U31146(.A(alu_logic_rs1_data_bf1[44]), .B(ecl_alu_casa_e), .Y(exu_n30547));
INVX1 exu_U31147(.A(exu_n30547), .Y(exu_n11195));
AND2X1 exu_U31148(.A(alu_logic_rs1_data_bf1[43]), .B(ecl_alu_casa_e), .Y(exu_n30549));
INVX1 exu_U31149(.A(exu_n30549), .Y(exu_n11196));
AND2X1 exu_U31150(.A(alu_logic_rs1_data_bf1[42]), .B(ecl_alu_casa_e), .Y(exu_n30551));
INVX1 exu_U31151(.A(exu_n30551), .Y(exu_n11197));
AND2X1 exu_U31152(.A(alu_logic_rs1_data_bf1[41]), .B(ecl_alu_casa_e), .Y(exu_n30553));
INVX1 exu_U31153(.A(exu_n30553), .Y(exu_n11198));
AND2X1 exu_U31154(.A(alu_logic_rs1_data_bf1[40]), .B(ecl_alu_casa_e), .Y(exu_n30555));
INVX1 exu_U31155(.A(exu_n30555), .Y(exu_n11199));
AND2X1 exu_U31156(.A(alu_logic_rs1_data_bf1[3]), .B(ecl_alu_casa_e), .Y(exu_n30557));
INVX1 exu_U31157(.A(exu_n30557), .Y(exu_n11200));
AND2X1 exu_U31158(.A(alu_logic_rs1_data_bf1[39]), .B(ecl_alu_casa_e), .Y(exu_n30559));
INVX1 exu_U31159(.A(exu_n30559), .Y(exu_n11201));
AND2X1 exu_U31160(.A(alu_logic_rs1_data_bf1[38]), .B(ecl_alu_casa_e), .Y(exu_n30561));
INVX1 exu_U31161(.A(exu_n30561), .Y(exu_n11202));
AND2X1 exu_U31162(.A(alu_logic_rs1_data_bf1[37]), .B(ecl_alu_casa_e), .Y(exu_n30563));
INVX1 exu_U31163(.A(exu_n30563), .Y(exu_n11203));
AND2X1 exu_U31164(.A(alu_logic_rs1_data_bf1[36]), .B(ecl_alu_casa_e), .Y(exu_n30565));
INVX1 exu_U31165(.A(exu_n30565), .Y(exu_n11204));
AND2X1 exu_U31166(.A(alu_logic_rs1_data_bf1[35]), .B(ecl_alu_casa_e), .Y(exu_n30567));
INVX1 exu_U31167(.A(exu_n30567), .Y(exu_n11205));
AND2X1 exu_U31168(.A(alu_logic_rs1_data_bf1[34]), .B(ecl_alu_casa_e), .Y(exu_n30569));
INVX1 exu_U31169(.A(exu_n30569), .Y(exu_n11206));
AND2X1 exu_U31170(.A(alu_logic_rs1_data_bf1[33]), .B(ecl_alu_casa_e), .Y(exu_n30571));
INVX1 exu_U31171(.A(exu_n30571), .Y(exu_n11207));
AND2X1 exu_U31172(.A(alu_logic_rs1_data_bf1[32]), .B(ecl_alu_casa_e), .Y(exu_n30573));
INVX1 exu_U31173(.A(exu_n30573), .Y(exu_n11208));
AND2X1 exu_U31174(.A(alu_logic_rs1_data_bf1[31]), .B(ecl_alu_casa_e), .Y(exu_n30575));
INVX1 exu_U31175(.A(exu_n30575), .Y(exu_n11209));
AND2X1 exu_U31176(.A(alu_logic_rs1_data_bf1[30]), .B(ecl_alu_casa_e), .Y(exu_n30577));
INVX1 exu_U31177(.A(exu_n30577), .Y(exu_n11210));
AND2X1 exu_U31178(.A(alu_logic_rs1_data_bf1[2]), .B(ecl_alu_casa_e), .Y(exu_n30579));
INVX1 exu_U31179(.A(exu_n30579), .Y(exu_n11211));
AND2X1 exu_U31180(.A(alu_logic_rs1_data_bf1[29]), .B(ecl_alu_casa_e), .Y(exu_n30581));
INVX1 exu_U31181(.A(exu_n30581), .Y(exu_n11212));
AND2X1 exu_U31182(.A(alu_logic_rs1_data_bf1[28]), .B(ecl_alu_casa_e), .Y(exu_n30583));
INVX1 exu_U31183(.A(exu_n30583), .Y(exu_n11213));
AND2X1 exu_U31184(.A(alu_logic_rs1_data_bf1[27]), .B(ecl_alu_casa_e), .Y(exu_n30585));
INVX1 exu_U31185(.A(exu_n30585), .Y(exu_n11214));
AND2X1 exu_U31186(.A(alu_logic_rs1_data_bf1[26]), .B(ecl_alu_casa_e), .Y(exu_n30587));
INVX1 exu_U31187(.A(exu_n30587), .Y(exu_n11215));
AND2X1 exu_U31188(.A(alu_logic_rs1_data_bf1[25]), .B(ecl_alu_casa_e), .Y(exu_n30589));
INVX1 exu_U31189(.A(exu_n30589), .Y(exu_n11216));
AND2X1 exu_U31190(.A(alu_logic_rs1_data_bf1[24]), .B(ecl_alu_casa_e), .Y(exu_n30591));
INVX1 exu_U31191(.A(exu_n30591), .Y(exu_n11217));
AND2X1 exu_U31192(.A(alu_logic_rs1_data_bf1[23]), .B(ecl_alu_casa_e), .Y(exu_n30593));
INVX1 exu_U31193(.A(exu_n30593), .Y(exu_n11218));
AND2X1 exu_U31194(.A(alu_logic_rs1_data_bf1[22]), .B(ecl_alu_casa_e), .Y(exu_n30595));
INVX1 exu_U31195(.A(exu_n30595), .Y(exu_n11219));
AND2X1 exu_U31196(.A(alu_logic_rs1_data_bf1[21]), .B(ecl_alu_casa_e), .Y(exu_n30597));
INVX1 exu_U31197(.A(exu_n30597), .Y(exu_n11220));
AND2X1 exu_U31198(.A(alu_logic_rs1_data_bf1[20]), .B(ecl_alu_casa_e), .Y(exu_n30599));
INVX1 exu_U31199(.A(exu_n30599), .Y(exu_n11221));
AND2X1 exu_U31200(.A(alu_logic_rs1_data_bf1[1]), .B(ecl_alu_casa_e), .Y(exu_n30601));
INVX1 exu_U31201(.A(exu_n30601), .Y(exu_n11222));
AND2X1 exu_U31202(.A(alu_logic_rs1_data_bf1[19]), .B(ecl_alu_casa_e), .Y(exu_n30603));
INVX1 exu_U31203(.A(exu_n30603), .Y(exu_n11223));
AND2X1 exu_U31204(.A(alu_logic_rs1_data_bf1[18]), .B(ecl_alu_casa_e), .Y(exu_n30605));
INVX1 exu_U31205(.A(exu_n30605), .Y(exu_n11224));
AND2X1 exu_U31206(.A(alu_logic_rs1_data_bf1[17]), .B(ecl_alu_casa_e), .Y(exu_n30607));
INVX1 exu_U31207(.A(exu_n30607), .Y(exu_n11225));
AND2X1 exu_U31208(.A(alu_logic_rs1_data_bf1[16]), .B(ecl_alu_casa_e), .Y(exu_n30609));
INVX1 exu_U31209(.A(exu_n30609), .Y(exu_n11226));
AND2X1 exu_U31210(.A(alu_logic_rs1_data_bf1[15]), .B(ecl_alu_casa_e), .Y(exu_n30611));
INVX1 exu_U31211(.A(exu_n30611), .Y(exu_n11227));
AND2X1 exu_U31212(.A(alu_logic_rs1_data_bf1[14]), .B(ecl_alu_casa_e), .Y(exu_n30613));
INVX1 exu_U31213(.A(exu_n30613), .Y(exu_n11228));
AND2X1 exu_U31214(.A(alu_logic_rs1_data_bf1[13]), .B(ecl_alu_casa_e), .Y(exu_n30615));
INVX1 exu_U31215(.A(exu_n30615), .Y(exu_n11229));
AND2X1 exu_U31216(.A(alu_logic_rs1_data_bf1[12]), .B(ecl_alu_casa_e), .Y(exu_n30617));
INVX1 exu_U31217(.A(exu_n30617), .Y(exu_n11230));
AND2X1 exu_U31218(.A(alu_logic_rs1_data_bf1[11]), .B(ecl_alu_casa_e), .Y(exu_n30619));
INVX1 exu_U31219(.A(exu_n30619), .Y(exu_n11231));
AND2X1 exu_U31220(.A(alu_logic_rs1_data_bf1[10]), .B(ecl_alu_casa_e), .Y(exu_n30621));
INVX1 exu_U31221(.A(exu_n30621), .Y(exu_n11232));
AND2X1 exu_U31222(.A(alu_logic_rs1_data_bf1[0]), .B(ecl_alu_casa_e), .Y(exu_n30623));
INVX1 exu_U31223(.A(exu_n30623), .Y(exu_n11233));
AND2X1 exu_U31224(.A(ecl_shft_lshift_e_l), .B(shft_rshift1[9]), .Y(exu_n30753));
INVX1 exu_U31225(.A(exu_n30753), .Y(exu_n11234));
INVX1 exu_U31226(.A(shft_alu_shift_out_e[8]), .Y(exu_n11235));
AND2X1 exu_U31227(.A(shft_rshift1[8]), .B(ecl_shft_lshift_e_l), .Y(exu_n30755));
INVX1 exu_U31228(.A(exu_n30755), .Y(exu_n11236));
INVX1 exu_U31229(.A(shft_alu_shift_out_e[7]), .Y(exu_n11237));
AND2X1 exu_U31230(.A(shft_rshift1[7]), .B(ecl_shft_lshift_e_l), .Y(exu_n30757));
INVX1 exu_U31231(.A(exu_n30757), .Y(exu_n11238));
INVX1 exu_U31232(.A(shft_alu_shift_out_e[6]), .Y(exu_n11239));
AND2X1 exu_U31233(.A(shft_rshift1[6]), .B(ecl_shft_lshift_e_l), .Y(exu_n30759));
INVX1 exu_U31234(.A(exu_n30759), .Y(exu_n11240));
INVX1 exu_U31235(.A(shft_alu_shift_out_e[63]), .Y(exu_n11241));
AND2X1 exu_U31236(.A(shft_rshift1[63]), .B(ecl_shft_lshift_e_l), .Y(exu_n30761));
INVX1 exu_U31237(.A(exu_n30761), .Y(exu_n11242));
INVX1 exu_U31238(.A(shft_alu_shift_out_e[62]), .Y(exu_n11243));
AND2X1 exu_U31239(.A(shft_rshift1[62]), .B(ecl_shft_lshift_e_l), .Y(exu_n30763));
INVX1 exu_U31240(.A(exu_n30763), .Y(exu_n11244));
INVX1 exu_U31241(.A(shft_alu_shift_out_e[61]), .Y(exu_n11245));
AND2X1 exu_U31242(.A(shft_rshift1[61]), .B(ecl_shft_lshift_e_l), .Y(exu_n30765));
INVX1 exu_U31243(.A(exu_n30765), .Y(exu_n11246));
INVX1 exu_U31244(.A(shft_alu_shift_out_e[60]), .Y(exu_n11247));
AND2X1 exu_U31245(.A(shft_rshift1[60]), .B(ecl_shft_lshift_e_l), .Y(exu_n30767));
INVX1 exu_U31246(.A(exu_n30767), .Y(exu_n11248));
INVX1 exu_U31247(.A(shft_alu_shift_out_e[5]), .Y(exu_n11249));
AND2X1 exu_U31248(.A(shft_rshift1[5]), .B(ecl_shft_lshift_e_l), .Y(exu_n30769));
INVX1 exu_U31249(.A(exu_n30769), .Y(exu_n11250));
INVX1 exu_U31250(.A(shft_alu_shift_out_e[59]), .Y(exu_n11251));
AND2X1 exu_U31251(.A(shft_rshift1[59]), .B(ecl_shft_lshift_e_l), .Y(exu_n30771));
INVX1 exu_U31252(.A(exu_n30771), .Y(exu_n11252));
INVX1 exu_U31253(.A(shft_alu_shift_out_e[58]), .Y(exu_n11253));
AND2X1 exu_U31254(.A(shft_rshift1[58]), .B(ecl_shft_lshift_e_l), .Y(exu_n30773));
INVX1 exu_U31255(.A(exu_n30773), .Y(exu_n11254));
INVX1 exu_U31256(.A(shft_alu_shift_out_e[57]), .Y(exu_n11255));
AND2X1 exu_U31257(.A(shft_rshift1[57]), .B(ecl_shft_lshift_e_l), .Y(exu_n30775));
INVX1 exu_U31258(.A(exu_n30775), .Y(exu_n11256));
INVX1 exu_U31259(.A(shft_alu_shift_out_e[56]), .Y(exu_n11257));
AND2X1 exu_U31260(.A(shft_rshift1[56]), .B(ecl_shft_lshift_e_l), .Y(exu_n30777));
INVX1 exu_U31261(.A(exu_n30777), .Y(exu_n11258));
INVX1 exu_U31262(.A(shft_alu_shift_out_e[55]), .Y(exu_n11259));
AND2X1 exu_U31263(.A(shft_rshift1[55]), .B(ecl_shft_lshift_e_l), .Y(exu_n30779));
INVX1 exu_U31264(.A(exu_n30779), .Y(exu_n11260));
INVX1 exu_U31265(.A(shft_alu_shift_out_e[54]), .Y(exu_n11261));
AND2X1 exu_U31266(.A(shft_rshift1[54]), .B(ecl_shft_lshift_e_l), .Y(exu_n30781));
INVX1 exu_U31267(.A(exu_n30781), .Y(exu_n11262));
INVX1 exu_U31268(.A(shft_alu_shift_out_e[53]), .Y(exu_n11263));
AND2X1 exu_U31269(.A(shft_rshift1[53]), .B(ecl_shft_lshift_e_l), .Y(exu_n30783));
INVX1 exu_U31270(.A(exu_n30783), .Y(exu_n11264));
INVX1 exu_U31271(.A(shft_alu_shift_out_e[52]), .Y(exu_n11265));
AND2X1 exu_U31272(.A(shft_rshift1[52]), .B(ecl_shft_lshift_e_l), .Y(exu_n30785));
INVX1 exu_U31273(.A(exu_n30785), .Y(exu_n11266));
INVX1 exu_U31274(.A(shft_alu_shift_out_e[51]), .Y(exu_n11267));
AND2X1 exu_U31275(.A(shft_rshift1[51]), .B(ecl_shft_lshift_e_l), .Y(exu_n30787));
INVX1 exu_U31276(.A(exu_n30787), .Y(exu_n11268));
INVX1 exu_U31277(.A(shft_alu_shift_out_e[50]), .Y(exu_n11269));
AND2X1 exu_U31278(.A(shft_rshift1[50]), .B(ecl_shft_lshift_e_l), .Y(exu_n30789));
INVX1 exu_U31279(.A(exu_n30789), .Y(exu_n11270));
INVX1 exu_U31280(.A(shft_alu_shift_out_e[4]), .Y(exu_n11271));
AND2X1 exu_U31281(.A(shft_rshift1[4]), .B(ecl_shft_lshift_e_l), .Y(exu_n30791));
INVX1 exu_U31282(.A(exu_n30791), .Y(exu_n11272));
INVX1 exu_U31283(.A(shft_alu_shift_out_e[49]), .Y(exu_n11273));
AND2X1 exu_U31284(.A(shft_rshift1[49]), .B(ecl_shft_lshift_e_l), .Y(exu_n30793));
INVX1 exu_U31285(.A(exu_n30793), .Y(exu_n11274));
INVX1 exu_U31286(.A(shft_alu_shift_out_e[48]), .Y(exu_n11275));
AND2X1 exu_U31287(.A(shft_rshift1[48]), .B(ecl_shft_lshift_e_l), .Y(exu_n30795));
INVX1 exu_U31288(.A(exu_n30795), .Y(exu_n11276));
INVX1 exu_U31289(.A(shft_alu_shift_out_e[47]), .Y(exu_n11277));
AND2X1 exu_U31290(.A(shft_rshift1[47]), .B(ecl_shft_lshift_e_l), .Y(exu_n30797));
INVX1 exu_U31291(.A(exu_n30797), .Y(exu_n11278));
INVX1 exu_U31292(.A(shft_alu_shift_out_e[46]), .Y(exu_n11279));
AND2X1 exu_U31293(.A(shft_rshift1[46]), .B(ecl_shft_lshift_e_l), .Y(exu_n30799));
INVX1 exu_U31294(.A(exu_n30799), .Y(exu_n11280));
INVX1 exu_U31295(.A(shft_alu_shift_out_e[45]), .Y(exu_n11281));
AND2X1 exu_U31296(.A(shft_rshift1[45]), .B(ecl_shft_lshift_e_l), .Y(exu_n30801));
INVX1 exu_U31297(.A(exu_n30801), .Y(exu_n11282));
INVX1 exu_U31298(.A(shft_alu_shift_out_e[44]), .Y(exu_n11283));
AND2X1 exu_U31299(.A(shft_rshift1[44]), .B(ecl_shft_lshift_e_l), .Y(exu_n30803));
INVX1 exu_U31300(.A(exu_n30803), .Y(exu_n11284));
INVX1 exu_U31301(.A(shft_alu_shift_out_e[43]), .Y(exu_n11285));
AND2X1 exu_U31302(.A(shft_rshift1[43]), .B(ecl_shft_lshift_e_l), .Y(exu_n30805));
INVX1 exu_U31303(.A(exu_n30805), .Y(exu_n11286));
INVX1 exu_U31304(.A(shft_alu_shift_out_e[42]), .Y(exu_n11287));
AND2X1 exu_U31305(.A(shft_rshift1[42]), .B(ecl_shft_lshift_e_l), .Y(exu_n30807));
INVX1 exu_U31306(.A(exu_n30807), .Y(exu_n11288));
INVX1 exu_U31307(.A(shft_alu_shift_out_e[41]), .Y(exu_n11289));
AND2X1 exu_U31308(.A(shft_rshift1[41]), .B(ecl_shft_lshift_e_l), .Y(exu_n30809));
INVX1 exu_U31309(.A(exu_n30809), .Y(exu_n11290));
INVX1 exu_U31310(.A(shft_alu_shift_out_e[40]), .Y(exu_n11291));
AND2X1 exu_U31311(.A(shft_rshift1[40]), .B(ecl_shft_lshift_e_l), .Y(exu_n30811));
INVX1 exu_U31312(.A(exu_n30811), .Y(exu_n11292));
INVX1 exu_U31313(.A(shft_alu_shift_out_e[3]), .Y(exu_n11293));
AND2X1 exu_U31314(.A(shft_rshift1[3]), .B(ecl_shft_lshift_e_l), .Y(exu_n30813));
INVX1 exu_U31315(.A(exu_n30813), .Y(exu_n11294));
INVX1 exu_U31316(.A(shft_alu_shift_out_e[39]), .Y(exu_n11295));
AND2X1 exu_U31317(.A(shft_rshift1[39]), .B(ecl_shft_lshift_e_l), .Y(exu_n30815));
INVX1 exu_U31318(.A(exu_n30815), .Y(exu_n11296));
INVX1 exu_U31319(.A(shft_alu_shift_out_e[38]), .Y(exu_n11297));
AND2X1 exu_U31320(.A(shft_rshift1[38]), .B(ecl_shft_lshift_e_l), .Y(exu_n30817));
INVX1 exu_U31321(.A(exu_n30817), .Y(exu_n11298));
INVX1 exu_U31322(.A(shft_alu_shift_out_e[37]), .Y(exu_n11299));
AND2X1 exu_U31323(.A(shft_rshift1[37]), .B(ecl_shft_lshift_e_l), .Y(exu_n30819));
INVX1 exu_U31324(.A(exu_n30819), .Y(exu_n11300));
INVX1 exu_U31325(.A(shft_alu_shift_out_e[36]), .Y(exu_n11301));
AND2X1 exu_U31326(.A(shft_rshift1[36]), .B(ecl_shft_lshift_e_l), .Y(exu_n30821));
INVX1 exu_U31327(.A(exu_n30821), .Y(exu_n11302));
INVX1 exu_U31328(.A(shft_alu_shift_out_e[35]), .Y(exu_n11303));
AND2X1 exu_U31329(.A(shft_rshift1[35]), .B(ecl_shft_lshift_e_l), .Y(exu_n30823));
INVX1 exu_U31330(.A(exu_n30823), .Y(exu_n11304));
INVX1 exu_U31331(.A(shft_alu_shift_out_e[34]), .Y(exu_n11305));
AND2X1 exu_U31332(.A(shft_rshift1[34]), .B(ecl_shft_lshift_e_l), .Y(exu_n30825));
INVX1 exu_U31333(.A(exu_n30825), .Y(exu_n11306));
INVX1 exu_U31334(.A(shft_alu_shift_out_e[33]), .Y(exu_n11307));
AND2X1 exu_U31335(.A(shft_rshift1[33]), .B(ecl_shft_lshift_e_l), .Y(exu_n30827));
INVX1 exu_U31336(.A(exu_n30827), .Y(exu_n11308));
INVX1 exu_U31337(.A(shft_alu_shift_out_e[32]), .Y(exu_n11309));
AND2X1 exu_U31338(.A(shft_rshift1[32]), .B(ecl_shft_lshift_e_l), .Y(exu_n30829));
INVX1 exu_U31339(.A(exu_n30829), .Y(exu_n11310));
INVX1 exu_U31340(.A(shft_alu_shift_out_e[31]), .Y(exu_n11311));
AND2X1 exu_U31341(.A(shft_rshift1[31]), .B(ecl_shft_lshift_e_l), .Y(exu_n30831));
INVX1 exu_U31342(.A(exu_n30831), .Y(exu_n11312));
INVX1 exu_U31343(.A(shft_alu_shift_out_e[30]), .Y(exu_n11313));
AND2X1 exu_U31344(.A(shft_rshift1[30]), .B(ecl_shft_lshift_e_l), .Y(exu_n30833));
INVX1 exu_U31345(.A(exu_n30833), .Y(exu_n11314));
INVX1 exu_U31346(.A(shft_alu_shift_out_e[2]), .Y(exu_n11315));
AND2X1 exu_U31347(.A(shft_rshift1[2]), .B(ecl_shft_lshift_e_l), .Y(exu_n30835));
INVX1 exu_U31348(.A(exu_n30835), .Y(exu_n11316));
INVX1 exu_U31349(.A(shft_alu_shift_out_e[29]), .Y(exu_n11317));
AND2X1 exu_U31350(.A(shft_rshift1[29]), .B(ecl_shft_lshift_e_l), .Y(exu_n30837));
INVX1 exu_U31351(.A(exu_n30837), .Y(exu_n11318));
INVX1 exu_U31352(.A(shft_alu_shift_out_e[28]), .Y(exu_n11319));
AND2X1 exu_U31353(.A(shft_rshift1[28]), .B(ecl_shft_lshift_e_l), .Y(exu_n30839));
INVX1 exu_U31354(.A(exu_n30839), .Y(exu_n11320));
INVX1 exu_U31355(.A(shft_alu_shift_out_e[27]), .Y(exu_n11321));
AND2X1 exu_U31356(.A(shft_rshift1[27]), .B(ecl_shft_lshift_e_l), .Y(exu_n30841));
INVX1 exu_U31357(.A(exu_n30841), .Y(exu_n11322));
INVX1 exu_U31358(.A(shft_alu_shift_out_e[26]), .Y(exu_n11323));
AND2X1 exu_U31359(.A(shft_rshift1[26]), .B(ecl_shft_lshift_e_l), .Y(exu_n30843));
INVX1 exu_U31360(.A(exu_n30843), .Y(exu_n11324));
INVX1 exu_U31361(.A(shft_alu_shift_out_e[25]), .Y(exu_n11325));
AND2X1 exu_U31362(.A(shft_rshift1[25]), .B(ecl_shft_lshift_e_l), .Y(exu_n30845));
INVX1 exu_U31363(.A(exu_n30845), .Y(exu_n11326));
INVX1 exu_U31364(.A(shft_alu_shift_out_e[24]), .Y(exu_n11327));
AND2X1 exu_U31365(.A(shft_rshift1[24]), .B(ecl_shft_lshift_e_l), .Y(exu_n30847));
INVX1 exu_U31366(.A(exu_n30847), .Y(exu_n11328));
INVX1 exu_U31367(.A(shft_alu_shift_out_e[23]), .Y(exu_n11329));
AND2X1 exu_U31368(.A(shft_rshift1[23]), .B(ecl_shft_lshift_e_l), .Y(exu_n30849));
INVX1 exu_U31369(.A(exu_n30849), .Y(exu_n11330));
INVX1 exu_U31370(.A(shft_alu_shift_out_e[22]), .Y(exu_n11331));
AND2X1 exu_U31371(.A(shft_rshift1[22]), .B(ecl_shft_lshift_e_l), .Y(exu_n30851));
INVX1 exu_U31372(.A(exu_n30851), .Y(exu_n11332));
INVX1 exu_U31373(.A(shft_alu_shift_out_e[21]), .Y(exu_n11333));
AND2X1 exu_U31374(.A(shft_rshift1[21]), .B(ecl_shft_lshift_e_l), .Y(exu_n30853));
INVX1 exu_U31375(.A(exu_n30853), .Y(exu_n11334));
INVX1 exu_U31376(.A(shft_alu_shift_out_e[20]), .Y(exu_n11335));
AND2X1 exu_U31377(.A(shft_rshift1[20]), .B(ecl_shft_lshift_e_l), .Y(exu_n30855));
INVX1 exu_U31378(.A(exu_n30855), .Y(exu_n11336));
INVX1 exu_U31379(.A(shft_alu_shift_out_e[1]), .Y(exu_n11337));
AND2X1 exu_U31380(.A(shft_rshift1[1]), .B(ecl_shft_lshift_e_l), .Y(exu_n30857));
INVX1 exu_U31381(.A(exu_n30857), .Y(exu_n11338));
INVX1 exu_U31382(.A(shft_alu_shift_out_e[19]), .Y(exu_n11339));
AND2X1 exu_U31383(.A(shft_rshift1[19]), .B(ecl_shft_lshift_e_l), .Y(exu_n30859));
INVX1 exu_U31384(.A(exu_n30859), .Y(exu_n11340));
INVX1 exu_U31385(.A(shft_alu_shift_out_e[18]), .Y(exu_n11341));
AND2X1 exu_U31386(.A(shft_rshift1[18]), .B(ecl_shft_lshift_e_l), .Y(exu_n30861));
INVX1 exu_U31387(.A(exu_n30861), .Y(exu_n11342));
INVX1 exu_U31388(.A(shft_alu_shift_out_e[17]), .Y(exu_n11343));
AND2X1 exu_U31389(.A(shft_rshift1[17]), .B(ecl_shft_lshift_e_l), .Y(exu_n30863));
INVX1 exu_U31390(.A(exu_n30863), .Y(exu_n11344));
INVX1 exu_U31391(.A(shft_alu_shift_out_e[16]), .Y(exu_n11345));
AND2X1 exu_U31392(.A(shft_rshift1[16]), .B(ecl_shft_lshift_e_l), .Y(exu_n30865));
INVX1 exu_U31393(.A(exu_n30865), .Y(exu_n11346));
INVX1 exu_U31394(.A(shft_alu_shift_out_e[15]), .Y(exu_n11347));
AND2X1 exu_U31395(.A(shft_rshift1[15]), .B(ecl_shft_lshift_e_l), .Y(exu_n30867));
INVX1 exu_U31396(.A(exu_n30867), .Y(exu_n11348));
INVX1 exu_U31397(.A(shft_alu_shift_out_e[14]), .Y(exu_n11349));
AND2X1 exu_U31398(.A(shft_rshift1[14]), .B(ecl_shft_lshift_e_l), .Y(exu_n30869));
INVX1 exu_U31399(.A(exu_n30869), .Y(exu_n11350));
INVX1 exu_U31400(.A(shft_alu_shift_out_e[13]), .Y(exu_n11351));
AND2X1 exu_U31401(.A(shft_rshift1[13]), .B(ecl_shft_lshift_e_l), .Y(exu_n30871));
INVX1 exu_U31402(.A(exu_n30871), .Y(exu_n11352));
INVX1 exu_U31403(.A(shft_alu_shift_out_e[12]), .Y(exu_n11353));
AND2X1 exu_U31404(.A(shft_rshift1[12]), .B(ecl_shft_lshift_e_l), .Y(exu_n30873));
INVX1 exu_U31405(.A(exu_n30873), .Y(exu_n11354));
INVX1 exu_U31406(.A(shft_alu_shift_out_e[11]), .Y(exu_n11355));
AND2X1 exu_U31407(.A(shft_rshift1[11]), .B(ecl_shft_lshift_e_l), .Y(exu_n30875));
INVX1 exu_U31408(.A(exu_n30875), .Y(exu_n11356));
INVX1 exu_U31409(.A(shft_alu_shift_out_e[10]), .Y(exu_n11357));
AND2X1 exu_U31410(.A(shft_rshift1[10]), .B(ecl_shft_lshift_e_l), .Y(exu_n30877));
INVX1 exu_U31411(.A(exu_n30877), .Y(exu_n11358));
INVX1 exu_U31412(.A(shft_alu_shift_out_e[0]), .Y(exu_n11359));
AND2X1 exu_U31413(.A(shft_rshift1[0]), .B(ecl_shft_lshift_e_l), .Y(exu_n30879));
INVX1 exu_U31414(.A(exu_n30879), .Y(exu_n11360));
AND2X1 exu_U31415(.A(exu_n16197), .B(div_d[9]), .Y(exu_n30881));
INVX1 exu_U31416(.A(exu_n30881), .Y(exu_n11361));
INVX1 exu_U31417(.A(div_byp_muldivout_g[8]), .Y(exu_n11362));
AND2X1 exu_U31418(.A(div_d[8]), .B(exu_n16197), .Y(exu_n30883));
INVX1 exu_U31419(.A(exu_n30883), .Y(exu_n11363));
INVX1 exu_U31420(.A(div_byp_muldivout_g[7]), .Y(exu_n11364));
AND2X1 exu_U31421(.A(div_d[7]), .B(exu_n16197), .Y(exu_n30884));
INVX1 exu_U31422(.A(exu_n30884), .Y(exu_n11365));
INVX1 exu_U31423(.A(div_byp_muldivout_g[6]), .Y(exu_n11366));
AND2X1 exu_U31424(.A(div_d[6]), .B(exu_n16197), .Y(exu_n30885));
INVX1 exu_U31425(.A(exu_n30885), .Y(exu_n11367));
INVX1 exu_U31426(.A(div_byp_muldivout_g[63]), .Y(exu_n11368));
AND2X1 exu_U31427(.A(div_d_63), .B(exu_n16197), .Y(exu_n30886));
INVX1 exu_U31428(.A(exu_n30886), .Y(exu_n11369));
INVX1 exu_U31429(.A(div_byp_muldivout_g[62]), .Y(exu_n11370));
AND2X1 exu_U31430(.A(div_ecl_d_62), .B(exu_n16197), .Y(exu_n30887));
INVX1 exu_U31431(.A(exu_n30887), .Y(exu_n11371));
INVX1 exu_U31432(.A(div_byp_muldivout_g[61]), .Y(exu_n11372));
AND2X1 exu_U31433(.A(div_d[61]), .B(exu_n16197), .Y(exu_n30888));
INVX1 exu_U31434(.A(exu_n30888), .Y(exu_n11373));
INVX1 exu_U31435(.A(div_byp_muldivout_g[60]), .Y(exu_n11374));
AND2X1 exu_U31436(.A(div_d[60]), .B(exu_n16197), .Y(exu_n30889));
INVX1 exu_U31437(.A(exu_n30889), .Y(exu_n11375));
INVX1 exu_U31438(.A(div_byp_muldivout_g[5]), .Y(exu_n11376));
AND2X1 exu_U31439(.A(div_d[5]), .B(exu_n16197), .Y(exu_n30890));
INVX1 exu_U31440(.A(exu_n30890), .Y(exu_n11377));
INVX1 exu_U31441(.A(div_byp_muldivout_g[59]), .Y(exu_n11378));
AND2X1 exu_U31442(.A(div_d[59]), .B(exu_n16195), .Y(exu_n30891));
INVX1 exu_U31443(.A(exu_n30891), .Y(exu_n11379));
INVX1 exu_U31444(.A(div_byp_muldivout_g[58]), .Y(exu_n11380));
AND2X1 exu_U31445(.A(div_d[58]), .B(exu_n16193), .Y(exu_n30892));
INVX1 exu_U31446(.A(exu_n30892), .Y(exu_n11381));
INVX1 exu_U31447(.A(div_byp_muldivout_g[57]), .Y(exu_n11382));
AND2X1 exu_U31448(.A(div_d[57]), .B(exu_n16194), .Y(exu_n30893));
INVX1 exu_U31449(.A(exu_n30893), .Y(exu_n11383));
INVX1 exu_U31450(.A(div_byp_muldivout_g[56]), .Y(exu_n11384));
AND2X1 exu_U31451(.A(div_d[56]), .B(exu_n16197), .Y(exu_n30894));
INVX1 exu_U31452(.A(exu_n30894), .Y(exu_n11385));
INVX1 exu_U31453(.A(div_byp_muldivout_g[55]), .Y(exu_n11386));
AND2X1 exu_U31454(.A(div_d[55]), .B(ecl_div_sel_div), .Y(exu_n30895));
INVX1 exu_U31455(.A(exu_n30895), .Y(exu_n11387));
INVX1 exu_U31456(.A(div_byp_muldivout_g[54]), .Y(exu_n11388));
AND2X1 exu_U31457(.A(div_d[54]), .B(exu_n16195), .Y(exu_n30896));
INVX1 exu_U31458(.A(exu_n30896), .Y(exu_n11389));
INVX1 exu_U31459(.A(div_byp_muldivout_g[53]), .Y(exu_n11390));
AND2X1 exu_U31460(.A(div_d[53]), .B(exu_n16193), .Y(exu_n30897));
INVX1 exu_U31461(.A(exu_n30897), .Y(exu_n11391));
INVX1 exu_U31462(.A(div_byp_muldivout_g[52]), .Y(exu_n11392));
AND2X1 exu_U31463(.A(div_d[52]), .B(exu_n16194), .Y(exu_n30898));
INVX1 exu_U31464(.A(exu_n30898), .Y(exu_n11393));
INVX1 exu_U31465(.A(div_byp_muldivout_g[51]), .Y(exu_n11394));
AND2X1 exu_U31466(.A(div_d[51]), .B(exu_n16197), .Y(exu_n30899));
INVX1 exu_U31467(.A(exu_n30899), .Y(exu_n11395));
INVX1 exu_U31468(.A(div_byp_muldivout_g[50]), .Y(exu_n11396));
AND2X1 exu_U31469(.A(div_d[50]), .B(ecl_div_sel_div), .Y(exu_n30900));
INVX1 exu_U31470(.A(exu_n30900), .Y(exu_n11397));
INVX1 exu_U31471(.A(div_byp_muldivout_g[4]), .Y(exu_n11398));
AND2X1 exu_U31472(.A(div_d[4]), .B(exu_n16195), .Y(exu_n30901));
INVX1 exu_U31473(.A(exu_n30901), .Y(exu_n11399));
INVX1 exu_U31474(.A(div_byp_muldivout_g[49]), .Y(exu_n11400));
AND2X1 exu_U31475(.A(div_d[49]), .B(exu_n16193), .Y(exu_n30902));
INVX1 exu_U31476(.A(exu_n30902), .Y(exu_n11401));
INVX1 exu_U31477(.A(div_byp_muldivout_g[48]), .Y(exu_n11402));
AND2X1 exu_U31478(.A(div_d[48]), .B(exu_n16194), .Y(exu_n30903));
INVX1 exu_U31479(.A(exu_n30903), .Y(exu_n11403));
INVX1 exu_U31480(.A(div_byp_muldivout_g[47]), .Y(exu_n11404));
AND2X1 exu_U31481(.A(div_d[47]), .B(ecl_div_sel_div), .Y(exu_n30904));
INVX1 exu_U31482(.A(exu_n30904), .Y(exu_n11405));
INVX1 exu_U31483(.A(div_byp_muldivout_g[46]), .Y(exu_n11406));
AND2X1 exu_U31484(.A(div_d[46]), .B(exu_n16194), .Y(exu_n30905));
INVX1 exu_U31485(.A(exu_n30905), .Y(exu_n11407));
INVX1 exu_U31486(.A(div_byp_muldivout_g[45]), .Y(exu_n11408));
AND2X1 exu_U31487(.A(div_d[45]), .B(ecl_div_sel_div), .Y(exu_n30906));
INVX1 exu_U31488(.A(exu_n30906), .Y(exu_n11409));
INVX1 exu_U31489(.A(div_byp_muldivout_g[44]), .Y(exu_n11410));
AND2X1 exu_U31490(.A(div_d[44]), .B(exu_n16194), .Y(exu_n30907));
INVX1 exu_U31491(.A(exu_n30907), .Y(exu_n11411));
INVX1 exu_U31492(.A(div_byp_muldivout_g[43]), .Y(exu_n11412));
AND2X1 exu_U31493(.A(div_d[43]), .B(ecl_div_sel_div), .Y(exu_n30908));
INVX1 exu_U31494(.A(exu_n30908), .Y(exu_n11413));
INVX1 exu_U31495(.A(div_byp_muldivout_g[42]), .Y(exu_n11414));
AND2X1 exu_U31496(.A(div_d[42]), .B(exu_n16194), .Y(exu_n30909));
INVX1 exu_U31497(.A(exu_n30909), .Y(exu_n11415));
INVX1 exu_U31498(.A(div_byp_muldivout_g[41]), .Y(exu_n11416));
AND2X1 exu_U31499(.A(div_d[41]), .B(ecl_div_sel_div), .Y(exu_n30910));
INVX1 exu_U31500(.A(exu_n30910), .Y(exu_n11417));
INVX1 exu_U31501(.A(div_byp_muldivout_g[40]), .Y(exu_n11418));
AND2X1 exu_U31502(.A(div_d[40]), .B(exu_n16194), .Y(exu_n30911));
INVX1 exu_U31503(.A(exu_n30911), .Y(exu_n11419));
INVX1 exu_U31504(.A(div_byp_muldivout_g[3]), .Y(exu_n11420));
AND2X1 exu_U31505(.A(div_d[3]), .B(ecl_div_sel_div), .Y(exu_n30912));
INVX1 exu_U31506(.A(exu_n30912), .Y(exu_n11421));
INVX1 exu_U31507(.A(div_byp_muldivout_g[39]), .Y(exu_n11422));
AND2X1 exu_U31508(.A(div_d[39]), .B(exu_n16194), .Y(exu_n30913));
INVX1 exu_U31509(.A(exu_n30913), .Y(exu_n11423));
INVX1 exu_U31510(.A(div_byp_muldivout_g[38]), .Y(exu_n11424));
AND2X1 exu_U31511(.A(div_d[38]), .B(exu_n16193), .Y(exu_n30914));
INVX1 exu_U31512(.A(exu_n30914), .Y(exu_n11425));
INVX1 exu_U31513(.A(div_byp_muldivout_g[37]), .Y(exu_n11426));
AND2X1 exu_U31514(.A(div_d[37]), .B(ecl_div_sel_div), .Y(exu_n30915));
INVX1 exu_U31515(.A(exu_n30915), .Y(exu_n11427));
INVX1 exu_U31516(.A(div_byp_muldivout_g[36]), .Y(exu_n11428));
AND2X1 exu_U31517(.A(div_d[36]), .B(ecl_div_sel_div), .Y(exu_n30916));
INVX1 exu_U31518(.A(exu_n30916), .Y(exu_n11429));
INVX1 exu_U31519(.A(div_byp_muldivout_g[35]), .Y(exu_n11430));
AND2X1 exu_U31520(.A(div_d[35]), .B(exu_n16194), .Y(exu_n30917));
INVX1 exu_U31521(.A(exu_n30917), .Y(exu_n11431));
INVX1 exu_U31522(.A(div_byp_muldivout_g[34]), .Y(exu_n11432));
AND2X1 exu_U31523(.A(div_d[34]), .B(ecl_div_sel_div), .Y(exu_n30918));
INVX1 exu_U31524(.A(exu_n30918), .Y(exu_n11433));
INVX1 exu_U31525(.A(div_byp_muldivout_g[33]), .Y(exu_n11434));
AND2X1 exu_U31526(.A(div_d[33]), .B(exu_n16194), .Y(exu_n30919));
INVX1 exu_U31527(.A(exu_n30919), .Y(exu_n11435));
INVX1 exu_U31528(.A(div_byp_muldivout_g[32]), .Y(exu_n11436));
AND2X1 exu_U31529(.A(div_d[32]), .B(exu_n16193), .Y(exu_n30920));
INVX1 exu_U31530(.A(exu_n30920), .Y(exu_n11437));
INVX1 exu_U31531(.A(div_byp_muldivout_g[31]), .Y(exu_n11438));
AND2X1 exu_U31532(.A(div_d[31]), .B(exu_n16197), .Y(exu_n30921));
INVX1 exu_U31533(.A(exu_n30921), .Y(exu_n11439));
INVX1 exu_U31534(.A(div_byp_muldivout_g[30]), .Y(exu_n11440));
AND2X1 exu_U31535(.A(div_d[30]), .B(exu_n16193), .Y(exu_n30922));
INVX1 exu_U31536(.A(exu_n30922), .Y(exu_n11441));
INVX1 exu_U31537(.A(div_byp_muldivout_g[2]), .Y(exu_n11442));
AND2X1 exu_U31538(.A(div_d[2]), .B(exu_n16193), .Y(exu_n30923));
INVX1 exu_U31539(.A(exu_n30923), .Y(exu_n11443));
INVX1 exu_U31540(.A(div_byp_muldivout_g[29]), .Y(exu_n11444));
AND2X1 exu_U31541(.A(div_d[29]), .B(exu_n16195), .Y(exu_n30924));
INVX1 exu_U31542(.A(exu_n30924), .Y(exu_n11445));
INVX1 exu_U31543(.A(div_byp_muldivout_g[28]), .Y(exu_n11446));
AND2X1 exu_U31544(.A(div_d[28]), .B(ecl_div_sel_div), .Y(exu_n30925));
INVX1 exu_U31545(.A(exu_n30925), .Y(exu_n11447));
INVX1 exu_U31546(.A(div_byp_muldivout_g[27]), .Y(exu_n11448));
AND2X1 exu_U31547(.A(div_d[27]), .B(exu_n16195), .Y(exu_n30926));
INVX1 exu_U31548(.A(exu_n30926), .Y(exu_n11449));
INVX1 exu_U31549(.A(div_byp_muldivout_g[26]), .Y(exu_n11450));
AND2X1 exu_U31550(.A(div_d[26]), .B(exu_n16194), .Y(exu_n30927));
INVX1 exu_U31551(.A(exu_n30927), .Y(exu_n11451));
INVX1 exu_U31552(.A(div_byp_muldivout_g[25]), .Y(exu_n11452));
AND2X1 exu_U31553(.A(div_d[25]), .B(exu_n16194), .Y(exu_n30928));
INVX1 exu_U31554(.A(exu_n30928), .Y(exu_n11453));
INVX1 exu_U31555(.A(div_byp_muldivout_g[24]), .Y(exu_n11454));
AND2X1 exu_U31556(.A(div_d[24]), .B(exu_n16197), .Y(exu_n30929));
INVX1 exu_U31557(.A(exu_n30929), .Y(exu_n11455));
INVX1 exu_U31558(.A(div_byp_muldivout_g[23]), .Y(exu_n11456));
AND2X1 exu_U31559(.A(div_d[23]), .B(exu_n16193), .Y(exu_n30930));
INVX1 exu_U31560(.A(exu_n30930), .Y(exu_n11457));
INVX1 exu_U31561(.A(div_byp_muldivout_g[22]), .Y(exu_n11458));
AND2X1 exu_U31562(.A(div_d[22]), .B(exu_n16194), .Y(exu_n30931));
INVX1 exu_U31563(.A(exu_n30931), .Y(exu_n11459));
INVX1 exu_U31564(.A(div_byp_muldivout_g[21]), .Y(exu_n11460));
AND2X1 exu_U31565(.A(div_d[21]), .B(exu_n16195), .Y(exu_n30932));
INVX1 exu_U31566(.A(exu_n30932), .Y(exu_n11461));
INVX1 exu_U31567(.A(div_byp_muldivout_g[20]), .Y(exu_n11462));
AND2X1 exu_U31568(.A(div_d[20]), .B(exu_n16197), .Y(exu_n30933));
INVX1 exu_U31569(.A(exu_n30933), .Y(exu_n11463));
INVX1 exu_U31570(.A(div_byp_muldivout_g[1]), .Y(exu_n11464));
AND2X1 exu_U31571(.A(div_d[1]), .B(exu_n16194), .Y(exu_n30934));
INVX1 exu_U31572(.A(exu_n30934), .Y(exu_n11465));
INVX1 exu_U31573(.A(div_byp_muldivout_g[19]), .Y(exu_n11466));
AND2X1 exu_U31574(.A(div_d[19]), .B(exu_n16195), .Y(exu_n30935));
INVX1 exu_U31575(.A(exu_n30935), .Y(exu_n11467));
INVX1 exu_U31576(.A(div_byp_muldivout_g[18]), .Y(exu_n11468));
AND2X1 exu_U31577(.A(div_d[18]), .B(exu_n16193), .Y(exu_n30936));
INVX1 exu_U31578(.A(exu_n30936), .Y(exu_n11469));
INVX1 exu_U31579(.A(div_byp_muldivout_g[17]), .Y(exu_n11470));
AND2X1 exu_U31580(.A(div_d[17]), .B(exu_n16195), .Y(exu_n30937));
INVX1 exu_U31581(.A(exu_n30937), .Y(exu_n11471));
INVX1 exu_U31582(.A(div_byp_muldivout_g[16]), .Y(exu_n11472));
AND2X1 exu_U31583(.A(div_d[16]), .B(ecl_div_sel_div), .Y(exu_n30938));
INVX1 exu_U31584(.A(exu_n30938), .Y(exu_n11473));
INVX1 exu_U31585(.A(div_byp_muldivout_g[15]), .Y(exu_n11474));
AND2X1 exu_U31586(.A(div_d[15]), .B(ecl_div_sel_div), .Y(exu_n30939));
INVX1 exu_U31587(.A(exu_n30939), .Y(exu_n11475));
INVX1 exu_U31588(.A(div_byp_muldivout_g[14]), .Y(exu_n11476));
AND2X1 exu_U31589(.A(div_d[14]), .B(exu_n16194), .Y(exu_n30940));
INVX1 exu_U31590(.A(exu_n30940), .Y(exu_n11477));
INVX1 exu_U31591(.A(div_byp_muldivout_g[13]), .Y(exu_n11478));
AND2X1 exu_U31592(.A(div_d[13]), .B(exu_n16193), .Y(exu_n30941));
INVX1 exu_U31593(.A(exu_n30941), .Y(exu_n11479));
INVX1 exu_U31594(.A(div_byp_muldivout_g[12]), .Y(exu_n11480));
AND2X1 exu_U31595(.A(div_d[12]), .B(exu_n16197), .Y(exu_n30942));
INVX1 exu_U31596(.A(exu_n30942), .Y(exu_n11481));
INVX1 exu_U31597(.A(div_byp_muldivout_g[11]), .Y(exu_n11482));
AND2X1 exu_U31598(.A(div_d[11]), .B(ecl_div_sel_div), .Y(exu_n30943));
INVX1 exu_U31599(.A(exu_n30943), .Y(exu_n11483));
INVX1 exu_U31600(.A(div_byp_muldivout_g[10]), .Y(exu_n11484));
AND2X1 exu_U31601(.A(div_d[10]), .B(ecl_div_sel_div), .Y(exu_n30944));
INVX1 exu_U31602(.A(exu_n30944), .Y(exu_n11485));
INVX1 exu_U31603(.A(div_byp_muldivout_g[0]), .Y(exu_n11486));
AND2X1 exu_U31604(.A(div_d[0]), .B(exu_n16193), .Y(exu_n30945));
INVX1 exu_U31605(.A(exu_n30945), .Y(exu_n11487));
AND2X1 exu_U31606(.A(ecl_div_mul_wen), .B(mul_data_out[9]), .Y(exu_n31329));
INVX1 exu_U31607(.A(exu_n31329), .Y(exu_n11488));
AND2X1 exu_U31608(.A(mul_data_out[8]), .B(ecl_div_mul_wen), .Y(exu_n31331));
INVX1 exu_U31609(.A(exu_n31331), .Y(exu_n11489));
AND2X1 exu_U31610(.A(mul_data_out[7]), .B(ecl_div_mul_wen), .Y(exu_n31333));
INVX1 exu_U31611(.A(exu_n31333), .Y(exu_n11490));
AND2X1 exu_U31612(.A(mul_data_out[6]), .B(ecl_div_mul_wen), .Y(exu_n31335));
INVX1 exu_U31613(.A(exu_n31335), .Y(exu_n11491));
AND2X1 exu_U31614(.A(mul_data_out[63]), .B(ecl_div_mul_wen), .Y(exu_n31337));
INVX1 exu_U31615(.A(exu_n31337), .Y(exu_n11492));
AND2X1 exu_U31616(.A(mul_data_out[62]), .B(ecl_div_mul_wen), .Y(exu_n31339));
INVX1 exu_U31617(.A(exu_n31339), .Y(exu_n11493));
AND2X1 exu_U31618(.A(mul_data_out[61]), .B(ecl_div_mul_wen), .Y(exu_n31341));
INVX1 exu_U31619(.A(exu_n31341), .Y(exu_n11494));
AND2X1 exu_U31620(.A(mul_data_out[60]), .B(ecl_div_mul_wen), .Y(exu_n31343));
INVX1 exu_U31621(.A(exu_n31343), .Y(exu_n11495));
AND2X1 exu_U31622(.A(mul_data_out[5]), .B(ecl_div_mul_wen), .Y(exu_n31345));
INVX1 exu_U31623(.A(exu_n31345), .Y(exu_n11496));
AND2X1 exu_U31624(.A(mul_data_out[59]), .B(ecl_div_mul_wen), .Y(exu_n31347));
INVX1 exu_U31625(.A(exu_n31347), .Y(exu_n11497));
AND2X1 exu_U31626(.A(mul_data_out[58]), .B(ecl_div_mul_wen), .Y(exu_n31349));
INVX1 exu_U31627(.A(exu_n31349), .Y(exu_n11498));
AND2X1 exu_U31628(.A(mul_data_out[57]), .B(ecl_div_mul_wen), .Y(exu_n31351));
INVX1 exu_U31629(.A(exu_n31351), .Y(exu_n11499));
AND2X1 exu_U31630(.A(mul_data_out[56]), .B(ecl_div_mul_wen), .Y(exu_n31353));
INVX1 exu_U31631(.A(exu_n31353), .Y(exu_n11500));
AND2X1 exu_U31632(.A(mul_data_out[55]), .B(ecl_div_mul_wen), .Y(exu_n31355));
INVX1 exu_U31633(.A(exu_n31355), .Y(exu_n11501));
AND2X1 exu_U31634(.A(mul_data_out[54]), .B(ecl_div_mul_wen), .Y(exu_n31357));
INVX1 exu_U31635(.A(exu_n31357), .Y(exu_n11502));
AND2X1 exu_U31636(.A(mul_data_out[53]), .B(ecl_div_mul_wen), .Y(exu_n31359));
INVX1 exu_U31637(.A(exu_n31359), .Y(exu_n11503));
AND2X1 exu_U31638(.A(mul_data_out[52]), .B(ecl_div_mul_wen), .Y(exu_n31361));
INVX1 exu_U31639(.A(exu_n31361), .Y(exu_n11504));
AND2X1 exu_U31640(.A(mul_data_out[51]), .B(ecl_div_mul_wen), .Y(exu_n31363));
INVX1 exu_U31641(.A(exu_n31363), .Y(exu_n11505));
AND2X1 exu_U31642(.A(mul_data_out[50]), .B(ecl_div_mul_wen), .Y(exu_n31365));
INVX1 exu_U31643(.A(exu_n31365), .Y(exu_n11506));
AND2X1 exu_U31644(.A(mul_data_out[4]), .B(ecl_div_mul_wen), .Y(exu_n31367));
INVX1 exu_U31645(.A(exu_n31367), .Y(exu_n11507));
AND2X1 exu_U31646(.A(mul_data_out[49]), .B(ecl_div_mul_wen), .Y(exu_n31369));
INVX1 exu_U31647(.A(exu_n31369), .Y(exu_n11508));
AND2X1 exu_U31648(.A(mul_data_out[48]), .B(ecl_div_mul_wen), .Y(exu_n31371));
INVX1 exu_U31649(.A(exu_n31371), .Y(exu_n11509));
AND2X1 exu_U31650(.A(mul_data_out[47]), .B(ecl_div_mul_wen), .Y(exu_n31373));
INVX1 exu_U31651(.A(exu_n31373), .Y(exu_n11510));
AND2X1 exu_U31652(.A(mul_data_out[46]), .B(ecl_div_mul_wen), .Y(exu_n31375));
INVX1 exu_U31653(.A(exu_n31375), .Y(exu_n11511));
AND2X1 exu_U31654(.A(mul_data_out[45]), .B(ecl_div_mul_wen), .Y(exu_n31377));
INVX1 exu_U31655(.A(exu_n31377), .Y(exu_n11512));
AND2X1 exu_U31656(.A(mul_data_out[44]), .B(ecl_div_mul_wen), .Y(exu_n31379));
INVX1 exu_U31657(.A(exu_n31379), .Y(exu_n11513));
AND2X1 exu_U31658(.A(mul_data_out[43]), .B(ecl_div_mul_wen), .Y(exu_n31381));
INVX1 exu_U31659(.A(exu_n31381), .Y(exu_n11514));
AND2X1 exu_U31660(.A(mul_data_out[42]), .B(ecl_div_mul_wen), .Y(exu_n31383));
INVX1 exu_U31661(.A(exu_n31383), .Y(exu_n11515));
AND2X1 exu_U31662(.A(mul_data_out[41]), .B(ecl_div_mul_wen), .Y(exu_n31385));
INVX1 exu_U31663(.A(exu_n31385), .Y(exu_n11516));
AND2X1 exu_U31664(.A(mul_data_out[40]), .B(ecl_div_mul_wen), .Y(exu_n31387));
INVX1 exu_U31665(.A(exu_n31387), .Y(exu_n11517));
AND2X1 exu_U31666(.A(mul_data_out[3]), .B(ecl_div_mul_wen), .Y(exu_n31389));
INVX1 exu_U31667(.A(exu_n31389), .Y(exu_n11518));
AND2X1 exu_U31668(.A(mul_data_out[39]), .B(ecl_div_mul_wen), .Y(exu_n31391));
INVX1 exu_U31669(.A(exu_n31391), .Y(exu_n11519));
AND2X1 exu_U31670(.A(mul_data_out[38]), .B(ecl_div_mul_wen), .Y(exu_n31393));
INVX1 exu_U31671(.A(exu_n31393), .Y(exu_n11520));
AND2X1 exu_U31672(.A(mul_data_out[37]), .B(ecl_div_mul_wen), .Y(exu_n31395));
INVX1 exu_U31673(.A(exu_n31395), .Y(exu_n11521));
AND2X1 exu_U31674(.A(mul_data_out[36]), .B(ecl_div_mul_wen), .Y(exu_n31397));
INVX1 exu_U31675(.A(exu_n31397), .Y(exu_n11522));
AND2X1 exu_U31676(.A(mul_data_out[35]), .B(ecl_div_mul_wen), .Y(exu_n31399));
INVX1 exu_U31677(.A(exu_n31399), .Y(exu_n11523));
AND2X1 exu_U31678(.A(mul_data_out[34]), .B(ecl_div_mul_wen), .Y(exu_n31401));
INVX1 exu_U31679(.A(exu_n31401), .Y(exu_n11524));
AND2X1 exu_U31680(.A(mul_data_out[33]), .B(ecl_div_mul_wen), .Y(exu_n31403));
INVX1 exu_U31681(.A(exu_n31403), .Y(exu_n11525));
AND2X1 exu_U31682(.A(mul_data_out[32]), .B(ecl_div_mul_wen), .Y(exu_n31405));
INVX1 exu_U31683(.A(exu_n31405), .Y(exu_n11526));
AND2X1 exu_U31684(.A(mul_data_out[31]), .B(ecl_div_mul_wen), .Y(exu_n31407));
INVX1 exu_U31685(.A(exu_n31407), .Y(exu_n11527));
AND2X1 exu_U31686(.A(mul_data_out[30]), .B(ecl_div_mul_wen), .Y(exu_n31409));
INVX1 exu_U31687(.A(exu_n31409), .Y(exu_n11528));
AND2X1 exu_U31688(.A(mul_data_out[2]), .B(ecl_div_mul_wen), .Y(exu_n31411));
INVX1 exu_U31689(.A(exu_n31411), .Y(exu_n11529));
AND2X1 exu_U31690(.A(mul_data_out[29]), .B(ecl_div_mul_wen), .Y(exu_n31413));
INVX1 exu_U31691(.A(exu_n31413), .Y(exu_n11530));
AND2X1 exu_U31692(.A(mul_data_out[28]), .B(ecl_div_mul_wen), .Y(exu_n31415));
INVX1 exu_U31693(.A(exu_n31415), .Y(exu_n11531));
AND2X1 exu_U31694(.A(mul_data_out[27]), .B(ecl_div_mul_wen), .Y(exu_n31417));
INVX1 exu_U31695(.A(exu_n31417), .Y(exu_n11532));
AND2X1 exu_U31696(.A(mul_data_out[26]), .B(ecl_div_mul_wen), .Y(exu_n31419));
INVX1 exu_U31697(.A(exu_n31419), .Y(exu_n11533));
AND2X1 exu_U31698(.A(mul_data_out[25]), .B(ecl_div_mul_wen), .Y(exu_n31421));
INVX1 exu_U31699(.A(exu_n31421), .Y(exu_n11534));
AND2X1 exu_U31700(.A(mul_data_out[24]), .B(ecl_div_mul_wen), .Y(exu_n31423));
INVX1 exu_U31701(.A(exu_n31423), .Y(exu_n11535));
AND2X1 exu_U31702(.A(mul_data_out[23]), .B(ecl_div_mul_wen), .Y(exu_n31425));
INVX1 exu_U31703(.A(exu_n31425), .Y(exu_n11536));
AND2X1 exu_U31704(.A(mul_data_out[22]), .B(ecl_div_mul_wen), .Y(exu_n31427));
INVX1 exu_U31705(.A(exu_n31427), .Y(exu_n11537));
AND2X1 exu_U31706(.A(mul_data_out[21]), .B(ecl_div_mul_wen), .Y(exu_n31429));
INVX1 exu_U31707(.A(exu_n31429), .Y(exu_n11538));
AND2X1 exu_U31708(.A(mul_data_out[20]), .B(ecl_div_mul_wen), .Y(exu_n31431));
INVX1 exu_U31709(.A(exu_n31431), .Y(exu_n11539));
AND2X1 exu_U31710(.A(mul_data_out[1]), .B(ecl_div_mul_wen), .Y(exu_n31433));
INVX1 exu_U31711(.A(exu_n31433), .Y(exu_n11540));
AND2X1 exu_U31712(.A(mul_data_out[19]), .B(ecl_div_mul_wen), .Y(exu_n31435));
INVX1 exu_U31713(.A(exu_n31435), .Y(exu_n11541));
AND2X1 exu_U31714(.A(mul_data_out[18]), .B(ecl_div_mul_wen), .Y(exu_n31437));
INVX1 exu_U31715(.A(exu_n31437), .Y(exu_n11542));
AND2X1 exu_U31716(.A(mul_data_out[17]), .B(ecl_div_mul_wen), .Y(exu_n31439));
INVX1 exu_U31717(.A(exu_n31439), .Y(exu_n11543));
AND2X1 exu_U31718(.A(mul_data_out[16]), .B(ecl_div_mul_wen), .Y(exu_n31441));
INVX1 exu_U31719(.A(exu_n31441), .Y(exu_n11544));
AND2X1 exu_U31720(.A(mul_data_out[15]), .B(ecl_div_mul_wen), .Y(exu_n31443));
INVX1 exu_U31721(.A(exu_n31443), .Y(exu_n11545));
AND2X1 exu_U31722(.A(mul_data_out[14]), .B(ecl_div_mul_wen), .Y(exu_n31445));
INVX1 exu_U31723(.A(exu_n31445), .Y(exu_n11546));
AND2X1 exu_U31724(.A(mul_data_out[13]), .B(ecl_div_mul_wen), .Y(exu_n31447));
INVX1 exu_U31725(.A(exu_n31447), .Y(exu_n11547));
AND2X1 exu_U31726(.A(mul_data_out[12]), .B(ecl_div_mul_wen), .Y(exu_n31449));
INVX1 exu_U31727(.A(exu_n31449), .Y(exu_n11548));
AND2X1 exu_U31728(.A(mul_data_out[11]), .B(ecl_div_mul_wen), .Y(exu_n31451));
INVX1 exu_U31729(.A(exu_n31451), .Y(exu_n11549));
AND2X1 exu_U31730(.A(mul_data_out[10]), .B(ecl_div_mul_wen), .Y(exu_n31453));
INVX1 exu_U31731(.A(exu_n31453), .Y(exu_n11550));
AND2X1 exu_U31732(.A(mul_data_out[0]), .B(ecl_div_mul_wen), .Y(exu_n31455));
INVX1 exu_U31733(.A(exu_n31455), .Y(exu_n11551));
AND2X1 exu_U31734(.A(rml_cwp_cwp_output_queue_pv[3]), .B(exu_n15027), .Y(rml_cwp_cwp_output_queue_n10));
INVX1 exu_U31735(.A(rml_cwp_cwp_output_queue_n10), .Y(exu_n11552));
AND2X1 exu_U31736(.A(rml_cwp_cwp_output_queue_pv[2]), .B(exu_n15027), .Y(rml_cwp_cwp_output_queue_n12));
INVX1 exu_U31737(.A(rml_cwp_cwp_output_queue_n12), .Y(exu_n11553));
AND2X1 exu_U31738(.A(rml_cwp_cwp_output_queue_pv[1]), .B(exu_n15027), .Y(rml_cwp_cwp_output_queue_n14));
INVX1 exu_U31739(.A(rml_cwp_cwp_output_queue_n14), .Y(exu_n11554));
AND2X1 exu_U31740(.A(rml_cwp_cwp_output_queue_pv[0]), .B(exu_n15027), .Y(rml_cwp_cwp_output_queue_n16));
INVX1 exu_U31741(.A(rml_cwp_cwp_output_queue_n16), .Y(exu_n11555));
INVX1 exu_U31742(.A(rml_cwp_cwp_output_queue_n25), .Y(exu_n11556));
INVX1 exu_U31743(.A(rml_cwp_cwp_output_queue_n35), .Y(exu_n11557));
AND2X1 exu_U31744(.A(exu_n16626), .B(exu_n16625), .Y(rml_cwp_cwp_output_queue_n36));
INVX1 exu_U31745(.A(rml_cwp_cwp_output_queue_n36), .Y(exu_n11558));
AND2X1 exu_U31746(.A(rml_cwp_n74), .B(rml_ecl_wtype_e[0]), .Y(rml_cwp_slot0_data_mux_n4));
INVX1 exu_U31747(.A(rml_cwp_slot0_data_mux_n4), .Y(exu_n11559));
AND2X1 exu_U31748(.A(rml_ecl_other_e), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n8));
INVX1 exu_U31749(.A(rml_cwp_slot0_data_mux_n8), .Y(exu_n11560));
AND2X1 exu_U31750(.A(exu_n15940), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n16));
INVX1 exu_U31751(.A(rml_cwp_slot0_data_mux_n16), .Y(exu_n11561));
AND2X1 exu_U31752(.A(rml_cwp_tlu_swap_data[12]), .B(rml_cwp_swap_sel_tlu[0]), .Y(rml_cwp_slot0_data_mux_n39));
INVX1 exu_U31753(.A(rml_cwp_slot0_data_mux_n39), .Y(exu_n11562));
AND2X1 exu_U31754(.A(rml_ecl_wtype_e[2]), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n44));
INVX1 exu_U31755(.A(rml_cwp_slot0_data_mux_n44), .Y(exu_n11563));
AND2X1 exu_U31756(.A(rml_ecl_wtype_e[1]), .B(rml_cwp_n74), .Y(rml_cwp_slot0_data_mux_n48));
INVX1 exu_U31757(.A(rml_cwp_slot0_data_mux_n48), .Y(exu_n11564));
AND2X1 exu_U31758(.A(ecl_tid_d[0]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n2));
INVX1 exu_U31759(.A(ecl_mdqctl_div_data_mux_n2), .Y(exu_n11565));
AND2X1 exu_U31760(.A(ecl_tid_d[1]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n4));
INVX1 exu_U31761(.A(ecl_mdqctl_div_data_mux_n4), .Y(exu_n11566));
AND2X1 exu_U31762(.A(ifu_exu_rd_d[0]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n6));
INVX1 exu_U31763(.A(ecl_mdqctl_div_data_mux_n6), .Y(exu_n11567));
AND2X1 exu_U31764(.A(ifu_exu_rd_d[1]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n8));
INVX1 exu_U31765(.A(ecl_mdqctl_div_data_mux_n8), .Y(exu_n11568));
AND2X1 exu_U31766(.A(ifu_exu_rd_d[2]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n10));
INVX1 exu_U31767(.A(ecl_mdqctl_div_data_mux_n10), .Y(exu_n11569));
AND2X1 exu_U31768(.A(ifu_exu_rd_d[3]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n12));
INVX1 exu_U31769(.A(ecl_mdqctl_div_data_mux_n12), .Y(exu_n11570));
AND2X1 exu_U31770(.A(ifu_exu_rd_d[4]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n14));
INVX1 exu_U31771(.A(ecl_mdqctl_div_data_mux_n14), .Y(exu_n11571));
AND2X1 exu_U31772(.A(ifu_exu_muldivop_d[0]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n16));
INVX1 exu_U31773(.A(ecl_mdqctl_div_data_mux_n16), .Y(exu_n11572));
AND2X1 exu_U31774(.A(ifu_exu_muldivop_d[1]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n18));
INVX1 exu_U31775(.A(ecl_mdqctl_div_data_mux_n18), .Y(exu_n11573));
AND2X1 exu_U31776(.A(ifu_exu_muldivop_d[2]), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n20));
INVX1 exu_U31777(.A(ecl_mdqctl_div_data_mux_n20), .Y(exu_n11574));
AND2X1 exu_U31778(.A(ifu_exu_muls_d), .B(ecl_mdqctl_new_div_vld), .Y(ecl_mdqctl_div_data_mux_n22));
INVX1 exu_U31779(.A(ecl_mdqctl_div_data_mux_n22), .Y(exu_n11575));
AND2X1 exu_U31780(.A(ecl_divcntl_inputs_neg_q), .B(exu_n16370), .Y(ecl_divcntl_inputs_neg_dff_n3));
INVX1 exu_U31781(.A(ecl_divcntl_inputs_neg_dff_n3), .Y(exu_n11576));
INVX1 exu_U31782(.A(ecl_divcntl_qnext_cout_mux_n2), .Y(exu_n11577));
INVX1 exu_U31783(.A(ecl_divcntl_cnt6_n14), .Y(exu_n11578));
AND2X1 exu_U31784(.A(ecl_divcntl_cntr[3]), .B(exu_n15366), .Y(ecl_divcntl_cnt6_n21));
INVX1 exu_U31785(.A(ecl_divcntl_cnt6_n21), .Y(exu_n11579));
AND2X1 exu_U31786(.A(ecl_divcntl_cntr[2]), .B(exu_n15367), .Y(ecl_divcntl_cnt6_n27));
INVX1 exu_U31787(.A(ecl_divcntl_cnt6_n27), .Y(exu_n11580));
INVX1 exu_U31788(.A(ecl_eccctl_wb_rd_m[3]), .Y(exu_n11581));
INVX1 exu_U31789(.A(ecl_eccctl_wb_rd_m[2]), .Y(exu_n11582));
INVX1 exu_U31790(.A(ecl_eccctl_wb_rd_m[1]), .Y(exu_n11583));
INVX1 exu_U31791(.A(ecl_eccctl_wb_rd_m[0]), .Y(exu_n11584));
AND2X1 exu_U31792(.A(ecl_rd_m[0]), .B(exu_n15816), .Y(ecl_writeback_restore_rd_dff_n5));
INVX1 exu_U31793(.A(ecl_writeback_restore_rd_dff_n5), .Y(exu_n11585));
AND2X1 exu_U31794(.A(ecl_rd_m[1]), .B(exu_n15816), .Y(ecl_writeback_restore_rd_dff_n10));
INVX1 exu_U31795(.A(ecl_writeback_restore_rd_dff_n10), .Y(exu_n11586));
AND2X1 exu_U31796(.A(ecl_rd_m[2]), .B(exu_n15816), .Y(ecl_writeback_restore_rd_dff_n14));
INVX1 exu_U31797(.A(ecl_writeback_restore_rd_dff_n14), .Y(exu_n11587));
AND2X1 exu_U31798(.A(ecl_rd_m[3]), .B(exu_n15816), .Y(ecl_writeback_restore_rd_dff_n18));
INVX1 exu_U31799(.A(ecl_writeback_restore_rd_dff_n18), .Y(exu_n11588));
AND2X1 exu_U31800(.A(ecl_rd_m[4]), .B(exu_n15816), .Y(ecl_writeback_restore_rd_dff_n22));
INVX1 exu_U31801(.A(ecl_writeback_restore_rd_dff_n22), .Y(exu_n11589));
AND2X1 exu_U31802(.A(ecl_writeback_restore_tid[0]), .B(exu_n15839), .Y(ecl_writeback_restore_tid_dff_n3));
INVX1 exu_U31803(.A(ecl_writeback_restore_tid_dff_n3), .Y(exu_n11590));
AND2X1 exu_U31804(.A(ecl_writeback_restore_tid[1]), .B(exu_n15839), .Y(ecl_writeback_restore_tid_dff_n9));
INVX1 exu_U31805(.A(ecl_writeback_restore_tid_dff_n9), .Y(exu_n11591));
AND2X1 exu_U31806(.A(ecl_mdqctl_wb_divsetcc_g), .B(ecl_div_sel_div), .Y(ecl_writeback_setcc_g_mux_n2));
INVX1 exu_U31807(.A(ecl_writeback_setcc_g_mux_n2), .Y(exu_n11592));
AND2X1 exu_U31808(.A(exu_n15701), .B(ecl_ccr_wen_thr0_w), .Y(ecl_ccr_mux_ccrin0_n12));
INVX1 exu_U31809(.A(ecl_ccr_mux_ccrin0_n12), .Y(exu_n11593));
AND2X1 exu_U31810(.A(exu_n15700), .B(ecl_ccr_wen_thr0_w), .Y(ecl_ccr_mux_ccrin0_n16));
INVX1 exu_U31811(.A(ecl_ccr_mux_ccrin0_n16), .Y(exu_n11594));
AND2X1 exu_U31812(.A(tlu_exu_ccr_m[0]), .B(tlu_exu_cwpccr_update_m), .Y(ecl_ccr_mux_ccr_m_n2));
INVX1 exu_U31813(.A(ecl_ccr_mux_ccr_m_n2), .Y(exu_n11595));
AND2X1 exu_U31814(.A(tlu_exu_ccr_m[1]), .B(tlu_exu_cwpccr_update_m), .Y(ecl_ccr_mux_ccr_m_n4));
INVX1 exu_U31815(.A(ecl_ccr_mux_ccr_m_n4), .Y(exu_n11596));
AND2X1 exu_U31816(.A(tlu_exu_ccr_m[2]), .B(tlu_exu_cwpccr_update_m), .Y(ecl_ccr_mux_ccr_m_n6));
INVX1 exu_U31817(.A(ecl_ccr_mux_ccr_m_n6), .Y(exu_n11597));
AND2X1 exu_U31818(.A(tlu_exu_ccr_m[3]), .B(tlu_exu_cwpccr_update_m), .Y(ecl_ccr_mux_ccr_m_n8));
INVX1 exu_U31819(.A(ecl_ccr_mux_ccr_m_n8), .Y(exu_n11598));
AND2X1 exu_U31820(.A(tlu_exu_ccr_m[4]), .B(tlu_exu_cwpccr_update_m), .Y(ecl_ccr_mux_ccr_m_n10));
INVX1 exu_U31821(.A(ecl_ccr_mux_ccr_m_n10), .Y(exu_n11599));
AND2X1 exu_U31822(.A(tlu_exu_ccr_m[5]), .B(tlu_exu_cwpccr_update_m), .Y(ecl_ccr_mux_ccr_m_n12));
INVX1 exu_U31823(.A(ecl_ccr_mux_ccr_m_n12), .Y(exu_n11600));
AND2X1 exu_U31824(.A(tlu_exu_ccr_m[6]), .B(tlu_exu_cwpccr_update_m), .Y(ecl_ccr_mux_ccr_m_n14));
INVX1 exu_U31825(.A(ecl_ccr_mux_ccr_m_n14), .Y(exu_n11601));
AND2X1 exu_U31826(.A(tlu_exu_ccr_m[7]), .B(tlu_exu_cwpccr_update_m), .Y(ecl_ccr_mux_ccr_m_n16));
INVX1 exu_U31827(.A(ecl_ccr_mux_ccr_m_n16), .Y(exu_n11602));
AND2X1 exu_U31828(.A(rml_new_agp[0]), .B(exu_n15486), .Y(rml_agp_next0_mux_n2));
INVX1 exu_U31829(.A(rml_agp_next0_mux_n2), .Y(exu_n11603));
AND2X1 exu_U31830(.A(rml_new_agp[1]), .B(exu_n15486), .Y(rml_agp_next0_mux_n4));
INVX1 exu_U31831(.A(rml_agp_next0_mux_n4), .Y(exu_n11604));
AND2X1 exu_U31832(.A(exu_n16589), .B(rml_cansave_wen_e), .Y(rml_next_cansave_mux_n2));
INVX1 exu_U31833(.A(rml_next_cansave_mux_n2), .Y(exu_n11605));
AND2X1 exu_U31834(.A(rml_rml_next_cansave_e[1]), .B(rml_cansave_wen_e), .Y(rml_next_cansave_mux_n4));
INVX1 exu_U31835(.A(rml_next_cansave_mux_n4), .Y(exu_n11606));
AND2X1 exu_U31836(.A(rml_rml_next_cansave_e[2]), .B(rml_cansave_wen_e), .Y(rml_next_cansave_mux_n6));
INVX1 exu_U31837(.A(rml_next_cansave_mux_n6), .Y(exu_n11607));
OR2X1 exu_U31838(.A(rml_cwp_n96), .B(rml_swap_locals_ins), .Y(rml_cwp_n25));
INVX1 exu_U31839(.A(rml_cwp_n25), .Y(exu_n11608));
OR2X1 exu_U31840(.A(exu_n15417), .B(exu_n15340), .Y(rml_cwp_swap_next_state[3]));
INVX1 exu_U31841(.A(rml_cwp_swap_next_state[3]), .Y(exu_n11609));
OR2X1 exu_U31842(.A(exu_n15416), .B(exu_n15341), .Y(rml_cwp_swap_next_state[2]));
INVX1 exu_U31843(.A(rml_cwp_swap_next_state[2]), .Y(exu_n11610));
OR2X1 exu_U31844(.A(exu_n15415), .B(exu_n15342), .Y(rml_cwp_swap_next_state[1]));
INVX1 exu_U31845(.A(rml_cwp_swap_next_state[1]), .Y(exu_n11611));
AND2X1 exu_U31846(.A(rml_rml_ecl_cwp_e[2]), .B(exu_n15027), .Y(rml_cwp_n53));
INVX1 exu_U31847(.A(rml_cwp_n53), .Y(exu_n11612));
AND2X1 exu_U31848(.A(rml_rml_ecl_cwp_e[1]), .B(exu_n15027), .Y(rml_cwp_n55));
INVX1 exu_U31849(.A(rml_cwp_n55), .Y(exu_n11613));
AND2X1 exu_U31850(.A(rml_rml_ecl_cwp_e[0]), .B(exu_n15027), .Y(rml_cwp_n57));
INVX1 exu_U31851(.A(rml_cwp_n57), .Y(exu_n11614));
AND2X1 exu_U31852(.A(exu_n15851), .B(exu_n15027), .Y(rml_cwp_n59));
INVX1 exu_U31853(.A(rml_cwp_n59), .Y(exu_n11615));
AND2X1 exu_U31854(.A(exu_n15852), .B(exu_n15027), .Y(rml_cwp_n61));
INVX1 exu_U31855(.A(rml_cwp_n61), .Y(exu_n11616));
AND2X1 exu_U31856(.A(exu_n15853), .B(exu_n15027), .Y(rml_cwp_n63));
INVX1 exu_U31857(.A(rml_cwp_n63), .Y(exu_n11617));
OR2X1 exu_U31858(.A(ecl_alu_sethi_inst_e), .B(exu_n16551), .Y(alu_logic_mov_data[63]));
INVX1 exu_U31859(.A(alu_logic_mov_data[63]), .Y(exu_n11618));
OR2X1 exu_U31860(.A(ecl_alu_sethi_inst_e), .B(exu_n16550), .Y(alu_logic_mov_data[62]));
INVX1 exu_U31861(.A(alu_logic_mov_data[62]), .Y(exu_n11619));
OR2X1 exu_U31862(.A(ecl_alu_sethi_inst_e), .B(exu_n16549), .Y(alu_logic_mov_data[61]));
INVX1 exu_U31863(.A(alu_logic_mov_data[61]), .Y(exu_n11620));
OR2X1 exu_U31864(.A(ecl_alu_sethi_inst_e), .B(exu_n16548), .Y(alu_logic_mov_data[60]));
INVX1 exu_U31865(.A(alu_logic_mov_data[60]), .Y(exu_n11621));
OR2X1 exu_U31866(.A(ecl_alu_sethi_inst_e), .B(exu_n16547), .Y(alu_logic_mov_data[59]));
INVX1 exu_U31867(.A(alu_logic_mov_data[59]), .Y(exu_n11622));
OR2X1 exu_U31868(.A(ecl_alu_sethi_inst_e), .B(exu_n16546), .Y(alu_logic_mov_data[58]));
INVX1 exu_U31869(.A(alu_logic_mov_data[58]), .Y(exu_n11623));
OR2X1 exu_U31870(.A(ecl_alu_sethi_inst_e), .B(exu_n16545), .Y(alu_logic_mov_data[57]));
INVX1 exu_U31871(.A(alu_logic_mov_data[57]), .Y(exu_n11624));
OR2X1 exu_U31872(.A(ecl_alu_sethi_inst_e), .B(exu_n16544), .Y(alu_logic_mov_data[56]));
INVX1 exu_U31873(.A(alu_logic_mov_data[56]), .Y(exu_n11625));
OR2X1 exu_U31874(.A(ecl_alu_sethi_inst_e), .B(exu_n16543), .Y(alu_logic_mov_data[55]));
INVX1 exu_U31875(.A(alu_logic_mov_data[55]), .Y(exu_n11626));
OR2X1 exu_U31876(.A(ecl_alu_sethi_inst_e), .B(exu_n16542), .Y(alu_logic_mov_data[54]));
INVX1 exu_U31877(.A(alu_logic_mov_data[54]), .Y(exu_n11627));
OR2X1 exu_U31878(.A(ecl_alu_sethi_inst_e), .B(exu_n16541), .Y(alu_logic_mov_data[53]));
INVX1 exu_U31879(.A(alu_logic_mov_data[53]), .Y(exu_n11628));
OR2X1 exu_U31880(.A(ecl_alu_sethi_inst_e), .B(exu_n16540), .Y(alu_logic_mov_data[52]));
INVX1 exu_U31881(.A(alu_logic_mov_data[52]), .Y(exu_n11629));
OR2X1 exu_U31882(.A(ecl_alu_sethi_inst_e), .B(exu_n16539), .Y(alu_logic_mov_data[51]));
INVX1 exu_U31883(.A(alu_logic_mov_data[51]), .Y(exu_n11630));
OR2X1 exu_U31884(.A(ecl_alu_sethi_inst_e), .B(exu_n16538), .Y(alu_logic_mov_data[50]));
INVX1 exu_U31885(.A(alu_logic_mov_data[50]), .Y(exu_n11631));
OR2X1 exu_U31886(.A(ecl_alu_sethi_inst_e), .B(exu_n16537), .Y(alu_logic_mov_data[49]));
INVX1 exu_U31887(.A(alu_logic_mov_data[49]), .Y(exu_n11632));
OR2X1 exu_U31888(.A(ecl_alu_sethi_inst_e), .B(exu_n16536), .Y(alu_logic_mov_data[48]));
INVX1 exu_U31889(.A(alu_logic_mov_data[48]), .Y(exu_n11633));
OR2X1 exu_U31890(.A(ecl_alu_sethi_inst_e), .B(exu_n16535), .Y(alu_logic_mov_data[47]));
INVX1 exu_U31891(.A(alu_logic_mov_data[47]), .Y(exu_n11634));
OR2X1 exu_U31892(.A(ecl_alu_sethi_inst_e), .B(exu_n16534), .Y(alu_logic_mov_data[46]));
INVX1 exu_U31893(.A(alu_logic_mov_data[46]), .Y(exu_n11635));
OR2X1 exu_U31894(.A(ecl_alu_sethi_inst_e), .B(exu_n16533), .Y(alu_logic_mov_data[45]));
INVX1 exu_U31895(.A(alu_logic_mov_data[45]), .Y(exu_n11636));
OR2X1 exu_U31896(.A(ecl_alu_sethi_inst_e), .B(exu_n16532), .Y(alu_logic_mov_data[44]));
INVX1 exu_U31897(.A(alu_logic_mov_data[44]), .Y(exu_n11637));
OR2X1 exu_U31898(.A(ecl_alu_sethi_inst_e), .B(exu_n16531), .Y(alu_logic_mov_data[43]));
INVX1 exu_U31899(.A(alu_logic_mov_data[43]), .Y(exu_n11638));
OR2X1 exu_U31900(.A(ecl_alu_sethi_inst_e), .B(exu_n16530), .Y(alu_logic_mov_data[42]));
INVX1 exu_U31901(.A(alu_logic_mov_data[42]), .Y(exu_n11639));
OR2X1 exu_U31902(.A(ecl_alu_sethi_inst_e), .B(exu_n16529), .Y(alu_logic_mov_data[41]));
INVX1 exu_U31903(.A(alu_logic_mov_data[41]), .Y(exu_n11640));
OR2X1 exu_U31904(.A(ecl_alu_sethi_inst_e), .B(exu_n16528), .Y(alu_logic_mov_data[40]));
INVX1 exu_U31905(.A(alu_logic_mov_data[40]), .Y(exu_n11641));
OR2X1 exu_U31906(.A(ecl_alu_sethi_inst_e), .B(exu_n16527), .Y(alu_logic_mov_data[39]));
INVX1 exu_U31907(.A(alu_logic_mov_data[39]), .Y(exu_n11642));
OR2X1 exu_U31908(.A(ecl_alu_sethi_inst_e), .B(exu_n16526), .Y(alu_logic_mov_data[38]));
INVX1 exu_U31909(.A(alu_logic_mov_data[38]), .Y(exu_n11643));
OR2X1 exu_U31910(.A(ecl_alu_sethi_inst_e), .B(exu_n16525), .Y(alu_logic_mov_data[37]));
INVX1 exu_U31911(.A(alu_logic_mov_data[37]), .Y(exu_n11644));
OR2X1 exu_U31912(.A(ecl_alu_sethi_inst_e), .B(exu_n16524), .Y(alu_logic_mov_data[36]));
INVX1 exu_U31913(.A(alu_logic_mov_data[36]), .Y(exu_n11645));
OR2X1 exu_U31914(.A(ecl_alu_sethi_inst_e), .B(exu_n16523), .Y(alu_logic_mov_data[35]));
INVX1 exu_U31915(.A(alu_logic_mov_data[35]), .Y(exu_n11646));
OR2X1 exu_U31916(.A(ecl_alu_sethi_inst_e), .B(exu_n16522), .Y(alu_logic_mov_data[34]));
INVX1 exu_U31917(.A(alu_logic_mov_data[34]), .Y(exu_n11647));
OR2X1 exu_U31918(.A(ecl_alu_sethi_inst_e), .B(exu_n16521), .Y(alu_logic_mov_data[33]));
INVX1 exu_U31919(.A(alu_logic_mov_data[33]), .Y(exu_n11648));
OR2X1 exu_U31920(.A(ecl_alu_sethi_inst_e), .B(exu_n16520), .Y(alu_logic_mov_data[32]));
INVX1 exu_U31921(.A(alu_logic_mov_data[32]), .Y(exu_n11649));
AND2X1 exu_U31922(.A(ecl_mdqctl_mul_data[9]), .B(exu_n16388), .Y(ecl_mdqctl_n26));
INVX1 exu_U31923(.A(ecl_mdqctl_n26), .Y(exu_n11650));
AND2X1 exu_U31924(.A(ecl_mdqctl_mul_data[8]), .B(exu_n16388), .Y(ecl_mdqctl_n28));
INVX1 exu_U31925(.A(ecl_mdqctl_n28), .Y(exu_n11651));
AND2X1 exu_U31926(.A(ecl_mdqctl_wb_mulsetcc_g), .B(exu_n16388), .Y(ecl_mdqctl_n30));
INVX1 exu_U31927(.A(ecl_mdqctl_n30), .Y(exu_n11652));
AND2X1 exu_U31928(.A(ifu_exu_rd_d[4]), .B(ifu_exu_muldivop_d[4]), .Y(ecl_mdqctl_n32));
INVX1 exu_U31929(.A(ecl_mdqctl_n32), .Y(exu_n11653));
AND2X1 exu_U31930(.A(ifu_exu_rd_d[3]), .B(ifu_exu_muldivop_d[4]), .Y(ecl_mdqctl_n34));
INVX1 exu_U31931(.A(ecl_mdqctl_n34), .Y(exu_n11654));
AND2X1 exu_U31932(.A(ifu_exu_rd_d[2]), .B(ifu_exu_muldivop_d[4]), .Y(ecl_mdqctl_n36));
INVX1 exu_U31933(.A(ecl_mdqctl_n36), .Y(exu_n11655));
AND2X1 exu_U31934(.A(ifu_exu_rd_d[1]), .B(ifu_exu_muldivop_d[4]), .Y(ecl_mdqctl_n38));
INVX1 exu_U31935(.A(ecl_mdqctl_n38), .Y(exu_n11656));
AND2X1 exu_U31936(.A(ifu_exu_rd_d[0]), .B(ifu_exu_muldivop_d[4]), .Y(ecl_mdqctl_n40));
INVX1 exu_U31937(.A(ecl_mdqctl_n40), .Y(exu_n11657));
AND2X1 exu_U31938(.A(ecl_tid_d[1]), .B(ifu_exu_muldivop_d[4]), .Y(ecl_mdqctl_n42));
INVX1 exu_U31939(.A(ecl_mdqctl_n42), .Y(exu_n11658));
AND2X1 exu_U31940(.A(ecl_tid_d[0]), .B(ifu_exu_muldivop_d[4]), .Y(ecl_mdqctl_n44));
INVX1 exu_U31941(.A(ecl_mdqctl_n44), .Y(exu_n11659));
OR2X1 exu_U31942(.A(exu_n16607), .B(ecl_mdqctl_n50), .Y(ecl_mdqctl_n48));
INVX1 exu_U31943(.A(ecl_mdqctl_n48), .Y(exu_n11660));
OR2X1 exu_U31944(.A(ecl_mdqctl_n46), .B(ecl_mdqctl_n54), .Y(ecl_mdqctl_curr_div_vld));
INVX1 exu_U31945(.A(ecl_mdqctl_curr_div_vld), .Y(exu_n11661));
INVX1 exu_U31946(.A(ecl_ccr_n35), .Y(exu_n11662));
OR2X1 exu_U31947(.A(ecl_ifu_tlu_flush_w), .B(ecl_rml_early_flush_w), .Y(ecl_ccr_n35));
OR2X1 exu_U31948(.A(exu_n16607), .B(ecl_mdqctl_n62), .Y(ecl_mdqctl_n60));
INVX1 exu_U31949(.A(ecl_mdqctl_n60), .Y(exu_n11663));
AND2X1 exu_U31950(.A(ecl_divcntl_div_state_0), .B(exu_n16213), .Y(ecl_divcntl_n32));
INVX1 exu_U31951(.A(ecl_divcntl_n32), .Y(exu_n11664));
AND2X1 exu_U31952(.A(exu_n11666), .B(ecl_divcntl_div_adder_out_31_w), .Y(ecl_divcntl_n41));
INVX1 exu_U31953(.A(ecl_divcntl_n41), .Y(exu_n11665));
OR2X1 exu_U31954(.A(ecl_divcntl_rs2_data_31_w), .B(ecl_divcntl_muls_rs1_data_31_w), .Y(ecl_divcntl_n44));
INVX1 exu_U31955(.A(ecl_divcntl_n44), .Y(exu_n11666));
AND2X1 exu_U31956(.A(ecl_divcntl_muls_v), .B(exu_n16504), .Y(ecl_divcntl_n38));
INVX1 exu_U31957(.A(ecl_divcntl_n38), .Y(exu_n11667));
AND2X1 exu_U31958(.A(ecl_divcntl_muls_c), .B(exu_n16438), .Y(ecl_divcntl_n45));
INVX1 exu_U31959(.A(ecl_divcntl_n45), .Y(exu_n11668));
OR2X1 exu_U31960(.A(ecl_ifu_exu_rs2_d[1]), .B(ecl_ifu_exu_rs2_d[0]), .Y(ecl_byplog_rs2_n49));
INVX1 exu_U31961(.A(ecl_byplog_rs2_n49), .Y(exu_n11669));
OR2X1 exu_U31962(.A(exu_n15769), .B(ecl_byplog_rs1_n24), .Y(ecl_byplog_rs1_n16));
INVX1 exu_U31963(.A(ecl_byplog_rs1_n16), .Y(exu_n11670));
AND2X1 exu_U31964(.A(ecl_eccctl_gl_m[1]), .B(exu_n15481), .Y(ecl_eccctl_n23));
INVX1 exu_U31965(.A(ecl_eccctl_n23), .Y(exu_n11671));
AND2X1 exu_U31966(.A(ecl_eccctl_gl_m[0]), .B(exu_n15481), .Y(ecl_eccctl_n26));
INVX1 exu_U31967(.A(ecl_eccctl_n26), .Y(exu_n11672));
OR2X1 exu_U31968(.A(ecl_eccctl_rs3_ue_m), .B(ecl_eccctl_rs1_ce_m), .Y(ecl_eccctl_n33));
INVX1 exu_U31969(.A(ecl_eccctl_n33), .Y(exu_n11673));
INVX1 exu_U31970(.A(ecl_writeback_n47), .Y(exu_n11674));
AND2X1 exu_U31971(.A(ecl_writeback_n167), .B(ecl_writeback_n51), .Y(ecl_writeback_n48));
INVX1 exu_U31972(.A(ecl_writeback_n48), .Y(exu_n11675));
AND2X1 exu_U31973(.A(sehold), .B(exu_n15031), .Y(ecl_writeback_n45));
INVX1 exu_U31974(.A(ecl_writeback_n45), .Y(exu_n11676));
OR2X1 exu_U31975(.A(ecl_writeback_restore_tid[0]), .B(exu_n15545), .Y(ecl_writeback_n109));
INVX1 exu_U31976(.A(ecl_writeback_n109), .Y(exu_n11677));
OR2X1 exu_U31977(.A(ecl_writeback_restore_tid[1]), .B(exu_n15545), .Y(ecl_writeback_n117));
INVX1 exu_U31978(.A(ecl_writeback_n117), .Y(exu_n11678));
OR2X1 exu_U31979(.A(ecl_writeback_restore_tid[1]), .B(ecl_writeback_restore_tid[0]), .Y(ecl_writeback_n128));
INVX1 exu_U31980(.A(ecl_writeback_n128), .Y(exu_n11679));
OR2X1 exu_U31981(.A(ecl_writeback_n148), .B(ecl_writeback_wen_no_inst_vld_w), .Y(ecl_writeback_n146));
INVX1 exu_U31982(.A(ecl_writeback_n146), .Y(exu_n11680));
INVX1 exu_U31983(.A(ecl_writeback_n152), .Y(exu_n11681));
OR2X1 exu_U31984(.A(exu_n16398), .B(exu_n15395), .Y(ecl_writeback_n162));
INVX1 exu_U31985(.A(ecl_writeback_n162), .Y(exu_n11682));
AND2X1 exu_U31986(.A(ecl_wb_byplog_wen_w2), .B(sehold), .Y(ecl_writeback_n150));
INVX1 exu_U31987(.A(ecl_writeback_n150), .Y(exu_n11683));
INVX1 exu_U31988(.A(ecl_writeback_n166), .Y(exu_n11684));
AND2X1 exu_U31989(.A(ecl_tid_m[1]), .B(exu_n15761), .Y(ecl_writeback_n168));
INVX1 exu_U31990(.A(ecl_writeback_n168), .Y(exu_n11685));
AND2X1 exu_U31991(.A(exu_n15764), .B(ecl_writeback_dfill_tid_g2[1]), .Y(ecl_writeback_n164));
INVX1 exu_U31992(.A(ecl_writeback_n164), .Y(exu_n11686));
INVX1 exu_U31993(.A(ecl_writeback_n172), .Y(exu_n11687));
AND2X1 exu_U31994(.A(ecl_tid_m[0]), .B(exu_n15761), .Y(ecl_writeback_n173));
INVX1 exu_U31995(.A(ecl_writeback_n173), .Y(exu_n11688));
AND2X1 exu_U31996(.A(ecl_writeback_n167), .B(ecl_writeback_dfill_tid_g2[0]), .Y(ecl_writeback_n170));
INVX1 exu_U31997(.A(ecl_writeback_n170), .Y(exu_n11689));
OR2X1 exu_U31998(.A(ecc_rs1_err_e[0]), .B(ecc_chk_rs1_n9), .Y(ecc_chk_rs1_n5));
INVX1 exu_U31999(.A(ecc_chk_rs1_n5), .Y(exu_n11690));
INVX1 exu_U32000(.A(bypass_full_rd_data_m[8]), .Y(exu_n11691));
INVX1 exu_U32001(.A(bypass_full_rd_data_m[7]), .Y(exu_n11692));
INVX1 exu_U32002(.A(bypass_full_rd_data_m[6]), .Y(exu_n11693));
INVX1 exu_U32003(.A(bypass_full_rd_data_m[63]), .Y(exu_n11694));
INVX1 exu_U32004(.A(bypass_full_rd_data_m[62]), .Y(exu_n11695));
INVX1 exu_U32005(.A(bypass_full_rd_data_m[61]), .Y(exu_n11696));
INVX1 exu_U32006(.A(bypass_full_rd_data_m[60]), .Y(exu_n11697));
INVX1 exu_U32007(.A(bypass_full_rd_data_m[5]), .Y(exu_n11698));
INVX1 exu_U32008(.A(bypass_full_rd_data_m[59]), .Y(exu_n11699));
INVX1 exu_U32009(.A(bypass_full_rd_data_m[58]), .Y(exu_n11700));
INVX1 exu_U32010(.A(bypass_full_rd_data_m[57]), .Y(exu_n11701));
INVX1 exu_U32011(.A(bypass_full_rd_data_m[56]), .Y(exu_n11702));
INVX1 exu_U32012(.A(bypass_full_rd_data_m[55]), .Y(exu_n11703));
INVX1 exu_U32013(.A(bypass_full_rd_data_m[54]), .Y(exu_n11704));
INVX1 exu_U32014(.A(bypass_full_rd_data_m[53]), .Y(exu_n11705));
INVX1 exu_U32015(.A(bypass_full_rd_data_m[52]), .Y(exu_n11706));
INVX1 exu_U32016(.A(bypass_full_rd_data_m[51]), .Y(exu_n11707));
INVX1 exu_U32017(.A(bypass_full_rd_data_m[50]), .Y(exu_n11708));
INVX1 exu_U32018(.A(bypass_full_rd_data_m[4]), .Y(exu_n11709));
INVX1 exu_U32019(.A(bypass_full_rd_data_m[49]), .Y(exu_n11710));
INVX1 exu_U32020(.A(bypass_full_rd_data_m[48]), .Y(exu_n11711));
INVX1 exu_U32021(.A(bypass_full_rd_data_m[47]), .Y(exu_n11712));
INVX1 exu_U32022(.A(bypass_full_rd_data_m[46]), .Y(exu_n11713));
INVX1 exu_U32023(.A(bypass_full_rd_data_m[45]), .Y(exu_n11714));
INVX1 exu_U32024(.A(bypass_full_rd_data_m[44]), .Y(exu_n11715));
INVX1 exu_U32025(.A(bypass_full_rd_data_m[43]), .Y(exu_n11716));
INVX1 exu_U32026(.A(bypass_full_rd_data_m[42]), .Y(exu_n11717));
INVX1 exu_U32027(.A(bypass_full_rd_data_m[41]), .Y(exu_n11718));
INVX1 exu_U32028(.A(bypass_full_rd_data_m[40]), .Y(exu_n11719));
INVX1 exu_U32029(.A(bypass_full_rd_data_m[3]), .Y(exu_n11720));
INVX1 exu_U32030(.A(bypass_full_rd_data_m[39]), .Y(exu_n11721));
INVX1 exu_U32031(.A(bypass_full_rd_data_m[38]), .Y(exu_n11722));
INVX1 exu_U32032(.A(bypass_full_rd_data_m[37]), .Y(exu_n11723));
INVX1 exu_U32033(.A(bypass_full_rd_data_m[36]), .Y(exu_n11724));
INVX1 exu_U32034(.A(bypass_full_rd_data_m[35]), .Y(exu_n11725));
INVX1 exu_U32035(.A(bypass_full_rd_data_m[34]), .Y(exu_n11726));
INVX1 exu_U32036(.A(bypass_full_rd_data_m[33]), .Y(exu_n11727));
INVX1 exu_U32037(.A(bypass_full_rd_data_m[32]), .Y(exu_n11728));
INVX1 exu_U32038(.A(bypass_full_rd_data_m[31]), .Y(exu_n11729));
INVX1 exu_U32039(.A(bypass_full_rd_data_m[30]), .Y(exu_n11730));
INVX1 exu_U32040(.A(bypass_full_rd_data_m[2]), .Y(exu_n11731));
INVX1 exu_U32041(.A(bypass_full_rd_data_m[29]), .Y(exu_n11732));
INVX1 exu_U32042(.A(bypass_full_rd_data_m[28]), .Y(exu_n11733));
INVX1 exu_U32043(.A(bypass_full_rd_data_m[27]), .Y(exu_n11734));
INVX1 exu_U32044(.A(bypass_full_rd_data_m[26]), .Y(exu_n11735));
INVX1 exu_U32045(.A(bypass_full_rd_data_m[25]), .Y(exu_n11736));
INVX1 exu_U32046(.A(bypass_full_rd_data_m[24]), .Y(exu_n11737));
INVX1 exu_U32047(.A(bypass_full_rd_data_m[23]), .Y(exu_n11738));
INVX1 exu_U32048(.A(bypass_full_rd_data_m[22]), .Y(exu_n11739));
INVX1 exu_U32049(.A(bypass_full_rd_data_m[21]), .Y(exu_n11740));
INVX1 exu_U32050(.A(bypass_full_rd_data_m[20]), .Y(exu_n11741));
INVX1 exu_U32051(.A(bypass_full_rd_data_m[1]), .Y(exu_n11742));
INVX1 exu_U32052(.A(bypass_full_rd_data_m[19]), .Y(exu_n11743));
INVX1 exu_U32053(.A(bypass_full_rd_data_m[18]), .Y(exu_n11744));
INVX1 exu_U32054(.A(bypass_full_rd_data_m[17]), .Y(exu_n11745));
INVX1 exu_U32055(.A(bypass_full_rd_data_m[16]), .Y(exu_n11746));
INVX1 exu_U32056(.A(bypass_full_rd_data_m[15]), .Y(exu_n11747));
INVX1 exu_U32057(.A(bypass_full_rd_data_m[14]), .Y(exu_n11748));
INVX1 exu_U32058(.A(bypass_full_rd_data_m[13]), .Y(exu_n11749));
INVX1 exu_U32059(.A(bypass_full_rd_data_m[12]), .Y(exu_n11750));
INVX1 exu_U32060(.A(bypass_full_rd_data_m[11]), .Y(exu_n11751));
INVX1 exu_U32061(.A(bypass_full_rd_data_m[10]), .Y(exu_n11752));
INVX1 exu_U32062(.A(bypass_full_rd_data_m[0]), .Y(exu_n11753));
AND2X1 exu_U32063(.A(alu_byp_rd_data_e[63]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n27));
INVX1 exu_U32064(.A(bypass_ifu_exu_sr_mux_n27), .Y(exu_n11754));
AND2X1 exu_U32065(.A(alu_byp_rd_data_e[62]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n33));
INVX1 exu_U32066(.A(bypass_ifu_exu_sr_mux_n33), .Y(exu_n11755));
AND2X1 exu_U32067(.A(alu_byp_rd_data_e[61]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n39));
INVX1 exu_U32068(.A(bypass_ifu_exu_sr_mux_n39), .Y(exu_n11756));
AND2X1 exu_U32069(.A(alu_byp_rd_data_e[60]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n45));
INVX1 exu_U32070(.A(bypass_ifu_exu_sr_mux_n45), .Y(exu_n11757));
AND2X1 exu_U32071(.A(alu_byp_rd_data_e[59]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n57));
INVX1 exu_U32072(.A(bypass_ifu_exu_sr_mux_n57), .Y(exu_n11758));
AND2X1 exu_U32073(.A(alu_byp_rd_data_e[58]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n63));
INVX1 exu_U32074(.A(bypass_ifu_exu_sr_mux_n63), .Y(exu_n11759));
AND2X1 exu_U32075(.A(alu_byp_rd_data_e[57]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n69));
INVX1 exu_U32076(.A(bypass_ifu_exu_sr_mux_n69), .Y(exu_n11760));
AND2X1 exu_U32077(.A(alu_byp_rd_data_e[56]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n75));
INVX1 exu_U32078(.A(bypass_ifu_exu_sr_mux_n75), .Y(exu_n11761));
AND2X1 exu_U32079(.A(alu_byp_rd_data_e[55]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n81));
INVX1 exu_U32080(.A(bypass_ifu_exu_sr_mux_n81), .Y(exu_n11762));
AND2X1 exu_U32081(.A(alu_byp_rd_data_e[54]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n87));
INVX1 exu_U32082(.A(bypass_ifu_exu_sr_mux_n87), .Y(exu_n11763));
AND2X1 exu_U32083(.A(alu_byp_rd_data_e[53]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n93));
INVX1 exu_U32084(.A(bypass_ifu_exu_sr_mux_n93), .Y(exu_n11764));
AND2X1 exu_U32085(.A(alu_byp_rd_data_e[52]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n99));
INVX1 exu_U32086(.A(bypass_ifu_exu_sr_mux_n99), .Y(exu_n11765));
AND2X1 exu_U32087(.A(alu_byp_rd_data_e[51]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n105));
INVX1 exu_U32088(.A(bypass_ifu_exu_sr_mux_n105), .Y(exu_n11766));
AND2X1 exu_U32089(.A(alu_byp_rd_data_e[50]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n111));
INVX1 exu_U32090(.A(bypass_ifu_exu_sr_mux_n111), .Y(exu_n11767));
AND2X1 exu_U32091(.A(alu_byp_rd_data_e[49]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n123));
INVX1 exu_U32092(.A(bypass_ifu_exu_sr_mux_n123), .Y(exu_n11768));
AND2X1 exu_U32093(.A(alu_byp_rd_data_e[48]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n129));
INVX1 exu_U32094(.A(bypass_ifu_exu_sr_mux_n129), .Y(exu_n11769));
AND2X1 exu_U32095(.A(alu_byp_rd_data_e[47]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n135));
INVX1 exu_U32096(.A(bypass_ifu_exu_sr_mux_n135), .Y(exu_n11770));
AND2X1 exu_U32097(.A(alu_byp_rd_data_e[46]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n141));
INVX1 exu_U32098(.A(bypass_ifu_exu_sr_mux_n141), .Y(exu_n11771));
AND2X1 exu_U32099(.A(alu_byp_rd_data_e[45]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n147));
INVX1 exu_U32100(.A(bypass_ifu_exu_sr_mux_n147), .Y(exu_n11772));
AND2X1 exu_U32101(.A(alu_byp_rd_data_e[44]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n153));
INVX1 exu_U32102(.A(bypass_ifu_exu_sr_mux_n153), .Y(exu_n11773));
AND2X1 exu_U32103(.A(alu_byp_rd_data_e[43]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n159));
INVX1 exu_U32104(.A(bypass_ifu_exu_sr_mux_n159), .Y(exu_n11774));
AND2X1 exu_U32105(.A(alu_byp_rd_data_e[42]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n165));
INVX1 exu_U32106(.A(bypass_ifu_exu_sr_mux_n165), .Y(exu_n11775));
AND2X1 exu_U32107(.A(alu_byp_rd_data_e[41]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n171));
INVX1 exu_U32108(.A(bypass_ifu_exu_sr_mux_n171), .Y(exu_n11776));
AND2X1 exu_U32109(.A(alu_byp_rd_data_e[40]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n177));
INVX1 exu_U32110(.A(bypass_ifu_exu_sr_mux_n177), .Y(exu_n11777));
AND2X1 exu_U32111(.A(alu_byp_rd_data_e[39]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n189));
INVX1 exu_U32112(.A(bypass_ifu_exu_sr_mux_n189), .Y(exu_n11778));
AND2X1 exu_U32113(.A(alu_byp_rd_data_e[38]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n195));
INVX1 exu_U32114(.A(bypass_ifu_exu_sr_mux_n195), .Y(exu_n11779));
AND2X1 exu_U32115(.A(alu_byp_rd_data_e[37]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n201));
INVX1 exu_U32116(.A(bypass_ifu_exu_sr_mux_n201), .Y(exu_n11780));
AND2X1 exu_U32117(.A(alu_byp_rd_data_e[36]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n207));
INVX1 exu_U32118(.A(bypass_ifu_exu_sr_mux_n207), .Y(exu_n11781));
AND2X1 exu_U32119(.A(alu_byp_rd_data_e[35]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n213));
INVX1 exu_U32120(.A(bypass_ifu_exu_sr_mux_n213), .Y(exu_n11782));
AND2X1 exu_U32121(.A(alu_byp_rd_data_e[34]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n219));
INVX1 exu_U32122(.A(bypass_ifu_exu_sr_mux_n219), .Y(exu_n11783));
AND2X1 exu_U32123(.A(alu_byp_rd_data_e[33]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n225));
INVX1 exu_U32124(.A(bypass_ifu_exu_sr_mux_n225), .Y(exu_n11784));
AND2X1 exu_U32125(.A(alu_byp_rd_data_e[32]), .B(ecl_byp_sel_alu_e), .Y(bypass_ifu_exu_sr_mux_n231));
INVX1 exu_U32126(.A(bypass_ifu_exu_sr_mux_n231), .Y(exu_n11785));
AND2X1 exu_U32127(.A(exu_n16269), .B(lsu_exu_ldxa_data_g[9]), .Y(bypass_dfill_data_mux_n2));
INVX1 exu_U32128(.A(bypass_dfill_data_mux_n2), .Y(exu_n11786));
AND2X1 exu_U32129(.A(lsu_exu_ldxa_data_g[8]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n4));
INVX1 exu_U32130(.A(bypass_dfill_data_mux_n4), .Y(exu_n11787));
AND2X1 exu_U32131(.A(lsu_exu_ldxa_data_g[7]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n6));
INVX1 exu_U32132(.A(bypass_dfill_data_mux_n6), .Y(exu_n11788));
AND2X1 exu_U32133(.A(lsu_exu_ldxa_data_g[6]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n8));
INVX1 exu_U32134(.A(bypass_dfill_data_mux_n8), .Y(exu_n11789));
AND2X1 exu_U32135(.A(lsu_exu_ldxa_data_g[63]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n10));
INVX1 exu_U32136(.A(bypass_dfill_data_mux_n10), .Y(exu_n11790));
AND2X1 exu_U32137(.A(lsu_exu_ldxa_data_g[62]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n12));
INVX1 exu_U32138(.A(bypass_dfill_data_mux_n12), .Y(exu_n11791));
AND2X1 exu_U32139(.A(lsu_exu_ldxa_data_g[61]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n14));
INVX1 exu_U32140(.A(bypass_dfill_data_mux_n14), .Y(exu_n11792));
AND2X1 exu_U32141(.A(lsu_exu_ldxa_data_g[60]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n16));
INVX1 exu_U32142(.A(bypass_dfill_data_mux_n16), .Y(exu_n11793));
AND2X1 exu_U32143(.A(lsu_exu_ldxa_data_g[5]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n18));
INVX1 exu_U32144(.A(bypass_dfill_data_mux_n18), .Y(exu_n11794));
AND2X1 exu_U32145(.A(lsu_exu_ldxa_data_g[59]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n20));
INVX1 exu_U32146(.A(bypass_dfill_data_mux_n20), .Y(exu_n11795));
AND2X1 exu_U32147(.A(lsu_exu_ldxa_data_g[58]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n22));
INVX1 exu_U32148(.A(bypass_dfill_data_mux_n22), .Y(exu_n11796));
AND2X1 exu_U32149(.A(lsu_exu_ldxa_data_g[57]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n24));
INVX1 exu_U32150(.A(bypass_dfill_data_mux_n24), .Y(exu_n11797));
AND2X1 exu_U32151(.A(lsu_exu_ldxa_data_g[56]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n26));
INVX1 exu_U32152(.A(bypass_dfill_data_mux_n26), .Y(exu_n11798));
AND2X1 exu_U32153(.A(lsu_exu_ldxa_data_g[55]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n28));
INVX1 exu_U32154(.A(bypass_dfill_data_mux_n28), .Y(exu_n11799));
AND2X1 exu_U32155(.A(lsu_exu_ldxa_data_g[54]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n30));
INVX1 exu_U32156(.A(bypass_dfill_data_mux_n30), .Y(exu_n11800));
AND2X1 exu_U32157(.A(lsu_exu_ldxa_data_g[53]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n32));
INVX1 exu_U32158(.A(bypass_dfill_data_mux_n32), .Y(exu_n11801));
AND2X1 exu_U32159(.A(lsu_exu_ldxa_data_g[52]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n34));
INVX1 exu_U32160(.A(bypass_dfill_data_mux_n34), .Y(exu_n11802));
AND2X1 exu_U32161(.A(lsu_exu_ldxa_data_g[51]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n36));
INVX1 exu_U32162(.A(bypass_dfill_data_mux_n36), .Y(exu_n11803));
AND2X1 exu_U32163(.A(lsu_exu_ldxa_data_g[50]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n38));
INVX1 exu_U32164(.A(bypass_dfill_data_mux_n38), .Y(exu_n11804));
AND2X1 exu_U32165(.A(lsu_exu_ldxa_data_g[4]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n40));
INVX1 exu_U32166(.A(bypass_dfill_data_mux_n40), .Y(exu_n11805));
AND2X1 exu_U32167(.A(lsu_exu_ldxa_data_g[49]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n42));
INVX1 exu_U32168(.A(bypass_dfill_data_mux_n42), .Y(exu_n11806));
AND2X1 exu_U32169(.A(lsu_exu_ldxa_data_g[48]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n44));
INVX1 exu_U32170(.A(bypass_dfill_data_mux_n44), .Y(exu_n11807));
AND2X1 exu_U32171(.A(lsu_exu_ldxa_data_g[47]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n46));
INVX1 exu_U32172(.A(bypass_dfill_data_mux_n46), .Y(exu_n11808));
AND2X1 exu_U32173(.A(lsu_exu_ldxa_data_g[46]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n48));
INVX1 exu_U32174(.A(bypass_dfill_data_mux_n48), .Y(exu_n11809));
AND2X1 exu_U32175(.A(lsu_exu_ldxa_data_g[45]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n50));
INVX1 exu_U32176(.A(bypass_dfill_data_mux_n50), .Y(exu_n11810));
AND2X1 exu_U32177(.A(lsu_exu_ldxa_data_g[44]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n52));
INVX1 exu_U32178(.A(bypass_dfill_data_mux_n52), .Y(exu_n11811));
AND2X1 exu_U32179(.A(lsu_exu_ldxa_data_g[43]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n54));
INVX1 exu_U32180(.A(bypass_dfill_data_mux_n54), .Y(exu_n11812));
AND2X1 exu_U32181(.A(lsu_exu_ldxa_data_g[42]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n56));
INVX1 exu_U32182(.A(bypass_dfill_data_mux_n56), .Y(exu_n11813));
AND2X1 exu_U32183(.A(lsu_exu_ldxa_data_g[41]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n58));
INVX1 exu_U32184(.A(bypass_dfill_data_mux_n58), .Y(exu_n11814));
AND2X1 exu_U32185(.A(lsu_exu_ldxa_data_g[40]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n60));
INVX1 exu_U32186(.A(bypass_dfill_data_mux_n60), .Y(exu_n11815));
AND2X1 exu_U32187(.A(lsu_exu_ldxa_data_g[3]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n62));
INVX1 exu_U32188(.A(bypass_dfill_data_mux_n62), .Y(exu_n11816));
AND2X1 exu_U32189(.A(lsu_exu_ldxa_data_g[39]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n64));
INVX1 exu_U32190(.A(bypass_dfill_data_mux_n64), .Y(exu_n11817));
AND2X1 exu_U32191(.A(lsu_exu_ldxa_data_g[38]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n66));
INVX1 exu_U32192(.A(bypass_dfill_data_mux_n66), .Y(exu_n11818));
AND2X1 exu_U32193(.A(lsu_exu_ldxa_data_g[37]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n68));
INVX1 exu_U32194(.A(bypass_dfill_data_mux_n68), .Y(exu_n11819));
AND2X1 exu_U32195(.A(lsu_exu_ldxa_data_g[36]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n70));
INVX1 exu_U32196(.A(bypass_dfill_data_mux_n70), .Y(exu_n11820));
AND2X1 exu_U32197(.A(lsu_exu_ldxa_data_g[35]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n72));
INVX1 exu_U32198(.A(bypass_dfill_data_mux_n72), .Y(exu_n11821));
AND2X1 exu_U32199(.A(lsu_exu_ldxa_data_g[34]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n74));
INVX1 exu_U32200(.A(bypass_dfill_data_mux_n74), .Y(exu_n11822));
AND2X1 exu_U32201(.A(lsu_exu_ldxa_data_g[33]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n76));
INVX1 exu_U32202(.A(bypass_dfill_data_mux_n76), .Y(exu_n11823));
AND2X1 exu_U32203(.A(lsu_exu_ldxa_data_g[32]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n78));
INVX1 exu_U32204(.A(bypass_dfill_data_mux_n78), .Y(exu_n11824));
AND2X1 exu_U32205(.A(lsu_exu_ldxa_data_g[31]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n80));
INVX1 exu_U32206(.A(bypass_dfill_data_mux_n80), .Y(exu_n11825));
AND2X1 exu_U32207(.A(lsu_exu_ldxa_data_g[30]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n82));
INVX1 exu_U32208(.A(bypass_dfill_data_mux_n82), .Y(exu_n11826));
AND2X1 exu_U32209(.A(lsu_exu_ldxa_data_g[2]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n84));
INVX1 exu_U32210(.A(bypass_dfill_data_mux_n84), .Y(exu_n11827));
AND2X1 exu_U32211(.A(lsu_exu_ldxa_data_g[29]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n86));
INVX1 exu_U32212(.A(bypass_dfill_data_mux_n86), .Y(exu_n11828));
AND2X1 exu_U32213(.A(lsu_exu_ldxa_data_g[28]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n88));
INVX1 exu_U32214(.A(bypass_dfill_data_mux_n88), .Y(exu_n11829));
AND2X1 exu_U32215(.A(lsu_exu_ldxa_data_g[27]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n90));
INVX1 exu_U32216(.A(bypass_dfill_data_mux_n90), .Y(exu_n11830));
AND2X1 exu_U32217(.A(lsu_exu_ldxa_data_g[26]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n92));
INVX1 exu_U32218(.A(bypass_dfill_data_mux_n92), .Y(exu_n11831));
AND2X1 exu_U32219(.A(lsu_exu_ldxa_data_g[25]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n94));
INVX1 exu_U32220(.A(bypass_dfill_data_mux_n94), .Y(exu_n11832));
AND2X1 exu_U32221(.A(lsu_exu_ldxa_data_g[24]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n96));
INVX1 exu_U32222(.A(bypass_dfill_data_mux_n96), .Y(exu_n11833));
AND2X1 exu_U32223(.A(lsu_exu_ldxa_data_g[23]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n98));
INVX1 exu_U32224(.A(bypass_dfill_data_mux_n98), .Y(exu_n11834));
AND2X1 exu_U32225(.A(lsu_exu_ldxa_data_g[22]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n100));
INVX1 exu_U32226(.A(bypass_dfill_data_mux_n100), .Y(exu_n11835));
AND2X1 exu_U32227(.A(lsu_exu_ldxa_data_g[21]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n102));
INVX1 exu_U32228(.A(bypass_dfill_data_mux_n102), .Y(exu_n11836));
AND2X1 exu_U32229(.A(lsu_exu_ldxa_data_g[20]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n104));
INVX1 exu_U32230(.A(bypass_dfill_data_mux_n104), .Y(exu_n11837));
AND2X1 exu_U32231(.A(lsu_exu_ldxa_data_g[1]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n106));
INVX1 exu_U32232(.A(bypass_dfill_data_mux_n106), .Y(exu_n11838));
AND2X1 exu_U32233(.A(lsu_exu_ldxa_data_g[19]), .B(exu_n16269), .Y(bypass_dfill_data_mux_n108));
INVX1 exu_U32234(.A(bypass_dfill_data_mux_n108), .Y(exu_n11839));
AND2X1 exu_U32235(.A(lsu_exu_ldxa_data_g[18]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n110));
INVX1 exu_U32236(.A(bypass_dfill_data_mux_n110), .Y(exu_n11840));
AND2X1 exu_U32237(.A(lsu_exu_ldxa_data_g[17]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n112));
INVX1 exu_U32238(.A(bypass_dfill_data_mux_n112), .Y(exu_n11841));
AND2X1 exu_U32239(.A(lsu_exu_ldxa_data_g[16]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n114));
INVX1 exu_U32240(.A(bypass_dfill_data_mux_n114), .Y(exu_n11842));
AND2X1 exu_U32241(.A(lsu_exu_ldxa_data_g[15]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n116));
INVX1 exu_U32242(.A(bypass_dfill_data_mux_n116), .Y(exu_n11843));
AND2X1 exu_U32243(.A(lsu_exu_ldxa_data_g[14]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n118));
INVX1 exu_U32244(.A(bypass_dfill_data_mux_n118), .Y(exu_n11844));
AND2X1 exu_U32245(.A(lsu_exu_ldxa_data_g[13]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n120));
INVX1 exu_U32246(.A(bypass_dfill_data_mux_n120), .Y(exu_n11845));
AND2X1 exu_U32247(.A(lsu_exu_ldxa_data_g[12]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n122));
INVX1 exu_U32248(.A(bypass_dfill_data_mux_n122), .Y(exu_n11846));
AND2X1 exu_U32249(.A(lsu_exu_ldxa_data_g[11]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n124));
INVX1 exu_U32250(.A(bypass_dfill_data_mux_n124), .Y(exu_n11847));
AND2X1 exu_U32251(.A(lsu_exu_ldxa_data_g[10]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n126));
INVX1 exu_U32252(.A(bypass_dfill_data_mux_n126), .Y(exu_n11848));
AND2X1 exu_U32253(.A(lsu_exu_ldxa_data_g[0]), .B(ecl_byp_ldxa_g), .Y(bypass_dfill_data_mux_n128));
INVX1 exu_U32254(.A(bypass_dfill_data_mux_n128), .Y(exu_n11849));
OR2X1 exu_U32255(.A(exu_n16590), .B(exu_n15683), .Y(rml_n40));
INVX1 exu_U32256(.A(rml_n40), .Y(exu_n11850));
OR2X1 exu_U32257(.A(rml_rml_ecl_cwp_e[1]), .B(rml_rml_ecl_cansave_e[1]), .Y(rml_n42));
INVX1 exu_U32258(.A(rml_n42), .Y(exu_n11851));
INVX1 exu_U32259(.A(rml_rml_next_cleanwin_e[2]), .Y(exu_n11852));
AND2X1 exu_U32260(.A(exu_n15857), .B(rml_n49), .Y(rml_n46));
INVX1 exu_U32261(.A(rml_n46), .Y(exu_n11853));
AND2X1 exu_U32262(.A(rml_n49), .B(exu_n15856), .Y(rml_n53));
INVX1 exu_U32263(.A(rml_n53), .Y(exu_n11854));
AND2X1 exu_U32264(.A(rml_n84), .B(exu_n15921), .Y(rml_n81));
INVX1 exu_U32265(.A(rml_n81), .Y(exu_n11855));
AND2X1 exu_U32266(.A(exu_n15922), .B(rml_n84), .Y(rml_n85));
INVX1 exu_U32267(.A(rml_n85), .Y(exu_n11856));
AND2X1 exu_U32268(.A(exu_n15923), .B(rml_n84), .Y(rml_n88));
INVX1 exu_U32269(.A(rml_n88), .Y(exu_n11857));
AND2X1 exu_U32270(.A(exu_n15924), .B(rml_n84), .Y(rml_n91));
INVX1 exu_U32271(.A(rml_n91), .Y(exu_n11858));
OR2X1 exu_U32272(.A(rml_ecl_clean_window_e), .B(exu_n15343), .Y(rml_n113));
INVX1 exu_U32273(.A(rml_n113), .Y(exu_n11859));
OR2X1 exu_U32274(.A(rml_rml_ecl_cansave_e[0]), .B(exu_n16590), .Y(rml_n120));
INVX1 exu_U32275(.A(rml_n120), .Y(exu_n11860));
AND2X1 exu_U32276(.A(ecl_divcntl_n70), .B(exu_n16412), .Y(div_u32[8]));
INVX1 exu_U32277(.A(div_u32[8]), .Y(exu_n11861));
AND2X1 exu_U32278(.A(ecl_divcntl_n70), .B(exu_n16411), .Y(div_u32[7]));
INVX1 exu_U32279(.A(div_u32[7]), .Y(exu_n11862));
AND2X1 exu_U32280(.A(ecl_divcntl_n70), .B(exu_n16410), .Y(div_u32[6]));
INVX1 exu_U32281(.A(div_u32[6]), .Y(exu_n11863));
AND2X1 exu_U32282(.A(ecl_divcntl_n70), .B(exu_n16409), .Y(div_u32[5]));
INVX1 exu_U32283(.A(div_u32[5]), .Y(exu_n11864));
AND2X1 exu_U32284(.A(ecl_divcntl_n70), .B(exu_n16408), .Y(div_u32[4]));
INVX1 exu_U32285(.A(div_u32[4]), .Y(exu_n11865));
AND2X1 exu_U32286(.A(ecl_divcntl_n70), .B(exu_n16407), .Y(div_u32[3]));
INVX1 exu_U32287(.A(div_u32[3]), .Y(exu_n11866));
AND2X1 exu_U32288(.A(exu_n16435), .B(ecl_divcntl_n70), .Y(div_u32[31]));
INVX1 exu_U32289(.A(div_u32[31]), .Y(exu_n11867));
AND2X1 exu_U32290(.A(ecl_divcntl_n70), .B(exu_n16434), .Y(div_u32[30]));
INVX1 exu_U32291(.A(div_u32[30]), .Y(exu_n11868));
AND2X1 exu_U32292(.A(ecl_divcntl_n70), .B(exu_n16406), .Y(div_u32[2]));
INVX1 exu_U32293(.A(div_u32[2]), .Y(exu_n11869));
AND2X1 exu_U32294(.A(ecl_divcntl_n70), .B(exu_n16433), .Y(div_u32[29]));
INVX1 exu_U32295(.A(div_u32[29]), .Y(exu_n11870));
AND2X1 exu_U32296(.A(ecl_divcntl_n70), .B(exu_n16432), .Y(div_u32[28]));
INVX1 exu_U32297(.A(div_u32[28]), .Y(exu_n11871));
AND2X1 exu_U32298(.A(ecl_divcntl_n70), .B(exu_n16431), .Y(div_u32[27]));
INVX1 exu_U32299(.A(div_u32[27]), .Y(exu_n11872));
AND2X1 exu_U32300(.A(ecl_divcntl_n70), .B(exu_n16430), .Y(div_u32[26]));
INVX1 exu_U32301(.A(div_u32[26]), .Y(exu_n11873));
AND2X1 exu_U32302(.A(ecl_divcntl_n70), .B(exu_n16429), .Y(div_u32[25]));
INVX1 exu_U32303(.A(div_u32[25]), .Y(exu_n11874));
AND2X1 exu_U32304(.A(ecl_divcntl_n70), .B(exu_n16428), .Y(div_u32[24]));
INVX1 exu_U32305(.A(div_u32[24]), .Y(exu_n11875));
AND2X1 exu_U32306(.A(ecl_divcntl_n70), .B(exu_n16427), .Y(div_u32[23]));
INVX1 exu_U32307(.A(div_u32[23]), .Y(exu_n11876));
AND2X1 exu_U32308(.A(ecl_divcntl_n70), .B(exu_n16426), .Y(div_u32[22]));
INVX1 exu_U32309(.A(div_u32[22]), .Y(exu_n11877));
AND2X1 exu_U32310(.A(ecl_divcntl_n70), .B(exu_n16425), .Y(div_u32[21]));
INVX1 exu_U32311(.A(div_u32[21]), .Y(exu_n11878));
AND2X1 exu_U32312(.A(ecl_divcntl_n70), .B(exu_n16424), .Y(div_u32[20]));
INVX1 exu_U32313(.A(div_u32[20]), .Y(exu_n11879));
AND2X1 exu_U32314(.A(ecl_divcntl_n70), .B(exu_n16405), .Y(div_u32[1]));
INVX1 exu_U32315(.A(div_u32[1]), .Y(exu_n11880));
AND2X1 exu_U32316(.A(ecl_divcntl_n70), .B(exu_n16423), .Y(div_u32[19]));
INVX1 exu_U32317(.A(div_u32[19]), .Y(exu_n11881));
AND2X1 exu_U32318(.A(ecl_divcntl_n70), .B(exu_n16422), .Y(div_u32[18]));
INVX1 exu_U32319(.A(div_u32[18]), .Y(exu_n11882));
AND2X1 exu_U32320(.A(ecl_divcntl_n70), .B(exu_n16421), .Y(div_u32[17]));
INVX1 exu_U32321(.A(div_u32[17]), .Y(exu_n11883));
AND2X1 exu_U32322(.A(ecl_divcntl_n70), .B(exu_n16420), .Y(div_u32[16]));
INVX1 exu_U32323(.A(div_u32[16]), .Y(exu_n11884));
AND2X1 exu_U32324(.A(ecl_divcntl_n70), .B(exu_n16419), .Y(div_u32[15]));
INVX1 exu_U32325(.A(div_u32[15]), .Y(exu_n11885));
AND2X1 exu_U32326(.A(ecl_divcntl_n70), .B(exu_n16418), .Y(div_u32[14]));
INVX1 exu_U32327(.A(div_u32[14]), .Y(exu_n11886));
AND2X1 exu_U32328(.A(ecl_divcntl_n70), .B(exu_n16417), .Y(div_u32[13]));
INVX1 exu_U32329(.A(div_u32[13]), .Y(exu_n11887));
AND2X1 exu_U32330(.A(ecl_divcntl_n70), .B(exu_n16416), .Y(div_u32[12]));
INVX1 exu_U32331(.A(div_u32[12]), .Y(exu_n11888));
AND2X1 exu_U32332(.A(ecl_divcntl_n70), .B(exu_n16415), .Y(div_u32[11]));
INVX1 exu_U32333(.A(div_u32[11]), .Y(exu_n11889));
AND2X1 exu_U32334(.A(ecl_divcntl_n70), .B(exu_n16414), .Y(div_u32[10]));
INVX1 exu_U32335(.A(div_u32[10]), .Y(exu_n11890));
AND2X1 exu_U32336(.A(ecl_divcntl_n70), .B(exu_n16404), .Y(div_u32[0]));
INVX1 exu_U32337(.A(div_u32[0]), .Y(exu_n11891));
AND2X1 exu_U32338(.A(exu_n16246), .B(exu_n16412), .Y(div_pos32[8]));
INVX1 exu_U32339(.A(div_pos32[8]), .Y(exu_n11892));
AND2X1 exu_U32340(.A(exu_n16246), .B(exu_n16411), .Y(div_pos32[7]));
INVX1 exu_U32341(.A(div_pos32[7]), .Y(exu_n11893));
AND2X1 exu_U32342(.A(exu_n16246), .B(exu_n16410), .Y(div_pos32[6]));
INVX1 exu_U32343(.A(div_pos32[6]), .Y(exu_n11894));
AND2X1 exu_U32344(.A(exu_n16246), .B(exu_n16409), .Y(div_pos32[5]));
INVX1 exu_U32345(.A(div_pos32[5]), .Y(exu_n11895));
AND2X1 exu_U32346(.A(exu_n16246), .B(exu_n16408), .Y(div_pos32[4]));
INVX1 exu_U32347(.A(div_pos32[4]), .Y(exu_n11896));
AND2X1 exu_U32348(.A(exu_n16246), .B(exu_n16407), .Y(div_pos32[3]));
INVX1 exu_U32349(.A(div_pos32[3]), .Y(exu_n11897));
AND2X1 exu_U32350(.A(exu_n16246), .B(exu_n16434), .Y(div_pos32[30]));
INVX1 exu_U32351(.A(div_pos32[30]), .Y(exu_n11898));
AND2X1 exu_U32352(.A(exu_n16246), .B(exu_n16406), .Y(div_pos32[2]));
INVX1 exu_U32353(.A(div_pos32[2]), .Y(exu_n11899));
AND2X1 exu_U32354(.A(exu_n16246), .B(exu_n16433), .Y(div_pos32[29]));
INVX1 exu_U32355(.A(div_pos32[29]), .Y(exu_n11900));
AND2X1 exu_U32356(.A(exu_n16246), .B(exu_n16432), .Y(div_pos32[28]));
INVX1 exu_U32357(.A(div_pos32[28]), .Y(exu_n11901));
AND2X1 exu_U32358(.A(exu_n16246), .B(exu_n16431), .Y(div_pos32[27]));
INVX1 exu_U32359(.A(div_pos32[27]), .Y(exu_n11902));
AND2X1 exu_U32360(.A(exu_n16246), .B(exu_n16430), .Y(div_pos32[26]));
INVX1 exu_U32361(.A(div_pos32[26]), .Y(exu_n11903));
AND2X1 exu_U32362(.A(exu_n16246), .B(exu_n16429), .Y(div_pos32[25]));
INVX1 exu_U32363(.A(div_pos32[25]), .Y(exu_n11904));
AND2X1 exu_U32364(.A(exu_n16246), .B(exu_n16428), .Y(div_pos32[24]));
INVX1 exu_U32365(.A(div_pos32[24]), .Y(exu_n11905));
AND2X1 exu_U32366(.A(exu_n16246), .B(exu_n16427), .Y(div_pos32[23]));
INVX1 exu_U32367(.A(div_pos32[23]), .Y(exu_n11906));
AND2X1 exu_U32368(.A(exu_n16246), .B(exu_n16426), .Y(div_pos32[22]));
INVX1 exu_U32369(.A(div_pos32[22]), .Y(exu_n11907));
AND2X1 exu_U32370(.A(exu_n16246), .B(exu_n16425), .Y(div_pos32[21]));
INVX1 exu_U32371(.A(div_pos32[21]), .Y(exu_n11908));
AND2X1 exu_U32372(.A(exu_n16246), .B(exu_n16424), .Y(div_pos32[20]));
INVX1 exu_U32373(.A(div_pos32[20]), .Y(exu_n11909));
AND2X1 exu_U32374(.A(exu_n16246), .B(exu_n16405), .Y(div_pos32[1]));
INVX1 exu_U32375(.A(div_pos32[1]), .Y(exu_n11910));
AND2X1 exu_U32376(.A(exu_n16246), .B(exu_n16423), .Y(div_pos32[19]));
INVX1 exu_U32377(.A(div_pos32[19]), .Y(exu_n11911));
AND2X1 exu_U32378(.A(exu_n16246), .B(exu_n16422), .Y(div_pos32[18]));
INVX1 exu_U32379(.A(div_pos32[18]), .Y(exu_n11912));
AND2X1 exu_U32380(.A(exu_n16246), .B(exu_n16421), .Y(div_pos32[17]));
INVX1 exu_U32381(.A(div_pos32[17]), .Y(exu_n11913));
AND2X1 exu_U32382(.A(exu_n16246), .B(exu_n16420), .Y(div_pos32[16]));
INVX1 exu_U32383(.A(div_pos32[16]), .Y(exu_n11914));
AND2X1 exu_U32384(.A(exu_n16246), .B(exu_n16419), .Y(div_pos32[15]));
INVX1 exu_U32385(.A(div_pos32[15]), .Y(exu_n11915));
AND2X1 exu_U32386(.A(exu_n16246), .B(exu_n16418), .Y(div_pos32[14]));
INVX1 exu_U32387(.A(div_pos32[14]), .Y(exu_n11916));
AND2X1 exu_U32388(.A(exu_n16246), .B(exu_n16417), .Y(div_pos32[13]));
INVX1 exu_U32389(.A(div_pos32[13]), .Y(exu_n11917));
AND2X1 exu_U32390(.A(exu_n16246), .B(exu_n16416), .Y(div_pos32[12]));
INVX1 exu_U32391(.A(div_pos32[12]), .Y(exu_n11918));
AND2X1 exu_U32392(.A(exu_n16246), .B(exu_n16415), .Y(div_pos32[11]));
INVX1 exu_U32393(.A(div_pos32[11]), .Y(exu_n11919));
AND2X1 exu_U32394(.A(exu_n16246), .B(exu_n16414), .Y(div_pos32[10]));
INVX1 exu_U32395(.A(div_pos32[10]), .Y(exu_n11920));
AND2X1 exu_U32396(.A(exu_n16246), .B(exu_n16404), .Y(div_pos32[0]));
INVX1 exu_U32397(.A(div_pos32[0]), .Y(exu_n11921));
AND2X1 exu_U32398(.A(lsu_exu_st_dtlb_perr_g), .B(ecl_rml_thr_w[3]), .Y(ecl_n49));
INVX1 exu_U32399(.A(ecl_n49), .Y(exu_n11922));
AND2X1 exu_U32400(.A(ecl_rml_thr_w[2]), .B(lsu_exu_st_dtlb_perr_g), .Y(ecl_n52));
INVX1 exu_U32401(.A(ecl_n52), .Y(exu_n11923));
AND2X1 exu_U32402(.A(exu_n15958), .B(lsu_exu_st_dtlb_perr_g), .Y(ecl_n55));
INVX1 exu_U32403(.A(ecl_n55), .Y(exu_n11924));
AND2X1 exu_U32404(.A(exu_n15960), .B(lsu_exu_st_dtlb_perr_g), .Y(ecl_n58));
INVX1 exu_U32405(.A(ecl_n58), .Y(exu_n11925));
OR2X1 exu_U32406(.A(exu_tlu_ttype_vld_m), .B(exu_tlu_va_oor_jl_ret_m), .Y(ecl_n61));
INVX1 exu_U32407(.A(ecl_n61), .Y(exu_n11926));
AND2X1 exu_U32408(.A(ecl_div_yreg_data_31_g), .B(exu_n16614), .Y(ecl_n63));
INVX1 exu_U32409(.A(ecl_n63), .Y(exu_n11927));
INVX1 exu_U32410(.A(ecl_early1_ttype_e[5]), .Y(exu_n11928));
AND2X1 exu_U32411(.A(rml_ecl_other_e), .B(exu_n15030), .Y(ecl_n114));
INVX1 exu_U32412(.A(ecl_n114), .Y(exu_n11929));
INVX1 exu_U32413(.A(ecl_early1_ttype_e[3]), .Y(exu_n11930));
OR2X1 exu_U32414(.A(exu_n15030), .B(exu_n15493), .Y(ecl_n119));
INVX1 exu_U32415(.A(ecl_n119), .Y(exu_n11931));
AND2X1 exu_U32416(.A(rml_ecl_wtype_e[1]), .B(exu_n15030), .Y(ecl_n117));
INVX1 exu_U32417(.A(ecl_n117), .Y(exu_n11932));
INVX1 exu_U32418(.A(ecl_early1_ttype_e[2]), .Y(exu_n11933));
AND2X1 exu_U32419(.A(rml_ecl_wtype_e[0]), .B(exu_n15030), .Y(ecl_n121));
INVX1 exu_U32420(.A(ecl_n121), .Y(exu_n11934));
OR2X1 exu_U32421(.A(alu_ecl_add_n64_e), .B(exu_n16552), .Y(ecl_n133));
INVX1 exu_U32422(.A(ecl_n133), .Y(exu_n11935));
AND2X1 exu_U32423(.A(exu_n11937), .B(alu_ecl_add_n64_e), .Y(ecl_n131));
INVX1 exu_U32424(.A(ecl_n131), .Y(exu_n11936));
OR2X1 exu_U32425(.A(alu_logic_rs1_data_bf1[63]), .B(alu_ecl_adderin2_63_e), .Y(ecl_n134));
INVX1 exu_U32426(.A(ecl_n134), .Y(exu_n11937));
OR2X1 exu_U32427(.A(alu_logic_rs1_data_bf1[1]), .B(alu_logic_rs1_data_bf1[0]), .Y(ecl_n140));
INVX1 exu_U32428(.A(ecl_n140), .Y(exu_n11938));
OR2X1 exu_U32429(.A(ecl_n141), .B(exu_n14997), .Y(ecl_n137));
INVX1 exu_U32430(.A(ecl_n137), .Y(exu_n11939));
AND2X1 exu_U32431(.A(exu_n16636), .B(exu_n16635), .Y(exu_n16640));
INVX1 exu_U32432(.A(exu_n16640), .Y(exu_n11940));
AND2X1 exu_U32433(.A(exu_n16664), .B(exu_n16663), .Y(exu_n16668));
INVX1 exu_U32434(.A(exu_n16668), .Y(exu_n11941));
AND2X1 exu_U32435(.A(exu_n16678), .B(exu_n16677), .Y(exu_n16682));
INVX1 exu_U32436(.A(exu_n16682), .Y(exu_n11942));
AND2X1 exu_U32437(.A(exu_n16692), .B(exu_n16691), .Y(exu_n16696));
INVX1 exu_U32438(.A(exu_n16696), .Y(exu_n11943));
AND2X1 exu_U32439(.A(exu_n16720), .B(exu_n16719), .Y(exu_n16724));
INVX1 exu_U32440(.A(exu_n16724), .Y(exu_n11944));
AND2X1 exu_U32441(.A(exu_n16734), .B(exu_n16733), .Y(exu_n16738));
INVX1 exu_U32442(.A(exu_n16738), .Y(exu_n11945));
AND2X1 exu_U32443(.A(exu_n17377), .B(exu_n17376), .Y(exu_n17381));
INVX1 exu_U32444(.A(exu_n17381), .Y(exu_n11946));
AND2X1 exu_U32445(.A(exu_n17391), .B(exu_n17390), .Y(exu_n17395));
INVX1 exu_U32446(.A(exu_n17395), .Y(exu_n11947));
AND2X1 exu_U32447(.A(exu_n17398), .B(exu_n17397), .Y(exu_n17402));
INVX1 exu_U32448(.A(exu_n17402), .Y(exu_n11948));
AND2X1 exu_U32449(.A(exu_n17412), .B(exu_n17411), .Y(exu_n17416));
INVX1 exu_U32450(.A(exu_n17416), .Y(exu_n11949));
AND2X1 exu_U32451(.A(exu_n17440), .B(exu_n17439), .Y(exu_n17444));
INVX1 exu_U32452(.A(exu_n17444), .Y(exu_n11950));
AND2X1 exu_U32453(.A(exu_n17454), .B(exu_n17453), .Y(exu_n17458));
INVX1 exu_U32454(.A(exu_n17458), .Y(exu_n11951));
AND2X1 exu_U32455(.A(exu_n17632), .B(exu_n17633), .Y(exu_n17628));
INVX1 exu_U32456(.A(exu_n17628), .Y(exu_n11952));
AND2X1 exu_U32457(.A(exu_n17644), .B(exu_n17645), .Y(exu_n17640));
INVX1 exu_U32458(.A(exu_n17640), .Y(exu_n11953));
AND2X1 exu_U32459(.A(exu_n17656), .B(exu_n17657), .Y(exu_n17652));
INVX1 exu_U32460(.A(exu_n17652), .Y(exu_n11954));
AND2X1 exu_U32461(.A(exu_n17668), .B(exu_n17669), .Y(exu_n17664));
INVX1 exu_U32462(.A(exu_n17664), .Y(exu_n11955));
AND2X1 exu_U32463(.A(exu_n17680), .B(exu_n17681), .Y(exu_n17676));
INVX1 exu_U32464(.A(exu_n17676), .Y(exu_n11956));
AND2X1 exu_U32465(.A(ecl_ecl_irf_rd_w[0]), .B(exu_n17692), .Y(exu_n17688));
INVX1 exu_U32466(.A(exu_n17688), .Y(exu_n11957));
AND2X1 exu_U32467(.A(ecl_wb_byplog_rd_w2[0]), .B(exu_n17703), .Y(exu_n17699));
INVX1 exu_U32468(.A(exu_n17699), .Y(exu_n11958));
INVX1 exu_U32469(.A(alu_zcomp_in[9]), .Y(exu_n11959));
INVX1 exu_U32470(.A(alu_zcomp_in[7]), .Y(exu_n11960));
INVX1 exu_U32471(.A(alu_zcomp_in[63]), .Y(exu_n11961));
INVX1 exu_U32472(.A(alu_zcomp_in[61]), .Y(exu_n11962));
INVX1 exu_U32473(.A(alu_zcomp_in[5]), .Y(exu_n11963));
INVX1 exu_U32474(.A(alu_zcomp_in[59]), .Y(exu_n11964));
INVX1 exu_U32475(.A(alu_zcomp_in[57]), .Y(exu_n11965));
INVX1 exu_U32476(.A(alu_zcomp_in[55]), .Y(exu_n11966));
INVX1 exu_U32477(.A(alu_zcomp_in[53]), .Y(exu_n11967));
INVX1 exu_U32478(.A(alu_zcomp_in[51]), .Y(exu_n11968));
INVX1 exu_U32479(.A(alu_zcomp_in[49]), .Y(exu_n11969));
INVX1 exu_U32480(.A(alu_zcomp_in[47]), .Y(exu_n11970));
INVX1 exu_U32481(.A(alu_zcomp_in[45]), .Y(exu_n11971));
INVX1 exu_U32482(.A(alu_zcomp_in[43]), .Y(exu_n11972));
INVX1 exu_U32483(.A(alu_zcomp_in[41]), .Y(exu_n11973));
INVX1 exu_U32484(.A(alu_zcomp_in[3]), .Y(exu_n11974));
INVX1 exu_U32485(.A(alu_zcomp_in[39]), .Y(exu_n11975));
INVX1 exu_U32486(.A(alu_zcomp_in[37]), .Y(exu_n11976));
INVX1 exu_U32487(.A(alu_zcomp_in[35]), .Y(exu_n11977));
INVX1 exu_U32488(.A(alu_zcomp_in[33]), .Y(exu_n11978));
INVX1 exu_U32489(.A(alu_zcomp_in[30]), .Y(exu_n11979));
INVX1 exu_U32490(.A(alu_zcomp_in[29]), .Y(exu_n11980));
INVX1 exu_U32491(.A(alu_zcomp_in[27]), .Y(exu_n11981));
INVX1 exu_U32492(.A(alu_zcomp_in[25]), .Y(exu_n11982));
INVX1 exu_U32493(.A(alu_zcomp_in[23]), .Y(exu_n11983));
INVX1 exu_U32494(.A(alu_zcomp_in[21]), .Y(exu_n11984));
INVX1 exu_U32495(.A(alu_zcomp_in[1]), .Y(exu_n11985));
INVX1 exu_U32496(.A(alu_zcomp_in[18]), .Y(exu_n11986));
INVX1 exu_U32497(.A(alu_zcomp_in[16]), .Y(exu_n11987));
INVX1 exu_U32498(.A(alu_zcomp_in[14]), .Y(exu_n11988));
INVX1 exu_U32499(.A(alu_zcomp_in[12]), .Y(exu_n11989));
INVX1 exu_U32500(.A(alu_zcomp_in[10]), .Y(exu_n11990));
INVX1 exu_U32501(.A(div_gencc_in_9), .Y(exu_n11991));
INVX1 exu_U32502(.A(div_gencc_in_7), .Y(exu_n11992));
INVX1 exu_U32503(.A(div_gencc_in_5), .Y(exu_n11993));
INVX1 exu_U32504(.A(div_gencc_in_3), .Y(exu_n11994));
INVX1 exu_U32505(.A(div_gencc_in_30), .Y(exu_n11995));
INVX1 exu_U32506(.A(div_gencc_in_29), .Y(exu_n11996));
INVX1 exu_U32507(.A(div_gencc_in_27), .Y(exu_n11997));
INVX1 exu_U32508(.A(div_gencc_in_25), .Y(exu_n11998));
INVX1 exu_U32509(.A(div_gencc_in_23), .Y(exu_n11999));
INVX1 exu_U32510(.A(div_gencc_in_21), .Y(exu_n12000));
INVX1 exu_U32511(.A(div_gencc_in_1), .Y(exu_n12001));
INVX1 exu_U32512(.A(div_gencc_in_18), .Y(exu_n12002));
INVX1 exu_U32513(.A(div_gencc_in_16), .Y(exu_n12003));
INVX1 exu_U32514(.A(div_gencc_in_14), .Y(exu_n12004));
INVX1 exu_U32515(.A(div_gencc_in_12), .Y(exu_n12005));
INVX1 exu_U32516(.A(div_gencc_in_10), .Y(exu_n12006));
INVX1 exu_U32517(.A(div_z_in[9]), .Y(exu_n12007));
INVX1 exu_U32518(.A(div_z_in[7]), .Y(exu_n12008));
INVX1 exu_U32519(.A(div_z_in[63]), .Y(exu_n12009));
INVX1 exu_U32520(.A(div_z_in[61]), .Y(exu_n12010));
INVX1 exu_U32521(.A(div_z_in[5]), .Y(exu_n12011));
INVX1 exu_U32522(.A(div_z_in[59]), .Y(exu_n12012));
INVX1 exu_U32523(.A(div_z_in[57]), .Y(exu_n12013));
INVX1 exu_U32524(.A(div_z_in[55]), .Y(exu_n12014));
INVX1 exu_U32525(.A(div_z_in[53]), .Y(exu_n12015));
INVX1 exu_U32526(.A(div_z_in[51]), .Y(exu_n12016));
INVX1 exu_U32527(.A(div_z_in[49]), .Y(exu_n12017));
INVX1 exu_U32528(.A(div_z_in[47]), .Y(exu_n12018));
INVX1 exu_U32529(.A(div_z_in[45]), .Y(exu_n12019));
INVX1 exu_U32530(.A(div_z_in[43]), .Y(exu_n12020));
INVX1 exu_U32531(.A(div_z_in[41]), .Y(exu_n12021));
INVX1 exu_U32532(.A(div_z_in[3]), .Y(exu_n12022));
INVX1 exu_U32533(.A(div_z_in[39]), .Y(exu_n12023));
INVX1 exu_U32534(.A(div_z_in[37]), .Y(exu_n12024));
INVX1 exu_U32535(.A(div_z_in[35]), .Y(exu_n12025));
INVX1 exu_U32536(.A(div_z_in[33]), .Y(exu_n12026));
INVX1 exu_U32537(.A(div_z_in[30]), .Y(exu_n12027));
INVX1 exu_U32538(.A(div_z_in[29]), .Y(exu_n12028));
INVX1 exu_U32539(.A(div_z_in[27]), .Y(exu_n12029));
INVX1 exu_U32540(.A(div_z_in[25]), .Y(exu_n12030));
INVX1 exu_U32541(.A(div_z_in[23]), .Y(exu_n12031));
INVX1 exu_U32542(.A(div_z_in[21]), .Y(exu_n12032));
INVX1 exu_U32543(.A(div_z_in[1]), .Y(exu_n12033));
INVX1 exu_U32544(.A(div_z_in[18]), .Y(exu_n12034));
INVX1 exu_U32545(.A(div_z_in[16]), .Y(exu_n12035));
INVX1 exu_U32546(.A(div_z_in[14]), .Y(exu_n12036));
INVX1 exu_U32547(.A(div_z_in[12]), .Y(exu_n12037));
INVX1 exu_U32548(.A(div_z_in[10]), .Y(exu_n12038));
INVX1 exu_U32549(.A(exu_n31620), .Y(exu_n12039));
INVX1 exu_U32550(.A(exu_n31626), .Y(exu_n12040));
INVX1 exu_U32551(.A(exu_n31634), .Y(exu_n12041));
INVX1 exu_U32552(.A(exu_n31640), .Y(exu_n12042));
INVX1 exu_U32553(.A(exu_n31650), .Y(exu_n12043));
INVX1 exu_U32554(.A(exu_n31656), .Y(exu_n12044));
INVX1 exu_U32555(.A(exu_n31664), .Y(exu_n12045));
INVX1 exu_U32556(.A(exu_n31670), .Y(exu_n12046));
INVX1 exu_U32557(.A(exu_n31680), .Y(exu_n12047));
INVX1 exu_U32558(.A(exu_n31686), .Y(exu_n12048));
INVX1 exu_U32559(.A(exu_n31693), .Y(exu_n12049));
INVX1 exu_U32560(.A(exu_n31699), .Y(exu_n12050));
AND2X1 exu_U32561(.A(ecl_byplog_rs1_w_comp7_n7), .B(ecl_byplog_rs1_w_comp7_n8), .Y(ecl_byplog_rs1_w_comp7_n3));
INVX1 exu_U32562(.A(ecl_byplog_rs1_w_comp7_n3), .Y(exu_n12051));
AND2X1 exu_U32563(.A(rml_cwp_n101), .B(tlu_exu_cwpccr_update_m), .Y(rml_cwp_n97));
INVX1 exu_U32564(.A(rml_cwp_n97), .Y(exu_n12052));
OR2X1 exu_U32565(.A(rml_rml_ecl_other_d), .B(rml_ecl_wstate_d[0]), .Y(rml_wtype_mux_n7));
INVX1 exu_U32566(.A(rml_wtype_mux_n7), .Y(exu_n12053));
OR2X1 exu_U32567(.A(rml_rml_ecl_other_d), .B(rml_ecl_wstate_d[1]), .Y(rml_wtype_mux_n9));
INVX1 exu_U32568(.A(rml_wtype_mux_n9), .Y(exu_n12054));
OR2X1 exu_U32569(.A(rml_rml_ecl_other_d), .B(rml_ecl_wstate_d[2]), .Y(rml_wtype_mux_n11));
INVX1 exu_U32570(.A(rml_wtype_mux_n11), .Y(exu_n12055));
INVX1 exu_U32571(.A(div_low32or_n5), .Y(exu_n12056));
INVX1 exu_U32572(.A(div_low32or_n11), .Y(exu_n12057));
INVX1 exu_U32573(.A(div_low32or_n19), .Y(exu_n12058));
INVX1 exu_U32574(.A(div_low32or_n25), .Y(exu_n12059));
AND2X1 exu_U32575(.A(alu_chk_mem_addr_n9), .B(alu_chk_mem_addr_n10), .Y(alu_chk_mem_addr_n5));
INVX1 exu_U32576(.A(alu_chk_mem_addr_n5), .Y(exu_n12060));
AND2X1 exu_U32577(.A(alu_chk_mem_addr_n15), .B(alu_chk_mem_addr_n16), .Y(alu_chk_mem_addr_n11));
INVX1 exu_U32578(.A(alu_chk_mem_addr_n11), .Y(exu_n12061));
INVX1 exu_U32579(.A(alu_chk_mem_addr_n1), .Y(exu_n12062));
AND2X1 exu_U32580(.A(alu_chk_mem_addr_n23), .B(alu_chk_mem_addr_n24), .Y(alu_chk_mem_addr_n19));
INVX1 exu_U32581(.A(alu_chk_mem_addr_n19), .Y(exu_n12063));
AND2X1 exu_U32582(.A(alu_chk_mem_addr_n29), .B(alu_chk_mem_addr_n30), .Y(alu_chk_mem_addr_n25));
INVX1 exu_U32583(.A(alu_chk_mem_addr_n25), .Y(exu_n12064));
AND2X1 exu_U32584(.A(exu_mul_input_vld), .B(exu_n15425), .Y(ecl_mdqctl_n24));
INVX1 exu_U32585(.A(ecl_mdqctl_n24), .Y(exu_n12065));
AND2X1 exu_U32586(.A(ecl_div_ld_inputs), .B(exu_n16185), .Y(ecl_mdqctl_n52));
INVX1 exu_U32587(.A(ecl_mdqctl_n52), .Y(exu_n12066));
INVX1 exu_U32588(.A(ecl_writeback_n59), .Y(exu_n12067));
AND2X1 exu_U32589(.A(exu_n16389), .B(exu_n16611), .Y(ecl_writeback_n63));
INVX1 exu_U32590(.A(ecl_writeback_n63), .Y(exu_n12068));
INVX1 exu_U32591(.A(div_n41), .Y(exu_n12069));
INVX1 exu_U32592(.A(div_n47), .Y(exu_n12070));
INVX1 exu_U32593(.A(div_n55), .Y(exu_n12071));
INVX1 exu_U32594(.A(div_n61), .Y(exu_n12072));
INVX1 exu_U32595(.A(div_n71), .Y(exu_n12073));
INVX1 exu_U32596(.A(div_n77), .Y(exu_n12074));
INVX1 exu_U32597(.A(div_n85), .Y(exu_n12075));
INVX1 exu_U32598(.A(div_n91), .Y(exu_n12076));
INVX1 exu_U32599(.A(alu_n73), .Y(exu_n12077));
INVX1 exu_U32600(.A(alu_n79), .Y(exu_n12078));
INVX1 exu_U32601(.A(alu_n87), .Y(exu_n12079));
INVX1 exu_U32602(.A(alu_n93), .Y(exu_n12080));
INVX1 exu_U32603(.A(alu_n103), .Y(exu_n12081));
INVX1 exu_U32604(.A(alu_n109), .Y(exu_n12082));
INVX1 exu_U32605(.A(alu_n99), .Y(exu_n12083));
INVX1 exu_U32606(.A(alu_n117), .Y(exu_n12084));
INVX1 exu_U32607(.A(alu_n123), .Y(exu_n12085));
AND2X1 exu_U32608(.A(exu_n16650), .B(exu_n16649), .Y(exu_n16654));
INVX1 exu_U32609(.A(exu_n16654), .Y(exu_n12086));
AND2X1 exu_U32610(.A(exu_n16706), .B(exu_n16705), .Y(exu_n16710));
INVX1 exu_U32611(.A(exu_n16710), .Y(exu_n12087));
AND2X1 exu_U32612(.A(exu_n17384), .B(exu_n17383), .Y(exu_n17388));
INVX1 exu_U32613(.A(exu_n17388), .Y(exu_n12088));
AND2X1 exu_U32614(.A(exu_n17426), .B(exu_n17425), .Y(exu_n17430));
INVX1 exu_U32615(.A(exu_n17430), .Y(exu_n12089));
INVX1 exu_U32616(.A(exu_n17728), .Y(exu_n12090));
INVX1 exu_U32617(.A(exu_n17734), .Y(exu_n12091));
INVX1 exu_U32618(.A(exu_n17740), .Y(exu_n12092));
INVX1 exu_U32619(.A(exu_n17746), .Y(exu_n12093));
INVX1 exu_U32620(.A(exu_n17752), .Y(exu_n12094));
INVX1 exu_U32621(.A(exu_n17758), .Y(exu_n12095));
INVX1 exu_U32622(.A(exu_n17764), .Y(exu_n12096));
INVX1 exu_U32623(.A(exu_n17770), .Y(exu_n12097));
INVX1 exu_U32624(.A(exu_n17776), .Y(exu_n12098));
INVX1 exu_U32625(.A(exu_n17782), .Y(exu_n12099));
INVX1 exu_U32626(.A(exu_n17788), .Y(exu_n12100));
INVX1 exu_U32627(.A(exu_n17794), .Y(exu_n12101));
INVX1 exu_U32628(.A(exu_n17800), .Y(exu_n12102));
INVX1 exu_U32629(.A(exu_n17806), .Y(exu_n12103));
INVX1 exu_U32630(.A(exu_n17812), .Y(exu_n12104));
INVX1 exu_U32631(.A(exu_n17818), .Y(exu_n12105));
INVX1 exu_U32632(.A(exu_n17824), .Y(exu_n12106));
INVX1 exu_U32633(.A(exu_n17830), .Y(exu_n12107));
INVX1 exu_U32634(.A(exu_n17836), .Y(exu_n12108));
INVX1 exu_U32635(.A(exu_n17842), .Y(exu_n12109));
INVX1 exu_U32636(.A(exu_n17848), .Y(exu_n12110));
INVX1 exu_U32637(.A(exu_n17854), .Y(exu_n12111));
INVX1 exu_U32638(.A(exu_n17860), .Y(exu_n12112));
INVX1 exu_U32639(.A(exu_n17866), .Y(exu_n12113));
INVX1 exu_U32640(.A(exu_n17872), .Y(exu_n12114));
INVX1 exu_U32641(.A(exu_n17878), .Y(exu_n12115));
INVX1 exu_U32642(.A(exu_n17884), .Y(exu_n12116));
INVX1 exu_U32643(.A(exu_n17890), .Y(exu_n12117));
INVX1 exu_U32644(.A(exu_n17896), .Y(exu_n12118));
INVX1 exu_U32645(.A(exu_n17902), .Y(exu_n12119));
INVX1 exu_U32646(.A(exu_n17908), .Y(exu_n12120));
INVX1 exu_U32647(.A(exu_n17914), .Y(exu_n12121));
INVX1 exu_U32648(.A(exu_n17920), .Y(exu_n12122));
INVX1 exu_U32649(.A(exu_n17926), .Y(exu_n12123));
INVX1 exu_U32650(.A(exu_n17932), .Y(exu_n12124));
INVX1 exu_U32651(.A(exu_n17938), .Y(exu_n12125));
INVX1 exu_U32652(.A(exu_n17944), .Y(exu_n12126));
INVX1 exu_U32653(.A(exu_n17950), .Y(exu_n12127));
INVX1 exu_U32654(.A(exu_n17956), .Y(exu_n12128));
INVX1 exu_U32655(.A(exu_n17962), .Y(exu_n12129));
INVX1 exu_U32656(.A(exu_n17968), .Y(exu_n12130));
INVX1 exu_U32657(.A(exu_n17974), .Y(exu_n12131));
INVX1 exu_U32658(.A(exu_n17981), .Y(exu_n12132));
INVX1 exu_U32659(.A(exu_n17987), .Y(exu_n12133));
INVX1 exu_U32660(.A(exu_n17993), .Y(exu_n12134));
INVX1 exu_U32661(.A(exu_n17999), .Y(exu_n12135));
INVX1 exu_U32662(.A(exu_n18005), .Y(exu_n12136));
INVX1 exu_U32663(.A(exu_n18019), .Y(exu_n12137));
INVX1 exu_U32664(.A(exu_n18025), .Y(exu_n12138));
INVX1 exu_U32665(.A(exu_n18031), .Y(exu_n12139));
AND2X1 exu_U32666(.A(exu_n15210), .B(exu_n16270), .Y(exu_n19198));
INVX1 exu_U32667(.A(exu_n19198), .Y(exu_n12140));
INVX1 exu_U32668(.A(exu_n19212), .Y(exu_n12141));
INVX1 exu_U32669(.A(exu_n19213), .Y(exu_n12142));
AND2X1 exu_U32670(.A(exu_n15209), .B(exu_n16270), .Y(exu_n19234));
INVX1 exu_U32671(.A(exu_n19234), .Y(exu_n12143));
INVX1 exu_U32672(.A(exu_n19248), .Y(exu_n12144));
INVX1 exu_U32673(.A(exu_n19249), .Y(exu_n12145));
INVX1 exu_U32674(.A(exu_n20476), .Y(exu_n12146));
INVX1 exu_U32675(.A(exu_n20482), .Y(exu_n12147));
INVX1 exu_U32676(.A(exu_n20488), .Y(exu_n12148));
INVX1 exu_U32677(.A(exu_n20494), .Y(exu_n12149));
INVX1 exu_U32678(.A(exu_n20500), .Y(exu_n12150));
INVX1 exu_U32679(.A(exu_n20506), .Y(exu_n12151));
INVX1 exu_U32680(.A(exu_n20512), .Y(exu_n12152));
INVX1 exu_U32681(.A(exu_n20518), .Y(exu_n12153));
INVX1 exu_U32682(.A(exu_n20524), .Y(exu_n12154));
INVX1 exu_U32683(.A(exu_n20530), .Y(exu_n12155));
INVX1 exu_U32684(.A(exu_n20536), .Y(exu_n12156));
INVX1 exu_U32685(.A(exu_n20542), .Y(exu_n12157));
INVX1 exu_U32686(.A(exu_n20548), .Y(exu_n12158));
INVX1 exu_U32687(.A(exu_n20554), .Y(exu_n12159));
INVX1 exu_U32688(.A(exu_n20560), .Y(exu_n12160));
INVX1 exu_U32689(.A(exu_n20566), .Y(exu_n12161));
INVX1 exu_U32690(.A(exu_n20572), .Y(exu_n12162));
INVX1 exu_U32691(.A(exu_n20578), .Y(exu_n12163));
INVX1 exu_U32692(.A(exu_n20584), .Y(exu_n12164));
INVX1 exu_U32693(.A(exu_n20590), .Y(exu_n12165));
INVX1 exu_U32694(.A(exu_n20596), .Y(exu_n12166));
INVX1 exu_U32695(.A(exu_n20602), .Y(exu_n12167));
INVX1 exu_U32696(.A(exu_n20608), .Y(exu_n12168));
INVX1 exu_U32697(.A(exu_n20614), .Y(exu_n12169));
INVX1 exu_U32698(.A(exu_n20620), .Y(exu_n12170));
INVX1 exu_U32699(.A(exu_n20626), .Y(exu_n12171));
INVX1 exu_U32700(.A(exu_n20632), .Y(exu_n12172));
INVX1 exu_U32701(.A(exu_n20638), .Y(exu_n12173));
INVX1 exu_U32702(.A(exu_n20644), .Y(exu_n12174));
INVX1 exu_U32703(.A(exu_n20650), .Y(exu_n12175));
INVX1 exu_U32704(.A(exu_n20656), .Y(exu_n12176));
INVX1 exu_U32705(.A(exu_n20662), .Y(exu_n12177));
INVX1 exu_U32706(.A(exu_n20668), .Y(exu_n12178));
INVX1 exu_U32707(.A(exu_n20674), .Y(exu_n12179));
INVX1 exu_U32708(.A(exu_n20680), .Y(exu_n12180));
INVX1 exu_U32709(.A(exu_n20686), .Y(exu_n12181));
INVX1 exu_U32710(.A(exu_n20692), .Y(exu_n12182));
INVX1 exu_U32711(.A(exu_n20698), .Y(exu_n12183));
INVX1 exu_U32712(.A(exu_n20704), .Y(exu_n12184));
INVX1 exu_U32713(.A(exu_n20710), .Y(exu_n12185));
INVX1 exu_U32714(.A(exu_n20716), .Y(exu_n12186));
INVX1 exu_U32715(.A(exu_n20722), .Y(exu_n12187));
INVX1 exu_U32716(.A(exu_n20728), .Y(exu_n12188));
INVX1 exu_U32717(.A(exu_n20734), .Y(exu_n12189));
INVX1 exu_U32718(.A(exu_n20740), .Y(exu_n12190));
INVX1 exu_U32719(.A(exu_n20746), .Y(exu_n12191));
INVX1 exu_U32720(.A(exu_n20752), .Y(exu_n12192));
INVX1 exu_U32721(.A(exu_n20758), .Y(exu_n12193));
INVX1 exu_U32722(.A(exu_n20764), .Y(exu_n12194));
INVX1 exu_U32723(.A(exu_n20770), .Y(exu_n12195));
INVX1 exu_U32724(.A(exu_n20776), .Y(exu_n12196));
INVX1 exu_U32725(.A(exu_n20782), .Y(exu_n12197));
INVX1 exu_U32726(.A(exu_n20788), .Y(exu_n12198));
INVX1 exu_U32727(.A(exu_n20794), .Y(exu_n12199));
INVX1 exu_U32728(.A(exu_n20800), .Y(exu_n12200));
INVX1 exu_U32729(.A(exu_n20806), .Y(exu_n12201));
INVX1 exu_U32730(.A(exu_n20812), .Y(exu_n12202));
INVX1 exu_U32731(.A(exu_n20818), .Y(exu_n12203));
INVX1 exu_U32732(.A(exu_n20824), .Y(exu_n12204));
INVX1 exu_U32733(.A(exu_n20830), .Y(exu_n12205));
INVX1 exu_U32734(.A(exu_n20836), .Y(exu_n12206));
INVX1 exu_U32735(.A(exu_n20842), .Y(exu_n12207));
INVX1 exu_U32736(.A(exu_n20848), .Y(exu_n12208));
INVX1 exu_U32737(.A(exu_n20854), .Y(exu_n12209));
INVX1 exu_U32738(.A(exu_n20860), .Y(exu_n12210));
INVX1 exu_U32739(.A(exu_n20866), .Y(exu_n12211));
INVX1 exu_U32740(.A(exu_n20872), .Y(exu_n12212));
INVX1 exu_U32741(.A(exu_n20878), .Y(exu_n12213));
INVX1 exu_U32742(.A(exu_n20884), .Y(exu_n12214));
INVX1 exu_U32743(.A(exu_n20890), .Y(exu_n12215));
INVX1 exu_U32744(.A(exu_n20896), .Y(exu_n12216));
INVX1 exu_U32745(.A(exu_n20902), .Y(exu_n12217));
INVX1 exu_U32746(.A(exu_n20908), .Y(exu_n12218));
INVX1 exu_U32747(.A(exu_n20914), .Y(exu_n12219));
INVX1 exu_U32748(.A(exu_n20920), .Y(exu_n12220));
INVX1 exu_U32749(.A(exu_n20926), .Y(exu_n12221));
INVX1 exu_U32750(.A(exu_n20932), .Y(exu_n12222));
INVX1 exu_U32751(.A(exu_n20938), .Y(exu_n12223));
INVX1 exu_U32752(.A(exu_n20944), .Y(exu_n12224));
INVX1 exu_U32753(.A(exu_n20950), .Y(exu_n12225));
INVX1 exu_U32754(.A(exu_n20956), .Y(exu_n12226));
INVX1 exu_U32755(.A(exu_n20962), .Y(exu_n12227));
INVX1 exu_U32756(.A(exu_n20968), .Y(exu_n12228));
INVX1 exu_U32757(.A(exu_n20974), .Y(exu_n12229));
INVX1 exu_U32758(.A(exu_n20980), .Y(exu_n12230));
INVX1 exu_U32759(.A(exu_n20986), .Y(exu_n12231));
INVX1 exu_U32760(.A(exu_n20992), .Y(exu_n12232));
INVX1 exu_U32761(.A(exu_n20998), .Y(exu_n12233));
INVX1 exu_U32762(.A(exu_n21004), .Y(exu_n12234));
INVX1 exu_U32763(.A(exu_n21010), .Y(exu_n12235));
INVX1 exu_U32764(.A(exu_n21016), .Y(exu_n12236));
INVX1 exu_U32765(.A(exu_n21022), .Y(exu_n12237));
INVX1 exu_U32766(.A(exu_n21028), .Y(exu_n12238));
INVX1 exu_U32767(.A(exu_n21034), .Y(exu_n12239));
INVX1 exu_U32768(.A(exu_n21040), .Y(exu_n12240));
INVX1 exu_U32769(.A(exu_n21046), .Y(exu_n12241));
INVX1 exu_U32770(.A(exu_n21052), .Y(exu_n12242));
INVX1 exu_U32771(.A(exu_n21058), .Y(exu_n12243));
INVX1 exu_U32772(.A(exu_n21064), .Y(exu_n12244));
INVX1 exu_U32773(.A(exu_n21070), .Y(exu_n12245));
INVX1 exu_U32774(.A(exu_n21076), .Y(exu_n12246));
INVX1 exu_U32775(.A(exu_n21082), .Y(exu_n12247));
INVX1 exu_U32776(.A(exu_n21088), .Y(exu_n12248));
INVX1 exu_U32777(.A(exu_n21094), .Y(exu_n12249));
INVX1 exu_U32778(.A(exu_n21100), .Y(exu_n12250));
INVX1 exu_U32779(.A(exu_n21106), .Y(exu_n12251));
INVX1 exu_U32780(.A(exu_n21112), .Y(exu_n12252));
INVX1 exu_U32781(.A(exu_n21118), .Y(exu_n12253));
INVX1 exu_U32782(.A(exu_n21124), .Y(exu_n12254));
INVX1 exu_U32783(.A(exu_n21130), .Y(exu_n12255));
INVX1 exu_U32784(.A(exu_n21136), .Y(exu_n12256));
INVX1 exu_U32785(.A(exu_n21142), .Y(exu_n12257));
INVX1 exu_U32786(.A(exu_n21148), .Y(exu_n12258));
INVX1 exu_U32787(.A(exu_n21154), .Y(exu_n12259));
INVX1 exu_U32788(.A(exu_n21160), .Y(exu_n12260));
INVX1 exu_U32789(.A(exu_n21166), .Y(exu_n12261));
INVX1 exu_U32790(.A(exu_n21172), .Y(exu_n12262));
INVX1 exu_U32791(.A(exu_n21178), .Y(exu_n12263));
INVX1 exu_U32792(.A(exu_n21184), .Y(exu_n12264));
INVX1 exu_U32793(.A(exu_n21190), .Y(exu_n12265));
INVX1 exu_U32794(.A(exu_n21196), .Y(exu_n12266));
INVX1 exu_U32795(.A(exu_n21202), .Y(exu_n12267));
INVX1 exu_U32796(.A(exu_n21208), .Y(exu_n12268));
INVX1 exu_U32797(.A(exu_n21214), .Y(exu_n12269));
INVX1 exu_U32798(.A(exu_n21220), .Y(exu_n12270));
INVX1 exu_U32799(.A(exu_n21226), .Y(exu_n12271));
INVX1 exu_U32800(.A(exu_n21232), .Y(exu_n12272));
INVX1 exu_U32801(.A(exu_n21238), .Y(exu_n12273));
INVX1 exu_U32802(.A(exu_n21244), .Y(exu_n12274));
INVX1 exu_U32803(.A(exu_n21250), .Y(exu_n12275));
INVX1 exu_U32804(.A(exu_n21256), .Y(exu_n12276));
INVX1 exu_U32805(.A(exu_n21262), .Y(exu_n12277));
INVX1 exu_U32806(.A(exu_n21268), .Y(exu_n12278));
INVX1 exu_U32807(.A(exu_n21274), .Y(exu_n12279));
INVX1 exu_U32808(.A(exu_n21280), .Y(exu_n12280));
INVX1 exu_U32809(.A(exu_n21286), .Y(exu_n12281));
INVX1 exu_U32810(.A(exu_n21292), .Y(exu_n12282));
INVX1 exu_U32811(.A(exu_n21298), .Y(exu_n12283));
INVX1 exu_U32812(.A(exu_n21304), .Y(exu_n12284));
INVX1 exu_U32813(.A(exu_n21310), .Y(exu_n12285));
INVX1 exu_U32814(.A(exu_n21316), .Y(exu_n12286));
INVX1 exu_U32815(.A(exu_n21322), .Y(exu_n12287));
INVX1 exu_U32816(.A(exu_n21328), .Y(exu_n12288));
INVX1 exu_U32817(.A(exu_n21334), .Y(exu_n12289));
INVX1 exu_U32818(.A(exu_n21340), .Y(exu_n12290));
INVX1 exu_U32819(.A(exu_n21346), .Y(exu_n12291));
INVX1 exu_U32820(.A(exu_n21352), .Y(exu_n12292));
INVX1 exu_U32821(.A(exu_n21358), .Y(exu_n12293));
INVX1 exu_U32822(.A(exu_n21364), .Y(exu_n12294));
INVX1 exu_U32823(.A(exu_n21370), .Y(exu_n12295));
INVX1 exu_U32824(.A(exu_n21376), .Y(exu_n12296));
INVX1 exu_U32825(.A(exu_n21382), .Y(exu_n12297));
INVX1 exu_U32826(.A(exu_n21388), .Y(exu_n12298));
INVX1 exu_U32827(.A(exu_n21394), .Y(exu_n12299));
INVX1 exu_U32828(.A(exu_n21400), .Y(exu_n12300));
INVX1 exu_U32829(.A(exu_n21406), .Y(exu_n12301));
INVX1 exu_U32830(.A(exu_n21412), .Y(exu_n12302));
INVX1 exu_U32831(.A(exu_n21418), .Y(exu_n12303));
INVX1 exu_U32832(.A(exu_n21424), .Y(exu_n12304));
INVX1 exu_U32833(.A(exu_n21430), .Y(exu_n12305));
INVX1 exu_U32834(.A(exu_n21436), .Y(exu_n12306));
INVX1 exu_U32835(.A(exu_n21442), .Y(exu_n12307));
INVX1 exu_U32836(.A(exu_n21448), .Y(exu_n12308));
INVX1 exu_U32837(.A(exu_n21454), .Y(exu_n12309));
INVX1 exu_U32838(.A(exu_n21460), .Y(exu_n12310));
INVX1 exu_U32839(.A(exu_n21466), .Y(exu_n12311));
INVX1 exu_U32840(.A(exu_n21472), .Y(exu_n12312));
INVX1 exu_U32841(.A(exu_n21478), .Y(exu_n12313));
INVX1 exu_U32842(.A(exu_n21484), .Y(exu_n12314));
INVX1 exu_U32843(.A(exu_n21490), .Y(exu_n12315));
INVX1 exu_U32844(.A(exu_n21496), .Y(exu_n12316));
INVX1 exu_U32845(.A(exu_n21502), .Y(exu_n12317));
INVX1 exu_U32846(.A(exu_n21508), .Y(exu_n12318));
INVX1 exu_U32847(.A(exu_n21514), .Y(exu_n12319));
INVX1 exu_U32848(.A(exu_n21520), .Y(exu_n12320));
INVX1 exu_U32849(.A(exu_n21526), .Y(exu_n12321));
INVX1 exu_U32850(.A(exu_n21532), .Y(exu_n12322));
INVX1 exu_U32851(.A(exu_n21538), .Y(exu_n12323));
INVX1 exu_U32852(.A(exu_n21544), .Y(exu_n12324));
INVX1 exu_U32853(.A(exu_n21550), .Y(exu_n12325));
INVX1 exu_U32854(.A(exu_n21556), .Y(exu_n12326));
INVX1 exu_U32855(.A(exu_n21562), .Y(exu_n12327));
INVX1 exu_U32856(.A(exu_n21568), .Y(exu_n12328));
INVX1 exu_U32857(.A(exu_n21574), .Y(exu_n12329));
INVX1 exu_U32858(.A(exu_n21580), .Y(exu_n12330));
INVX1 exu_U32859(.A(exu_n21586), .Y(exu_n12331));
INVX1 exu_U32860(.A(exu_n21592), .Y(exu_n12332));
INVX1 exu_U32861(.A(exu_n21598), .Y(exu_n12333));
INVX1 exu_U32862(.A(exu_n21604), .Y(exu_n12334));
INVX1 exu_U32863(.A(exu_n21610), .Y(exu_n12335));
INVX1 exu_U32864(.A(exu_n21616), .Y(exu_n12336));
INVX1 exu_U32865(.A(exu_n21622), .Y(exu_n12337));
INVX1 exu_U32866(.A(exu_n23201), .Y(exu_n12338));
INVX1 exu_U32867(.A(exu_n23207), .Y(exu_n12339));
INVX1 exu_U32868(.A(exu_n23213), .Y(exu_n12340));
INVX1 exu_U32869(.A(exu_n23219), .Y(exu_n12341));
INVX1 exu_U32870(.A(exu_n23225), .Y(exu_n12342));
INVX1 exu_U32871(.A(exu_n23231), .Y(exu_n12343));
INVX1 exu_U32872(.A(exu_n23237), .Y(exu_n12344));
INVX1 exu_U32873(.A(exu_n23243), .Y(exu_n12345));
INVX1 exu_U32874(.A(exu_n23249), .Y(exu_n12346));
INVX1 exu_U32875(.A(exu_n23255), .Y(exu_n12347));
INVX1 exu_U32876(.A(exu_n23261), .Y(exu_n12348));
INVX1 exu_U32877(.A(exu_n23267), .Y(exu_n12349));
INVX1 exu_U32878(.A(exu_n23273), .Y(exu_n12350));
INVX1 exu_U32879(.A(exu_n23279), .Y(exu_n12351));
INVX1 exu_U32880(.A(exu_n23285), .Y(exu_n12352));
INVX1 exu_U32881(.A(exu_n23291), .Y(exu_n12353));
INVX1 exu_U32882(.A(exu_n23297), .Y(exu_n12354));
INVX1 exu_U32883(.A(exu_n23303), .Y(exu_n12355));
INVX1 exu_U32884(.A(exu_n23309), .Y(exu_n12356));
INVX1 exu_U32885(.A(exu_n23315), .Y(exu_n12357));
INVX1 exu_U32886(.A(exu_n23321), .Y(exu_n12358));
INVX1 exu_U32887(.A(exu_n23327), .Y(exu_n12359));
INVX1 exu_U32888(.A(exu_n23333), .Y(exu_n12360));
INVX1 exu_U32889(.A(exu_n23339), .Y(exu_n12361));
INVX1 exu_U32890(.A(exu_n23345), .Y(exu_n12362));
INVX1 exu_U32891(.A(exu_n23351), .Y(exu_n12363));
INVX1 exu_U32892(.A(exu_n23357), .Y(exu_n12364));
INVX1 exu_U32893(.A(exu_n23363), .Y(exu_n12365));
INVX1 exu_U32894(.A(exu_n23369), .Y(exu_n12366));
INVX1 exu_U32895(.A(exu_n23375), .Y(exu_n12367));
INVX1 exu_U32896(.A(exu_n23381), .Y(exu_n12368));
INVX1 exu_U32897(.A(exu_n23387), .Y(exu_n12369));
INVX1 exu_U32898(.A(exu_n23393), .Y(exu_n12370));
INVX1 exu_U32899(.A(exu_n23399), .Y(exu_n12371));
INVX1 exu_U32900(.A(exu_n23405), .Y(exu_n12372));
INVX1 exu_U32901(.A(exu_n23411), .Y(exu_n12373));
INVX1 exu_U32902(.A(exu_n23417), .Y(exu_n12374));
INVX1 exu_U32903(.A(exu_n23423), .Y(exu_n12375));
INVX1 exu_U32904(.A(exu_n23429), .Y(exu_n12376));
INVX1 exu_U32905(.A(exu_n23435), .Y(exu_n12377));
INVX1 exu_U32906(.A(exu_n23441), .Y(exu_n12378));
INVX1 exu_U32907(.A(exu_n23447), .Y(exu_n12379));
INVX1 exu_U32908(.A(exu_n23453), .Y(exu_n12380));
INVX1 exu_U32909(.A(exu_n23459), .Y(exu_n12381));
INVX1 exu_U32910(.A(exu_n23465), .Y(exu_n12382));
INVX1 exu_U32911(.A(exu_n23471), .Y(exu_n12383));
INVX1 exu_U32912(.A(exu_n23477), .Y(exu_n12384));
INVX1 exu_U32913(.A(exu_n23483), .Y(exu_n12385));
INVX1 exu_U32914(.A(exu_n23489), .Y(exu_n12386));
INVX1 exu_U32915(.A(exu_n23495), .Y(exu_n12387));
INVX1 exu_U32916(.A(exu_n23501), .Y(exu_n12388));
INVX1 exu_U32917(.A(exu_n23507), .Y(exu_n12389));
INVX1 exu_U32918(.A(exu_n23513), .Y(exu_n12390));
INVX1 exu_U32919(.A(exu_n23519), .Y(exu_n12391));
INVX1 exu_U32920(.A(exu_n23525), .Y(exu_n12392));
INVX1 exu_U32921(.A(exu_n23531), .Y(exu_n12393));
INVX1 exu_U32922(.A(exu_n23537), .Y(exu_n12394));
INVX1 exu_U32923(.A(exu_n23543), .Y(exu_n12395));
INVX1 exu_U32924(.A(exu_n23549), .Y(exu_n12396));
INVX1 exu_U32925(.A(exu_n23555), .Y(exu_n12397));
INVX1 exu_U32926(.A(exu_n23561), .Y(exu_n12398));
INVX1 exu_U32927(.A(exu_n23567), .Y(exu_n12399));
INVX1 exu_U32928(.A(exu_n23573), .Y(exu_n12400));
INVX1 exu_U32929(.A(exu_n23579), .Y(exu_n12401));
INVX1 exu_U32930(.A(exu_n23585), .Y(exu_n12402));
INVX1 exu_U32931(.A(exu_n23591), .Y(exu_n12403));
INVX1 exu_U32932(.A(exu_n23597), .Y(exu_n12404));
INVX1 exu_U32933(.A(exu_n23603), .Y(exu_n12405));
INVX1 exu_U32934(.A(exu_n23609), .Y(exu_n12406));
INVX1 exu_U32935(.A(exu_n23614), .Y(exu_n12407));
INVX1 exu_U32936(.A(exu_n23619), .Y(exu_n12408));
INVX1 exu_U32937(.A(exu_n23624), .Y(exu_n12409));
INVX1 exu_U32938(.A(exu_n23629), .Y(exu_n12410));
INVX1 exu_U32939(.A(exu_n23635), .Y(exu_n12411));
INVX1 exu_U32940(.A(exu_n23640), .Y(exu_n12412));
INVX1 exu_U32941(.A(exu_n23645), .Y(exu_n12413));
INVX1 exu_U32942(.A(exu_n23650), .Y(exu_n12414));
INVX1 exu_U32943(.A(exu_n23655), .Y(exu_n12415));
INVX1 exu_U32944(.A(exu_n23660), .Y(exu_n12416));
INVX1 exu_U32945(.A(exu_n23665), .Y(exu_n12417));
INVX1 exu_U32946(.A(exu_n23670), .Y(exu_n12418));
INVX1 exu_U32947(.A(exu_n23675), .Y(exu_n12419));
INVX1 exu_U32948(.A(exu_n23680), .Y(exu_n12420));
INVX1 exu_U32949(.A(exu_n23685), .Y(exu_n12421));
INVX1 exu_U32950(.A(exu_n23691), .Y(exu_n12422));
INVX1 exu_U32951(.A(exu_n23696), .Y(exu_n12423));
INVX1 exu_U32952(.A(exu_n23701), .Y(exu_n12424));
INVX1 exu_U32953(.A(exu_n23707), .Y(exu_n12425));
INVX1 exu_U32954(.A(exu_n23713), .Y(exu_n12426));
INVX1 exu_U32955(.A(exu_n23719), .Y(exu_n12427));
INVX1 exu_U32956(.A(exu_n23725), .Y(exu_n12428));
INVX1 exu_U32957(.A(exu_n23731), .Y(exu_n12429));
INVX1 exu_U32958(.A(exu_n23737), .Y(exu_n12430));
INVX1 exu_U32959(.A(exu_n23743), .Y(exu_n12431));
INVX1 exu_U32960(.A(exu_n23749), .Y(exu_n12432));
INVX1 exu_U32961(.A(exu_n23755), .Y(exu_n12433));
INVX1 exu_U32962(.A(exu_n23761), .Y(exu_n12434));
INVX1 exu_U32963(.A(exu_n23767), .Y(exu_n12435));
INVX1 exu_U32964(.A(exu_n23773), .Y(exu_n12436));
INVX1 exu_U32965(.A(exu_n23779), .Y(exu_n12437));
INVX1 exu_U32966(.A(exu_n23785), .Y(exu_n12438));
INVX1 exu_U32967(.A(exu_n23791), .Y(exu_n12439));
INVX1 exu_U32968(.A(exu_n23797), .Y(exu_n12440));
INVX1 exu_U32969(.A(exu_n23803), .Y(exu_n12441));
INVX1 exu_U32970(.A(exu_n23809), .Y(exu_n12442));
INVX1 exu_U32971(.A(exu_n23815), .Y(exu_n12443));
INVX1 exu_U32972(.A(exu_n23821), .Y(exu_n12444));
INVX1 exu_U32973(.A(exu_n23827), .Y(exu_n12445));
INVX1 exu_U32974(.A(exu_n23833), .Y(exu_n12446));
INVX1 exu_U32975(.A(exu_n23839), .Y(exu_n12447));
INVX1 exu_U32976(.A(exu_n23845), .Y(exu_n12448));
INVX1 exu_U32977(.A(exu_n23851), .Y(exu_n12449));
INVX1 exu_U32978(.A(exu_n23857), .Y(exu_n12450));
INVX1 exu_U32979(.A(exu_n23863), .Y(exu_n12451));
INVX1 exu_U32980(.A(exu_n23869), .Y(exu_n12452));
INVX1 exu_U32981(.A(exu_n23875), .Y(exu_n12453));
INVX1 exu_U32982(.A(exu_n23881), .Y(exu_n12454));
INVX1 exu_U32983(.A(exu_n23887), .Y(exu_n12455));
INVX1 exu_U32984(.A(exu_n23893), .Y(exu_n12456));
INVX1 exu_U32985(.A(exu_n23899), .Y(exu_n12457));
INVX1 exu_U32986(.A(exu_n23905), .Y(exu_n12458));
INVX1 exu_U32987(.A(exu_n23911), .Y(exu_n12459));
INVX1 exu_U32988(.A(exu_n23917), .Y(exu_n12460));
INVX1 exu_U32989(.A(exu_n23923), .Y(exu_n12461));
INVX1 exu_U32990(.A(exu_n23929), .Y(exu_n12462));
INVX1 exu_U32991(.A(exu_n23935), .Y(exu_n12463));
INVX1 exu_U32992(.A(exu_n23941), .Y(exu_n12464));
INVX1 exu_U32993(.A(exu_n23947), .Y(exu_n12465));
INVX1 exu_U32994(.A(exu_n23953), .Y(exu_n12466));
INVX1 exu_U32995(.A(exu_n23959), .Y(exu_n12467));
INVX1 exu_U32996(.A(exu_n23965), .Y(exu_n12468));
INVX1 exu_U32997(.A(exu_n23971), .Y(exu_n12469));
INVX1 exu_U32998(.A(exu_n23977), .Y(exu_n12470));
INVX1 exu_U32999(.A(exu_n23983), .Y(exu_n12471));
INVX1 exu_U33000(.A(exu_n23989), .Y(exu_n12472));
INVX1 exu_U33001(.A(exu_n23995), .Y(exu_n12473));
INVX1 exu_U33002(.A(exu_n24001), .Y(exu_n12474));
INVX1 exu_U33003(.A(exu_n24007), .Y(exu_n12475));
INVX1 exu_U33004(.A(exu_n24013), .Y(exu_n12476));
INVX1 exu_U33005(.A(exu_n24019), .Y(exu_n12477));
INVX1 exu_U33006(.A(exu_n24025), .Y(exu_n12478));
INVX1 exu_U33007(.A(exu_n24031), .Y(exu_n12479));
INVX1 exu_U33008(.A(exu_n24037), .Y(exu_n12480));
INVX1 exu_U33009(.A(exu_n24043), .Y(exu_n12481));
INVX1 exu_U33010(.A(exu_n24049), .Y(exu_n12482));
INVX1 exu_U33011(.A(exu_n24055), .Y(exu_n12483));
INVX1 exu_U33012(.A(exu_n24061), .Y(exu_n12484));
INVX1 exu_U33013(.A(exu_n24067), .Y(exu_n12485));
INVX1 exu_U33014(.A(exu_n24073), .Y(exu_n12486));
INVX1 exu_U33015(.A(exu_n24079), .Y(exu_n12487));
INVX1 exu_U33016(.A(exu_n24085), .Y(exu_n12488));
INVX1 exu_U33017(.A(exu_n24091), .Y(exu_n12489));
INVX1 exu_U33018(.A(exu_n24097), .Y(exu_n12490));
INVX1 exu_U33019(.A(exu_n24103), .Y(exu_n12491));
INVX1 exu_U33020(.A(exu_n24109), .Y(exu_n12492));
INVX1 exu_U33021(.A(exu_n24115), .Y(exu_n12493));
INVX1 exu_U33022(.A(exu_n24121), .Y(exu_n12494));
INVX1 exu_U33023(.A(exu_n24127), .Y(exu_n12495));
INVX1 exu_U33024(.A(exu_n24133), .Y(exu_n12496));
INVX1 exu_U33025(.A(exu_n24139), .Y(exu_n12497));
INVX1 exu_U33026(.A(exu_n24145), .Y(exu_n12498));
INVX1 exu_U33027(.A(exu_n24151), .Y(exu_n12499));
INVX1 exu_U33028(.A(exu_n24157), .Y(exu_n12500));
INVX1 exu_U33029(.A(exu_n24163), .Y(exu_n12501));
INVX1 exu_U33030(.A(exu_n24169), .Y(exu_n12502));
INVX1 exu_U33031(.A(exu_n24175), .Y(exu_n12503));
INVX1 exu_U33032(.A(exu_n24181), .Y(exu_n12504));
INVX1 exu_U33033(.A(exu_n24187), .Y(exu_n12505));
INVX1 exu_U33034(.A(exu_n24193), .Y(exu_n12506));
INVX1 exu_U33035(.A(exu_n24199), .Y(exu_n12507));
INVX1 exu_U33036(.A(exu_n24205), .Y(exu_n12508));
INVX1 exu_U33037(.A(exu_n24211), .Y(exu_n12509));
INVX1 exu_U33038(.A(exu_n24217), .Y(exu_n12510));
INVX1 exu_U33039(.A(exu_n24223), .Y(exu_n12511));
INVX1 exu_U33040(.A(exu_n24229), .Y(exu_n12512));
INVX1 exu_U33041(.A(exu_n24235), .Y(exu_n12513));
INVX1 exu_U33042(.A(exu_n24241), .Y(exu_n12514));
INVX1 exu_U33043(.A(exu_n24247), .Y(exu_n12515));
INVX1 exu_U33044(.A(exu_n24253), .Y(exu_n12516));
INVX1 exu_U33045(.A(exu_n24259), .Y(exu_n12517));
INVX1 exu_U33046(.A(exu_n24265), .Y(exu_n12518));
INVX1 exu_U33047(.A(exu_n24271), .Y(exu_n12519));
INVX1 exu_U33048(.A(exu_n24277), .Y(exu_n12520));
INVX1 exu_U33049(.A(exu_n24283), .Y(exu_n12521));
INVX1 exu_U33050(.A(exu_n24289), .Y(exu_n12522));
INVX1 exu_U33051(.A(exu_n24295), .Y(exu_n12523));
INVX1 exu_U33052(.A(exu_n24301), .Y(exu_n12524));
INVX1 exu_U33053(.A(exu_n24307), .Y(exu_n12525));
INVX1 exu_U33054(.A(exu_n24313), .Y(exu_n12526));
INVX1 exu_U33055(.A(exu_n24319), .Y(exu_n12527));
INVX1 exu_U33056(.A(exu_n24325), .Y(exu_n12528));
INVX1 exu_U33057(.A(exu_n24331), .Y(exu_n12529));
INVX1 exu_U33058(.A(exu_n24337), .Y(exu_n12530));
INVX1 exu_U33059(.A(exu_n24341), .Y(exu_n12531));
INVX1 exu_U33060(.A(exu_n24345), .Y(exu_n12532));
INVX1 exu_U33061(.A(exu_n24349), .Y(exu_n12533));
INVX1 exu_U33062(.A(exu_n24353), .Y(exu_n12534));
INVX1 exu_U33063(.A(exu_n24357), .Y(exu_n12535));
INVX1 exu_U33064(.A(exu_n24361), .Y(exu_n12536));
INVX1 exu_U33065(.A(exu_n24365), .Y(exu_n12537));
INVX1 exu_U33066(.A(exu_n24369), .Y(exu_n12538));
INVX1 exu_U33067(.A(exu_n24373), .Y(exu_n12539));
INVX1 exu_U33068(.A(exu_n24377), .Y(exu_n12540));
INVX1 exu_U33069(.A(exu_n24381), .Y(exu_n12541));
INVX1 exu_U33070(.A(exu_n24385), .Y(exu_n12542));
INVX1 exu_U33071(.A(exu_n24389), .Y(exu_n12543));
INVX1 exu_U33072(.A(exu_n24393), .Y(exu_n12544));
INVX1 exu_U33073(.A(exu_n24397), .Y(exu_n12545));
INVX1 exu_U33074(.A(exu_n24401), .Y(exu_n12546));
INVX1 exu_U33075(.A(exu_n24405), .Y(exu_n12547));
INVX1 exu_U33076(.A(exu_n24409), .Y(exu_n12548));
INVX1 exu_U33077(.A(exu_n24413), .Y(exu_n12549));
INVX1 exu_U33078(.A(exu_n24417), .Y(exu_n12550));
INVX1 exu_U33079(.A(exu_n24421), .Y(exu_n12551));
INVX1 exu_U33080(.A(exu_n24425), .Y(exu_n12552));
INVX1 exu_U33081(.A(exu_n24429), .Y(exu_n12553));
INVX1 exu_U33082(.A(exu_n24433), .Y(exu_n12554));
INVX1 exu_U33083(.A(exu_n24437), .Y(exu_n12555));
INVX1 exu_U33084(.A(exu_n24441), .Y(exu_n12556));
INVX1 exu_U33085(.A(exu_n24445), .Y(exu_n12557));
INVX1 exu_U33086(.A(exu_n24449), .Y(exu_n12558));
INVX1 exu_U33087(.A(exu_n24453), .Y(exu_n12559));
INVX1 exu_U33088(.A(exu_n24457), .Y(exu_n12560));
INVX1 exu_U33089(.A(exu_n24461), .Y(exu_n12561));
INVX1 exu_U33090(.A(exu_n24465), .Y(exu_n12562));
INVX1 exu_U33091(.A(exu_n24469), .Y(exu_n12563));
INVX1 exu_U33092(.A(exu_n24473), .Y(exu_n12564));
INVX1 exu_U33093(.A(exu_n24477), .Y(exu_n12565));
INVX1 exu_U33094(.A(exu_n24481), .Y(exu_n12566));
INVX1 exu_U33095(.A(exu_n24485), .Y(exu_n12567));
INVX1 exu_U33096(.A(exu_n24489), .Y(exu_n12568));
INVX1 exu_U33097(.A(exu_n24493), .Y(exu_n12569));
INVX1 exu_U33098(.A(exu_n24497), .Y(exu_n12570));
INVX1 exu_U33099(.A(exu_n24501), .Y(exu_n12571));
INVX1 exu_U33100(.A(exu_n24505), .Y(exu_n12572));
INVX1 exu_U33101(.A(exu_n24509), .Y(exu_n12573));
INVX1 exu_U33102(.A(exu_n24513), .Y(exu_n12574));
INVX1 exu_U33103(.A(exu_n24517), .Y(exu_n12575));
INVX1 exu_U33104(.A(exu_n24521), .Y(exu_n12576));
INVX1 exu_U33105(.A(exu_n24525), .Y(exu_n12577));
INVX1 exu_U33106(.A(exu_n24529), .Y(exu_n12578));
INVX1 exu_U33107(.A(exu_n24533), .Y(exu_n12579));
INVX1 exu_U33108(.A(exu_n24537), .Y(exu_n12580));
INVX1 exu_U33109(.A(exu_n24541), .Y(exu_n12581));
INVX1 exu_U33110(.A(exu_n24545), .Y(exu_n12582));
INVX1 exu_U33111(.A(exu_n24549), .Y(exu_n12583));
INVX1 exu_U33112(.A(exu_n24553), .Y(exu_n12584));
INVX1 exu_U33113(.A(exu_n24557), .Y(exu_n12585));
INVX1 exu_U33114(.A(exu_n24561), .Y(exu_n12586));
INVX1 exu_U33115(.A(exu_n24565), .Y(exu_n12587));
INVX1 exu_U33116(.A(exu_n24569), .Y(exu_n12588));
INVX1 exu_U33117(.A(exu_n24573), .Y(exu_n12589));
INVX1 exu_U33118(.A(exu_n24577), .Y(exu_n12590));
INVX1 exu_U33119(.A(exu_n24581), .Y(exu_n12591));
INVX1 exu_U33120(.A(exu_n24585), .Y(exu_n12592));
INVX1 exu_U33121(.A(exu_n24589), .Y(exu_n12593));
INVX1 exu_U33122(.A(exu_n24593), .Y(exu_n12594));
INVX1 exu_U33123(.A(exu_n24599), .Y(exu_n12595));
INVX1 exu_U33124(.A(exu_n24605), .Y(exu_n12596));
INVX1 exu_U33125(.A(exu_n24611), .Y(exu_n12597));
INVX1 exu_U33126(.A(exu_n24617), .Y(exu_n12598));
INVX1 exu_U33127(.A(exu_n24623), .Y(exu_n12599));
INVX1 exu_U33128(.A(exu_n24629), .Y(exu_n12600));
INVX1 exu_U33129(.A(exu_n24635), .Y(exu_n12601));
INVX1 exu_U33130(.A(exu_n24641), .Y(exu_n12602));
INVX1 exu_U33131(.A(exu_n24647), .Y(exu_n12603));
INVX1 exu_U33132(.A(exu_n24653), .Y(exu_n12604));
INVX1 exu_U33133(.A(exu_n24659), .Y(exu_n12605));
INVX1 exu_U33134(.A(exu_n24665), .Y(exu_n12606));
INVX1 exu_U33135(.A(exu_n24671), .Y(exu_n12607));
INVX1 exu_U33136(.A(exu_n24677), .Y(exu_n12608));
INVX1 exu_U33137(.A(exu_n24683), .Y(exu_n12609));
INVX1 exu_U33138(.A(exu_n24689), .Y(exu_n12610));
INVX1 exu_U33139(.A(exu_n24695), .Y(exu_n12611));
INVX1 exu_U33140(.A(exu_n24701), .Y(exu_n12612));
INVX1 exu_U33141(.A(exu_n24707), .Y(exu_n12613));
INVX1 exu_U33142(.A(exu_n24713), .Y(exu_n12614));
INVX1 exu_U33143(.A(exu_n24719), .Y(exu_n12615));
INVX1 exu_U33144(.A(exu_n24725), .Y(exu_n12616));
INVX1 exu_U33145(.A(exu_n24731), .Y(exu_n12617));
INVX1 exu_U33146(.A(exu_n24737), .Y(exu_n12618));
INVX1 exu_U33147(.A(exu_n24743), .Y(exu_n12619));
INVX1 exu_U33148(.A(exu_n24749), .Y(exu_n12620));
INVX1 exu_U33149(.A(exu_n24755), .Y(exu_n12621));
INVX1 exu_U33150(.A(exu_n24761), .Y(exu_n12622));
INVX1 exu_U33151(.A(exu_n24767), .Y(exu_n12623));
INVX1 exu_U33152(.A(exu_n24773), .Y(exu_n12624));
INVX1 exu_U33153(.A(exu_n24779), .Y(exu_n12625));
INVX1 exu_U33154(.A(exu_n24785), .Y(exu_n12626));
INVX1 exu_U33155(.A(exu_n24791), .Y(exu_n12627));
INVX1 exu_U33156(.A(exu_n24797), .Y(exu_n12628));
INVX1 exu_U33157(.A(exu_n24803), .Y(exu_n12629));
INVX1 exu_U33158(.A(exu_n24809), .Y(exu_n12630));
INVX1 exu_U33159(.A(exu_n24815), .Y(exu_n12631));
INVX1 exu_U33160(.A(exu_n24821), .Y(exu_n12632));
INVX1 exu_U33161(.A(exu_n24827), .Y(exu_n12633));
INVX1 exu_U33162(.A(exu_n24833), .Y(exu_n12634));
INVX1 exu_U33163(.A(exu_n24839), .Y(exu_n12635));
INVX1 exu_U33164(.A(exu_n24845), .Y(exu_n12636));
INVX1 exu_U33165(.A(exu_n24851), .Y(exu_n12637));
INVX1 exu_U33166(.A(exu_n24857), .Y(exu_n12638));
INVX1 exu_U33167(.A(exu_n24863), .Y(exu_n12639));
INVX1 exu_U33168(.A(exu_n24869), .Y(exu_n12640));
INVX1 exu_U33169(.A(exu_n24875), .Y(exu_n12641));
INVX1 exu_U33170(.A(exu_n24881), .Y(exu_n12642));
INVX1 exu_U33171(.A(exu_n24887), .Y(exu_n12643));
INVX1 exu_U33172(.A(exu_n24893), .Y(exu_n12644));
INVX1 exu_U33173(.A(exu_n24899), .Y(exu_n12645));
INVX1 exu_U33174(.A(exu_n24905), .Y(exu_n12646));
INVX1 exu_U33175(.A(exu_n24911), .Y(exu_n12647));
INVX1 exu_U33176(.A(exu_n24917), .Y(exu_n12648));
INVX1 exu_U33177(.A(exu_n24923), .Y(exu_n12649));
INVX1 exu_U33178(.A(exu_n24929), .Y(exu_n12650));
INVX1 exu_U33179(.A(exu_n24935), .Y(exu_n12651));
INVX1 exu_U33180(.A(exu_n24941), .Y(exu_n12652));
INVX1 exu_U33181(.A(exu_n24947), .Y(exu_n12653));
INVX1 exu_U33182(.A(exu_n24953), .Y(exu_n12654));
INVX1 exu_U33183(.A(exu_n24959), .Y(exu_n12655));
INVX1 exu_U33184(.A(exu_n24965), .Y(exu_n12656));
INVX1 exu_U33185(.A(exu_n24971), .Y(exu_n12657));
INVX1 exu_U33186(.A(exu_n24977), .Y(exu_n12658));
INVX1 exu_U33187(.A(exu_n24983), .Y(exu_n12659));
INVX1 exu_U33188(.A(exu_n24989), .Y(exu_n12660));
INVX1 exu_U33189(.A(exu_n24995), .Y(exu_n12661));
INVX1 exu_U33190(.A(exu_n25001), .Y(exu_n12662));
INVX1 exu_U33191(.A(exu_n25006), .Y(exu_n12663));
INVX1 exu_U33192(.A(exu_n25011), .Y(exu_n12664));
INVX1 exu_U33193(.A(exu_n25016), .Y(exu_n12665));
INVX1 exu_U33194(.A(exu_n25021), .Y(exu_n12666));
INVX1 exu_U33195(.A(exu_n25027), .Y(exu_n12667));
INVX1 exu_U33196(.A(exu_n25032), .Y(exu_n12668));
INVX1 exu_U33197(.A(exu_n25037), .Y(exu_n12669));
INVX1 exu_U33198(.A(exu_n25042), .Y(exu_n12670));
INVX1 exu_U33199(.A(exu_n25047), .Y(exu_n12671));
INVX1 exu_U33200(.A(exu_n25052), .Y(exu_n12672));
INVX1 exu_U33201(.A(exu_n25057), .Y(exu_n12673));
INVX1 exu_U33202(.A(exu_n25062), .Y(exu_n12674));
INVX1 exu_U33203(.A(exu_n25067), .Y(exu_n12675));
INVX1 exu_U33204(.A(exu_n25072), .Y(exu_n12676));
INVX1 exu_U33205(.A(exu_n25077), .Y(exu_n12677));
INVX1 exu_U33206(.A(exu_n25083), .Y(exu_n12678));
INVX1 exu_U33207(.A(exu_n25088), .Y(exu_n12679));
INVX1 exu_U33208(.A(exu_n25093), .Y(exu_n12680));
INVX1 exu_U33209(.A(exu_n25098), .Y(exu_n12681));
INVX1 exu_U33210(.A(exu_n25103), .Y(exu_n12682));
INVX1 exu_U33211(.A(exu_n25108), .Y(exu_n12683));
INVX1 exu_U33212(.A(exu_n25113), .Y(exu_n12684));
INVX1 exu_U33213(.A(exu_n25118), .Y(exu_n12685));
INVX1 exu_U33214(.A(exu_n25123), .Y(exu_n12686));
INVX1 exu_U33215(.A(exu_n25128), .Y(exu_n12687));
INVX1 exu_U33216(.A(exu_n25133), .Y(exu_n12688));
INVX1 exu_U33217(.A(exu_n25139), .Y(exu_n12689));
INVX1 exu_U33218(.A(exu_n25144), .Y(exu_n12690));
INVX1 exu_U33219(.A(exu_n25149), .Y(exu_n12691));
INVX1 exu_U33220(.A(exu_n25154), .Y(exu_n12692));
INVX1 exu_U33221(.A(exu_n25159), .Y(exu_n12693));
INVX1 exu_U33222(.A(exu_n25164), .Y(exu_n12694));
INVX1 exu_U33223(.A(exu_n25169), .Y(exu_n12695));
INVX1 exu_U33224(.A(exu_n25174), .Y(exu_n12696));
INVX1 exu_U33225(.A(exu_n25179), .Y(exu_n12697));
INVX1 exu_U33226(.A(exu_n25185), .Y(exu_n12698));
INVX1 exu_U33227(.A(exu_n25191), .Y(exu_n12699));
INVX1 exu_U33228(.A(exu_n25197), .Y(exu_n12700));
INVX1 exu_U33229(.A(exu_n25203), .Y(exu_n12701));
INVX1 exu_U33230(.A(exu_n25209), .Y(exu_n12702));
INVX1 exu_U33231(.A(exu_n25215), .Y(exu_n12703));
INVX1 exu_U33232(.A(exu_n25221), .Y(exu_n12704));
INVX1 exu_U33233(.A(exu_n25227), .Y(exu_n12705));
INVX1 exu_U33234(.A(exu_n25233), .Y(exu_n12706));
INVX1 exu_U33235(.A(exu_n25239), .Y(exu_n12707));
INVX1 exu_U33236(.A(exu_n25245), .Y(exu_n12708));
INVX1 exu_U33237(.A(exu_n25251), .Y(exu_n12709));
INVX1 exu_U33238(.A(exu_n25257), .Y(exu_n12710));
INVX1 exu_U33239(.A(exu_n25263), .Y(exu_n12711));
INVX1 exu_U33240(.A(exu_n25269), .Y(exu_n12712));
INVX1 exu_U33241(.A(exu_n25275), .Y(exu_n12713));
INVX1 exu_U33242(.A(exu_n25281), .Y(exu_n12714));
INVX1 exu_U33243(.A(exu_n25287), .Y(exu_n12715));
INVX1 exu_U33244(.A(exu_n25293), .Y(exu_n12716));
INVX1 exu_U33245(.A(exu_n25299), .Y(exu_n12717));
INVX1 exu_U33246(.A(exu_n25305), .Y(exu_n12718));
INVX1 exu_U33247(.A(exu_n25311), .Y(exu_n12719));
INVX1 exu_U33248(.A(exu_n25317), .Y(exu_n12720));
INVX1 exu_U33249(.A(exu_n25323), .Y(exu_n12721));
INVX1 exu_U33250(.A(exu_n25329), .Y(exu_n12722));
INVX1 exu_U33251(.A(exu_n25335), .Y(exu_n12723));
INVX1 exu_U33252(.A(exu_n25341), .Y(exu_n12724));
INVX1 exu_U33253(.A(exu_n25347), .Y(exu_n12725));
INVX1 exu_U33254(.A(exu_n25353), .Y(exu_n12726));
INVX1 exu_U33255(.A(exu_n25359), .Y(exu_n12727));
INVX1 exu_U33256(.A(exu_n25365), .Y(exu_n12728));
INVX1 exu_U33257(.A(exu_n25371), .Y(exu_n12729));
INVX1 exu_U33258(.A(exu_n25377), .Y(exu_n12730));
INVX1 exu_U33259(.A(exu_n25383), .Y(exu_n12731));
INVX1 exu_U33260(.A(exu_n25389), .Y(exu_n12732));
INVX1 exu_U33261(.A(exu_n25395), .Y(exu_n12733));
INVX1 exu_U33262(.A(exu_n25401), .Y(exu_n12734));
INVX1 exu_U33263(.A(exu_n25407), .Y(exu_n12735));
INVX1 exu_U33264(.A(exu_n25413), .Y(exu_n12736));
INVX1 exu_U33265(.A(exu_n25419), .Y(exu_n12737));
INVX1 exu_U33266(.A(exu_n25425), .Y(exu_n12738));
INVX1 exu_U33267(.A(exu_n25431), .Y(exu_n12739));
INVX1 exu_U33268(.A(exu_n25437), .Y(exu_n12740));
INVX1 exu_U33269(.A(exu_n25443), .Y(exu_n12741));
INVX1 exu_U33270(.A(exu_n25449), .Y(exu_n12742));
INVX1 exu_U33271(.A(exu_n25455), .Y(exu_n12743));
INVX1 exu_U33272(.A(exu_n25461), .Y(exu_n12744));
INVX1 exu_U33273(.A(exu_n25467), .Y(exu_n12745));
INVX1 exu_U33274(.A(exu_n25473), .Y(exu_n12746));
INVX1 exu_U33275(.A(exu_n25479), .Y(exu_n12747));
INVX1 exu_U33276(.A(exu_n25485), .Y(exu_n12748));
INVX1 exu_U33277(.A(exu_n25491), .Y(exu_n12749));
INVX1 exu_U33278(.A(exu_n25497), .Y(exu_n12750));
INVX1 exu_U33279(.A(exu_n25503), .Y(exu_n12751));
INVX1 exu_U33280(.A(exu_n25509), .Y(exu_n12752));
INVX1 exu_U33281(.A(exu_n25515), .Y(exu_n12753));
INVX1 exu_U33282(.A(exu_n25521), .Y(exu_n12754));
INVX1 exu_U33283(.A(exu_n25527), .Y(exu_n12755));
INVX1 exu_U33284(.A(exu_n25533), .Y(exu_n12756));
INVX1 exu_U33285(.A(exu_n25539), .Y(exu_n12757));
INVX1 exu_U33286(.A(exu_n25545), .Y(exu_n12758));
INVX1 exu_U33287(.A(exu_n25551), .Y(exu_n12759));
INVX1 exu_U33288(.A(exu_n25557), .Y(exu_n12760));
INVX1 exu_U33289(.A(exu_n25563), .Y(exu_n12761));
INVX1 exu_U33290(.A(exu_n25569), .Y(exu_n12762));
INVX1 exu_U33291(.A(exu_n25575), .Y(exu_n12763));
INVX1 exu_U33292(.A(exu_n25581), .Y(exu_n12764));
INVX1 exu_U33293(.A(exu_n25587), .Y(exu_n12765));
INVX1 exu_U33294(.A(exu_n25593), .Y(exu_n12766));
INVX1 exu_U33295(.A(exu_n25599), .Y(exu_n12767));
INVX1 exu_U33296(.A(exu_n25605), .Y(exu_n12768));
INVX1 exu_U33297(.A(exu_n25611), .Y(exu_n12769));
INVX1 exu_U33298(.A(exu_n25617), .Y(exu_n12770));
INVX1 exu_U33299(.A(exu_n25623), .Y(exu_n12771));
INVX1 exu_U33300(.A(exu_n25629), .Y(exu_n12772));
INVX1 exu_U33301(.A(exu_n25635), .Y(exu_n12773));
INVX1 exu_U33302(.A(exu_n25641), .Y(exu_n12774));
INVX1 exu_U33303(.A(exu_n25647), .Y(exu_n12775));
INVX1 exu_U33304(.A(exu_n25653), .Y(exu_n12776));
INVX1 exu_U33305(.A(exu_n25659), .Y(exu_n12777));
INVX1 exu_U33306(.A(exu_n25665), .Y(exu_n12778));
INVX1 exu_U33307(.A(exu_n25671), .Y(exu_n12779));
INVX1 exu_U33308(.A(exu_n25677), .Y(exu_n12780));
INVX1 exu_U33309(.A(exu_n25683), .Y(exu_n12781));
INVX1 exu_U33310(.A(exu_n25689), .Y(exu_n12782));
INVX1 exu_U33311(.A(exu_n25695), .Y(exu_n12783));
INVX1 exu_U33312(.A(exu_n25701), .Y(exu_n12784));
INVX1 exu_U33313(.A(exu_n25707), .Y(exu_n12785));
INVX1 exu_U33314(.A(exu_n25713), .Y(exu_n12786));
INVX1 exu_U33315(.A(exu_n25717), .Y(exu_n12787));
INVX1 exu_U33316(.A(exu_n25721), .Y(exu_n12788));
INVX1 exu_U33317(.A(exu_n25725), .Y(exu_n12789));
INVX1 exu_U33318(.A(exu_n25729), .Y(exu_n12790));
INVX1 exu_U33319(.A(exu_n25733), .Y(exu_n12791));
INVX1 exu_U33320(.A(exu_n25737), .Y(exu_n12792));
INVX1 exu_U33321(.A(exu_n25741), .Y(exu_n12793));
INVX1 exu_U33322(.A(exu_n25745), .Y(exu_n12794));
INVX1 exu_U33323(.A(exu_n25749), .Y(exu_n12795));
INVX1 exu_U33324(.A(exu_n25753), .Y(exu_n12796));
INVX1 exu_U33325(.A(exu_n25757), .Y(exu_n12797));
INVX1 exu_U33326(.A(exu_n25761), .Y(exu_n12798));
INVX1 exu_U33327(.A(exu_n25765), .Y(exu_n12799));
INVX1 exu_U33328(.A(exu_n25769), .Y(exu_n12800));
INVX1 exu_U33329(.A(exu_n25773), .Y(exu_n12801));
INVX1 exu_U33330(.A(exu_n25777), .Y(exu_n12802));
INVX1 exu_U33331(.A(exu_n25781), .Y(exu_n12803));
INVX1 exu_U33332(.A(exu_n25785), .Y(exu_n12804));
INVX1 exu_U33333(.A(exu_n25789), .Y(exu_n12805));
INVX1 exu_U33334(.A(exu_n25793), .Y(exu_n12806));
INVX1 exu_U33335(.A(exu_n25797), .Y(exu_n12807));
INVX1 exu_U33336(.A(exu_n25801), .Y(exu_n12808));
INVX1 exu_U33337(.A(exu_n25805), .Y(exu_n12809));
INVX1 exu_U33338(.A(exu_n25809), .Y(exu_n12810));
INVX1 exu_U33339(.A(exu_n25813), .Y(exu_n12811));
INVX1 exu_U33340(.A(exu_n25817), .Y(exu_n12812));
INVX1 exu_U33341(.A(exu_n25821), .Y(exu_n12813));
INVX1 exu_U33342(.A(exu_n25825), .Y(exu_n12814));
INVX1 exu_U33343(.A(exu_n25829), .Y(exu_n12815));
INVX1 exu_U33344(.A(exu_n25833), .Y(exu_n12816));
INVX1 exu_U33345(.A(exu_n25837), .Y(exu_n12817));
INVX1 exu_U33346(.A(exu_n25841), .Y(exu_n12818));
INVX1 exu_U33347(.A(exu_n25845), .Y(exu_n12819));
INVX1 exu_U33348(.A(exu_n25849), .Y(exu_n12820));
INVX1 exu_U33349(.A(exu_n25853), .Y(exu_n12821));
INVX1 exu_U33350(.A(exu_n25857), .Y(exu_n12822));
INVX1 exu_U33351(.A(exu_n25861), .Y(exu_n12823));
INVX1 exu_U33352(.A(exu_n25865), .Y(exu_n12824));
INVX1 exu_U33353(.A(exu_n25869), .Y(exu_n12825));
INVX1 exu_U33354(.A(exu_n25873), .Y(exu_n12826));
INVX1 exu_U33355(.A(exu_n25877), .Y(exu_n12827));
INVX1 exu_U33356(.A(exu_n25881), .Y(exu_n12828));
INVX1 exu_U33357(.A(exu_n25885), .Y(exu_n12829));
INVX1 exu_U33358(.A(exu_n25889), .Y(exu_n12830));
INVX1 exu_U33359(.A(exu_n25893), .Y(exu_n12831));
INVX1 exu_U33360(.A(exu_n25897), .Y(exu_n12832));
INVX1 exu_U33361(.A(exu_n25901), .Y(exu_n12833));
INVX1 exu_U33362(.A(exu_n25905), .Y(exu_n12834));
INVX1 exu_U33363(.A(exu_n25909), .Y(exu_n12835));
INVX1 exu_U33364(.A(exu_n25913), .Y(exu_n12836));
INVX1 exu_U33365(.A(exu_n25917), .Y(exu_n12837));
INVX1 exu_U33366(.A(exu_n25921), .Y(exu_n12838));
INVX1 exu_U33367(.A(exu_n25925), .Y(exu_n12839));
INVX1 exu_U33368(.A(exu_n25929), .Y(exu_n12840));
INVX1 exu_U33369(.A(exu_n25933), .Y(exu_n12841));
INVX1 exu_U33370(.A(exu_n25937), .Y(exu_n12842));
INVX1 exu_U33371(.A(exu_n25941), .Y(exu_n12843));
INVX1 exu_U33372(.A(exu_n25945), .Y(exu_n12844));
INVX1 exu_U33373(.A(exu_n25949), .Y(exu_n12845));
INVX1 exu_U33374(.A(exu_n25953), .Y(exu_n12846));
INVX1 exu_U33375(.A(exu_n25957), .Y(exu_n12847));
INVX1 exu_U33376(.A(exu_n25961), .Y(exu_n12848));
INVX1 exu_U33377(.A(exu_n25965), .Y(exu_n12849));
INVX1 exu_U33378(.A(exu_n25969), .Y(exu_n12850));
INVX1 exu_U33379(.A(exu_n25975), .Y(exu_n12851));
INVX1 exu_U33380(.A(exu_n25981), .Y(exu_n12852));
INVX1 exu_U33381(.A(exu_n25987), .Y(exu_n12853));
INVX1 exu_U33382(.A(exu_n25993), .Y(exu_n12854));
INVX1 exu_U33383(.A(exu_n25999), .Y(exu_n12855));
INVX1 exu_U33384(.A(exu_n26005), .Y(exu_n12856));
INVX1 exu_U33385(.A(exu_n26011), .Y(exu_n12857));
INVX1 exu_U33386(.A(exu_n26017), .Y(exu_n12858));
INVX1 exu_U33387(.A(exu_n26023), .Y(exu_n12859));
INVX1 exu_U33388(.A(exu_n26029), .Y(exu_n12860));
INVX1 exu_U33389(.A(exu_n26035), .Y(exu_n12861));
INVX1 exu_U33390(.A(exu_n26041), .Y(exu_n12862));
INVX1 exu_U33391(.A(exu_n26047), .Y(exu_n12863));
INVX1 exu_U33392(.A(exu_n26053), .Y(exu_n12864));
INVX1 exu_U33393(.A(exu_n26059), .Y(exu_n12865));
INVX1 exu_U33394(.A(exu_n26065), .Y(exu_n12866));
INVX1 exu_U33395(.A(exu_n26071), .Y(exu_n12867));
INVX1 exu_U33396(.A(exu_n26077), .Y(exu_n12868));
INVX1 exu_U33397(.A(exu_n26083), .Y(exu_n12869));
INVX1 exu_U33398(.A(exu_n26089), .Y(exu_n12870));
INVX1 exu_U33399(.A(exu_n26095), .Y(exu_n12871));
INVX1 exu_U33400(.A(exu_n26101), .Y(exu_n12872));
INVX1 exu_U33401(.A(exu_n26107), .Y(exu_n12873));
INVX1 exu_U33402(.A(exu_n26113), .Y(exu_n12874));
INVX1 exu_U33403(.A(exu_n26119), .Y(exu_n12875));
INVX1 exu_U33404(.A(exu_n26125), .Y(exu_n12876));
INVX1 exu_U33405(.A(exu_n26131), .Y(exu_n12877));
INVX1 exu_U33406(.A(exu_n26137), .Y(exu_n12878));
INVX1 exu_U33407(.A(exu_n26143), .Y(exu_n12879));
INVX1 exu_U33408(.A(exu_n26149), .Y(exu_n12880));
INVX1 exu_U33409(.A(exu_n26155), .Y(exu_n12881));
INVX1 exu_U33410(.A(exu_n26161), .Y(exu_n12882));
INVX1 exu_U33411(.A(exu_n26167), .Y(exu_n12883));
INVX1 exu_U33412(.A(exu_n26173), .Y(exu_n12884));
INVX1 exu_U33413(.A(exu_n26179), .Y(exu_n12885));
INVX1 exu_U33414(.A(exu_n26185), .Y(exu_n12886));
INVX1 exu_U33415(.A(exu_n26191), .Y(exu_n12887));
INVX1 exu_U33416(.A(exu_n26197), .Y(exu_n12888));
INVX1 exu_U33417(.A(exu_n26203), .Y(exu_n12889));
INVX1 exu_U33418(.A(exu_n26209), .Y(exu_n12890));
INVX1 exu_U33419(.A(exu_n26215), .Y(exu_n12891));
INVX1 exu_U33420(.A(exu_n26221), .Y(exu_n12892));
INVX1 exu_U33421(.A(exu_n26227), .Y(exu_n12893));
INVX1 exu_U33422(.A(exu_n26233), .Y(exu_n12894));
INVX1 exu_U33423(.A(exu_n26239), .Y(exu_n12895));
INVX1 exu_U33424(.A(exu_n26245), .Y(exu_n12896));
INVX1 exu_U33425(.A(exu_n26251), .Y(exu_n12897));
INVX1 exu_U33426(.A(exu_n26257), .Y(exu_n12898));
INVX1 exu_U33427(.A(exu_n26263), .Y(exu_n12899));
INVX1 exu_U33428(.A(exu_n26269), .Y(exu_n12900));
INVX1 exu_U33429(.A(exu_n26275), .Y(exu_n12901));
INVX1 exu_U33430(.A(exu_n26281), .Y(exu_n12902));
INVX1 exu_U33431(.A(exu_n26287), .Y(exu_n12903));
INVX1 exu_U33432(.A(exu_n26293), .Y(exu_n12904));
INVX1 exu_U33433(.A(exu_n26299), .Y(exu_n12905));
INVX1 exu_U33434(.A(exu_n26305), .Y(exu_n12906));
INVX1 exu_U33435(.A(exu_n26311), .Y(exu_n12907));
INVX1 exu_U33436(.A(exu_n26317), .Y(exu_n12908));
INVX1 exu_U33437(.A(exu_n26323), .Y(exu_n12909));
INVX1 exu_U33438(.A(exu_n26329), .Y(exu_n12910));
INVX1 exu_U33439(.A(exu_n26335), .Y(exu_n12911));
INVX1 exu_U33440(.A(exu_n26341), .Y(exu_n12912));
INVX1 exu_U33441(.A(exu_n26347), .Y(exu_n12913));
INVX1 exu_U33442(.A(exu_n26353), .Y(exu_n12914));
INVX1 exu_U33443(.A(exu_n26359), .Y(exu_n12915));
INVX1 exu_U33444(.A(exu_n26365), .Y(exu_n12916));
INVX1 exu_U33445(.A(exu_n26371), .Y(exu_n12917));
INVX1 exu_U33446(.A(exu_n26377), .Y(exu_n12918));
INVX1 exu_U33447(.A(exu_n26382), .Y(exu_n12919));
INVX1 exu_U33448(.A(exu_n26388), .Y(exu_n12920));
INVX1 exu_U33449(.A(exu_n26394), .Y(exu_n12921));
INVX1 exu_U33450(.A(exu_n26400), .Y(exu_n12922));
INVX1 exu_U33451(.A(exu_n26406), .Y(exu_n12923));
INVX1 exu_U33452(.A(exu_n26412), .Y(exu_n12924));
INVX1 exu_U33453(.A(exu_n26418), .Y(exu_n12925));
INVX1 exu_U33454(.A(exu_n26424), .Y(exu_n12926));
INVX1 exu_U33455(.A(exu_n26430), .Y(exu_n12927));
INVX1 exu_U33456(.A(exu_n26436), .Y(exu_n12928));
INVX1 exu_U33457(.A(exu_n26442), .Y(exu_n12929));
INVX1 exu_U33458(.A(exu_n26448), .Y(exu_n12930));
INVX1 exu_U33459(.A(exu_n26454), .Y(exu_n12931));
INVX1 exu_U33460(.A(exu_n26460), .Y(exu_n12932));
INVX1 exu_U33461(.A(exu_n26466), .Y(exu_n12933));
INVX1 exu_U33462(.A(exu_n26472), .Y(exu_n12934));
INVX1 exu_U33463(.A(exu_n26478), .Y(exu_n12935));
INVX1 exu_U33464(.A(exu_n26484), .Y(exu_n12936));
INVX1 exu_U33465(.A(exu_n26490), .Y(exu_n12937));
INVX1 exu_U33466(.A(exu_n26496), .Y(exu_n12938));
INVX1 exu_U33467(.A(exu_n26502), .Y(exu_n12939));
INVX1 exu_U33468(.A(exu_n26508), .Y(exu_n12940));
INVX1 exu_U33469(.A(exu_n26514), .Y(exu_n12941));
INVX1 exu_U33470(.A(exu_n26520), .Y(exu_n12942));
INVX1 exu_U33471(.A(exu_n26526), .Y(exu_n12943));
INVX1 exu_U33472(.A(exu_n26532), .Y(exu_n12944));
INVX1 exu_U33473(.A(exu_n26538), .Y(exu_n12945));
INVX1 exu_U33474(.A(exu_n26544), .Y(exu_n12946));
INVX1 exu_U33475(.A(exu_n26550), .Y(exu_n12947));
INVX1 exu_U33476(.A(exu_n26556), .Y(exu_n12948));
INVX1 exu_U33477(.A(exu_n26562), .Y(exu_n12949));
INVX1 exu_U33478(.A(exu_n26568), .Y(exu_n12950));
INVX1 exu_U33479(.A(exu_n26574), .Y(exu_n12951));
INVX1 exu_U33480(.A(exu_n26580), .Y(exu_n12952));
INVX1 exu_U33481(.A(exu_n26586), .Y(exu_n12953));
INVX1 exu_U33482(.A(exu_n26591), .Y(exu_n12954));
INVX1 exu_U33483(.A(exu_n26597), .Y(exu_n12955));
INVX1 exu_U33484(.A(exu_n26603), .Y(exu_n12956));
INVX1 exu_U33485(.A(exu_n26609), .Y(exu_n12957));
INVX1 exu_U33486(.A(exu_n26615), .Y(exu_n12958));
INVX1 exu_U33487(.A(exu_n26621), .Y(exu_n12959));
INVX1 exu_U33488(.A(exu_n26627), .Y(exu_n12960));
INVX1 exu_U33489(.A(exu_n26633), .Y(exu_n12961));
INVX1 exu_U33490(.A(exu_n26639), .Y(exu_n12962));
INVX1 exu_U33491(.A(exu_n26645), .Y(exu_n12963));
INVX1 exu_U33492(.A(exu_n26651), .Y(exu_n12964));
INVX1 exu_U33493(.A(exu_n26657), .Y(exu_n12965));
INVX1 exu_U33494(.A(exu_n26663), .Y(exu_n12966));
INVX1 exu_U33495(.A(exu_n26669), .Y(exu_n12967));
INVX1 exu_U33496(.A(exu_n26675), .Y(exu_n12968));
INVX1 exu_U33497(.A(exu_n26681), .Y(exu_n12969));
INVX1 exu_U33498(.A(exu_n26687), .Y(exu_n12970));
INVX1 exu_U33499(.A(exu_n26693), .Y(exu_n12971));
INVX1 exu_U33500(.A(exu_n26699), .Y(exu_n12972));
INVX1 exu_U33501(.A(exu_n26705), .Y(exu_n12973));
INVX1 exu_U33502(.A(exu_n26711), .Y(exu_n12974));
INVX1 exu_U33503(.A(exu_n26717), .Y(exu_n12975));
INVX1 exu_U33504(.A(exu_n26723), .Y(exu_n12976));
INVX1 exu_U33505(.A(exu_n26729), .Y(exu_n12977));
INVX1 exu_U33506(.A(exu_n26735), .Y(exu_n12978));
INVX1 exu_U33507(.A(exu_n26740), .Y(exu_n12979));
INVX1 exu_U33508(.A(exu_n26744), .Y(exu_n12980));
INVX1 exu_U33509(.A(exu_n26748), .Y(exu_n12981));
INVX1 exu_U33510(.A(exu_n26752), .Y(exu_n12982));
INVX1 exu_U33511(.A(exu_n26756), .Y(exu_n12983));
INVX1 exu_U33512(.A(exu_n26760), .Y(exu_n12984));
INVX1 exu_U33513(.A(exu_n26764), .Y(exu_n12985));
INVX1 exu_U33514(.A(exu_n26768), .Y(exu_n12986));
INVX1 exu_U33515(.A(exu_n26772), .Y(exu_n12987));
INVX1 exu_U33516(.A(exu_n26776), .Y(exu_n12988));
INVX1 exu_U33517(.A(exu_n26780), .Y(exu_n12989));
INVX1 exu_U33518(.A(exu_n26784), .Y(exu_n12990));
INVX1 exu_U33519(.A(exu_n26788), .Y(exu_n12991));
INVX1 exu_U33520(.A(exu_n26792), .Y(exu_n12992));
INVX1 exu_U33521(.A(exu_n26796), .Y(exu_n12993));
INVX1 exu_U33522(.A(exu_n26800), .Y(exu_n12994));
INVX1 exu_U33523(.A(exu_n26804), .Y(exu_n12995));
INVX1 exu_U33524(.A(exu_n26808), .Y(exu_n12996));
INVX1 exu_U33525(.A(exu_n26812), .Y(exu_n12997));
INVX1 exu_U33526(.A(exu_n26816), .Y(exu_n12998));
INVX1 exu_U33527(.A(exu_n26820), .Y(exu_n12999));
INVX1 exu_U33528(.A(exu_n26825), .Y(exu_n13000));
INVX1 exu_U33529(.A(exu_n26830), .Y(exu_n13001));
INVX1 exu_U33530(.A(exu_n26835), .Y(exu_n13002));
INVX1 exu_U33531(.A(exu_n26840), .Y(exu_n13003));
INVX1 exu_U33532(.A(exu_n26845), .Y(exu_n13004));
INVX1 exu_U33533(.A(exu_n26850), .Y(exu_n13005));
INVX1 exu_U33534(.A(exu_n26855), .Y(exu_n13006));
INVX1 exu_U33535(.A(exu_n26860), .Y(exu_n13007));
INVX1 exu_U33536(.A(exu_n26865), .Y(exu_n13008));
INVX1 exu_U33537(.A(exu_n26869), .Y(exu_n13009));
INVX1 exu_U33538(.A(exu_n26874), .Y(exu_n13010));
INVX1 exu_U33539(.A(exu_n26879), .Y(exu_n13011));
INVX1 exu_U33540(.A(exu_n26884), .Y(exu_n13012));
INVX1 exu_U33541(.A(exu_n26889), .Y(exu_n13013));
INVX1 exu_U33542(.A(exu_n26894), .Y(exu_n13014));
INVX1 exu_U33543(.A(exu_n26899), .Y(exu_n13015));
INVX1 exu_U33544(.A(exu_n26904), .Y(exu_n13016));
INVX1 exu_U33545(.A(exu_n26910), .Y(exu_n13017));
INVX1 exu_U33546(.A(exu_n26914), .Y(exu_n13018));
INVX1 exu_U33547(.A(exu_n26918), .Y(exu_n13019));
INVX1 exu_U33548(.A(exu_n26922), .Y(exu_n13020));
INVX1 exu_U33549(.A(exu_n26926), .Y(exu_n13021));
INVX1 exu_U33550(.A(exu_n26930), .Y(exu_n13022));
INVX1 exu_U33551(.A(exu_n26934), .Y(exu_n13023));
INVX1 exu_U33552(.A(exu_n26938), .Y(exu_n13024));
INVX1 exu_U33553(.A(exu_n26942), .Y(exu_n13025));
INVX1 exu_U33554(.A(exu_n26946), .Y(exu_n13026));
INVX1 exu_U33555(.A(exu_n26950), .Y(exu_n13027));
INVX1 exu_U33556(.A(exu_n26954), .Y(exu_n13028));
INVX1 exu_U33557(.A(exu_n26958), .Y(exu_n13029));
INVX1 exu_U33558(.A(exu_n26962), .Y(exu_n13030));
INVX1 exu_U33559(.A(exu_n26966), .Y(exu_n13031));
INVX1 exu_U33560(.A(exu_n26970), .Y(exu_n13032));
INVX1 exu_U33561(.A(exu_n26974), .Y(exu_n13033));
INVX1 exu_U33562(.A(exu_n26978), .Y(exu_n13034));
INVX1 exu_U33563(.A(exu_n26983), .Y(exu_n13035));
INVX1 exu_U33564(.A(exu_n26987), .Y(exu_n13036));
INVX1 exu_U33565(.A(exu_n26991), .Y(exu_n13037));
INVX1 exu_U33566(.A(exu_n26995), .Y(exu_n13038));
INVX1 exu_U33567(.A(exu_n26999), .Y(exu_n13039));
INVX1 exu_U33568(.A(exu_n27003), .Y(exu_n13040));
INVX1 exu_U33569(.A(exu_n27007), .Y(exu_n13041));
INVX1 exu_U33570(.A(exu_n27011), .Y(exu_n13042));
INVX1 exu_U33571(.A(exu_n27017), .Y(exu_n13043));
INVX1 exu_U33572(.A(exu_n27023), .Y(exu_n13044));
INVX1 exu_U33573(.A(exu_n27029), .Y(exu_n13045));
INVX1 exu_U33574(.A(exu_n27037), .Y(exu_n13046));
INVX1 exu_U33575(.A(exu_n27040), .Y(exu_n13047));
INVX1 exu_U33576(.A(exu_n27043), .Y(exu_n13048));
INVX1 exu_U33577(.A(exu_n27048), .Y(exu_n13049));
INVX1 exu_U33578(.A(exu_n27054), .Y(exu_n13050));
INVX1 exu_U33579(.A(exu_n27059), .Y(exu_n13051));
INVX1 exu_U33580(.A(exu_n27067), .Y(exu_n13052));
INVX1 exu_U33581(.A(exu_n27072), .Y(exu_n13053));
INVX1 exu_U33582(.A(exu_n27077), .Y(exu_n13054));
INVX1 exu_U33583(.A(exu_n27082), .Y(exu_n13055));
INVX1 exu_U33584(.A(exu_n27087), .Y(exu_n13056));
INVX1 exu_U33585(.A(exu_n27092), .Y(exu_n13057));
INVX1 exu_U33586(.A(exu_n27098), .Y(exu_n13058));
INVX1 exu_U33587(.A(exu_n27104), .Y(exu_n13059));
INVX1 exu_U33588(.A(exu_n27110), .Y(exu_n13060));
INVX1 exu_U33589(.A(exu_n27116), .Y(exu_n13061));
INVX1 exu_U33590(.A(exu_n27122), .Y(exu_n13062));
INVX1 exu_U33591(.A(exu_n27128), .Y(exu_n13063));
INVX1 exu_U33592(.A(exu_n27134), .Y(exu_n13064));
INVX1 exu_U33593(.A(exu_n27140), .Y(exu_n13065));
INVX1 exu_U33594(.A(exu_n27146), .Y(exu_n13066));
INVX1 exu_U33595(.A(exu_n27152), .Y(exu_n13067));
INVX1 exu_U33596(.A(exu_n27158), .Y(exu_n13068));
INVX1 exu_U33597(.A(exu_n27164), .Y(exu_n13069));
INVX1 exu_U33598(.A(exu_n27170), .Y(exu_n13070));
INVX1 exu_U33599(.A(exu_n27176), .Y(exu_n13071));
INVX1 exu_U33600(.A(exu_n27182), .Y(exu_n13072));
INVX1 exu_U33601(.A(exu_n27188), .Y(exu_n13073));
INVX1 exu_U33602(.A(exu_n27194), .Y(exu_n13074));
INVX1 exu_U33603(.A(exu_n27200), .Y(exu_n13075));
INVX1 exu_U33604(.A(exu_n27206), .Y(exu_n13076));
INVX1 exu_U33605(.A(exu_n27212), .Y(exu_n13077));
INVX1 exu_U33606(.A(exu_n27218), .Y(exu_n13078));
INVX1 exu_U33607(.A(exu_n27224), .Y(exu_n13079));
INVX1 exu_U33608(.A(exu_n27230), .Y(exu_n13080));
INVX1 exu_U33609(.A(exu_n27236), .Y(exu_n13081));
INVX1 exu_U33610(.A(exu_n27242), .Y(exu_n13082));
INVX1 exu_U33611(.A(exu_n27248), .Y(exu_n13083));
INVX1 exu_U33612(.A(exu_n27254), .Y(exu_n13084));
INVX1 exu_U33613(.A(exu_n27260), .Y(exu_n13085));
INVX1 exu_U33614(.A(exu_n27266), .Y(exu_n13086));
INVX1 exu_U33615(.A(exu_n27272), .Y(exu_n13087));
INVX1 exu_U33616(.A(exu_n27278), .Y(exu_n13088));
INVX1 exu_U33617(.A(exu_n27284), .Y(exu_n13089));
INVX1 exu_U33618(.A(exu_n27290), .Y(exu_n13090));
INVX1 exu_U33619(.A(exu_n27296), .Y(exu_n13091));
INVX1 exu_U33620(.A(exu_n27302), .Y(exu_n13092));
INVX1 exu_U33621(.A(exu_n27308), .Y(exu_n13093));
INVX1 exu_U33622(.A(exu_n27314), .Y(exu_n13094));
INVX1 exu_U33623(.A(exu_n27320), .Y(exu_n13095));
INVX1 exu_U33624(.A(exu_n27326), .Y(exu_n13096));
INVX1 exu_U33625(.A(exu_n27332), .Y(exu_n13097));
INVX1 exu_U33626(.A(exu_n27338), .Y(exu_n13098));
INVX1 exu_U33627(.A(exu_n27344), .Y(exu_n13099));
INVX1 exu_U33628(.A(exu_n27350), .Y(exu_n13100));
INVX1 exu_U33629(.A(exu_n27356), .Y(exu_n13101));
INVX1 exu_U33630(.A(exu_n27362), .Y(exu_n13102));
INVX1 exu_U33631(.A(exu_n27368), .Y(exu_n13103));
INVX1 exu_U33632(.A(exu_n27374), .Y(exu_n13104));
INVX1 exu_U33633(.A(exu_n27380), .Y(exu_n13105));
INVX1 exu_U33634(.A(exu_n27386), .Y(exu_n13106));
INVX1 exu_U33635(.A(exu_n27392), .Y(exu_n13107));
INVX1 exu_U33636(.A(exu_n27398), .Y(exu_n13108));
INVX1 exu_U33637(.A(exu_n27407), .Y(exu_n13109));
INVX1 exu_U33638(.A(exu_n27412), .Y(exu_n13110));
INVX1 exu_U33639(.A(exu_n27418), .Y(exu_n13111));
INVX1 exu_U33640(.A(exu_n27424), .Y(exu_n13112));
INVX1 exu_U33641(.A(exu_n27430), .Y(exu_n13113));
INVX1 exu_U33642(.A(exu_n27436), .Y(exu_n13114));
INVX1 exu_U33643(.A(exu_n27442), .Y(exu_n13115));
INVX1 exu_U33644(.A(exu_n27448), .Y(exu_n13116));
INVX1 exu_U33645(.A(exu_n27454), .Y(exu_n13117));
INVX1 exu_U33646(.A(exu_n27460), .Y(exu_n13118));
INVX1 exu_U33647(.A(exu_n27466), .Y(exu_n13119));
INVX1 exu_U33648(.A(exu_n27472), .Y(exu_n13120));
INVX1 exu_U33649(.A(exu_n27478), .Y(exu_n13121));
INVX1 exu_U33650(.A(exu_n27484), .Y(exu_n13122));
INVX1 exu_U33651(.A(exu_n27490), .Y(exu_n13123));
INVX1 exu_U33652(.A(exu_n27496), .Y(exu_n13124));
INVX1 exu_U33653(.A(exu_n27502), .Y(exu_n13125));
INVX1 exu_U33654(.A(exu_n27508), .Y(exu_n13126));
INVX1 exu_U33655(.A(exu_n27514), .Y(exu_n13127));
INVX1 exu_U33656(.A(exu_n27520), .Y(exu_n13128));
INVX1 exu_U33657(.A(exu_n27526), .Y(exu_n13129));
INVX1 exu_U33658(.A(exu_n27532), .Y(exu_n13130));
INVX1 exu_U33659(.A(exu_n27538), .Y(exu_n13131));
INVX1 exu_U33660(.A(exu_n27544), .Y(exu_n13132));
INVX1 exu_U33661(.A(exu_n27550), .Y(exu_n13133));
INVX1 exu_U33662(.A(exu_n27556), .Y(exu_n13134));
INVX1 exu_U33663(.A(exu_n27562), .Y(exu_n13135));
INVX1 exu_U33664(.A(exu_n27568), .Y(exu_n13136));
INVX1 exu_U33665(.A(exu_n27574), .Y(exu_n13137));
INVX1 exu_U33666(.A(exu_n27580), .Y(exu_n13138));
INVX1 exu_U33667(.A(exu_n27586), .Y(exu_n13139));
INVX1 exu_U33668(.A(exu_n27592), .Y(exu_n13140));
INVX1 exu_U33669(.A(exu_n27598), .Y(exu_n13141));
INVX1 exu_U33670(.A(exu_n27604), .Y(exu_n13142));
INVX1 exu_U33671(.A(exu_n27610), .Y(exu_n13143));
INVX1 exu_U33672(.A(exu_n27616), .Y(exu_n13144));
INVX1 exu_U33673(.A(exu_n27622), .Y(exu_n13145));
INVX1 exu_U33674(.A(exu_n27628), .Y(exu_n13146));
INVX1 exu_U33675(.A(exu_n27634), .Y(exu_n13147));
INVX1 exu_U33676(.A(exu_n27640), .Y(exu_n13148));
INVX1 exu_U33677(.A(exu_n27646), .Y(exu_n13149));
INVX1 exu_U33678(.A(exu_n27652), .Y(exu_n13150));
INVX1 exu_U33679(.A(exu_n27658), .Y(exu_n13151));
INVX1 exu_U33680(.A(exu_n27664), .Y(exu_n13152));
INVX1 exu_U33681(.A(exu_n27670), .Y(exu_n13153));
INVX1 exu_U33682(.A(exu_n27676), .Y(exu_n13154));
INVX1 exu_U33683(.A(exu_n27682), .Y(exu_n13155));
INVX1 exu_U33684(.A(exu_n27688), .Y(exu_n13156));
INVX1 exu_U33685(.A(exu_n27694), .Y(exu_n13157));
INVX1 exu_U33686(.A(exu_n27700), .Y(exu_n13158));
INVX1 exu_U33687(.A(exu_n27706), .Y(exu_n13159));
INVX1 exu_U33688(.A(exu_n27712), .Y(exu_n13160));
INVX1 exu_U33689(.A(exu_n27718), .Y(exu_n13161));
INVX1 exu_U33690(.A(exu_n27724), .Y(exu_n13162));
INVX1 exu_U33691(.A(exu_n27730), .Y(exu_n13163));
INVX1 exu_U33692(.A(exu_n27736), .Y(exu_n13164));
INVX1 exu_U33693(.A(exu_n27742), .Y(exu_n13165));
INVX1 exu_U33694(.A(exu_n27748), .Y(exu_n13166));
INVX1 exu_U33695(.A(exu_n27758), .Y(exu_n13167));
INVX1 exu_U33696(.A(exu_n27764), .Y(exu_n13168));
INVX1 exu_U33697(.A(exu_n27770), .Y(exu_n13169));
INVX1 exu_U33698(.A(exu_n27776), .Y(exu_n13170));
INVX1 exu_U33699(.A(exu_n27783), .Y(exu_n13171));
INVX1 exu_U33700(.A(exu_n27789), .Y(exu_n13172));
INVX1 exu_U33701(.A(exu_n27795), .Y(exu_n13173));
INVX1 exu_U33702(.A(exu_n27801), .Y(exu_n13174));
INVX1 exu_U33703(.A(exu_n27807), .Y(exu_n13175));
INVX1 exu_U33704(.A(exu_n27813), .Y(exu_n13176));
INVX1 exu_U33705(.A(exu_n27819), .Y(exu_n13177));
INVX1 exu_U33706(.A(exu_n27825), .Y(exu_n13178));
INVX1 exu_U33707(.A(exu_n27831), .Y(exu_n13179));
INVX1 exu_U33708(.A(exu_n27837), .Y(exu_n13180));
INVX1 exu_U33709(.A(exu_n27844), .Y(exu_n13181));
INVX1 exu_U33710(.A(exu_n27850), .Y(exu_n13182));
INVX1 exu_U33711(.A(exu_n27992), .Y(exu_n13183));
INVX1 exu_U33712(.A(exu_n27998), .Y(exu_n13184));
INVX1 exu_U33713(.A(exu_n28004), .Y(exu_n13185));
INVX1 exu_U33714(.A(exu_n28010), .Y(exu_n13186));
INVX1 exu_U33715(.A(exu_n28019), .Y(exu_n13187));
INVX1 exu_U33716(.A(exu_n28025), .Y(exu_n13188));
INVX1 exu_U33717(.A(exu_n28031), .Y(exu_n13189));
INVX1 exu_U33718(.A(exu_n28037), .Y(exu_n13190));
INVX1 exu_U33719(.A(exu_n28043), .Y(exu_n13191));
INVX1 exu_U33720(.A(exu_n28049), .Y(exu_n13192));
INVX1 exu_U33721(.A(exu_n28055), .Y(exu_n13193));
INVX1 exu_U33722(.A(exu_n28061), .Y(exu_n13194));
INVX1 exu_U33723(.A(exu_n28067), .Y(exu_n13195));
INVX1 exu_U33724(.A(exu_n28073), .Y(exu_n13196));
INVX1 exu_U33725(.A(exu_n28082), .Y(exu_n13197));
INVX1 exu_U33726(.A(exu_n28088), .Y(exu_n13198));
INVX1 exu_U33727(.A(exu_n28094), .Y(exu_n13199));
INVX1 exu_U33728(.A(exu_n28100), .Y(exu_n13200));
INVX1 exu_U33729(.A(exu_n28106), .Y(exu_n13201));
INVX1 exu_U33730(.A(exu_n28112), .Y(exu_n13202));
INVX1 exu_U33731(.A(exu_n28118), .Y(exu_n13203));
INVX1 exu_U33732(.A(exu_n28124), .Y(exu_n13204));
INVX1 exu_U33733(.A(exu_n28130), .Y(exu_n13205));
INVX1 exu_U33734(.A(exu_n28136), .Y(exu_n13206));
INVX1 exu_U33735(.A(exu_n28143), .Y(exu_n13207));
INVX1 exu_U33736(.A(exu_n28149), .Y(exu_n13208));
INVX1 exu_U33737(.A(exu_n28155), .Y(exu_n13209));
INVX1 exu_U33738(.A(exu_n28161), .Y(exu_n13210));
INVX1 exu_U33739(.A(exu_n28167), .Y(exu_n13211));
INVX1 exu_U33740(.A(exu_n28173), .Y(exu_n13212));
INVX1 exu_U33741(.A(exu_n28179), .Y(exu_n13213));
INVX1 exu_U33742(.A(exu_n28185), .Y(exu_n13214));
INVX1 exu_U33743(.A(exu_n28191), .Y(exu_n13215));
INVX1 exu_U33744(.A(exu_n28197), .Y(exu_n13216));
INVX1 exu_U33745(.A(exu_n28204), .Y(exu_n13217));
INVX1 exu_U33746(.A(exu_n28210), .Y(exu_n13218));
INVX1 exu_U33747(.A(exu_n28216), .Y(exu_n13219));
INVX1 exu_U33748(.A(exu_n28222), .Y(exu_n13220));
INVX1 exu_U33749(.A(exu_n28228), .Y(exu_n13221));
INVX1 exu_U33750(.A(exu_n28234), .Y(exu_n13222));
INVX1 exu_U33751(.A(exu_n28240), .Y(exu_n13223));
INVX1 exu_U33752(.A(exu_n28246), .Y(exu_n13224));
INVX1 exu_U33753(.A(exu_n28252), .Y(exu_n13225));
INVX1 exu_U33754(.A(exu_n28258), .Y(exu_n13226));
INVX1 exu_U33755(.A(exu_n28265), .Y(exu_n13227));
INVX1 exu_U33756(.A(exu_n28271), .Y(exu_n13228));
INVX1 exu_U33757(.A(exu_n28277), .Y(exu_n13229));
INVX1 exu_U33758(.A(exu_n28283), .Y(exu_n13230));
INVX1 exu_U33759(.A(exu_n28289), .Y(exu_n13231));
INVX1 exu_U33760(.A(exu_n28295), .Y(exu_n13232));
INVX1 exu_U33761(.A(exu_n28301), .Y(exu_n13233));
INVX1 exu_U33762(.A(exu_n28307), .Y(exu_n13234));
INVX1 exu_U33763(.A(exu_n28322), .Y(exu_n13235));
INVX1 exu_U33764(.A(exu_n28328), .Y(exu_n13236));
INVX1 exu_U33765(.A(exu_n28334), .Y(exu_n13237));
INVX1 exu_U33766(.A(exu_n28340), .Y(exu_n13238));
INVX1 exu_U33767(.A(exu_n28346), .Y(exu_n13239));
INVX1 exu_U33768(.A(exu_n28352), .Y(exu_n13240));
INVX1 exu_U33769(.A(exu_n28358), .Y(exu_n13241));
INVX1 exu_U33770(.A(exu_n28364), .Y(exu_n13242));
INVX1 exu_U33771(.A(exu_n28370), .Y(exu_n13243));
INVX1 exu_U33772(.A(exu_n28376), .Y(exu_n13244));
INVX1 exu_U33773(.A(exu_n28382), .Y(exu_n13245));
INVX1 exu_U33774(.A(exu_n28388), .Y(exu_n13246));
INVX1 exu_U33775(.A(exu_n28394), .Y(exu_n13247));
INVX1 exu_U33776(.A(exu_n28400), .Y(exu_n13248));
INVX1 exu_U33777(.A(exu_n28406), .Y(exu_n13249));
INVX1 exu_U33778(.A(exu_n28412), .Y(exu_n13250));
INVX1 exu_U33779(.A(exu_n28418), .Y(exu_n13251));
INVX1 exu_U33780(.A(exu_n28424), .Y(exu_n13252));
INVX1 exu_U33781(.A(exu_n28430), .Y(exu_n13253));
INVX1 exu_U33782(.A(exu_n28436), .Y(exu_n13254));
INVX1 exu_U33783(.A(exu_n28442), .Y(exu_n13255));
INVX1 exu_U33784(.A(exu_n28448), .Y(exu_n13256));
INVX1 exu_U33785(.A(exu_n28454), .Y(exu_n13257));
INVX1 exu_U33786(.A(exu_n28460), .Y(exu_n13258));
INVX1 exu_U33787(.A(exu_n28466), .Y(exu_n13259));
INVX1 exu_U33788(.A(exu_n28472), .Y(exu_n13260));
INVX1 exu_U33789(.A(exu_n28478), .Y(exu_n13261));
INVX1 exu_U33790(.A(exu_n28484), .Y(exu_n13262));
INVX1 exu_U33791(.A(exu_n28490), .Y(exu_n13263));
INVX1 exu_U33792(.A(exu_n28496), .Y(exu_n13264));
INVX1 exu_U33793(.A(exu_n28502), .Y(exu_n13265));
INVX1 exu_U33794(.A(exu_n28508), .Y(exu_n13266));
INVX1 exu_U33795(.A(exu_n28514), .Y(exu_n13267));
INVX1 exu_U33796(.A(exu_n28520), .Y(exu_n13268));
INVX1 exu_U33797(.A(exu_n28526), .Y(exu_n13269));
INVX1 exu_U33798(.A(exu_n28532), .Y(exu_n13270));
INVX1 exu_U33799(.A(exu_n28538), .Y(exu_n13271));
INVX1 exu_U33800(.A(exu_n28544), .Y(exu_n13272));
INVX1 exu_U33801(.A(exu_n28550), .Y(exu_n13273));
INVX1 exu_U33802(.A(exu_n28556), .Y(exu_n13274));
INVX1 exu_U33803(.A(exu_n28562), .Y(exu_n13275));
INVX1 exu_U33804(.A(exu_n28572), .Y(exu_n13276));
INVX1 exu_U33805(.A(exu_n28578), .Y(exu_n13277));
INVX1 exu_U33806(.A(exu_n28584), .Y(exu_n13278));
INVX1 exu_U33807(.A(exu_n28590), .Y(exu_n13279));
INVX1 exu_U33808(.A(exu_n28596), .Y(exu_n13280));
INVX1 exu_U33809(.A(exu_n28602), .Y(exu_n13281));
INVX1 exu_U33810(.A(exu_n28608), .Y(exu_n13282));
INVX1 exu_U33811(.A(exu_n28614), .Y(exu_n13283));
INVX1 exu_U33812(.A(exu_n28620), .Y(exu_n13284));
INVX1 exu_U33813(.A(exu_n28626), .Y(exu_n13285));
INVX1 exu_U33814(.A(exu_n28635), .Y(exu_n13286));
INVX1 exu_U33815(.A(exu_n28641), .Y(exu_n13287));
INVX1 exu_U33816(.A(exu_n28647), .Y(exu_n13288));
INVX1 exu_U33817(.A(exu_n28653), .Y(exu_n13289));
INVX1 exu_U33818(.A(exu_n28659), .Y(exu_n13290));
INVX1 exu_U33819(.A(exu_n28665), .Y(exu_n13291));
INVX1 exu_U33820(.A(exu_n28671), .Y(exu_n13292));
INVX1 exu_U33821(.A(exu_n28677), .Y(exu_n13293));
INVX1 exu_U33822(.A(exu_n28683), .Y(exu_n13294));
INVX1 exu_U33823(.A(exu_n28689), .Y(exu_n13295));
INVX1 exu_U33824(.A(exu_n28696), .Y(exu_n13296));
INVX1 exu_U33825(.A(exu_n28702), .Y(exu_n13297));
INVX1 exu_U33826(.A(exu_n28708), .Y(exu_n13298));
INVX1 exu_U33827(.A(exu_n28714), .Y(exu_n13299));
INVX1 exu_U33828(.A(exu_n28724), .Y(exu_n13300));
INVX1 exu_U33829(.A(exu_n28740), .Y(exu_n13301));
INVX1 exu_U33830(.A(exu_n28756), .Y(exu_n13302));
INVX1 exu_U33831(.A(exu_n28770), .Y(exu_n13303));
INVX1 exu_U33832(.A(exu_n28773), .Y(exu_n13304));
INVX1 exu_U33833(.A(exu_n28779), .Y(exu_n13305));
INVX1 exu_U33834(.A(exu_n28785), .Y(exu_n13306));
INVX1 exu_U33835(.A(exu_n28791), .Y(exu_n13307));
INVX1 exu_U33836(.A(exu_n28797), .Y(exu_n13308));
INVX1 exu_U33837(.A(exu_n28803), .Y(exu_n13309));
INVX1 exu_U33838(.A(exu_n28809), .Y(exu_n13310));
INVX1 exu_U33839(.A(exu_n28815), .Y(exu_n13311));
INVX1 exu_U33840(.A(exu_n28821), .Y(exu_n13312));
INVX1 exu_U33841(.A(exu_n28827), .Y(exu_n13313));
INVX1 exu_U33842(.A(exu_n28833), .Y(exu_n13314));
INVX1 exu_U33843(.A(exu_n28839), .Y(exu_n13315));
INVX1 exu_U33844(.A(exu_n28845), .Y(exu_n13316));
INVX1 exu_U33845(.A(exu_n28851), .Y(exu_n13317));
INVX1 exu_U33846(.A(exu_n28857), .Y(exu_n13318));
INVX1 exu_U33847(.A(exu_n28863), .Y(exu_n13319));
INVX1 exu_U33848(.A(exu_n28869), .Y(exu_n13320));
INVX1 exu_U33849(.A(exu_n28875), .Y(exu_n13321));
INVX1 exu_U33850(.A(exu_n28881), .Y(exu_n13322));
INVX1 exu_U33851(.A(exu_n28887), .Y(exu_n13323));
INVX1 exu_U33852(.A(exu_n28893), .Y(exu_n13324));
INVX1 exu_U33853(.A(exu_n28899), .Y(exu_n13325));
INVX1 exu_U33854(.A(exu_n28905), .Y(exu_n13326));
INVX1 exu_U33855(.A(exu_n28911), .Y(exu_n13327));
INVX1 exu_U33856(.A(exu_n28917), .Y(exu_n13328));
INVX1 exu_U33857(.A(exu_n28923), .Y(exu_n13329));
INVX1 exu_U33858(.A(exu_n28929), .Y(exu_n13330));
INVX1 exu_U33859(.A(exu_n28935), .Y(exu_n13331));
INVX1 exu_U33860(.A(exu_n28941), .Y(exu_n13332));
INVX1 exu_U33861(.A(exu_n28947), .Y(exu_n13333));
INVX1 exu_U33862(.A(exu_n28953), .Y(exu_n13334));
INVX1 exu_U33863(.A(exu_n28959), .Y(exu_n13335));
INVX1 exu_U33864(.A(exu_n28965), .Y(exu_n13336));
INVX1 exu_U33865(.A(exu_n28971), .Y(exu_n13337));
INVX1 exu_U33866(.A(exu_n28977), .Y(exu_n13338));
INVX1 exu_U33867(.A(exu_n28983), .Y(exu_n13339));
INVX1 exu_U33868(.A(exu_n28989), .Y(exu_n13340));
INVX1 exu_U33869(.A(exu_n28995), .Y(exu_n13341));
INVX1 exu_U33870(.A(exu_n29001), .Y(exu_n13342));
INVX1 exu_U33871(.A(exu_n29007), .Y(exu_n13343));
INVX1 exu_U33872(.A(exu_n29013), .Y(exu_n13344));
INVX1 exu_U33873(.A(exu_n29019), .Y(exu_n13345));
INVX1 exu_U33874(.A(exu_n29025), .Y(exu_n13346));
INVX1 exu_U33875(.A(exu_n29031), .Y(exu_n13347));
INVX1 exu_U33876(.A(exu_n29037), .Y(exu_n13348));
INVX1 exu_U33877(.A(exu_n29043), .Y(exu_n13349));
INVX1 exu_U33878(.A(exu_n29049), .Y(exu_n13350));
INVX1 exu_U33879(.A(exu_n29055), .Y(exu_n13351));
INVX1 exu_U33880(.A(exu_n29061), .Y(exu_n13352));
INVX1 exu_U33881(.A(exu_n29067), .Y(exu_n13353));
INVX1 exu_U33882(.A(exu_n29073), .Y(exu_n13354));
INVX1 exu_U33883(.A(exu_n29079), .Y(exu_n13355));
INVX1 exu_U33884(.A(exu_n29085), .Y(exu_n13356));
INVX1 exu_U33885(.A(exu_n29091), .Y(exu_n13357));
INVX1 exu_U33886(.A(exu_n29097), .Y(exu_n13358));
INVX1 exu_U33887(.A(exu_n29103), .Y(exu_n13359));
INVX1 exu_U33888(.A(exu_n29109), .Y(exu_n13360));
INVX1 exu_U33889(.A(exu_n29115), .Y(exu_n13361));
INVX1 exu_U33890(.A(exu_n29121), .Y(exu_n13362));
INVX1 exu_U33891(.A(exu_n29127), .Y(exu_n13363));
INVX1 exu_U33892(.A(exu_n29133), .Y(exu_n13364));
INVX1 exu_U33893(.A(exu_n29139), .Y(exu_n13365));
INVX1 exu_U33894(.A(exu_n29145), .Y(exu_n13366));
INVX1 exu_U33895(.A(exu_n29151), .Y(exu_n13367));
INVX1 exu_U33896(.A(exu_n29157), .Y(exu_n13368));
INVX1 exu_U33897(.A(exu_n29163), .Y(exu_n13369));
INVX1 exu_U33898(.A(exu_n29169), .Y(exu_n13370));
INVX1 exu_U33899(.A(exu_n29175), .Y(exu_n13371));
INVX1 exu_U33900(.A(exu_n29181), .Y(exu_n13372));
INVX1 exu_U33901(.A(exu_n29187), .Y(exu_n13373));
INVX1 exu_U33902(.A(exu_n29193), .Y(exu_n13374));
INVX1 exu_U33903(.A(exu_n29199), .Y(exu_n13375));
INVX1 exu_U33904(.A(exu_n29205), .Y(exu_n13376));
INVX1 exu_U33905(.A(exu_n29211), .Y(exu_n13377));
INVX1 exu_U33906(.A(exu_n29217), .Y(exu_n13378));
INVX1 exu_U33907(.A(exu_n29223), .Y(exu_n13379));
INVX1 exu_U33908(.A(exu_n29229), .Y(exu_n13380));
INVX1 exu_U33909(.A(exu_n29235), .Y(exu_n13381));
INVX1 exu_U33910(.A(exu_n29241), .Y(exu_n13382));
INVX1 exu_U33911(.A(exu_n29247), .Y(exu_n13383));
INVX1 exu_U33912(.A(exu_n29253), .Y(exu_n13384));
INVX1 exu_U33913(.A(exu_n29259), .Y(exu_n13385));
INVX1 exu_U33914(.A(exu_n29265), .Y(exu_n13386));
INVX1 exu_U33915(.A(exu_n29271), .Y(exu_n13387));
INVX1 exu_U33916(.A(exu_n29277), .Y(exu_n13388));
INVX1 exu_U33917(.A(exu_n29283), .Y(exu_n13389));
INVX1 exu_U33918(.A(exu_n29289), .Y(exu_n13390));
INVX1 exu_U33919(.A(exu_n29295), .Y(exu_n13391));
INVX1 exu_U33920(.A(exu_n31457), .Y(exu_n13392));
INVX1 exu_U33921(.A(exu_n31463), .Y(exu_n13393));
INVX1 exu_U33922(.A(exu_n31616), .Y(exu_n13394));
INVX1 exu_U33923(.A(exu_n31646), .Y(exu_n13395));
INVX1 exu_U33924(.A(exu_n31676), .Y(exu_n13396));
INVX1 exu_U33925(.A(rml_cwp_cwp_output_mux_n1), .Y(exu_n13397));
INVX1 exu_U33926(.A(rml_cwp_cwp_output_mux_n7), .Y(exu_n13398));
INVX1 exu_U33927(.A(rml_cwp_cwp_output_mux_n13), .Y(exu_n13399));
INVX1 exu_U33928(.A(rml_cwp_cwp_output_mux_n19), .Y(exu_n13400));
INVX1 exu_U33929(.A(rml_cwp_cwp_output_mux_n25), .Y(exu_n13401));
INVX1 exu_U33930(.A(rml_cwp_cwp_output_mux_n31), .Y(exu_n13402));
INVX1 exu_U33931(.A(rml_cwp_cwp_output_mux_n37), .Y(exu_n13403));
INVX1 exu_U33932(.A(rml_cwp_cwp_output_mux_n43), .Y(exu_n13404));
INVX1 exu_U33933(.A(rml_cwp_cwp_output_mux_n49), .Y(exu_n13405));
INVX1 exu_U33934(.A(rml_cwp_cwp_output_mux_n55), .Y(exu_n13406));
INVX1 exu_U33935(.A(rml_cwp_cwp_output_mux_n61), .Y(exu_n13407));
INVX1 exu_U33936(.A(rml_cwp_cwp_output_mux_n67), .Y(exu_n13408));
INVX1 exu_U33937(.A(rml_cwp_cwp_output_mux_n73), .Y(exu_n13409));
INVX1 exu_U33938(.A(rml_cwp_cwp_output_mux_n79), .Y(exu_n13410));
INVX1 exu_U33939(.A(rml_cwp_cwp_output_mux_n85), .Y(exu_n13411));
INVX1 exu_U33940(.A(ecl_writeback_rdpr_mux1_n1), .Y(exu_n13412));
INVX1 exu_U33941(.A(ecl_writeback_rdpr_mux1_n7), .Y(exu_n13413));
INVX1 exu_U33942(.A(ecl_writeback_rdpr_mux1_n13), .Y(exu_n13414));
INVX1 exu_U33943(.A(ecl_writeback_rd_g_mux_n1), .Y(exu_n13415));
INVX1 exu_U33944(.A(ecl_writeback_rd_g_mux_n7), .Y(exu_n13416));
INVX1 exu_U33945(.A(ecl_writeback_rd_g_mux_n13), .Y(exu_n13417));
INVX1 exu_U33946(.A(ecl_writeback_rd_g_mux_n19), .Y(exu_n13418));
INVX1 exu_U33947(.A(ecl_writeback_rd_g_mux_n25), .Y(exu_n13419));
INVX1 exu_U33948(.A(ecl_ccr_mux_ccr_out_n1), .Y(exu_n13420));
INVX1 exu_U33949(.A(ecl_ccr_mux_ccr_out_n7), .Y(exu_n13421));
INVX1 exu_U33950(.A(ecl_ccr_mux_ccr_out_n13), .Y(exu_n13422));
INVX1 exu_U33951(.A(ecl_ccr_mux_ccr_out_n19), .Y(exu_n13423));
INVX1 exu_U33952(.A(ecl_ccr_mux_ccr_out_n25), .Y(exu_n13424));
INVX1 exu_U33953(.A(ecl_ccr_mux_ccr_out_n31), .Y(exu_n13425));
INVX1 exu_U33954(.A(ecl_ccr_mux_ccr_out_n37), .Y(exu_n13426));
INVX1 exu_U33955(.A(ecl_ccr_mux_ccr_out_n43), .Y(exu_n13427));
INVX1 exu_U33956(.A(rml_mux_agp_out1_n1), .Y(exu_n13428));
INVX1 exu_U33957(.A(rml_mux_agp_out1_n7), .Y(exu_n13429));
INVX1 exu_U33958(.A(div_low32or_n1), .Y(exu_n13430));
AND2X1 exu_U33959(.A(exu_n15425), .B(exu_n16371), .Y(ecl_mdqctl_n18));
INVX1 exu_U33960(.A(ecl_mdqctl_n18), .Y(exu_n13431));
AND2X1 exu_U33961(.A(exu_n16504), .B(exu_n16505), .Y(ecl_divcntl_n48));
INVX1 exu_U33962(.A(ecl_divcntl_n48), .Y(exu_n13432));
OR2X1 exu_U33963(.A(exu_n16508), .B(ecl_divcntl_n59), .Y(ecl_divcntl_n57));
INVX1 exu_U33964(.A(ecl_divcntl_n57), .Y(exu_n13433));
AND2X1 exu_U33965(.A(ecl_divcntl_n89), .B(ecl_divcntl_cntr[2]), .Y(ecl_divcntl_n86));
INVX1 exu_U33966(.A(ecl_divcntl_n86), .Y(exu_n13434));
AND2X1 exu_U33967(.A(exu_n15208), .B(exu_n16270), .Y(ecl_byplog_rs2_n27));
INVX1 exu_U33968(.A(ecl_byplog_rs2_n27), .Y(exu_n13435));
INVX1 exu_U33969(.A(ecl_byplog_rs2_n42), .Y(exu_n13436));
INVX1 exu_U33970(.A(ecl_byplog_rs2_n44), .Y(exu_n13437));
AND2X1 exu_U33971(.A(exu_n15207), .B(exu_n16270), .Y(ecl_byplog_rs1_n36));
INVX1 exu_U33972(.A(ecl_byplog_rs1_n36), .Y(exu_n13438));
AND2X1 exu_U33973(.A(exu_n15437), .B(exu_n15203), .Y(ecl_byplog_rs1_n33));
INVX1 exu_U33974(.A(ecl_byplog_rs1_n33), .Y(exu_n13439));
INVX1 exu_U33975(.A(ecl_byplog_rs1_n47), .Y(exu_n13440));
INVX1 exu_U33976(.A(ecl_byplog_rs1_n49), .Y(exu_n13441));
OR2X1 exu_U33977(.A(exu_n16611), .B(ecl_writeback_n68), .Y(ecl_writeback_n67));
INVX1 exu_U33978(.A(ecl_writeback_n67), .Y(exu_n13442));
OR2X1 exu_U33979(.A(exu_n16553), .B(ecl_writeback_n133), .Y(ecl_rml_otherwin_wen_w));
INVX1 exu_U33980(.A(ecl_rml_otherwin_wen_w), .Y(exu_n13443));
AND2X1 exu_U33981(.A(ecl_writeback_sraddr_e[0]), .B(exu_ffu_wsr_inst_e), .Y(ecl_writeback_n136));
INVX1 exu_U33982(.A(ecl_writeback_n136), .Y(exu_n13444));
INVX1 exu_U33983(.A(ecl_writeback_n134), .Y(exu_n13445));
OR2X1 exu_U33984(.A(ecl_writeback_n131), .B(exu_n14972), .Y(ecl_rml_cleanwin_wen_w));
INVX1 exu_U33985(.A(ecl_rml_cleanwin_wen_w), .Y(exu_n13446));
OR2X1 exu_U33986(.A(ecl_writeback_sraddr_w[0]), .B(ecl_writeback_n142), .Y(ecl_rml_cansave_wen_w));
INVX1 exu_U33987(.A(ecl_rml_cansave_wen_w), .Y(exu_n13447));
OR2X1 exu_U33988(.A(exu_n16553), .B(ecl_writeback_n142), .Y(ecl_rml_canrestore_wen_w));
INVX1 exu_U33989(.A(ecl_rml_canrestore_wen_w), .Y(exu_n13448));
AND2X1 exu_U33990(.A(ecl_mdqctl_wb_multhr_g[0]), .B(exu_n15741), .Y(ecl_writeback_n184));
INVX1 exu_U33991(.A(ecl_writeback_n184), .Y(exu_n13449));
AND2X1 exu_U33992(.A(exu_n15743), .B(exu_n16509), .Y(ecl_writeback_n186));
INVX1 exu_U33993(.A(ecl_writeback_n186), .Y(exu_n13450));
AND2X1 exu_U33994(.A(exu_n15744), .B(exu_n16510), .Y(ecl_writeback_n187));
INVX1 exu_U33995(.A(ecl_writeback_n187), .Y(exu_n13451));
AND2X1 exu_U33996(.A(exu_n16509), .B(exu_n16510), .Y(ecl_writeback_n189));
INVX1 exu_U33997(.A(ecl_writeback_n189), .Y(exu_n13452));
INVX1 exu_U33998(.A(ecl_yreg0_mux_n1), .Y(exu_n13453));
AND2X1 exu_U33999(.A(ecc_err_m[4]), .B(ecc_err_m[5]), .Y(ecc_decode_n25));
INVX1 exu_U34000(.A(ecc_decode_n25), .Y(exu_n13454));
INVX1 exu_U34001(.A(bypass_mux_rs3h_data_1_n1), .Y(exu_n13455));
INVX1 exu_U34002(.A(bypass_mux_rs3h_data_1_n7), .Y(exu_n13456));
INVX1 exu_U34003(.A(bypass_mux_rs3h_data_1_n13), .Y(exu_n13457));
INVX1 exu_U34004(.A(bypass_mux_rs3h_data_1_n19), .Y(exu_n13458));
INVX1 exu_U34005(.A(bypass_mux_rs3h_data_1_n25), .Y(exu_n13459));
INVX1 exu_U34006(.A(bypass_mux_rs3h_data_1_n31), .Y(exu_n13460));
INVX1 exu_U34007(.A(bypass_mux_rs3h_data_1_n37), .Y(exu_n13461));
INVX1 exu_U34008(.A(bypass_mux_rs3h_data_1_n43), .Y(exu_n13462));
INVX1 exu_U34009(.A(bypass_mux_rs3h_data_1_n49), .Y(exu_n13463));
INVX1 exu_U34010(.A(bypass_mux_rs3h_data_1_n55), .Y(exu_n13464));
INVX1 exu_U34011(.A(bypass_mux_rs3h_data_1_n61), .Y(exu_n13465));
INVX1 exu_U34012(.A(bypass_mux_rs3h_data_1_n67), .Y(exu_n13466));
INVX1 exu_U34013(.A(bypass_mux_rs3h_data_1_n73), .Y(exu_n13467));
INVX1 exu_U34014(.A(bypass_mux_rs3h_data_1_n79), .Y(exu_n13468));
INVX1 exu_U34015(.A(bypass_mux_rs3h_data_1_n85), .Y(exu_n13469));
INVX1 exu_U34016(.A(bypass_mux_rs3h_data_1_n91), .Y(exu_n13470));
INVX1 exu_U34017(.A(bypass_mux_rs3h_data_1_n97), .Y(exu_n13471));
INVX1 exu_U34018(.A(bypass_mux_rs3h_data_1_n103), .Y(exu_n13472));
INVX1 exu_U34019(.A(bypass_mux_rs3h_data_1_n109), .Y(exu_n13473));
INVX1 exu_U34020(.A(bypass_mux_rs3h_data_1_n115), .Y(exu_n13474));
INVX1 exu_U34021(.A(bypass_mux_rs3h_data_1_n121), .Y(exu_n13475));
INVX1 exu_U34022(.A(bypass_mux_rs3h_data_1_n127), .Y(exu_n13476));
INVX1 exu_U34023(.A(bypass_mux_rs3h_data_1_n133), .Y(exu_n13477));
INVX1 exu_U34024(.A(bypass_mux_rs3h_data_1_n139), .Y(exu_n13478));
INVX1 exu_U34025(.A(bypass_mux_rs3h_data_1_n145), .Y(exu_n13479));
INVX1 exu_U34026(.A(bypass_mux_rs3h_data_1_n151), .Y(exu_n13480));
INVX1 exu_U34027(.A(bypass_mux_rs3h_data_1_n157), .Y(exu_n13481));
INVX1 exu_U34028(.A(bypass_mux_rs3h_data_1_n163), .Y(exu_n13482));
INVX1 exu_U34029(.A(bypass_mux_rs3h_data_1_n169), .Y(exu_n13483));
INVX1 exu_U34030(.A(bypass_mux_rs3h_data_1_n175), .Y(exu_n13484));
INVX1 exu_U34031(.A(bypass_mux_rs3h_data_1_n181), .Y(exu_n13485));
INVX1 exu_U34032(.A(bypass_mux_rs3h_data_1_n187), .Y(exu_n13486));
INVX1 exu_U34033(.A(bypass_ifu_exu_sr_mux_n13), .Y(exu_n13487));
INVX1 exu_U34034(.A(bypass_ifu_exu_sr_mux_n19), .Y(exu_n13488));
INVX1 exu_U34035(.A(bypass_ifu_exu_sr_mux_n49), .Y(exu_n13489));
INVX1 exu_U34036(.A(bypass_ifu_exu_sr_mux_n115), .Y(exu_n13490));
INVX1 exu_U34037(.A(bypass_ifu_exu_sr_mux_n181), .Y(exu_n13491));
INVX1 exu_U34038(.A(bypass_ifu_exu_sr_mux_n247), .Y(exu_n13492));
INVX1 exu_U34039(.A(bypass_ifu_exu_sr_mux_n313), .Y(exu_n13493));
INVX1 exu_U34040(.A(bypass_ifu_exu_sr_mux_n379), .Y(exu_n13494));
INVX1 exu_U34041(.A(rml_n62), .Y(exu_n13495));
INVX1 exu_U34042(.A(rml_n71), .Y(exu_n13496));
INVX1 exu_U34043(.A(div_n37), .Y(exu_n13497));
INVX1 exu_U34044(.A(div_n67), .Y(exu_n13498));
INVX1 exu_U34045(.A(alu_n69), .Y(exu_n13499));
INVX1 exu_U34046(.A(ecl_n82), .Y(exu_n13500));
AND2X1 exu_U34047(.A(exu_n16381), .B(rml_ecl_fill_e), .Y(ecl_n110));
INVX1 exu_U34048(.A(ecl_n110), .Y(exu_n13501));
AND2X1 exu_U34049(.A(exu_n16652), .B(exu_n16651), .Y(exu_n16653));
INVX1 exu_U34050(.A(exu_n16653), .Y(exu_n13502));
AND2X1 exu_U34051(.A(exu_n16708), .B(exu_n16707), .Y(exu_n16709));
INVX1 exu_U34052(.A(exu_n16709), .Y(exu_n13503));
AND2X1 exu_U34053(.A(exu_n17386), .B(exu_n17385), .Y(exu_n17387));
INVX1 exu_U34054(.A(exu_n17387), .Y(exu_n13504));
AND2X1 exu_U34055(.A(exu_n17428), .B(exu_n17427), .Y(exu_n17429));
INVX1 exu_U34056(.A(exu_n17429), .Y(exu_n13505));
INVX1 exu_U34057(.A(exu_n17729), .Y(exu_n13506));
INVX1 exu_U34058(.A(exu_n17735), .Y(exu_n13507));
INVX1 exu_U34059(.A(exu_n17741), .Y(exu_n13508));
INVX1 exu_U34060(.A(exu_n17747), .Y(exu_n13509));
INVX1 exu_U34061(.A(exu_n17753), .Y(exu_n13510));
INVX1 exu_U34062(.A(exu_n17759), .Y(exu_n13511));
INVX1 exu_U34063(.A(exu_n17765), .Y(exu_n13512));
INVX1 exu_U34064(.A(exu_n17771), .Y(exu_n13513));
INVX1 exu_U34065(.A(exu_n17777), .Y(exu_n13514));
INVX1 exu_U34066(.A(exu_n17783), .Y(exu_n13515));
INVX1 exu_U34067(.A(exu_n17789), .Y(exu_n13516));
INVX1 exu_U34068(.A(exu_n17795), .Y(exu_n13517));
INVX1 exu_U34069(.A(exu_n17801), .Y(exu_n13518));
INVX1 exu_U34070(.A(exu_n17807), .Y(exu_n13519));
INVX1 exu_U34071(.A(exu_n17813), .Y(exu_n13520));
INVX1 exu_U34072(.A(exu_n17819), .Y(exu_n13521));
INVX1 exu_U34073(.A(exu_n17825), .Y(exu_n13522));
INVX1 exu_U34074(.A(exu_n17831), .Y(exu_n13523));
INVX1 exu_U34075(.A(exu_n17837), .Y(exu_n13524));
INVX1 exu_U34076(.A(exu_n17843), .Y(exu_n13525));
INVX1 exu_U34077(.A(exu_n17849), .Y(exu_n13526));
INVX1 exu_U34078(.A(exu_n17855), .Y(exu_n13527));
INVX1 exu_U34079(.A(exu_n17861), .Y(exu_n13528));
INVX1 exu_U34080(.A(exu_n17867), .Y(exu_n13529));
INVX1 exu_U34081(.A(exu_n17873), .Y(exu_n13530));
INVX1 exu_U34082(.A(exu_n17879), .Y(exu_n13531));
INVX1 exu_U34083(.A(exu_n17885), .Y(exu_n13532));
INVX1 exu_U34084(.A(exu_n17891), .Y(exu_n13533));
INVX1 exu_U34085(.A(exu_n17897), .Y(exu_n13534));
INVX1 exu_U34086(.A(exu_n17903), .Y(exu_n13535));
INVX1 exu_U34087(.A(exu_n17909), .Y(exu_n13536));
INVX1 exu_U34088(.A(exu_n17915), .Y(exu_n13537));
INVX1 exu_U34089(.A(exu_n17921), .Y(exu_n13538));
INVX1 exu_U34090(.A(exu_n17927), .Y(exu_n13539));
INVX1 exu_U34091(.A(exu_n17933), .Y(exu_n13540));
INVX1 exu_U34092(.A(exu_n17939), .Y(exu_n13541));
INVX1 exu_U34093(.A(exu_n17945), .Y(exu_n13542));
INVX1 exu_U34094(.A(exu_n17951), .Y(exu_n13543));
INVX1 exu_U34095(.A(exu_n17957), .Y(exu_n13544));
INVX1 exu_U34096(.A(exu_n17963), .Y(exu_n13545));
INVX1 exu_U34097(.A(exu_n17969), .Y(exu_n13546));
INVX1 exu_U34098(.A(exu_n17975), .Y(exu_n13547));
INVX1 exu_U34099(.A(exu_n17982), .Y(exu_n13548));
INVX1 exu_U34100(.A(exu_n17988), .Y(exu_n13549));
INVX1 exu_U34101(.A(exu_n17994), .Y(exu_n13550));
INVX1 exu_U34102(.A(exu_n18000), .Y(exu_n13551));
INVX1 exu_U34103(.A(exu_n18006), .Y(exu_n13552));
INVX1 exu_U34104(.A(exu_n18020), .Y(exu_n13553));
INVX1 exu_U34105(.A(exu_n18026), .Y(exu_n13554));
INVX1 exu_U34106(.A(exu_n18032), .Y(exu_n13555));
AND2X1 exu_U34107(.A(exu_n19190), .B(exu_n19199), .Y(exu_n19193));
INVX1 exu_U34108(.A(exu_n19193), .Y(exu_n13556));
AND2X1 exu_U34109(.A(exu_n19226), .B(exu_n19235), .Y(exu_n19229));
INVX1 exu_U34110(.A(exu_n19229), .Y(exu_n13557));
INVX1 exu_U34111(.A(exu_n20477), .Y(exu_n13558));
INVX1 exu_U34112(.A(exu_n20483), .Y(exu_n13559));
INVX1 exu_U34113(.A(exu_n20489), .Y(exu_n13560));
INVX1 exu_U34114(.A(exu_n20495), .Y(exu_n13561));
INVX1 exu_U34115(.A(exu_n20501), .Y(exu_n13562));
INVX1 exu_U34116(.A(exu_n20507), .Y(exu_n13563));
INVX1 exu_U34117(.A(exu_n20513), .Y(exu_n13564));
INVX1 exu_U34118(.A(exu_n20519), .Y(exu_n13565));
INVX1 exu_U34119(.A(exu_n20525), .Y(exu_n13566));
INVX1 exu_U34120(.A(exu_n20531), .Y(exu_n13567));
INVX1 exu_U34121(.A(exu_n20537), .Y(exu_n13568));
INVX1 exu_U34122(.A(exu_n20543), .Y(exu_n13569));
INVX1 exu_U34123(.A(exu_n20549), .Y(exu_n13570));
INVX1 exu_U34124(.A(exu_n20555), .Y(exu_n13571));
INVX1 exu_U34125(.A(exu_n20561), .Y(exu_n13572));
INVX1 exu_U34126(.A(exu_n20567), .Y(exu_n13573));
INVX1 exu_U34127(.A(exu_n20573), .Y(exu_n13574));
INVX1 exu_U34128(.A(exu_n20579), .Y(exu_n13575));
INVX1 exu_U34129(.A(exu_n20585), .Y(exu_n13576));
INVX1 exu_U34130(.A(exu_n20591), .Y(exu_n13577));
INVX1 exu_U34131(.A(exu_n20597), .Y(exu_n13578));
INVX1 exu_U34132(.A(exu_n20603), .Y(exu_n13579));
INVX1 exu_U34133(.A(exu_n20609), .Y(exu_n13580));
INVX1 exu_U34134(.A(exu_n20615), .Y(exu_n13581));
INVX1 exu_U34135(.A(exu_n20621), .Y(exu_n13582));
INVX1 exu_U34136(.A(exu_n20627), .Y(exu_n13583));
INVX1 exu_U34137(.A(exu_n20633), .Y(exu_n13584));
INVX1 exu_U34138(.A(exu_n20639), .Y(exu_n13585));
INVX1 exu_U34139(.A(exu_n20645), .Y(exu_n13586));
INVX1 exu_U34140(.A(exu_n20651), .Y(exu_n13587));
INVX1 exu_U34141(.A(exu_n20657), .Y(exu_n13588));
INVX1 exu_U34142(.A(exu_n20663), .Y(exu_n13589));
INVX1 exu_U34143(.A(exu_n20669), .Y(exu_n13590));
INVX1 exu_U34144(.A(exu_n20675), .Y(exu_n13591));
INVX1 exu_U34145(.A(exu_n20681), .Y(exu_n13592));
INVX1 exu_U34146(.A(exu_n20687), .Y(exu_n13593));
INVX1 exu_U34147(.A(exu_n20693), .Y(exu_n13594));
INVX1 exu_U34148(.A(exu_n20699), .Y(exu_n13595));
INVX1 exu_U34149(.A(exu_n20705), .Y(exu_n13596));
INVX1 exu_U34150(.A(exu_n20711), .Y(exu_n13597));
INVX1 exu_U34151(.A(exu_n20717), .Y(exu_n13598));
INVX1 exu_U34152(.A(exu_n20723), .Y(exu_n13599));
INVX1 exu_U34153(.A(exu_n20729), .Y(exu_n13600));
INVX1 exu_U34154(.A(exu_n20735), .Y(exu_n13601));
INVX1 exu_U34155(.A(exu_n20741), .Y(exu_n13602));
INVX1 exu_U34156(.A(exu_n20747), .Y(exu_n13603));
INVX1 exu_U34157(.A(exu_n20753), .Y(exu_n13604));
INVX1 exu_U34158(.A(exu_n20759), .Y(exu_n13605));
INVX1 exu_U34159(.A(exu_n20765), .Y(exu_n13606));
INVX1 exu_U34160(.A(exu_n20771), .Y(exu_n13607));
INVX1 exu_U34161(.A(exu_n20777), .Y(exu_n13608));
INVX1 exu_U34162(.A(exu_n20783), .Y(exu_n13609));
INVX1 exu_U34163(.A(exu_n20789), .Y(exu_n13610));
INVX1 exu_U34164(.A(exu_n20795), .Y(exu_n13611));
INVX1 exu_U34165(.A(exu_n20801), .Y(exu_n13612));
INVX1 exu_U34166(.A(exu_n20807), .Y(exu_n13613));
INVX1 exu_U34167(.A(exu_n20813), .Y(exu_n13614));
INVX1 exu_U34168(.A(exu_n20819), .Y(exu_n13615));
INVX1 exu_U34169(.A(exu_n20825), .Y(exu_n13616));
INVX1 exu_U34170(.A(exu_n20831), .Y(exu_n13617));
INVX1 exu_U34171(.A(exu_n20837), .Y(exu_n13618));
INVX1 exu_U34172(.A(exu_n20843), .Y(exu_n13619));
INVX1 exu_U34173(.A(exu_n20849), .Y(exu_n13620));
INVX1 exu_U34174(.A(exu_n20855), .Y(exu_n13621));
INVX1 exu_U34175(.A(exu_n20861), .Y(exu_n13622));
INVX1 exu_U34176(.A(exu_n20867), .Y(exu_n13623));
INVX1 exu_U34177(.A(exu_n20873), .Y(exu_n13624));
INVX1 exu_U34178(.A(exu_n20879), .Y(exu_n13625));
INVX1 exu_U34179(.A(exu_n20885), .Y(exu_n13626));
INVX1 exu_U34180(.A(exu_n20891), .Y(exu_n13627));
INVX1 exu_U34181(.A(exu_n20897), .Y(exu_n13628));
INVX1 exu_U34182(.A(exu_n20903), .Y(exu_n13629));
INVX1 exu_U34183(.A(exu_n20909), .Y(exu_n13630));
INVX1 exu_U34184(.A(exu_n20915), .Y(exu_n13631));
INVX1 exu_U34185(.A(exu_n20921), .Y(exu_n13632));
INVX1 exu_U34186(.A(exu_n20927), .Y(exu_n13633));
INVX1 exu_U34187(.A(exu_n20933), .Y(exu_n13634));
INVX1 exu_U34188(.A(exu_n20939), .Y(exu_n13635));
INVX1 exu_U34189(.A(exu_n20945), .Y(exu_n13636));
INVX1 exu_U34190(.A(exu_n20951), .Y(exu_n13637));
INVX1 exu_U34191(.A(exu_n20957), .Y(exu_n13638));
INVX1 exu_U34192(.A(exu_n20963), .Y(exu_n13639));
INVX1 exu_U34193(.A(exu_n20969), .Y(exu_n13640));
INVX1 exu_U34194(.A(exu_n20975), .Y(exu_n13641));
INVX1 exu_U34195(.A(exu_n20981), .Y(exu_n13642));
INVX1 exu_U34196(.A(exu_n20987), .Y(exu_n13643));
INVX1 exu_U34197(.A(exu_n20993), .Y(exu_n13644));
INVX1 exu_U34198(.A(exu_n20999), .Y(exu_n13645));
INVX1 exu_U34199(.A(exu_n21005), .Y(exu_n13646));
INVX1 exu_U34200(.A(exu_n21011), .Y(exu_n13647));
INVX1 exu_U34201(.A(exu_n21017), .Y(exu_n13648));
INVX1 exu_U34202(.A(exu_n21023), .Y(exu_n13649));
INVX1 exu_U34203(.A(exu_n21029), .Y(exu_n13650));
INVX1 exu_U34204(.A(exu_n21035), .Y(exu_n13651));
INVX1 exu_U34205(.A(exu_n21041), .Y(exu_n13652));
INVX1 exu_U34206(.A(exu_n21047), .Y(exu_n13653));
INVX1 exu_U34207(.A(exu_n21053), .Y(exu_n13654));
INVX1 exu_U34208(.A(exu_n21059), .Y(exu_n13655));
INVX1 exu_U34209(.A(exu_n21065), .Y(exu_n13656));
INVX1 exu_U34210(.A(exu_n21071), .Y(exu_n13657));
INVX1 exu_U34211(.A(exu_n21077), .Y(exu_n13658));
INVX1 exu_U34212(.A(exu_n21083), .Y(exu_n13659));
INVX1 exu_U34213(.A(exu_n21089), .Y(exu_n13660));
INVX1 exu_U34214(.A(exu_n21095), .Y(exu_n13661));
INVX1 exu_U34215(.A(exu_n21101), .Y(exu_n13662));
INVX1 exu_U34216(.A(exu_n21107), .Y(exu_n13663));
INVX1 exu_U34217(.A(exu_n21113), .Y(exu_n13664));
INVX1 exu_U34218(.A(exu_n21119), .Y(exu_n13665));
INVX1 exu_U34219(.A(exu_n21125), .Y(exu_n13666));
INVX1 exu_U34220(.A(exu_n21131), .Y(exu_n13667));
INVX1 exu_U34221(.A(exu_n21137), .Y(exu_n13668));
INVX1 exu_U34222(.A(exu_n21143), .Y(exu_n13669));
INVX1 exu_U34223(.A(exu_n21149), .Y(exu_n13670));
INVX1 exu_U34224(.A(exu_n21155), .Y(exu_n13671));
INVX1 exu_U34225(.A(exu_n21161), .Y(exu_n13672));
INVX1 exu_U34226(.A(exu_n21167), .Y(exu_n13673));
INVX1 exu_U34227(.A(exu_n21173), .Y(exu_n13674));
INVX1 exu_U34228(.A(exu_n21179), .Y(exu_n13675));
INVX1 exu_U34229(.A(exu_n21185), .Y(exu_n13676));
INVX1 exu_U34230(.A(exu_n21191), .Y(exu_n13677));
INVX1 exu_U34231(.A(exu_n21197), .Y(exu_n13678));
INVX1 exu_U34232(.A(exu_n21203), .Y(exu_n13679));
INVX1 exu_U34233(.A(exu_n21209), .Y(exu_n13680));
INVX1 exu_U34234(.A(exu_n21215), .Y(exu_n13681));
INVX1 exu_U34235(.A(exu_n21221), .Y(exu_n13682));
INVX1 exu_U34236(.A(exu_n21227), .Y(exu_n13683));
INVX1 exu_U34237(.A(exu_n21233), .Y(exu_n13684));
INVX1 exu_U34238(.A(exu_n21239), .Y(exu_n13685));
INVX1 exu_U34239(.A(exu_n21245), .Y(exu_n13686));
INVX1 exu_U34240(.A(exu_n21251), .Y(exu_n13687));
INVX1 exu_U34241(.A(exu_n21257), .Y(exu_n13688));
INVX1 exu_U34242(.A(exu_n21263), .Y(exu_n13689));
INVX1 exu_U34243(.A(exu_n21269), .Y(exu_n13690));
INVX1 exu_U34244(.A(exu_n21275), .Y(exu_n13691));
INVX1 exu_U34245(.A(exu_n21281), .Y(exu_n13692));
INVX1 exu_U34246(.A(exu_n21287), .Y(exu_n13693));
INVX1 exu_U34247(.A(exu_n21293), .Y(exu_n13694));
INVX1 exu_U34248(.A(exu_n21299), .Y(exu_n13695));
INVX1 exu_U34249(.A(exu_n21305), .Y(exu_n13696));
INVX1 exu_U34250(.A(exu_n21311), .Y(exu_n13697));
INVX1 exu_U34251(.A(exu_n21317), .Y(exu_n13698));
INVX1 exu_U34252(.A(exu_n21323), .Y(exu_n13699));
INVX1 exu_U34253(.A(exu_n21329), .Y(exu_n13700));
INVX1 exu_U34254(.A(exu_n21335), .Y(exu_n13701));
INVX1 exu_U34255(.A(exu_n21341), .Y(exu_n13702));
INVX1 exu_U34256(.A(exu_n21347), .Y(exu_n13703));
INVX1 exu_U34257(.A(exu_n21353), .Y(exu_n13704));
INVX1 exu_U34258(.A(exu_n21359), .Y(exu_n13705));
INVX1 exu_U34259(.A(exu_n21365), .Y(exu_n13706));
INVX1 exu_U34260(.A(exu_n21371), .Y(exu_n13707));
INVX1 exu_U34261(.A(exu_n21377), .Y(exu_n13708));
INVX1 exu_U34262(.A(exu_n21383), .Y(exu_n13709));
INVX1 exu_U34263(.A(exu_n21389), .Y(exu_n13710));
INVX1 exu_U34264(.A(exu_n21395), .Y(exu_n13711));
INVX1 exu_U34265(.A(exu_n21401), .Y(exu_n13712));
INVX1 exu_U34266(.A(exu_n21407), .Y(exu_n13713));
INVX1 exu_U34267(.A(exu_n21413), .Y(exu_n13714));
INVX1 exu_U34268(.A(exu_n21419), .Y(exu_n13715));
INVX1 exu_U34269(.A(exu_n21425), .Y(exu_n13716));
INVX1 exu_U34270(.A(exu_n21431), .Y(exu_n13717));
INVX1 exu_U34271(.A(exu_n21437), .Y(exu_n13718));
INVX1 exu_U34272(.A(exu_n21443), .Y(exu_n13719));
INVX1 exu_U34273(.A(exu_n21449), .Y(exu_n13720));
INVX1 exu_U34274(.A(exu_n21455), .Y(exu_n13721));
INVX1 exu_U34275(.A(exu_n21461), .Y(exu_n13722));
INVX1 exu_U34276(.A(exu_n21467), .Y(exu_n13723));
INVX1 exu_U34277(.A(exu_n21473), .Y(exu_n13724));
INVX1 exu_U34278(.A(exu_n21479), .Y(exu_n13725));
INVX1 exu_U34279(.A(exu_n21485), .Y(exu_n13726));
INVX1 exu_U34280(.A(exu_n21491), .Y(exu_n13727));
INVX1 exu_U34281(.A(exu_n21497), .Y(exu_n13728));
INVX1 exu_U34282(.A(exu_n21503), .Y(exu_n13729));
INVX1 exu_U34283(.A(exu_n21509), .Y(exu_n13730));
INVX1 exu_U34284(.A(exu_n21515), .Y(exu_n13731));
INVX1 exu_U34285(.A(exu_n21521), .Y(exu_n13732));
INVX1 exu_U34286(.A(exu_n21527), .Y(exu_n13733));
INVX1 exu_U34287(.A(exu_n21533), .Y(exu_n13734));
INVX1 exu_U34288(.A(exu_n21539), .Y(exu_n13735));
INVX1 exu_U34289(.A(exu_n21545), .Y(exu_n13736));
INVX1 exu_U34290(.A(exu_n21551), .Y(exu_n13737));
INVX1 exu_U34291(.A(exu_n21557), .Y(exu_n13738));
INVX1 exu_U34292(.A(exu_n21563), .Y(exu_n13739));
INVX1 exu_U34293(.A(exu_n21569), .Y(exu_n13740));
INVX1 exu_U34294(.A(exu_n21575), .Y(exu_n13741));
INVX1 exu_U34295(.A(exu_n21581), .Y(exu_n13742));
INVX1 exu_U34296(.A(exu_n21587), .Y(exu_n13743));
INVX1 exu_U34297(.A(exu_n21593), .Y(exu_n13744));
INVX1 exu_U34298(.A(exu_n21599), .Y(exu_n13745));
INVX1 exu_U34299(.A(exu_n21605), .Y(exu_n13746));
INVX1 exu_U34300(.A(exu_n21611), .Y(exu_n13747));
INVX1 exu_U34301(.A(exu_n21617), .Y(exu_n13748));
INVX1 exu_U34302(.A(exu_n21623), .Y(exu_n13749));
INVX1 exu_U34303(.A(exu_n23202), .Y(exu_n13750));
INVX1 exu_U34304(.A(exu_n23208), .Y(exu_n13751));
INVX1 exu_U34305(.A(exu_n23214), .Y(exu_n13752));
INVX1 exu_U34306(.A(exu_n23220), .Y(exu_n13753));
INVX1 exu_U34307(.A(exu_n23226), .Y(exu_n13754));
INVX1 exu_U34308(.A(exu_n23232), .Y(exu_n13755));
INVX1 exu_U34309(.A(exu_n23238), .Y(exu_n13756));
INVX1 exu_U34310(.A(exu_n23244), .Y(exu_n13757));
INVX1 exu_U34311(.A(exu_n23250), .Y(exu_n13758));
INVX1 exu_U34312(.A(exu_n23256), .Y(exu_n13759));
INVX1 exu_U34313(.A(exu_n23262), .Y(exu_n13760));
INVX1 exu_U34314(.A(exu_n23268), .Y(exu_n13761));
INVX1 exu_U34315(.A(exu_n23274), .Y(exu_n13762));
INVX1 exu_U34316(.A(exu_n23280), .Y(exu_n13763));
INVX1 exu_U34317(.A(exu_n23286), .Y(exu_n13764));
INVX1 exu_U34318(.A(exu_n23292), .Y(exu_n13765));
INVX1 exu_U34319(.A(exu_n23298), .Y(exu_n13766));
INVX1 exu_U34320(.A(exu_n23304), .Y(exu_n13767));
INVX1 exu_U34321(.A(exu_n23310), .Y(exu_n13768));
INVX1 exu_U34322(.A(exu_n23316), .Y(exu_n13769));
INVX1 exu_U34323(.A(exu_n23322), .Y(exu_n13770));
INVX1 exu_U34324(.A(exu_n23328), .Y(exu_n13771));
INVX1 exu_U34325(.A(exu_n23334), .Y(exu_n13772));
INVX1 exu_U34326(.A(exu_n23340), .Y(exu_n13773));
INVX1 exu_U34327(.A(exu_n23346), .Y(exu_n13774));
INVX1 exu_U34328(.A(exu_n23352), .Y(exu_n13775));
INVX1 exu_U34329(.A(exu_n23358), .Y(exu_n13776));
INVX1 exu_U34330(.A(exu_n23364), .Y(exu_n13777));
INVX1 exu_U34331(.A(exu_n23370), .Y(exu_n13778));
INVX1 exu_U34332(.A(exu_n23376), .Y(exu_n13779));
INVX1 exu_U34333(.A(exu_n23382), .Y(exu_n13780));
INVX1 exu_U34334(.A(exu_n23388), .Y(exu_n13781));
INVX1 exu_U34335(.A(exu_n23394), .Y(exu_n13782));
INVX1 exu_U34336(.A(exu_n23400), .Y(exu_n13783));
INVX1 exu_U34337(.A(exu_n23406), .Y(exu_n13784));
INVX1 exu_U34338(.A(exu_n23412), .Y(exu_n13785));
INVX1 exu_U34339(.A(exu_n23418), .Y(exu_n13786));
INVX1 exu_U34340(.A(exu_n23424), .Y(exu_n13787));
INVX1 exu_U34341(.A(exu_n23430), .Y(exu_n13788));
INVX1 exu_U34342(.A(exu_n23436), .Y(exu_n13789));
INVX1 exu_U34343(.A(exu_n23442), .Y(exu_n13790));
INVX1 exu_U34344(.A(exu_n23448), .Y(exu_n13791));
INVX1 exu_U34345(.A(exu_n23454), .Y(exu_n13792));
INVX1 exu_U34346(.A(exu_n23460), .Y(exu_n13793));
INVX1 exu_U34347(.A(exu_n23466), .Y(exu_n13794));
INVX1 exu_U34348(.A(exu_n23472), .Y(exu_n13795));
INVX1 exu_U34349(.A(exu_n23478), .Y(exu_n13796));
INVX1 exu_U34350(.A(exu_n23484), .Y(exu_n13797));
INVX1 exu_U34351(.A(exu_n23490), .Y(exu_n13798));
INVX1 exu_U34352(.A(exu_n23496), .Y(exu_n13799));
INVX1 exu_U34353(.A(exu_n23502), .Y(exu_n13800));
INVX1 exu_U34354(.A(exu_n23508), .Y(exu_n13801));
INVX1 exu_U34355(.A(exu_n23514), .Y(exu_n13802));
INVX1 exu_U34356(.A(exu_n23520), .Y(exu_n13803));
INVX1 exu_U34357(.A(exu_n23526), .Y(exu_n13804));
INVX1 exu_U34358(.A(exu_n23532), .Y(exu_n13805));
INVX1 exu_U34359(.A(exu_n23538), .Y(exu_n13806));
INVX1 exu_U34360(.A(exu_n23544), .Y(exu_n13807));
INVX1 exu_U34361(.A(exu_n23550), .Y(exu_n13808));
INVX1 exu_U34362(.A(exu_n23556), .Y(exu_n13809));
INVX1 exu_U34363(.A(exu_n23562), .Y(exu_n13810));
INVX1 exu_U34364(.A(exu_n23568), .Y(exu_n13811));
INVX1 exu_U34365(.A(exu_n23574), .Y(exu_n13812));
INVX1 exu_U34366(.A(exu_n23580), .Y(exu_n13813));
INVX1 exu_U34367(.A(exu_n23586), .Y(exu_n13814));
INVX1 exu_U34368(.A(exu_n23592), .Y(exu_n13815));
INVX1 exu_U34369(.A(exu_n23598), .Y(exu_n13816));
INVX1 exu_U34370(.A(exu_n23604), .Y(exu_n13817));
INVX1 exu_U34371(.A(exu_n23610), .Y(exu_n13818));
INVX1 exu_U34372(.A(exu_n23615), .Y(exu_n13819));
INVX1 exu_U34373(.A(exu_n23620), .Y(exu_n13820));
INVX1 exu_U34374(.A(exu_n23625), .Y(exu_n13821));
INVX1 exu_U34375(.A(exu_n23630), .Y(exu_n13822));
INVX1 exu_U34376(.A(exu_n23636), .Y(exu_n13823));
INVX1 exu_U34377(.A(exu_n23641), .Y(exu_n13824));
INVX1 exu_U34378(.A(exu_n23646), .Y(exu_n13825));
INVX1 exu_U34379(.A(exu_n23651), .Y(exu_n13826));
INVX1 exu_U34380(.A(exu_n23656), .Y(exu_n13827));
INVX1 exu_U34381(.A(exu_n23661), .Y(exu_n13828));
INVX1 exu_U34382(.A(exu_n23666), .Y(exu_n13829));
INVX1 exu_U34383(.A(exu_n23671), .Y(exu_n13830));
INVX1 exu_U34384(.A(exu_n23676), .Y(exu_n13831));
INVX1 exu_U34385(.A(exu_n23681), .Y(exu_n13832));
INVX1 exu_U34386(.A(exu_n23686), .Y(exu_n13833));
INVX1 exu_U34387(.A(exu_n23692), .Y(exu_n13834));
INVX1 exu_U34388(.A(exu_n23697), .Y(exu_n13835));
INVX1 exu_U34389(.A(exu_n23702), .Y(exu_n13836));
INVX1 exu_U34390(.A(exu_n23708), .Y(exu_n13837));
INVX1 exu_U34391(.A(exu_n23714), .Y(exu_n13838));
INVX1 exu_U34392(.A(exu_n23720), .Y(exu_n13839));
INVX1 exu_U34393(.A(exu_n23726), .Y(exu_n13840));
INVX1 exu_U34394(.A(exu_n23732), .Y(exu_n13841));
INVX1 exu_U34395(.A(exu_n23738), .Y(exu_n13842));
INVX1 exu_U34396(.A(exu_n23744), .Y(exu_n13843));
INVX1 exu_U34397(.A(exu_n23750), .Y(exu_n13844));
INVX1 exu_U34398(.A(exu_n23756), .Y(exu_n13845));
INVX1 exu_U34399(.A(exu_n23762), .Y(exu_n13846));
INVX1 exu_U34400(.A(exu_n23768), .Y(exu_n13847));
INVX1 exu_U34401(.A(exu_n23774), .Y(exu_n13848));
INVX1 exu_U34402(.A(exu_n23780), .Y(exu_n13849));
INVX1 exu_U34403(.A(exu_n23786), .Y(exu_n13850));
INVX1 exu_U34404(.A(exu_n23792), .Y(exu_n13851));
INVX1 exu_U34405(.A(exu_n23798), .Y(exu_n13852));
INVX1 exu_U34406(.A(exu_n23804), .Y(exu_n13853));
INVX1 exu_U34407(.A(exu_n23810), .Y(exu_n13854));
INVX1 exu_U34408(.A(exu_n23816), .Y(exu_n13855));
INVX1 exu_U34409(.A(exu_n23822), .Y(exu_n13856));
INVX1 exu_U34410(.A(exu_n23828), .Y(exu_n13857));
INVX1 exu_U34411(.A(exu_n23834), .Y(exu_n13858));
INVX1 exu_U34412(.A(exu_n23840), .Y(exu_n13859));
INVX1 exu_U34413(.A(exu_n23846), .Y(exu_n13860));
INVX1 exu_U34414(.A(exu_n23852), .Y(exu_n13861));
INVX1 exu_U34415(.A(exu_n23858), .Y(exu_n13862));
INVX1 exu_U34416(.A(exu_n23864), .Y(exu_n13863));
INVX1 exu_U34417(.A(exu_n23870), .Y(exu_n13864));
INVX1 exu_U34418(.A(exu_n23876), .Y(exu_n13865));
INVX1 exu_U34419(.A(exu_n23882), .Y(exu_n13866));
INVX1 exu_U34420(.A(exu_n23888), .Y(exu_n13867));
INVX1 exu_U34421(.A(exu_n23894), .Y(exu_n13868));
INVX1 exu_U34422(.A(exu_n23900), .Y(exu_n13869));
INVX1 exu_U34423(.A(exu_n23906), .Y(exu_n13870));
INVX1 exu_U34424(.A(exu_n23912), .Y(exu_n13871));
INVX1 exu_U34425(.A(exu_n23918), .Y(exu_n13872));
INVX1 exu_U34426(.A(exu_n23924), .Y(exu_n13873));
INVX1 exu_U34427(.A(exu_n23930), .Y(exu_n13874));
INVX1 exu_U34428(.A(exu_n23936), .Y(exu_n13875));
INVX1 exu_U34429(.A(exu_n23942), .Y(exu_n13876));
INVX1 exu_U34430(.A(exu_n23948), .Y(exu_n13877));
INVX1 exu_U34431(.A(exu_n23954), .Y(exu_n13878));
INVX1 exu_U34432(.A(exu_n23960), .Y(exu_n13879));
INVX1 exu_U34433(.A(exu_n23966), .Y(exu_n13880));
INVX1 exu_U34434(.A(exu_n23972), .Y(exu_n13881));
INVX1 exu_U34435(.A(exu_n23978), .Y(exu_n13882));
INVX1 exu_U34436(.A(exu_n23984), .Y(exu_n13883));
INVX1 exu_U34437(.A(exu_n23990), .Y(exu_n13884));
INVX1 exu_U34438(.A(exu_n23996), .Y(exu_n13885));
INVX1 exu_U34439(.A(exu_n24002), .Y(exu_n13886));
INVX1 exu_U34440(.A(exu_n24008), .Y(exu_n13887));
INVX1 exu_U34441(.A(exu_n24014), .Y(exu_n13888));
INVX1 exu_U34442(.A(exu_n24020), .Y(exu_n13889));
INVX1 exu_U34443(.A(exu_n24026), .Y(exu_n13890));
INVX1 exu_U34444(.A(exu_n24032), .Y(exu_n13891));
INVX1 exu_U34445(.A(exu_n24038), .Y(exu_n13892));
INVX1 exu_U34446(.A(exu_n24044), .Y(exu_n13893));
INVX1 exu_U34447(.A(exu_n24050), .Y(exu_n13894));
INVX1 exu_U34448(.A(exu_n24056), .Y(exu_n13895));
INVX1 exu_U34449(.A(exu_n24062), .Y(exu_n13896));
INVX1 exu_U34450(.A(exu_n24068), .Y(exu_n13897));
INVX1 exu_U34451(.A(exu_n24074), .Y(exu_n13898));
INVX1 exu_U34452(.A(exu_n24080), .Y(exu_n13899));
INVX1 exu_U34453(.A(exu_n24086), .Y(exu_n13900));
INVX1 exu_U34454(.A(exu_n24092), .Y(exu_n13901));
INVX1 exu_U34455(.A(exu_n24098), .Y(exu_n13902));
INVX1 exu_U34456(.A(exu_n24104), .Y(exu_n13903));
INVX1 exu_U34457(.A(exu_n24110), .Y(exu_n13904));
INVX1 exu_U34458(.A(exu_n24116), .Y(exu_n13905));
INVX1 exu_U34459(.A(exu_n24122), .Y(exu_n13906));
INVX1 exu_U34460(.A(exu_n24128), .Y(exu_n13907));
INVX1 exu_U34461(.A(exu_n24134), .Y(exu_n13908));
INVX1 exu_U34462(.A(exu_n24140), .Y(exu_n13909));
INVX1 exu_U34463(.A(exu_n24146), .Y(exu_n13910));
INVX1 exu_U34464(.A(exu_n24152), .Y(exu_n13911));
INVX1 exu_U34465(.A(exu_n24158), .Y(exu_n13912));
INVX1 exu_U34466(.A(exu_n24164), .Y(exu_n13913));
INVX1 exu_U34467(.A(exu_n24170), .Y(exu_n13914));
INVX1 exu_U34468(.A(exu_n24176), .Y(exu_n13915));
INVX1 exu_U34469(.A(exu_n24182), .Y(exu_n13916));
INVX1 exu_U34470(.A(exu_n24188), .Y(exu_n13917));
INVX1 exu_U34471(.A(exu_n24194), .Y(exu_n13918));
INVX1 exu_U34472(.A(exu_n24200), .Y(exu_n13919));
INVX1 exu_U34473(.A(exu_n24206), .Y(exu_n13920));
INVX1 exu_U34474(.A(exu_n24212), .Y(exu_n13921));
INVX1 exu_U34475(.A(exu_n24218), .Y(exu_n13922));
INVX1 exu_U34476(.A(exu_n24224), .Y(exu_n13923));
INVX1 exu_U34477(.A(exu_n24230), .Y(exu_n13924));
INVX1 exu_U34478(.A(exu_n24236), .Y(exu_n13925));
INVX1 exu_U34479(.A(exu_n24242), .Y(exu_n13926));
INVX1 exu_U34480(.A(exu_n24248), .Y(exu_n13927));
INVX1 exu_U34481(.A(exu_n24254), .Y(exu_n13928));
INVX1 exu_U34482(.A(exu_n24260), .Y(exu_n13929));
INVX1 exu_U34483(.A(exu_n24266), .Y(exu_n13930));
INVX1 exu_U34484(.A(exu_n24272), .Y(exu_n13931));
INVX1 exu_U34485(.A(exu_n24278), .Y(exu_n13932));
INVX1 exu_U34486(.A(exu_n24284), .Y(exu_n13933));
INVX1 exu_U34487(.A(exu_n24290), .Y(exu_n13934));
INVX1 exu_U34488(.A(exu_n24296), .Y(exu_n13935));
INVX1 exu_U34489(.A(exu_n24302), .Y(exu_n13936));
INVX1 exu_U34490(.A(exu_n24308), .Y(exu_n13937));
INVX1 exu_U34491(.A(exu_n24314), .Y(exu_n13938));
INVX1 exu_U34492(.A(exu_n24320), .Y(exu_n13939));
INVX1 exu_U34493(.A(exu_n24326), .Y(exu_n13940));
INVX1 exu_U34494(.A(exu_n24332), .Y(exu_n13941));
INVX1 exu_U34495(.A(exu_n24594), .Y(exu_n13942));
INVX1 exu_U34496(.A(exu_n24600), .Y(exu_n13943));
INVX1 exu_U34497(.A(exu_n24606), .Y(exu_n13944));
INVX1 exu_U34498(.A(exu_n24612), .Y(exu_n13945));
INVX1 exu_U34499(.A(exu_n24618), .Y(exu_n13946));
INVX1 exu_U34500(.A(exu_n24624), .Y(exu_n13947));
INVX1 exu_U34501(.A(exu_n24630), .Y(exu_n13948));
INVX1 exu_U34502(.A(exu_n24636), .Y(exu_n13949));
INVX1 exu_U34503(.A(exu_n24642), .Y(exu_n13950));
INVX1 exu_U34504(.A(exu_n24648), .Y(exu_n13951));
INVX1 exu_U34505(.A(exu_n24654), .Y(exu_n13952));
INVX1 exu_U34506(.A(exu_n24660), .Y(exu_n13953));
INVX1 exu_U34507(.A(exu_n24666), .Y(exu_n13954));
INVX1 exu_U34508(.A(exu_n24672), .Y(exu_n13955));
INVX1 exu_U34509(.A(exu_n24678), .Y(exu_n13956));
INVX1 exu_U34510(.A(exu_n24684), .Y(exu_n13957));
INVX1 exu_U34511(.A(exu_n24690), .Y(exu_n13958));
INVX1 exu_U34512(.A(exu_n24696), .Y(exu_n13959));
INVX1 exu_U34513(.A(exu_n24702), .Y(exu_n13960));
INVX1 exu_U34514(.A(exu_n24708), .Y(exu_n13961));
INVX1 exu_U34515(.A(exu_n24714), .Y(exu_n13962));
INVX1 exu_U34516(.A(exu_n24720), .Y(exu_n13963));
INVX1 exu_U34517(.A(exu_n24726), .Y(exu_n13964));
INVX1 exu_U34518(.A(exu_n24732), .Y(exu_n13965));
INVX1 exu_U34519(.A(exu_n24738), .Y(exu_n13966));
INVX1 exu_U34520(.A(exu_n24744), .Y(exu_n13967));
INVX1 exu_U34521(.A(exu_n24750), .Y(exu_n13968));
INVX1 exu_U34522(.A(exu_n24756), .Y(exu_n13969));
INVX1 exu_U34523(.A(exu_n24762), .Y(exu_n13970));
INVX1 exu_U34524(.A(exu_n24768), .Y(exu_n13971));
INVX1 exu_U34525(.A(exu_n24774), .Y(exu_n13972));
INVX1 exu_U34526(.A(exu_n24780), .Y(exu_n13973));
INVX1 exu_U34527(.A(exu_n24786), .Y(exu_n13974));
INVX1 exu_U34528(.A(exu_n24792), .Y(exu_n13975));
INVX1 exu_U34529(.A(exu_n24798), .Y(exu_n13976));
INVX1 exu_U34530(.A(exu_n24804), .Y(exu_n13977));
INVX1 exu_U34531(.A(exu_n24810), .Y(exu_n13978));
INVX1 exu_U34532(.A(exu_n24816), .Y(exu_n13979));
INVX1 exu_U34533(.A(exu_n24822), .Y(exu_n13980));
INVX1 exu_U34534(.A(exu_n24828), .Y(exu_n13981));
INVX1 exu_U34535(.A(exu_n24834), .Y(exu_n13982));
INVX1 exu_U34536(.A(exu_n24840), .Y(exu_n13983));
INVX1 exu_U34537(.A(exu_n24846), .Y(exu_n13984));
INVX1 exu_U34538(.A(exu_n24852), .Y(exu_n13985));
INVX1 exu_U34539(.A(exu_n24858), .Y(exu_n13986));
INVX1 exu_U34540(.A(exu_n24864), .Y(exu_n13987));
INVX1 exu_U34541(.A(exu_n24870), .Y(exu_n13988));
INVX1 exu_U34542(.A(exu_n24876), .Y(exu_n13989));
INVX1 exu_U34543(.A(exu_n24882), .Y(exu_n13990));
INVX1 exu_U34544(.A(exu_n24888), .Y(exu_n13991));
INVX1 exu_U34545(.A(exu_n24894), .Y(exu_n13992));
INVX1 exu_U34546(.A(exu_n24900), .Y(exu_n13993));
INVX1 exu_U34547(.A(exu_n24906), .Y(exu_n13994));
INVX1 exu_U34548(.A(exu_n24912), .Y(exu_n13995));
INVX1 exu_U34549(.A(exu_n24918), .Y(exu_n13996));
INVX1 exu_U34550(.A(exu_n24924), .Y(exu_n13997));
INVX1 exu_U34551(.A(exu_n24930), .Y(exu_n13998));
INVX1 exu_U34552(.A(exu_n24936), .Y(exu_n13999));
INVX1 exu_U34553(.A(exu_n24942), .Y(exu_n14000));
INVX1 exu_U34554(.A(exu_n24948), .Y(exu_n14001));
INVX1 exu_U34555(.A(exu_n24954), .Y(exu_n14002));
INVX1 exu_U34556(.A(exu_n24960), .Y(exu_n14003));
INVX1 exu_U34557(.A(exu_n24966), .Y(exu_n14004));
INVX1 exu_U34558(.A(exu_n24972), .Y(exu_n14005));
INVX1 exu_U34559(.A(exu_n24978), .Y(exu_n14006));
INVX1 exu_U34560(.A(exu_n24984), .Y(exu_n14007));
INVX1 exu_U34561(.A(exu_n24990), .Y(exu_n14008));
INVX1 exu_U34562(.A(exu_n24996), .Y(exu_n14009));
INVX1 exu_U34563(.A(exu_n25002), .Y(exu_n14010));
INVX1 exu_U34564(.A(exu_n25007), .Y(exu_n14011));
INVX1 exu_U34565(.A(exu_n25012), .Y(exu_n14012));
INVX1 exu_U34566(.A(exu_n25017), .Y(exu_n14013));
INVX1 exu_U34567(.A(exu_n25022), .Y(exu_n14014));
INVX1 exu_U34568(.A(exu_n25028), .Y(exu_n14015));
INVX1 exu_U34569(.A(exu_n25033), .Y(exu_n14016));
INVX1 exu_U34570(.A(exu_n25038), .Y(exu_n14017));
INVX1 exu_U34571(.A(exu_n25043), .Y(exu_n14018));
INVX1 exu_U34572(.A(exu_n25048), .Y(exu_n14019));
INVX1 exu_U34573(.A(exu_n25053), .Y(exu_n14020));
INVX1 exu_U34574(.A(exu_n25058), .Y(exu_n14021));
INVX1 exu_U34575(.A(exu_n25063), .Y(exu_n14022));
INVX1 exu_U34576(.A(exu_n25068), .Y(exu_n14023));
INVX1 exu_U34577(.A(exu_n25073), .Y(exu_n14024));
INVX1 exu_U34578(.A(exu_n25078), .Y(exu_n14025));
INVX1 exu_U34579(.A(exu_n25084), .Y(exu_n14026));
INVX1 exu_U34580(.A(exu_n25089), .Y(exu_n14027));
INVX1 exu_U34581(.A(exu_n25094), .Y(exu_n14028));
INVX1 exu_U34582(.A(exu_n25099), .Y(exu_n14029));
INVX1 exu_U34583(.A(exu_n25104), .Y(exu_n14030));
INVX1 exu_U34584(.A(exu_n25109), .Y(exu_n14031));
INVX1 exu_U34585(.A(exu_n25114), .Y(exu_n14032));
INVX1 exu_U34586(.A(exu_n25119), .Y(exu_n14033));
INVX1 exu_U34587(.A(exu_n25124), .Y(exu_n14034));
INVX1 exu_U34588(.A(exu_n25129), .Y(exu_n14035));
INVX1 exu_U34589(.A(exu_n25134), .Y(exu_n14036));
INVX1 exu_U34590(.A(exu_n25140), .Y(exu_n14037));
INVX1 exu_U34591(.A(exu_n25145), .Y(exu_n14038));
INVX1 exu_U34592(.A(exu_n25150), .Y(exu_n14039));
INVX1 exu_U34593(.A(exu_n25155), .Y(exu_n14040));
INVX1 exu_U34594(.A(exu_n25160), .Y(exu_n14041));
INVX1 exu_U34595(.A(exu_n25165), .Y(exu_n14042));
INVX1 exu_U34596(.A(exu_n25170), .Y(exu_n14043));
INVX1 exu_U34597(.A(exu_n25175), .Y(exu_n14044));
INVX1 exu_U34598(.A(exu_n25180), .Y(exu_n14045));
INVX1 exu_U34599(.A(exu_n25186), .Y(exu_n14046));
INVX1 exu_U34600(.A(exu_n25192), .Y(exu_n14047));
INVX1 exu_U34601(.A(exu_n25198), .Y(exu_n14048));
INVX1 exu_U34602(.A(exu_n25204), .Y(exu_n14049));
INVX1 exu_U34603(.A(exu_n25210), .Y(exu_n14050));
INVX1 exu_U34604(.A(exu_n25216), .Y(exu_n14051));
INVX1 exu_U34605(.A(exu_n25222), .Y(exu_n14052));
INVX1 exu_U34606(.A(exu_n25228), .Y(exu_n14053));
INVX1 exu_U34607(.A(exu_n25234), .Y(exu_n14054));
INVX1 exu_U34608(.A(exu_n25240), .Y(exu_n14055));
INVX1 exu_U34609(.A(exu_n25246), .Y(exu_n14056));
INVX1 exu_U34610(.A(exu_n25252), .Y(exu_n14057));
INVX1 exu_U34611(.A(exu_n25258), .Y(exu_n14058));
INVX1 exu_U34612(.A(exu_n25264), .Y(exu_n14059));
INVX1 exu_U34613(.A(exu_n25270), .Y(exu_n14060));
INVX1 exu_U34614(.A(exu_n25276), .Y(exu_n14061));
INVX1 exu_U34615(.A(exu_n25282), .Y(exu_n14062));
INVX1 exu_U34616(.A(exu_n25288), .Y(exu_n14063));
INVX1 exu_U34617(.A(exu_n25294), .Y(exu_n14064));
INVX1 exu_U34618(.A(exu_n25300), .Y(exu_n14065));
INVX1 exu_U34619(.A(exu_n25306), .Y(exu_n14066));
INVX1 exu_U34620(.A(exu_n25312), .Y(exu_n14067));
INVX1 exu_U34621(.A(exu_n25318), .Y(exu_n14068));
INVX1 exu_U34622(.A(exu_n25324), .Y(exu_n14069));
INVX1 exu_U34623(.A(exu_n25330), .Y(exu_n14070));
INVX1 exu_U34624(.A(exu_n25336), .Y(exu_n14071));
INVX1 exu_U34625(.A(exu_n25342), .Y(exu_n14072));
INVX1 exu_U34626(.A(exu_n25348), .Y(exu_n14073));
INVX1 exu_U34627(.A(exu_n25354), .Y(exu_n14074));
INVX1 exu_U34628(.A(exu_n25360), .Y(exu_n14075));
INVX1 exu_U34629(.A(exu_n25366), .Y(exu_n14076));
INVX1 exu_U34630(.A(exu_n25372), .Y(exu_n14077));
INVX1 exu_U34631(.A(exu_n25378), .Y(exu_n14078));
INVX1 exu_U34632(.A(exu_n25384), .Y(exu_n14079));
INVX1 exu_U34633(.A(exu_n25390), .Y(exu_n14080));
INVX1 exu_U34634(.A(exu_n25396), .Y(exu_n14081));
INVX1 exu_U34635(.A(exu_n25402), .Y(exu_n14082));
INVX1 exu_U34636(.A(exu_n25408), .Y(exu_n14083));
INVX1 exu_U34637(.A(exu_n25414), .Y(exu_n14084));
INVX1 exu_U34638(.A(exu_n25420), .Y(exu_n14085));
INVX1 exu_U34639(.A(exu_n25426), .Y(exu_n14086));
INVX1 exu_U34640(.A(exu_n25432), .Y(exu_n14087));
INVX1 exu_U34641(.A(exu_n25438), .Y(exu_n14088));
INVX1 exu_U34642(.A(exu_n25444), .Y(exu_n14089));
INVX1 exu_U34643(.A(exu_n25450), .Y(exu_n14090));
INVX1 exu_U34644(.A(exu_n25456), .Y(exu_n14091));
INVX1 exu_U34645(.A(exu_n25462), .Y(exu_n14092));
INVX1 exu_U34646(.A(exu_n25468), .Y(exu_n14093));
INVX1 exu_U34647(.A(exu_n25474), .Y(exu_n14094));
INVX1 exu_U34648(.A(exu_n25480), .Y(exu_n14095));
INVX1 exu_U34649(.A(exu_n25486), .Y(exu_n14096));
INVX1 exu_U34650(.A(exu_n25492), .Y(exu_n14097));
INVX1 exu_U34651(.A(exu_n25498), .Y(exu_n14098));
INVX1 exu_U34652(.A(exu_n25504), .Y(exu_n14099));
INVX1 exu_U34653(.A(exu_n25510), .Y(exu_n14100));
INVX1 exu_U34654(.A(exu_n25516), .Y(exu_n14101));
INVX1 exu_U34655(.A(exu_n25522), .Y(exu_n14102));
INVX1 exu_U34656(.A(exu_n25528), .Y(exu_n14103));
INVX1 exu_U34657(.A(exu_n25534), .Y(exu_n14104));
INVX1 exu_U34658(.A(exu_n25540), .Y(exu_n14105));
INVX1 exu_U34659(.A(exu_n25546), .Y(exu_n14106));
INVX1 exu_U34660(.A(exu_n25552), .Y(exu_n14107));
INVX1 exu_U34661(.A(exu_n25558), .Y(exu_n14108));
INVX1 exu_U34662(.A(exu_n25564), .Y(exu_n14109));
INVX1 exu_U34663(.A(exu_n25570), .Y(exu_n14110));
INVX1 exu_U34664(.A(exu_n25576), .Y(exu_n14111));
INVX1 exu_U34665(.A(exu_n25582), .Y(exu_n14112));
INVX1 exu_U34666(.A(exu_n25588), .Y(exu_n14113));
INVX1 exu_U34667(.A(exu_n25594), .Y(exu_n14114));
INVX1 exu_U34668(.A(exu_n25600), .Y(exu_n14115));
INVX1 exu_U34669(.A(exu_n25606), .Y(exu_n14116));
INVX1 exu_U34670(.A(exu_n25612), .Y(exu_n14117));
INVX1 exu_U34671(.A(exu_n25618), .Y(exu_n14118));
INVX1 exu_U34672(.A(exu_n25624), .Y(exu_n14119));
INVX1 exu_U34673(.A(exu_n25630), .Y(exu_n14120));
INVX1 exu_U34674(.A(exu_n25636), .Y(exu_n14121));
INVX1 exu_U34675(.A(exu_n25642), .Y(exu_n14122));
INVX1 exu_U34676(.A(exu_n25648), .Y(exu_n14123));
INVX1 exu_U34677(.A(exu_n25654), .Y(exu_n14124));
INVX1 exu_U34678(.A(exu_n25660), .Y(exu_n14125));
INVX1 exu_U34679(.A(exu_n25666), .Y(exu_n14126));
INVX1 exu_U34680(.A(exu_n25672), .Y(exu_n14127));
INVX1 exu_U34681(.A(exu_n25678), .Y(exu_n14128));
INVX1 exu_U34682(.A(exu_n25684), .Y(exu_n14129));
INVX1 exu_U34683(.A(exu_n25690), .Y(exu_n14130));
INVX1 exu_U34684(.A(exu_n25696), .Y(exu_n14131));
INVX1 exu_U34685(.A(exu_n25702), .Y(exu_n14132));
INVX1 exu_U34686(.A(exu_n25708), .Y(exu_n14133));
INVX1 exu_U34687(.A(exu_n25970), .Y(exu_n14134));
INVX1 exu_U34688(.A(exu_n25976), .Y(exu_n14135));
INVX1 exu_U34689(.A(exu_n25982), .Y(exu_n14136));
INVX1 exu_U34690(.A(exu_n25988), .Y(exu_n14137));
INVX1 exu_U34691(.A(exu_n25994), .Y(exu_n14138));
INVX1 exu_U34692(.A(exu_n26000), .Y(exu_n14139));
INVX1 exu_U34693(.A(exu_n26006), .Y(exu_n14140));
INVX1 exu_U34694(.A(exu_n26012), .Y(exu_n14141));
INVX1 exu_U34695(.A(exu_n26018), .Y(exu_n14142));
INVX1 exu_U34696(.A(exu_n26024), .Y(exu_n14143));
INVX1 exu_U34697(.A(exu_n26030), .Y(exu_n14144));
INVX1 exu_U34698(.A(exu_n26036), .Y(exu_n14145));
INVX1 exu_U34699(.A(exu_n26042), .Y(exu_n14146));
INVX1 exu_U34700(.A(exu_n26048), .Y(exu_n14147));
INVX1 exu_U34701(.A(exu_n26054), .Y(exu_n14148));
INVX1 exu_U34702(.A(exu_n26060), .Y(exu_n14149));
INVX1 exu_U34703(.A(exu_n26066), .Y(exu_n14150));
INVX1 exu_U34704(.A(exu_n26072), .Y(exu_n14151));
INVX1 exu_U34705(.A(exu_n26078), .Y(exu_n14152));
INVX1 exu_U34706(.A(exu_n26084), .Y(exu_n14153));
INVX1 exu_U34707(.A(exu_n26090), .Y(exu_n14154));
INVX1 exu_U34708(.A(exu_n26096), .Y(exu_n14155));
INVX1 exu_U34709(.A(exu_n26102), .Y(exu_n14156));
INVX1 exu_U34710(.A(exu_n26108), .Y(exu_n14157));
INVX1 exu_U34711(.A(exu_n26114), .Y(exu_n14158));
INVX1 exu_U34712(.A(exu_n26120), .Y(exu_n14159));
INVX1 exu_U34713(.A(exu_n26126), .Y(exu_n14160));
INVX1 exu_U34714(.A(exu_n26132), .Y(exu_n14161));
INVX1 exu_U34715(.A(exu_n26138), .Y(exu_n14162));
INVX1 exu_U34716(.A(exu_n26144), .Y(exu_n14163));
INVX1 exu_U34717(.A(exu_n26150), .Y(exu_n14164));
INVX1 exu_U34718(.A(exu_n26156), .Y(exu_n14165));
INVX1 exu_U34719(.A(exu_n26162), .Y(exu_n14166));
INVX1 exu_U34720(.A(exu_n26168), .Y(exu_n14167));
INVX1 exu_U34721(.A(exu_n26174), .Y(exu_n14168));
INVX1 exu_U34722(.A(exu_n26180), .Y(exu_n14169));
INVX1 exu_U34723(.A(exu_n26186), .Y(exu_n14170));
INVX1 exu_U34724(.A(exu_n26192), .Y(exu_n14171));
INVX1 exu_U34725(.A(exu_n26198), .Y(exu_n14172));
INVX1 exu_U34726(.A(exu_n26204), .Y(exu_n14173));
INVX1 exu_U34727(.A(exu_n26210), .Y(exu_n14174));
INVX1 exu_U34728(.A(exu_n26216), .Y(exu_n14175));
INVX1 exu_U34729(.A(exu_n26222), .Y(exu_n14176));
INVX1 exu_U34730(.A(exu_n26228), .Y(exu_n14177));
INVX1 exu_U34731(.A(exu_n26234), .Y(exu_n14178));
INVX1 exu_U34732(.A(exu_n26240), .Y(exu_n14179));
INVX1 exu_U34733(.A(exu_n26246), .Y(exu_n14180));
INVX1 exu_U34734(.A(exu_n26252), .Y(exu_n14181));
INVX1 exu_U34735(.A(exu_n26258), .Y(exu_n14182));
INVX1 exu_U34736(.A(exu_n26264), .Y(exu_n14183));
INVX1 exu_U34737(.A(exu_n26270), .Y(exu_n14184));
INVX1 exu_U34738(.A(exu_n26276), .Y(exu_n14185));
INVX1 exu_U34739(.A(exu_n26282), .Y(exu_n14186));
INVX1 exu_U34740(.A(exu_n26288), .Y(exu_n14187));
INVX1 exu_U34741(.A(exu_n26294), .Y(exu_n14188));
INVX1 exu_U34742(.A(exu_n26300), .Y(exu_n14189));
INVX1 exu_U34743(.A(exu_n26306), .Y(exu_n14190));
INVX1 exu_U34744(.A(exu_n26312), .Y(exu_n14191));
INVX1 exu_U34745(.A(exu_n26318), .Y(exu_n14192));
INVX1 exu_U34746(.A(exu_n26324), .Y(exu_n14193));
INVX1 exu_U34747(.A(exu_n26330), .Y(exu_n14194));
INVX1 exu_U34748(.A(exu_n26336), .Y(exu_n14195));
INVX1 exu_U34749(.A(exu_n26342), .Y(exu_n14196));
INVX1 exu_U34750(.A(exu_n26348), .Y(exu_n14197));
INVX1 exu_U34751(.A(exu_n26354), .Y(exu_n14198));
INVX1 exu_U34752(.A(exu_n26360), .Y(exu_n14199));
INVX1 exu_U34753(.A(exu_n26366), .Y(exu_n14200));
INVX1 exu_U34754(.A(exu_n26372), .Y(exu_n14201));
INVX1 exu_U34755(.A(exu_n26378), .Y(exu_n14202));
INVX1 exu_U34756(.A(exu_n26383), .Y(exu_n14203));
INVX1 exu_U34757(.A(exu_n26389), .Y(exu_n14204));
INVX1 exu_U34758(.A(exu_n26395), .Y(exu_n14205));
INVX1 exu_U34759(.A(exu_n26401), .Y(exu_n14206));
INVX1 exu_U34760(.A(exu_n26407), .Y(exu_n14207));
INVX1 exu_U34761(.A(exu_n26413), .Y(exu_n14208));
INVX1 exu_U34762(.A(exu_n26419), .Y(exu_n14209));
INVX1 exu_U34763(.A(exu_n26425), .Y(exu_n14210));
INVX1 exu_U34764(.A(exu_n26431), .Y(exu_n14211));
INVX1 exu_U34765(.A(exu_n26437), .Y(exu_n14212));
INVX1 exu_U34766(.A(exu_n26443), .Y(exu_n14213));
INVX1 exu_U34767(.A(exu_n26449), .Y(exu_n14214));
INVX1 exu_U34768(.A(exu_n26455), .Y(exu_n14215));
INVX1 exu_U34769(.A(exu_n26461), .Y(exu_n14216));
INVX1 exu_U34770(.A(exu_n26467), .Y(exu_n14217));
INVX1 exu_U34771(.A(exu_n26473), .Y(exu_n14218));
INVX1 exu_U34772(.A(exu_n26479), .Y(exu_n14219));
INVX1 exu_U34773(.A(exu_n26485), .Y(exu_n14220));
INVX1 exu_U34774(.A(exu_n26491), .Y(exu_n14221));
INVX1 exu_U34775(.A(exu_n26497), .Y(exu_n14222));
INVX1 exu_U34776(.A(exu_n26503), .Y(exu_n14223));
INVX1 exu_U34777(.A(exu_n26509), .Y(exu_n14224));
INVX1 exu_U34778(.A(exu_n26515), .Y(exu_n14225));
INVX1 exu_U34779(.A(exu_n26521), .Y(exu_n14226));
INVX1 exu_U34780(.A(exu_n26527), .Y(exu_n14227));
INVX1 exu_U34781(.A(exu_n26533), .Y(exu_n14228));
INVX1 exu_U34782(.A(exu_n26539), .Y(exu_n14229));
INVX1 exu_U34783(.A(exu_n26545), .Y(exu_n14230));
INVX1 exu_U34784(.A(exu_n26551), .Y(exu_n14231));
INVX1 exu_U34785(.A(exu_n26557), .Y(exu_n14232));
INVX1 exu_U34786(.A(exu_n26563), .Y(exu_n14233));
INVX1 exu_U34787(.A(exu_n26569), .Y(exu_n14234));
INVX1 exu_U34788(.A(exu_n26575), .Y(exu_n14235));
INVX1 exu_U34789(.A(exu_n26581), .Y(exu_n14236));
INVX1 exu_U34790(.A(exu_n26587), .Y(exu_n14237));
INVX1 exu_U34791(.A(exu_n26592), .Y(exu_n14238));
INVX1 exu_U34792(.A(exu_n26598), .Y(exu_n14239));
INVX1 exu_U34793(.A(exu_n26604), .Y(exu_n14240));
INVX1 exu_U34794(.A(exu_n26610), .Y(exu_n14241));
INVX1 exu_U34795(.A(exu_n26616), .Y(exu_n14242));
INVX1 exu_U34796(.A(exu_n26622), .Y(exu_n14243));
INVX1 exu_U34797(.A(exu_n26628), .Y(exu_n14244));
INVX1 exu_U34798(.A(exu_n26634), .Y(exu_n14245));
INVX1 exu_U34799(.A(exu_n26640), .Y(exu_n14246));
INVX1 exu_U34800(.A(exu_n26646), .Y(exu_n14247));
INVX1 exu_U34801(.A(exu_n26652), .Y(exu_n14248));
INVX1 exu_U34802(.A(exu_n26658), .Y(exu_n14249));
INVX1 exu_U34803(.A(exu_n26664), .Y(exu_n14250));
INVX1 exu_U34804(.A(exu_n26670), .Y(exu_n14251));
INVX1 exu_U34805(.A(exu_n26676), .Y(exu_n14252));
INVX1 exu_U34806(.A(exu_n26682), .Y(exu_n14253));
INVX1 exu_U34807(.A(exu_n26688), .Y(exu_n14254));
INVX1 exu_U34808(.A(exu_n26694), .Y(exu_n14255));
INVX1 exu_U34809(.A(exu_n26700), .Y(exu_n14256));
INVX1 exu_U34810(.A(exu_n26706), .Y(exu_n14257));
INVX1 exu_U34811(.A(exu_n26712), .Y(exu_n14258));
INVX1 exu_U34812(.A(exu_n26718), .Y(exu_n14259));
INVX1 exu_U34813(.A(exu_n26724), .Y(exu_n14260));
INVX1 exu_U34814(.A(exu_n26730), .Y(exu_n14261));
INVX1 exu_U34815(.A(exu_n26736), .Y(exu_n14262));
INVX1 exu_U34816(.A(exu_n26741), .Y(exu_n14263));
INVX1 exu_U34817(.A(exu_n26745), .Y(exu_n14264));
INVX1 exu_U34818(.A(exu_n26749), .Y(exu_n14265));
INVX1 exu_U34819(.A(exu_n26753), .Y(exu_n14266));
INVX1 exu_U34820(.A(exu_n26757), .Y(exu_n14267));
INVX1 exu_U34821(.A(exu_n26761), .Y(exu_n14268));
INVX1 exu_U34822(.A(exu_n26765), .Y(exu_n14269));
INVX1 exu_U34823(.A(exu_n26769), .Y(exu_n14270));
INVX1 exu_U34824(.A(exu_n26773), .Y(exu_n14271));
INVX1 exu_U34825(.A(exu_n26777), .Y(exu_n14272));
INVX1 exu_U34826(.A(exu_n26781), .Y(exu_n14273));
INVX1 exu_U34827(.A(exu_n26785), .Y(exu_n14274));
INVX1 exu_U34828(.A(exu_n26789), .Y(exu_n14275));
INVX1 exu_U34829(.A(exu_n26793), .Y(exu_n14276));
INVX1 exu_U34830(.A(exu_n26797), .Y(exu_n14277));
INVX1 exu_U34831(.A(exu_n26801), .Y(exu_n14278));
INVX1 exu_U34832(.A(exu_n26805), .Y(exu_n14279));
INVX1 exu_U34833(.A(exu_n26809), .Y(exu_n14280));
INVX1 exu_U34834(.A(exu_n26813), .Y(exu_n14281));
INVX1 exu_U34835(.A(exu_n26817), .Y(exu_n14282));
INVX1 exu_U34836(.A(exu_n26821), .Y(exu_n14283));
INVX1 exu_U34837(.A(exu_n26826), .Y(exu_n14284));
INVX1 exu_U34838(.A(exu_n26831), .Y(exu_n14285));
INVX1 exu_U34839(.A(exu_n26836), .Y(exu_n14286));
INVX1 exu_U34840(.A(exu_n26841), .Y(exu_n14287));
INVX1 exu_U34841(.A(exu_n26846), .Y(exu_n14288));
INVX1 exu_U34842(.A(exu_n26851), .Y(exu_n14289));
INVX1 exu_U34843(.A(exu_n26856), .Y(exu_n14290));
INVX1 exu_U34844(.A(exu_n26861), .Y(exu_n14291));
INVX1 exu_U34845(.A(exu_n26866), .Y(exu_n14292));
INVX1 exu_U34846(.A(exu_n26870), .Y(exu_n14293));
INVX1 exu_U34847(.A(exu_n26875), .Y(exu_n14294));
INVX1 exu_U34848(.A(exu_n26880), .Y(exu_n14295));
INVX1 exu_U34849(.A(exu_n26885), .Y(exu_n14296));
INVX1 exu_U34850(.A(exu_n26890), .Y(exu_n14297));
INVX1 exu_U34851(.A(exu_n26895), .Y(exu_n14298));
INVX1 exu_U34852(.A(exu_n26900), .Y(exu_n14299));
INVX1 exu_U34853(.A(exu_n26905), .Y(exu_n14300));
INVX1 exu_U34854(.A(exu_n26911), .Y(exu_n14301));
INVX1 exu_U34855(.A(exu_n26915), .Y(exu_n14302));
INVX1 exu_U34856(.A(exu_n26919), .Y(exu_n14303));
INVX1 exu_U34857(.A(exu_n26923), .Y(exu_n14304));
INVX1 exu_U34858(.A(exu_n26927), .Y(exu_n14305));
INVX1 exu_U34859(.A(exu_n26931), .Y(exu_n14306));
INVX1 exu_U34860(.A(exu_n26935), .Y(exu_n14307));
INVX1 exu_U34861(.A(exu_n26939), .Y(exu_n14308));
INVX1 exu_U34862(.A(exu_n26943), .Y(exu_n14309));
INVX1 exu_U34863(.A(exu_n26947), .Y(exu_n14310));
INVX1 exu_U34864(.A(exu_n26951), .Y(exu_n14311));
INVX1 exu_U34865(.A(exu_n26955), .Y(exu_n14312));
INVX1 exu_U34866(.A(exu_n26959), .Y(exu_n14313));
INVX1 exu_U34867(.A(exu_n26963), .Y(exu_n14314));
INVX1 exu_U34868(.A(exu_n26967), .Y(exu_n14315));
INVX1 exu_U34869(.A(exu_n26971), .Y(exu_n14316));
INVX1 exu_U34870(.A(exu_n26975), .Y(exu_n14317));
INVX1 exu_U34871(.A(exu_n26979), .Y(exu_n14318));
INVX1 exu_U34872(.A(exu_n26984), .Y(exu_n14319));
INVX1 exu_U34873(.A(exu_n26988), .Y(exu_n14320));
INVX1 exu_U34874(.A(exu_n26992), .Y(exu_n14321));
INVX1 exu_U34875(.A(exu_n26996), .Y(exu_n14322));
INVX1 exu_U34876(.A(exu_n27000), .Y(exu_n14323));
INVX1 exu_U34877(.A(exu_n27004), .Y(exu_n14324));
INVX1 exu_U34878(.A(exu_n27008), .Y(exu_n14325));
INVX1 exu_U34879(.A(exu_n27012), .Y(exu_n14326));
INVX1 exu_U34880(.A(exu_n27018), .Y(exu_n14327));
INVX1 exu_U34881(.A(exu_n27024), .Y(exu_n14328));
INVX1 exu_U34882(.A(exu_n27030), .Y(exu_n14329));
INVX1 exu_U34883(.A(exu_n27035), .Y(exu_n14330));
INVX1 exu_U34884(.A(exu_n27038), .Y(exu_n14331));
INVX1 exu_U34885(.A(exu_n27041), .Y(exu_n14332));
INVX1 exu_U34886(.A(exu_n27044), .Y(exu_n14333));
INVX1 exu_U34887(.A(exu_n27049), .Y(exu_n14334));
INVX1 exu_U34888(.A(exu_n27055), .Y(exu_n14335));
INVX1 exu_U34889(.A(exu_n27060), .Y(exu_n14336));
INVX1 exu_U34890(.A(exu_n27064), .Y(exu_n14337));
INVX1 exu_U34891(.A(exu_n27068), .Y(exu_n14338));
INVX1 exu_U34892(.A(exu_n27073), .Y(exu_n14339));
INVX1 exu_U34893(.A(exu_n27078), .Y(exu_n14340));
INVX1 exu_U34894(.A(exu_n27083), .Y(exu_n14341));
INVX1 exu_U34895(.A(exu_n27088), .Y(exu_n14342));
INVX1 exu_U34896(.A(exu_n27093), .Y(exu_n14343));
INVX1 exu_U34897(.A(exu_n27099), .Y(exu_n14344));
INVX1 exu_U34898(.A(exu_n27105), .Y(exu_n14345));
INVX1 exu_U34899(.A(exu_n27111), .Y(exu_n14346));
INVX1 exu_U34900(.A(exu_n27117), .Y(exu_n14347));
INVX1 exu_U34901(.A(exu_n27123), .Y(exu_n14348));
INVX1 exu_U34902(.A(exu_n27129), .Y(exu_n14349));
INVX1 exu_U34903(.A(exu_n27135), .Y(exu_n14350));
INVX1 exu_U34904(.A(exu_n27141), .Y(exu_n14351));
INVX1 exu_U34905(.A(exu_n27147), .Y(exu_n14352));
INVX1 exu_U34906(.A(exu_n27153), .Y(exu_n14353));
INVX1 exu_U34907(.A(exu_n27159), .Y(exu_n14354));
INVX1 exu_U34908(.A(exu_n27165), .Y(exu_n14355));
INVX1 exu_U34909(.A(exu_n27171), .Y(exu_n14356));
INVX1 exu_U34910(.A(exu_n27177), .Y(exu_n14357));
INVX1 exu_U34911(.A(exu_n27183), .Y(exu_n14358));
INVX1 exu_U34912(.A(exu_n27189), .Y(exu_n14359));
INVX1 exu_U34913(.A(exu_n27195), .Y(exu_n14360));
INVX1 exu_U34914(.A(exu_n27201), .Y(exu_n14361));
INVX1 exu_U34915(.A(exu_n27207), .Y(exu_n14362));
INVX1 exu_U34916(.A(exu_n27213), .Y(exu_n14363));
INVX1 exu_U34917(.A(exu_n27219), .Y(exu_n14364));
INVX1 exu_U34918(.A(exu_n27225), .Y(exu_n14365));
INVX1 exu_U34919(.A(exu_n27231), .Y(exu_n14366));
INVX1 exu_U34920(.A(exu_n27237), .Y(exu_n14367));
INVX1 exu_U34921(.A(exu_n27243), .Y(exu_n14368));
INVX1 exu_U34922(.A(exu_n27249), .Y(exu_n14369));
INVX1 exu_U34923(.A(exu_n27255), .Y(exu_n14370));
INVX1 exu_U34924(.A(exu_n27261), .Y(exu_n14371));
INVX1 exu_U34925(.A(exu_n27267), .Y(exu_n14372));
INVX1 exu_U34926(.A(exu_n27273), .Y(exu_n14373));
INVX1 exu_U34927(.A(exu_n27279), .Y(exu_n14374));
INVX1 exu_U34928(.A(exu_n27285), .Y(exu_n14375));
INVX1 exu_U34929(.A(exu_n27291), .Y(exu_n14376));
INVX1 exu_U34930(.A(exu_n27297), .Y(exu_n14377));
INVX1 exu_U34931(.A(exu_n27303), .Y(exu_n14378));
INVX1 exu_U34932(.A(exu_n27309), .Y(exu_n14379));
INVX1 exu_U34933(.A(exu_n27315), .Y(exu_n14380));
INVX1 exu_U34934(.A(exu_n27321), .Y(exu_n14381));
INVX1 exu_U34935(.A(exu_n27327), .Y(exu_n14382));
INVX1 exu_U34936(.A(exu_n27333), .Y(exu_n14383));
INVX1 exu_U34937(.A(exu_n27339), .Y(exu_n14384));
INVX1 exu_U34938(.A(exu_n27345), .Y(exu_n14385));
INVX1 exu_U34939(.A(exu_n27351), .Y(exu_n14386));
INVX1 exu_U34940(.A(exu_n27357), .Y(exu_n14387));
INVX1 exu_U34941(.A(exu_n27363), .Y(exu_n14388));
INVX1 exu_U34942(.A(exu_n27369), .Y(exu_n14389));
INVX1 exu_U34943(.A(exu_n27375), .Y(exu_n14390));
INVX1 exu_U34944(.A(exu_n27381), .Y(exu_n14391));
INVX1 exu_U34945(.A(exu_n27387), .Y(exu_n14392));
INVX1 exu_U34946(.A(exu_n27393), .Y(exu_n14393));
INVX1 exu_U34947(.A(exu_n27399), .Y(exu_n14394));
INVX1 exu_U34948(.A(exu_n27402), .Y(exu_n14395));
INVX1 exu_U34949(.A(exu_n27408), .Y(exu_n14396));
INVX1 exu_U34950(.A(exu_n27413), .Y(exu_n14397));
INVX1 exu_U34951(.A(exu_n27419), .Y(exu_n14398));
INVX1 exu_U34952(.A(exu_n27425), .Y(exu_n14399));
INVX1 exu_U34953(.A(exu_n27431), .Y(exu_n14400));
INVX1 exu_U34954(.A(exu_n27437), .Y(exu_n14401));
INVX1 exu_U34955(.A(exu_n27443), .Y(exu_n14402));
INVX1 exu_U34956(.A(exu_n27449), .Y(exu_n14403));
INVX1 exu_U34957(.A(exu_n27455), .Y(exu_n14404));
INVX1 exu_U34958(.A(exu_n27461), .Y(exu_n14405));
INVX1 exu_U34959(.A(exu_n27467), .Y(exu_n14406));
INVX1 exu_U34960(.A(exu_n27473), .Y(exu_n14407));
INVX1 exu_U34961(.A(exu_n27479), .Y(exu_n14408));
INVX1 exu_U34962(.A(exu_n27485), .Y(exu_n14409));
INVX1 exu_U34963(.A(exu_n27491), .Y(exu_n14410));
INVX1 exu_U34964(.A(exu_n27497), .Y(exu_n14411));
INVX1 exu_U34965(.A(exu_n27503), .Y(exu_n14412));
INVX1 exu_U34966(.A(exu_n27509), .Y(exu_n14413));
INVX1 exu_U34967(.A(exu_n27515), .Y(exu_n14414));
INVX1 exu_U34968(.A(exu_n27521), .Y(exu_n14415));
INVX1 exu_U34969(.A(exu_n27527), .Y(exu_n14416));
INVX1 exu_U34970(.A(exu_n27533), .Y(exu_n14417));
INVX1 exu_U34971(.A(exu_n27539), .Y(exu_n14418));
INVX1 exu_U34972(.A(exu_n27545), .Y(exu_n14419));
INVX1 exu_U34973(.A(exu_n27551), .Y(exu_n14420));
INVX1 exu_U34974(.A(exu_n27557), .Y(exu_n14421));
INVX1 exu_U34975(.A(exu_n27563), .Y(exu_n14422));
INVX1 exu_U34976(.A(exu_n27569), .Y(exu_n14423));
INVX1 exu_U34977(.A(exu_n27575), .Y(exu_n14424));
INVX1 exu_U34978(.A(exu_n27581), .Y(exu_n14425));
INVX1 exu_U34979(.A(exu_n27587), .Y(exu_n14426));
INVX1 exu_U34980(.A(exu_n27593), .Y(exu_n14427));
INVX1 exu_U34981(.A(exu_n27599), .Y(exu_n14428));
INVX1 exu_U34982(.A(exu_n27605), .Y(exu_n14429));
INVX1 exu_U34983(.A(exu_n27611), .Y(exu_n14430));
INVX1 exu_U34984(.A(exu_n27617), .Y(exu_n14431));
INVX1 exu_U34985(.A(exu_n27623), .Y(exu_n14432));
INVX1 exu_U34986(.A(exu_n27629), .Y(exu_n14433));
INVX1 exu_U34987(.A(exu_n27635), .Y(exu_n14434));
INVX1 exu_U34988(.A(exu_n27641), .Y(exu_n14435));
INVX1 exu_U34989(.A(exu_n27647), .Y(exu_n14436));
INVX1 exu_U34990(.A(exu_n27653), .Y(exu_n14437));
INVX1 exu_U34991(.A(exu_n27659), .Y(exu_n14438));
INVX1 exu_U34992(.A(exu_n27665), .Y(exu_n14439));
INVX1 exu_U34993(.A(exu_n27671), .Y(exu_n14440));
INVX1 exu_U34994(.A(exu_n27677), .Y(exu_n14441));
INVX1 exu_U34995(.A(exu_n27683), .Y(exu_n14442));
INVX1 exu_U34996(.A(exu_n27689), .Y(exu_n14443));
INVX1 exu_U34997(.A(exu_n27695), .Y(exu_n14444));
INVX1 exu_U34998(.A(exu_n27701), .Y(exu_n14445));
INVX1 exu_U34999(.A(exu_n27707), .Y(exu_n14446));
INVX1 exu_U35000(.A(exu_n27713), .Y(exu_n14447));
INVX1 exu_U35001(.A(exu_n27719), .Y(exu_n14448));
INVX1 exu_U35002(.A(exu_n27725), .Y(exu_n14449));
INVX1 exu_U35003(.A(exu_n27731), .Y(exu_n14450));
INVX1 exu_U35004(.A(exu_n27737), .Y(exu_n14451));
INVX1 exu_U35005(.A(exu_n27743), .Y(exu_n14452));
INVX1 exu_U35006(.A(exu_n27749), .Y(exu_n14453));
INVX1 exu_U35007(.A(exu_n27759), .Y(exu_n14454));
INVX1 exu_U35008(.A(exu_n27765), .Y(exu_n14455));
INVX1 exu_U35009(.A(exu_n27771), .Y(exu_n14456));
INVX1 exu_U35010(.A(exu_n27777), .Y(exu_n14457));
INVX1 exu_U35011(.A(exu_n27784), .Y(exu_n14458));
INVX1 exu_U35012(.A(exu_n27790), .Y(exu_n14459));
INVX1 exu_U35013(.A(exu_n27796), .Y(exu_n14460));
INVX1 exu_U35014(.A(exu_n27802), .Y(exu_n14461));
INVX1 exu_U35015(.A(exu_n27808), .Y(exu_n14462));
INVX1 exu_U35016(.A(exu_n27814), .Y(exu_n14463));
INVX1 exu_U35017(.A(exu_n27820), .Y(exu_n14464));
INVX1 exu_U35018(.A(exu_n27826), .Y(exu_n14465));
INVX1 exu_U35019(.A(exu_n27832), .Y(exu_n14466));
INVX1 exu_U35020(.A(exu_n27838), .Y(exu_n14467));
INVX1 exu_U35021(.A(exu_n27845), .Y(exu_n14468));
INVX1 exu_U35022(.A(exu_n27851), .Y(exu_n14469));
INVX1 exu_U35023(.A(exu_n27856), .Y(exu_n14470));
INVX1 exu_U35024(.A(exu_n27860), .Y(exu_n14471));
INVX1 exu_U35025(.A(exu_n27864), .Y(exu_n14472));
INVX1 exu_U35026(.A(exu_n27868), .Y(exu_n14473));
INVX1 exu_U35027(.A(exu_n27872), .Y(exu_n14474));
INVX1 exu_U35028(.A(exu_n27876), .Y(exu_n14475));
INVX1 exu_U35029(.A(exu_n27880), .Y(exu_n14476));
INVX1 exu_U35030(.A(exu_n27884), .Y(exu_n14477));
INVX1 exu_U35031(.A(exu_n27889), .Y(exu_n14478));
INVX1 exu_U35032(.A(exu_n27893), .Y(exu_n14479));
INVX1 exu_U35033(.A(exu_n27897), .Y(exu_n14480));
INVX1 exu_U35034(.A(exu_n27901), .Y(exu_n14481));
INVX1 exu_U35035(.A(exu_n27905), .Y(exu_n14482));
INVX1 exu_U35036(.A(exu_n27909), .Y(exu_n14483));
INVX1 exu_U35037(.A(exu_n27913), .Y(exu_n14484));
INVX1 exu_U35038(.A(exu_n27917), .Y(exu_n14485));
INVX1 exu_U35039(.A(exu_n27978), .Y(exu_n14486));
INVX1 exu_U35040(.A(exu_n27982), .Y(exu_n14487));
INVX1 exu_U35041(.A(exu_n27993), .Y(exu_n14488));
INVX1 exu_U35042(.A(exu_n27999), .Y(exu_n14489));
INVX1 exu_U35043(.A(exu_n28005), .Y(exu_n14490));
INVX1 exu_U35044(.A(exu_n28011), .Y(exu_n14491));
INVX1 exu_U35045(.A(exu_n28020), .Y(exu_n14492));
INVX1 exu_U35046(.A(exu_n28026), .Y(exu_n14493));
INVX1 exu_U35047(.A(exu_n28032), .Y(exu_n14494));
INVX1 exu_U35048(.A(exu_n28038), .Y(exu_n14495));
INVX1 exu_U35049(.A(exu_n28044), .Y(exu_n14496));
INVX1 exu_U35050(.A(exu_n28050), .Y(exu_n14497));
INVX1 exu_U35051(.A(exu_n28056), .Y(exu_n14498));
INVX1 exu_U35052(.A(exu_n28062), .Y(exu_n14499));
INVX1 exu_U35053(.A(exu_n28068), .Y(exu_n14500));
INVX1 exu_U35054(.A(exu_n28074), .Y(exu_n14501));
INVX1 exu_U35055(.A(exu_n28083), .Y(exu_n14502));
INVX1 exu_U35056(.A(exu_n28089), .Y(exu_n14503));
INVX1 exu_U35057(.A(exu_n28095), .Y(exu_n14504));
INVX1 exu_U35058(.A(exu_n28101), .Y(exu_n14505));
INVX1 exu_U35059(.A(exu_n28107), .Y(exu_n14506));
INVX1 exu_U35060(.A(exu_n28113), .Y(exu_n14507));
INVX1 exu_U35061(.A(exu_n28119), .Y(exu_n14508));
INVX1 exu_U35062(.A(exu_n28125), .Y(exu_n14509));
INVX1 exu_U35063(.A(exu_n28131), .Y(exu_n14510));
INVX1 exu_U35064(.A(exu_n28137), .Y(exu_n14511));
INVX1 exu_U35065(.A(exu_n28144), .Y(exu_n14512));
INVX1 exu_U35066(.A(exu_n28150), .Y(exu_n14513));
INVX1 exu_U35067(.A(exu_n28156), .Y(exu_n14514));
INVX1 exu_U35068(.A(exu_n28162), .Y(exu_n14515));
INVX1 exu_U35069(.A(exu_n28168), .Y(exu_n14516));
INVX1 exu_U35070(.A(exu_n28174), .Y(exu_n14517));
INVX1 exu_U35071(.A(exu_n28180), .Y(exu_n14518));
INVX1 exu_U35072(.A(exu_n28186), .Y(exu_n14519));
INVX1 exu_U35073(.A(exu_n28192), .Y(exu_n14520));
INVX1 exu_U35074(.A(exu_n28198), .Y(exu_n14521));
INVX1 exu_U35075(.A(exu_n28205), .Y(exu_n14522));
INVX1 exu_U35076(.A(exu_n28211), .Y(exu_n14523));
INVX1 exu_U35077(.A(exu_n28217), .Y(exu_n14524));
INVX1 exu_U35078(.A(exu_n28223), .Y(exu_n14525));
INVX1 exu_U35079(.A(exu_n28229), .Y(exu_n14526));
INVX1 exu_U35080(.A(exu_n28235), .Y(exu_n14527));
INVX1 exu_U35081(.A(exu_n28241), .Y(exu_n14528));
INVX1 exu_U35082(.A(exu_n28247), .Y(exu_n14529));
INVX1 exu_U35083(.A(exu_n28253), .Y(exu_n14530));
INVX1 exu_U35084(.A(exu_n28259), .Y(exu_n14531));
INVX1 exu_U35085(.A(exu_n28266), .Y(exu_n14532));
INVX1 exu_U35086(.A(exu_n28272), .Y(exu_n14533));
INVX1 exu_U35087(.A(exu_n28278), .Y(exu_n14534));
INVX1 exu_U35088(.A(exu_n28284), .Y(exu_n14535));
INVX1 exu_U35089(.A(exu_n28290), .Y(exu_n14536));
INVX1 exu_U35090(.A(exu_n28296), .Y(exu_n14537));
INVX1 exu_U35091(.A(exu_n28302), .Y(exu_n14538));
INVX1 exu_U35092(.A(exu_n28308), .Y(exu_n14539));
INVX1 exu_U35093(.A(exu_n28313), .Y(exu_n14540));
INVX1 exu_U35094(.A(exu_n28317), .Y(exu_n14541));
INVX1 exu_U35095(.A(exu_n28323), .Y(exu_n14542));
INVX1 exu_U35096(.A(exu_n28329), .Y(exu_n14543));
INVX1 exu_U35097(.A(exu_n28335), .Y(exu_n14544));
INVX1 exu_U35098(.A(exu_n28341), .Y(exu_n14545));
INVX1 exu_U35099(.A(exu_n28347), .Y(exu_n14546));
INVX1 exu_U35100(.A(exu_n28353), .Y(exu_n14547));
INVX1 exu_U35101(.A(exu_n28359), .Y(exu_n14548));
INVX1 exu_U35102(.A(exu_n28365), .Y(exu_n14549));
INVX1 exu_U35103(.A(exu_n28371), .Y(exu_n14550));
INVX1 exu_U35104(.A(exu_n28377), .Y(exu_n14551));
INVX1 exu_U35105(.A(exu_n28383), .Y(exu_n14552));
INVX1 exu_U35106(.A(exu_n28389), .Y(exu_n14553));
INVX1 exu_U35107(.A(exu_n28395), .Y(exu_n14554));
INVX1 exu_U35108(.A(exu_n28401), .Y(exu_n14555));
INVX1 exu_U35109(.A(exu_n28407), .Y(exu_n14556));
INVX1 exu_U35110(.A(exu_n28413), .Y(exu_n14557));
INVX1 exu_U35111(.A(exu_n28419), .Y(exu_n14558));
INVX1 exu_U35112(.A(exu_n28425), .Y(exu_n14559));
INVX1 exu_U35113(.A(exu_n28431), .Y(exu_n14560));
INVX1 exu_U35114(.A(exu_n28437), .Y(exu_n14561));
INVX1 exu_U35115(.A(exu_n28443), .Y(exu_n14562));
INVX1 exu_U35116(.A(exu_n28449), .Y(exu_n14563));
INVX1 exu_U35117(.A(exu_n28455), .Y(exu_n14564));
INVX1 exu_U35118(.A(exu_n28461), .Y(exu_n14565));
INVX1 exu_U35119(.A(exu_n28467), .Y(exu_n14566));
INVX1 exu_U35120(.A(exu_n28473), .Y(exu_n14567));
INVX1 exu_U35121(.A(exu_n28479), .Y(exu_n14568));
INVX1 exu_U35122(.A(exu_n28485), .Y(exu_n14569));
INVX1 exu_U35123(.A(exu_n28491), .Y(exu_n14570));
INVX1 exu_U35124(.A(exu_n28497), .Y(exu_n14571));
INVX1 exu_U35125(.A(exu_n28503), .Y(exu_n14572));
INVX1 exu_U35126(.A(exu_n28509), .Y(exu_n14573));
INVX1 exu_U35127(.A(exu_n28515), .Y(exu_n14574));
INVX1 exu_U35128(.A(exu_n28521), .Y(exu_n14575));
INVX1 exu_U35129(.A(exu_n28527), .Y(exu_n14576));
INVX1 exu_U35130(.A(exu_n28533), .Y(exu_n14577));
INVX1 exu_U35131(.A(exu_n28539), .Y(exu_n14578));
INVX1 exu_U35132(.A(exu_n28545), .Y(exu_n14579));
INVX1 exu_U35133(.A(exu_n28551), .Y(exu_n14580));
INVX1 exu_U35134(.A(exu_n28557), .Y(exu_n14581));
INVX1 exu_U35135(.A(exu_n28563), .Y(exu_n14582));
INVX1 exu_U35136(.A(exu_n28568), .Y(exu_n14583));
INVX1 exu_U35137(.A(exu_n28573), .Y(exu_n14584));
INVX1 exu_U35138(.A(exu_n28579), .Y(exu_n14585));
INVX1 exu_U35139(.A(exu_n28585), .Y(exu_n14586));
INVX1 exu_U35140(.A(exu_n28591), .Y(exu_n14587));
INVX1 exu_U35141(.A(exu_n28597), .Y(exu_n14588));
INVX1 exu_U35142(.A(exu_n28603), .Y(exu_n14589));
INVX1 exu_U35143(.A(exu_n28609), .Y(exu_n14590));
INVX1 exu_U35144(.A(exu_n28615), .Y(exu_n14591));
INVX1 exu_U35145(.A(exu_n28621), .Y(exu_n14592));
INVX1 exu_U35146(.A(exu_n28627), .Y(exu_n14593));
INVX1 exu_U35147(.A(exu_n28636), .Y(exu_n14594));
INVX1 exu_U35148(.A(exu_n28642), .Y(exu_n14595));
INVX1 exu_U35149(.A(exu_n28648), .Y(exu_n14596));
INVX1 exu_U35150(.A(exu_n28654), .Y(exu_n14597));
INVX1 exu_U35151(.A(exu_n28660), .Y(exu_n14598));
INVX1 exu_U35152(.A(exu_n28666), .Y(exu_n14599));
INVX1 exu_U35153(.A(exu_n28672), .Y(exu_n14600));
INVX1 exu_U35154(.A(exu_n28678), .Y(exu_n14601));
INVX1 exu_U35155(.A(exu_n28684), .Y(exu_n14602));
INVX1 exu_U35156(.A(exu_n28690), .Y(exu_n14603));
INVX1 exu_U35157(.A(exu_n28697), .Y(exu_n14604));
INVX1 exu_U35158(.A(exu_n28703), .Y(exu_n14605));
INVX1 exu_U35159(.A(exu_n28709), .Y(exu_n14606));
INVX1 exu_U35160(.A(exu_n28715), .Y(exu_n14607));
INVX1 exu_U35161(.A(exu_n28725), .Y(exu_n14608));
INVX1 exu_U35162(.A(exu_n28741), .Y(exu_n14609));
INVX1 exu_U35163(.A(exu_n28757), .Y(exu_n14610));
INVX1 exu_U35164(.A(exu_n28774), .Y(exu_n14611));
INVX1 exu_U35165(.A(exu_n28780), .Y(exu_n14612));
INVX1 exu_U35166(.A(exu_n28786), .Y(exu_n14613));
INVX1 exu_U35167(.A(exu_n28792), .Y(exu_n14614));
INVX1 exu_U35168(.A(exu_n28798), .Y(exu_n14615));
INVX1 exu_U35169(.A(exu_n28804), .Y(exu_n14616));
INVX1 exu_U35170(.A(exu_n28810), .Y(exu_n14617));
INVX1 exu_U35171(.A(exu_n28816), .Y(exu_n14618));
INVX1 exu_U35172(.A(exu_n28822), .Y(exu_n14619));
INVX1 exu_U35173(.A(exu_n28828), .Y(exu_n14620));
INVX1 exu_U35174(.A(exu_n28834), .Y(exu_n14621));
INVX1 exu_U35175(.A(exu_n28840), .Y(exu_n14622));
INVX1 exu_U35176(.A(exu_n28846), .Y(exu_n14623));
INVX1 exu_U35177(.A(exu_n28852), .Y(exu_n14624));
INVX1 exu_U35178(.A(exu_n28858), .Y(exu_n14625));
INVX1 exu_U35179(.A(exu_n28864), .Y(exu_n14626));
INVX1 exu_U35180(.A(exu_n28870), .Y(exu_n14627));
INVX1 exu_U35181(.A(exu_n28876), .Y(exu_n14628));
INVX1 exu_U35182(.A(exu_n28882), .Y(exu_n14629));
INVX1 exu_U35183(.A(exu_n28888), .Y(exu_n14630));
INVX1 exu_U35184(.A(exu_n28894), .Y(exu_n14631));
INVX1 exu_U35185(.A(exu_n28900), .Y(exu_n14632));
INVX1 exu_U35186(.A(exu_n28906), .Y(exu_n14633));
INVX1 exu_U35187(.A(exu_n28912), .Y(exu_n14634));
INVX1 exu_U35188(.A(exu_n28918), .Y(exu_n14635));
INVX1 exu_U35189(.A(exu_n28924), .Y(exu_n14636));
INVX1 exu_U35190(.A(exu_n28930), .Y(exu_n14637));
INVX1 exu_U35191(.A(exu_n28936), .Y(exu_n14638));
INVX1 exu_U35192(.A(exu_n28942), .Y(exu_n14639));
INVX1 exu_U35193(.A(exu_n28948), .Y(exu_n14640));
INVX1 exu_U35194(.A(exu_n28954), .Y(exu_n14641));
INVX1 exu_U35195(.A(exu_n28960), .Y(exu_n14642));
INVX1 exu_U35196(.A(exu_n28966), .Y(exu_n14643));
INVX1 exu_U35197(.A(exu_n28972), .Y(exu_n14644));
INVX1 exu_U35198(.A(exu_n28978), .Y(exu_n14645));
INVX1 exu_U35199(.A(exu_n28984), .Y(exu_n14646));
INVX1 exu_U35200(.A(exu_n28990), .Y(exu_n14647));
INVX1 exu_U35201(.A(exu_n28996), .Y(exu_n14648));
INVX1 exu_U35202(.A(exu_n29002), .Y(exu_n14649));
INVX1 exu_U35203(.A(exu_n29008), .Y(exu_n14650));
INVX1 exu_U35204(.A(exu_n29014), .Y(exu_n14651));
INVX1 exu_U35205(.A(exu_n29020), .Y(exu_n14652));
INVX1 exu_U35206(.A(exu_n29026), .Y(exu_n14653));
INVX1 exu_U35207(.A(exu_n29032), .Y(exu_n14654));
INVX1 exu_U35208(.A(exu_n29038), .Y(exu_n14655));
INVX1 exu_U35209(.A(exu_n29044), .Y(exu_n14656));
INVX1 exu_U35210(.A(exu_n29050), .Y(exu_n14657));
INVX1 exu_U35211(.A(exu_n29056), .Y(exu_n14658));
INVX1 exu_U35212(.A(exu_n29062), .Y(exu_n14659));
INVX1 exu_U35213(.A(exu_n29068), .Y(exu_n14660));
INVX1 exu_U35214(.A(exu_n29074), .Y(exu_n14661));
INVX1 exu_U35215(.A(exu_n29080), .Y(exu_n14662));
INVX1 exu_U35216(.A(exu_n29086), .Y(exu_n14663));
INVX1 exu_U35217(.A(exu_n29092), .Y(exu_n14664));
INVX1 exu_U35218(.A(exu_n29098), .Y(exu_n14665));
INVX1 exu_U35219(.A(exu_n29104), .Y(exu_n14666));
INVX1 exu_U35220(.A(exu_n29110), .Y(exu_n14667));
INVX1 exu_U35221(.A(exu_n29116), .Y(exu_n14668));
INVX1 exu_U35222(.A(exu_n29122), .Y(exu_n14669));
INVX1 exu_U35223(.A(exu_n29128), .Y(exu_n14670));
INVX1 exu_U35224(.A(exu_n29134), .Y(exu_n14671));
INVX1 exu_U35225(.A(exu_n29140), .Y(exu_n14672));
INVX1 exu_U35226(.A(exu_n29146), .Y(exu_n14673));
INVX1 exu_U35227(.A(exu_n29152), .Y(exu_n14674));
INVX1 exu_U35228(.A(exu_n29158), .Y(exu_n14675));
INVX1 exu_U35229(.A(exu_n29164), .Y(exu_n14676));
INVX1 exu_U35230(.A(exu_n29170), .Y(exu_n14677));
INVX1 exu_U35231(.A(exu_n29176), .Y(exu_n14678));
INVX1 exu_U35232(.A(exu_n29182), .Y(exu_n14679));
INVX1 exu_U35233(.A(exu_n29188), .Y(exu_n14680));
INVX1 exu_U35234(.A(exu_n29194), .Y(exu_n14681));
INVX1 exu_U35235(.A(exu_n29200), .Y(exu_n14682));
INVX1 exu_U35236(.A(exu_n29206), .Y(exu_n14683));
INVX1 exu_U35237(.A(exu_n29212), .Y(exu_n14684));
INVX1 exu_U35238(.A(exu_n29218), .Y(exu_n14685));
INVX1 exu_U35239(.A(exu_n29224), .Y(exu_n14686));
INVX1 exu_U35240(.A(exu_n29230), .Y(exu_n14687));
INVX1 exu_U35241(.A(exu_n29236), .Y(exu_n14688));
INVX1 exu_U35242(.A(exu_n29242), .Y(exu_n14689));
INVX1 exu_U35243(.A(exu_n29248), .Y(exu_n14690));
INVX1 exu_U35244(.A(exu_n29254), .Y(exu_n14691));
INVX1 exu_U35245(.A(exu_n29260), .Y(exu_n14692));
INVX1 exu_U35246(.A(exu_n29266), .Y(exu_n14693));
INVX1 exu_U35247(.A(exu_n29272), .Y(exu_n14694));
INVX1 exu_U35248(.A(exu_n29278), .Y(exu_n14695));
INVX1 exu_U35249(.A(exu_n29284), .Y(exu_n14696));
INVX1 exu_U35250(.A(exu_n29290), .Y(exu_n14697));
INVX1 exu_U35251(.A(exu_n29296), .Y(exu_n14698));
INVX1 exu_U35252(.A(exu_n31458), .Y(exu_n14699));
INVX1 exu_U35253(.A(exu_n31464), .Y(exu_n14700));
INVX1 exu_U35254(.A(exu_n31469), .Y(exu_n14701));
INVX1 exu_U35255(.A(exu_n31474), .Y(exu_n14702));
INVX1 exu_U35256(.A(exu_n31479), .Y(exu_n14703));
INVX1 exu_U35257(.A(exu_n31484), .Y(exu_n14704));
INVX1 exu_U35258(.A(exu_n31617), .Y(exu_n14705));
INVX1 exu_U35259(.A(exu_n31647), .Y(exu_n14706));
INVX1 exu_U35260(.A(exu_n31677), .Y(exu_n14707));
INVX1 exu_U35261(.A(rml_cwp_cwp_output_mux_n2), .Y(exu_n14708));
INVX1 exu_U35262(.A(rml_cwp_cwp_output_mux_n8), .Y(exu_n14709));
INVX1 exu_U35263(.A(rml_cwp_cwp_output_mux_n14), .Y(exu_n14710));
INVX1 exu_U35264(.A(rml_cwp_cwp_output_mux_n20), .Y(exu_n14711));
INVX1 exu_U35265(.A(rml_cwp_cwp_output_mux_n26), .Y(exu_n14712));
INVX1 exu_U35266(.A(rml_cwp_cwp_output_mux_n32), .Y(exu_n14713));
INVX1 exu_U35267(.A(rml_cwp_cwp_output_mux_n38), .Y(exu_n14714));
INVX1 exu_U35268(.A(rml_cwp_cwp_output_mux_n44), .Y(exu_n14715));
INVX1 exu_U35269(.A(rml_cwp_cwp_output_mux_n50), .Y(exu_n14716));
INVX1 exu_U35270(.A(rml_cwp_cwp_output_mux_n56), .Y(exu_n14717));
INVX1 exu_U35271(.A(rml_cwp_cwp_output_mux_n62), .Y(exu_n14718));
INVX1 exu_U35272(.A(rml_cwp_cwp_output_mux_n68), .Y(exu_n14719));
INVX1 exu_U35273(.A(rml_cwp_cwp_output_mux_n74), .Y(exu_n14720));
INVX1 exu_U35274(.A(rml_cwp_cwp_output_mux_n80), .Y(exu_n14721));
INVX1 exu_U35275(.A(rml_cwp_cwp_output_mux_n86), .Y(exu_n14722));
AND2X1 exu_U35276(.A(ecl_divcntl_cnt6_n23), .B(ecl_divcntl_cntr[3]), .Y(ecl_divcntl_cnt6_n17));
INVX1 exu_U35277(.A(ecl_divcntl_cnt6_n17), .Y(exu_n14723));
AND2X1 exu_U35278(.A(ecl_divcntl_cntr[2]), .B(exu_n16623), .Y(ecl_divcntl_cnt6_n24));
INVX1 exu_U35279(.A(ecl_divcntl_cnt6_n24), .Y(exu_n14724));
INVX1 exu_U35280(.A(ecl_writeback_rdpr_mux1_n2), .Y(exu_n14725));
INVX1 exu_U35281(.A(ecl_writeback_rdpr_mux1_n8), .Y(exu_n14726));
INVX1 exu_U35282(.A(ecl_writeback_rdpr_mux1_n14), .Y(exu_n14727));
INVX1 exu_U35283(.A(ecl_writeback_rd_g_mux_n2), .Y(exu_n14728));
INVX1 exu_U35284(.A(ecl_writeback_rd_g_mux_n8), .Y(exu_n14729));
INVX1 exu_U35285(.A(ecl_writeback_rd_g_mux_n14), .Y(exu_n14730));
INVX1 exu_U35286(.A(ecl_writeback_rd_g_mux_n20), .Y(exu_n14731));
INVX1 exu_U35287(.A(ecl_writeback_rd_g_mux_n26), .Y(exu_n14732));
INVX1 exu_U35288(.A(ecl_ccr_mux_ccr_out_n2), .Y(exu_n14733));
INVX1 exu_U35289(.A(ecl_ccr_mux_ccr_out_n8), .Y(exu_n14734));
INVX1 exu_U35290(.A(ecl_ccr_mux_ccr_out_n14), .Y(exu_n14735));
INVX1 exu_U35291(.A(ecl_ccr_mux_ccr_out_n20), .Y(exu_n14736));
INVX1 exu_U35292(.A(ecl_ccr_mux_ccr_out_n26), .Y(exu_n14737));
INVX1 exu_U35293(.A(ecl_ccr_mux_ccr_out_n32), .Y(exu_n14738));
INVX1 exu_U35294(.A(ecl_ccr_mux_ccr_out_n38), .Y(exu_n14739));
INVX1 exu_U35295(.A(ecl_ccr_mux_ccr_out_n44), .Y(exu_n14740));
INVX1 exu_U35296(.A(rml_mux_agp_out1_n2), .Y(exu_n14741));
INVX1 exu_U35297(.A(rml_mux_agp_out1_n8), .Y(exu_n14742));
AND2X1 exu_U35298(.A(exu_n15472), .B(exu_n15368), .Y(rml_cwp_n78));
INVX1 exu_U35299(.A(rml_cwp_n78), .Y(exu_n14743));
AND2X1 exu_U35300(.A(exu_n15473), .B(exu_n15369), .Y(rml_cwp_n81));
INVX1 exu_U35301(.A(rml_cwp_n81), .Y(exu_n14744));
AND2X1 exu_U35302(.A(exu_n15474), .B(exu_n15370), .Y(rml_cwp_n84));
INVX1 exu_U35303(.A(rml_cwp_n84), .Y(exu_n14745));
AND2X1 exu_U35304(.A(exu_n15475), .B(exu_n15371), .Y(rml_cwp_n87));
INVX1 exu_U35305(.A(rml_cwp_n87), .Y(exu_n14746));
INVX1 exu_U35306(.A(div_low32or_n2), .Y(exu_n14747));
AND2X1 exu_U35307(.A(exu_mul_input_vld), .B(ecl_mdqctl_n20), .Y(ecl_mdqctl_n19));
INVX1 exu_U35308(.A(ecl_mdqctl_n19), .Y(exu_n14748));
AND2X1 exu_U35309(.A(ecl_divcntl_div_state_1), .B(exu_n16185), .Y(ecl_divcntl_n34));
INVX1 exu_U35310(.A(ecl_divcntl_n34), .Y(exu_n14749));
AND2X1 exu_U35311(.A(exu_n16257), .B(exu_n16205), .Y(ecl_divcntl_n47));
INVX1 exu_U35312(.A(ecl_divcntl_n47), .Y(exu_n14750));
AND2X1 exu_U35313(.A(ecl_mdqctl_divcntl_muldone), .B(exu_n16503), .Y(ecl_divcntl_n49));
INVX1 exu_U35314(.A(ecl_divcntl_n49), .Y(exu_n14751));
AND2X1 exu_U35315(.A(exu_n15424), .B(exu_n16185), .Y(ecl_divcntl_n58));
INVX1 exu_U35316(.A(ecl_divcntl_n58), .Y(exu_n14752));
AND2X1 exu_U35317(.A(exu_n15684), .B(exu_n16557), .Y(ecl_divcntl_n73));
INVX1 exu_U35318(.A(ecl_divcntl_n73), .Y(exu_n14753));
AND2X1 exu_U35319(.A(ecl_divcntl_n88), .B(ecl_divcntl_cntr[5]), .Y(ecl_divcntl_n87));
INVX1 exu_U35320(.A(ecl_divcntl_n87), .Y(exu_n14754));
AND2X1 exu_U35321(.A(ecl_byplog_rs2_n19), .B(ecl_byplog_rs2_n29), .Y(ecl_byplog_rs2_n22));
INVX1 exu_U35322(.A(ecl_byplog_rs2_n22), .Y(exu_n14755));
AND2X1 exu_U35323(.A(ecl_byplog_rs1_n17), .B(exu_n15767), .Y(ecl_byplog_rs1_n27));
INVX1 exu_U35324(.A(ecl_byplog_rs1_n27), .Y(exu_n14756));
AND2X1 exu_U35325(.A(exu_n15345), .B(ecl_byplog_rs1_n35), .Y(ecl_byplog_rs1_n34));
INVX1 exu_U35326(.A(ecl_byplog_rs1_n34), .Y(exu_n14757));
AND2X1 exu_U35327(.A(lsu_exu_dfill_vld_g), .B(ecl_ld_thr_match_dg), .Y(ecl_byplog_rs1_n37));
INVX1 exu_U35328(.A(ecl_byplog_rs1_n37), .Y(exu_n14758));
AND2X1 exu_U35329(.A(ecl_thr_match_dm), .B(ecl_bypass_m), .Y(ecl_byplog_rs1_n48));
INVX1 exu_U35330(.A(ecl_byplog_rs1_n48), .Y(exu_n14759));
AND2X1 exu_U35331(.A(ecl_wb_e), .B(ecl_thr_match_de), .Y(ecl_byplog_rs1_n50));
INVX1 exu_U35332(.A(ecl_byplog_rs1_n50), .Y(exu_n14760));
AND2X1 exu_U35333(.A(exu_n15692), .B(ifu_tlu_sraddr_d[3]), .Y(ecl_writeback_n69));
INVX1 exu_U35334(.A(ecl_writeback_n69), .Y(exu_n14761));
AND2X1 exu_U35335(.A(ifu_tlu_sraddr_d[3]), .B(exu_n16374), .Y(ecl_writeback_n71));
INVX1 exu_U35336(.A(ecl_writeback_n71), .Y(exu_n14762));
AND2X1 exu_U35337(.A(exu_n15741), .B(ecl_writeback_n77), .Y(ecl_writeback_n75));
INVX1 exu_U35338(.A(ecl_writeback_n75), .Y(exu_n14763));
AND2X1 exu_U35339(.A(exu_n15743), .B(ecl_writeback_n81), .Y(ecl_writeback_n79));
INVX1 exu_U35340(.A(ecl_writeback_n79), .Y(exu_n14764));
AND2X1 exu_U35341(.A(exu_n15744), .B(ecl_writeback_n85), .Y(ecl_writeback_n83));
INVX1 exu_U35342(.A(ecl_writeback_n83), .Y(exu_n14765));
AND2X1 exu_U35343(.A(ecl_writeback_sraddr_e[5]), .B(ecl_writeback_sraddr_e[3]), .Y(ecl_writeback_n137));
INVX1 exu_U35344(.A(ecl_writeback_n137), .Y(exu_n14766));
AND2X1 exu_U35345(.A(ecl_writeback_sraddr_w[1]), .B(exu_n16555), .Y(ecl_writeback_n143));
INVX1 exu_U35346(.A(ecl_writeback_n143), .Y(exu_n14767));
AND2X1 exu_U35347(.A(ecl_tid_w1[0]), .B(ecl_tid_w1[1]), .Y(ecl_writeback_n177));
INVX1 exu_U35348(.A(ecl_writeback_n177), .Y(exu_n14768));
AND2X1 exu_U35349(.A(ecl_tid_w1[1]), .B(exu_n16575), .Y(ecl_writeback_n179));
INVX1 exu_U35350(.A(ecl_writeback_n179), .Y(exu_n14769));
AND2X1 exu_U35351(.A(exu_n15457), .B(ecl_mdqctl_wb_multhr_g[0]), .Y(ecl_writeback_n188));
INVX1 exu_U35352(.A(ecl_writeback_n188), .Y(exu_n14770));
AND2X1 exu_U35353(.A(exu_n15457), .B(exu_n15374), .Y(ecl_writeback_n190));
INVX1 exu_U35354(.A(ecl_writeback_n190), .Y(exu_n14771));
INVX1 exu_U35355(.A(ecl_ccr_n36), .Y(exu_n14772));
INVX1 exu_U35356(.A(ecl_yreg0_mux_n2), .Y(exu_n14773));
AND2X1 exu_U35357(.A(exu_n15480), .B(ecc_err_m[3]), .Y(ecc_decode_n26));
INVX1 exu_U35358(.A(ecc_decode_n26), .Y(exu_n14774));
AND2X1 exu_U35359(.A(ecc_decode_n27), .B(ecc_decode_n34), .Y(ecc_decode_n33));
INVX1 exu_U35360(.A(ecc_decode_n33), .Y(exu_n14775));
INVX1 exu_U35361(.A(bypass_ifu_exu_sr_mux_n2), .Y(exu_n14776));
INVX1 exu_U35362(.A(bypass_ifu_exu_sr_mux_n8), .Y(exu_n14777));
INVX1 exu_U35363(.A(bypass_ifu_exu_sr_mux_n14), .Y(exu_n14778));
INVX1 exu_U35364(.A(bypass_ifu_exu_sr_mux_n20), .Y(exu_n14779));
INVX1 exu_U35365(.A(bypass_ifu_exu_sr_mux_n50), .Y(exu_n14780));
INVX1 exu_U35366(.A(bypass_ifu_exu_sr_mux_n116), .Y(exu_n14781));
INVX1 exu_U35367(.A(bypass_ifu_exu_sr_mux_n182), .Y(exu_n14782));
INVX1 exu_U35368(.A(bypass_ifu_exu_sr_mux_n236), .Y(exu_n14783));
INVX1 exu_U35369(.A(bypass_ifu_exu_sr_mux_n242), .Y(exu_n14784));
INVX1 exu_U35370(.A(bypass_ifu_exu_sr_mux_n248), .Y(exu_n14785));
INVX1 exu_U35371(.A(bypass_ifu_exu_sr_mux_n254), .Y(exu_n14786));
INVX1 exu_U35372(.A(bypass_ifu_exu_sr_mux_n260), .Y(exu_n14787));
INVX1 exu_U35373(.A(bypass_ifu_exu_sr_mux_n266), .Y(exu_n14788));
INVX1 exu_U35374(.A(bypass_ifu_exu_sr_mux_n272), .Y(exu_n14789));
INVX1 exu_U35375(.A(bypass_ifu_exu_sr_mux_n278), .Y(exu_n14790));
INVX1 exu_U35376(.A(bypass_ifu_exu_sr_mux_n284), .Y(exu_n14791));
INVX1 exu_U35377(.A(bypass_ifu_exu_sr_mux_n290), .Y(exu_n14792));
INVX1 exu_U35378(.A(bypass_ifu_exu_sr_mux_n296), .Y(exu_n14793));
INVX1 exu_U35379(.A(bypass_ifu_exu_sr_mux_n302), .Y(exu_n14794));
INVX1 exu_U35380(.A(bypass_ifu_exu_sr_mux_n308), .Y(exu_n14795));
INVX1 exu_U35381(.A(bypass_ifu_exu_sr_mux_n314), .Y(exu_n14796));
INVX1 exu_U35382(.A(bypass_ifu_exu_sr_mux_n320), .Y(exu_n14797));
INVX1 exu_U35383(.A(bypass_ifu_exu_sr_mux_n326), .Y(exu_n14798));
INVX1 exu_U35384(.A(bypass_ifu_exu_sr_mux_n332), .Y(exu_n14799));
INVX1 exu_U35385(.A(bypass_ifu_exu_sr_mux_n338), .Y(exu_n14800));
INVX1 exu_U35386(.A(bypass_ifu_exu_sr_mux_n344), .Y(exu_n14801));
INVX1 exu_U35387(.A(bypass_ifu_exu_sr_mux_n350), .Y(exu_n14802));
INVX1 exu_U35388(.A(bypass_ifu_exu_sr_mux_n356), .Y(exu_n14803));
INVX1 exu_U35389(.A(bypass_ifu_exu_sr_mux_n362), .Y(exu_n14804));
INVX1 exu_U35390(.A(bypass_ifu_exu_sr_mux_n368), .Y(exu_n14805));
INVX1 exu_U35391(.A(bypass_ifu_exu_sr_mux_n374), .Y(exu_n14806));
INVX1 exu_U35392(.A(bypass_ifu_exu_sr_mux_n380), .Y(exu_n14807));
AND2X1 exu_U35393(.A(exu_n15685), .B(ecl_rml_cwp_wen_e), .Y(rml_n56));
INVX1 exu_U35394(.A(rml_n56), .Y(exu_n14808));
INVX1 exu_U35395(.A(rml_ecl_rmlop_done_e), .Y(exu_n14809));
INVX1 exu_U35396(.A(rml_n63), .Y(exu_n14810));
INVX1 exu_U35397(.A(rml_n72), .Y(exu_n14811));
INVX1 exu_U35398(.A(rml_n104), .Y(exu_n14812));
INVX1 exu_U35399(.A(rml_n109), .Y(exu_n14813));
INVX1 exu_U35400(.A(div_n38), .Y(exu_n14814));
INVX1 exu_U35401(.A(div_n68), .Y(exu_n14815));
INVX1 exu_U35402(.A(alu_n70), .Y(exu_n14816));
AND2X1 exu_U35403(.A(ecl_misalign_addr_e), .B(exu_n16381), .Y(ecl_n48));
INVX1 exu_U35404(.A(ecl_n48), .Y(exu_n14817));
INVX1 exu_U35405(.A(ecl_n83), .Y(exu_n14818));
AND2X1 exu_U35406(.A(ecl_ifu_exu_aluop_e[0]), .B(exu_n16402), .Y(ecl_n106));
INVX1 exu_U35407(.A(ecl_n106), .Y(exu_n14819));
AND2X1 exu_U35408(.A(exu_n16400), .B(exu_n16402), .Y(ecl_n107));
INVX1 exu_U35409(.A(ecl_n107), .Y(exu_n14820));
AND2X1 exu_U35410(.A(exu_n16401), .B(exu_n16402), .Y(ecl_n109));
INVX1 exu_U35411(.A(ecl_n109), .Y(exu_n14821));
AND2X1 exu_U35412(.A(exu_n16638), .B(exu_n16637), .Y(exu_n16639));
INVX1 exu_U35413(.A(exu_n16639), .Y(exu_n14822));
AND2X1 exu_U35414(.A(exu_n16666), .B(exu_n16665), .Y(exu_n16667));
INVX1 exu_U35415(.A(exu_n16667), .Y(exu_n14823));
AND2X1 exu_U35416(.A(exu_n16680), .B(exu_n16679), .Y(exu_n16681));
INVX1 exu_U35417(.A(exu_n16681), .Y(exu_n14824));
AND2X1 exu_U35418(.A(exu_n16694), .B(exu_n16693), .Y(exu_n16695));
INVX1 exu_U35419(.A(exu_n16695), .Y(exu_n14825));
AND2X1 exu_U35420(.A(exu_n16722), .B(exu_n16721), .Y(exu_n16723));
INVX1 exu_U35421(.A(exu_n16723), .Y(exu_n14826));
AND2X1 exu_U35422(.A(exu_n16736), .B(exu_n16735), .Y(exu_n16737));
INVX1 exu_U35423(.A(exu_n16737), .Y(exu_n14827));
AND2X1 exu_U35424(.A(exu_n17379), .B(exu_n17378), .Y(exu_n17380));
INVX1 exu_U35425(.A(exu_n17380), .Y(exu_n14828));
AND2X1 exu_U35426(.A(exu_n17393), .B(exu_n17392), .Y(exu_n17394));
INVX1 exu_U35427(.A(exu_n17394), .Y(exu_n14829));
AND2X1 exu_U35428(.A(exu_n17400), .B(exu_n17399), .Y(exu_n17401));
INVX1 exu_U35429(.A(exu_n17401), .Y(exu_n14830));
AND2X1 exu_U35430(.A(exu_n17414), .B(exu_n17413), .Y(exu_n17415));
INVX1 exu_U35431(.A(exu_n17415), .Y(exu_n14831));
AND2X1 exu_U35432(.A(exu_n17442), .B(exu_n17441), .Y(exu_n17443));
INVX1 exu_U35433(.A(exu_n17443), .Y(exu_n14832));
AND2X1 exu_U35434(.A(exu_n17456), .B(exu_n17455), .Y(exu_n17457));
INVX1 exu_U35435(.A(exu_n17457), .Y(exu_n14833));
AND2X1 exu_U35436(.A(exu_n17630), .B(exu_n17631), .Y(exu_n17629));
INVX1 exu_U35437(.A(exu_n17629), .Y(exu_n14834));
AND2X1 exu_U35438(.A(exu_n17636), .B(exu_n17637), .Y(exu_n17635));
INVX1 exu_U35439(.A(exu_n17635), .Y(exu_n14835));
AND2X1 exu_U35440(.A(exu_n17642), .B(exu_n17643), .Y(exu_n17641));
INVX1 exu_U35441(.A(exu_n17641), .Y(exu_n14836));
AND2X1 exu_U35442(.A(exu_n17648), .B(exu_n17649), .Y(exu_n17647));
INVX1 exu_U35443(.A(exu_n17647), .Y(exu_n14837));
AND2X1 exu_U35444(.A(exu_n17654), .B(exu_n17655), .Y(exu_n17653));
INVX1 exu_U35445(.A(exu_n17653), .Y(exu_n14838));
AND2X1 exu_U35446(.A(exu_n17660), .B(exu_n17661), .Y(exu_n17659));
INVX1 exu_U35447(.A(exu_n17659), .Y(exu_n14839));
AND2X1 exu_U35448(.A(exu_n17666), .B(exu_n17667), .Y(exu_n17665));
INVX1 exu_U35449(.A(exu_n17665), .Y(exu_n14840));
AND2X1 exu_U35450(.A(exu_n17672), .B(exu_n17673), .Y(exu_n17671));
INVX1 exu_U35451(.A(exu_n17671), .Y(exu_n14841));
AND2X1 exu_U35452(.A(exu_n17678), .B(exu_n17679), .Y(exu_n17677));
INVX1 exu_U35453(.A(exu_n17677), .Y(exu_n14842));
AND2X1 exu_U35454(.A(exu_n17684), .B(exu_n17685), .Y(exu_n17683));
INVX1 exu_U35455(.A(exu_n17683), .Y(exu_n14843));
AND2X1 exu_U35456(.A(exu_n17690), .B(exu_n17691), .Y(exu_n17689));
INVX1 exu_U35457(.A(exu_n17689), .Y(exu_n14844));
AND2X1 exu_U35458(.A(exu_n17695), .B(exu_n17696), .Y(exu_n17694));
INVX1 exu_U35459(.A(exu_n17694), .Y(exu_n14845));
AND2X1 exu_U35460(.A(exu_n17701), .B(exu_n17702), .Y(exu_n17700));
INVX1 exu_U35461(.A(exu_n17700), .Y(exu_n14846));
AND2X1 exu_U35462(.A(exu_n17706), .B(exu_n17707), .Y(exu_n17705));
INVX1 exu_U35463(.A(exu_n17705), .Y(exu_n14847));
INVX1 exu_U35464(.A(alu_zcomp_in[8]), .Y(exu_n14848));
INVX1 exu_U35465(.A(alu_zcomp_in[6]), .Y(exu_n14849));
INVX1 exu_U35466(.A(alu_zcomp_in[62]), .Y(exu_n14850));
INVX1 exu_U35467(.A(alu_zcomp_in[60]), .Y(exu_n14851));
INVX1 exu_U35468(.A(alu_zcomp_in[58]), .Y(exu_n14852));
INVX1 exu_U35469(.A(alu_zcomp_in[56]), .Y(exu_n14853));
INVX1 exu_U35470(.A(alu_zcomp_in[54]), .Y(exu_n14854));
INVX1 exu_U35471(.A(alu_zcomp_in[52]), .Y(exu_n14855));
INVX1 exu_U35472(.A(alu_zcomp_in[50]), .Y(exu_n14856));
INVX1 exu_U35473(.A(alu_zcomp_in[4]), .Y(exu_n14857));
INVX1 exu_U35474(.A(alu_zcomp_in[48]), .Y(exu_n14858));
INVX1 exu_U35475(.A(alu_zcomp_in[46]), .Y(exu_n14859));
INVX1 exu_U35476(.A(alu_zcomp_in[44]), .Y(exu_n14860));
INVX1 exu_U35477(.A(alu_zcomp_in[42]), .Y(exu_n14861));
INVX1 exu_U35478(.A(alu_zcomp_in[40]), .Y(exu_n14862));
INVX1 exu_U35479(.A(alu_zcomp_in[38]), .Y(exu_n14863));
INVX1 exu_U35480(.A(alu_zcomp_in[36]), .Y(exu_n14864));
INVX1 exu_U35481(.A(alu_zcomp_in[34]), .Y(exu_n14865));
INVX1 exu_U35482(.A(alu_zcomp_in[32]), .Y(exu_n14866));
INVX1 exu_U35483(.A(alu_zcomp_in[31]), .Y(exu_n14867));
INVX1 exu_U35484(.A(alu_zcomp_in[2]), .Y(exu_n14868));
INVX1 exu_U35485(.A(alu_zcomp_in[28]), .Y(exu_n14869));
INVX1 exu_U35486(.A(alu_zcomp_in[26]), .Y(exu_n14870));
INVX1 exu_U35487(.A(alu_zcomp_in[24]), .Y(exu_n14871));
INVX1 exu_U35488(.A(alu_zcomp_in[22]), .Y(exu_n14872));
INVX1 exu_U35489(.A(alu_zcomp_in[20]), .Y(exu_n14873));
INVX1 exu_U35490(.A(alu_zcomp_in[19]), .Y(exu_n14874));
INVX1 exu_U35491(.A(alu_zcomp_in[17]), .Y(exu_n14875));
INVX1 exu_U35492(.A(alu_zcomp_in[15]), .Y(exu_n14876));
INVX1 exu_U35493(.A(alu_zcomp_in[13]), .Y(exu_n14877));
INVX1 exu_U35494(.A(alu_zcomp_in[11]), .Y(exu_n14878));
INVX1 exu_U35495(.A(alu_zcomp_in[0]), .Y(exu_n14879));
INVX1 exu_U35496(.A(div_gencc_in_8), .Y(exu_n14880));
INVX1 exu_U35497(.A(div_gencc_in_6), .Y(exu_n14881));
INVX1 exu_U35498(.A(div_gencc_in_4), .Y(exu_n14882));
INVX1 exu_U35499(.A(div_gencc_in_2), .Y(exu_n14883));
INVX1 exu_U35500(.A(div_gencc_in_28), .Y(exu_n14884));
INVX1 exu_U35501(.A(div_gencc_in_26), .Y(exu_n14885));
INVX1 exu_U35502(.A(div_gencc_in_24), .Y(exu_n14886));
INVX1 exu_U35503(.A(div_gencc_in_22), .Y(exu_n14887));
INVX1 exu_U35504(.A(div_gencc_in_20), .Y(exu_n14888));
INVX1 exu_U35505(.A(div_gencc_in_19), .Y(exu_n14889));
INVX1 exu_U35506(.A(div_gencc_in_17), .Y(exu_n14890));
INVX1 exu_U35507(.A(div_gencc_in_15), .Y(exu_n14891));
INVX1 exu_U35508(.A(div_gencc_in_13), .Y(exu_n14892));
INVX1 exu_U35509(.A(div_gencc_in_11), .Y(exu_n14893));
INVX1 exu_U35510(.A(div_gencc_in_0), .Y(exu_n14894));
INVX1 exu_U35511(.A(div_z_in[8]), .Y(exu_n14895));
INVX1 exu_U35512(.A(div_z_in[6]), .Y(exu_n14896));
INVX1 exu_U35513(.A(div_z_in[62]), .Y(exu_n14897));
INVX1 exu_U35514(.A(div_z_in[60]), .Y(exu_n14898));
INVX1 exu_U35515(.A(div_z_in[58]), .Y(exu_n14899));
INVX1 exu_U35516(.A(div_z_in[56]), .Y(exu_n14900));
INVX1 exu_U35517(.A(div_z_in[54]), .Y(exu_n14901));
INVX1 exu_U35518(.A(div_z_in[52]), .Y(exu_n14902));
INVX1 exu_U35519(.A(div_z_in[50]), .Y(exu_n14903));
INVX1 exu_U35520(.A(div_z_in[4]), .Y(exu_n14904));
INVX1 exu_U35521(.A(div_z_in[48]), .Y(exu_n14905));
INVX1 exu_U35522(.A(div_z_in[46]), .Y(exu_n14906));
INVX1 exu_U35523(.A(div_z_in[44]), .Y(exu_n14907));
INVX1 exu_U35524(.A(div_z_in[42]), .Y(exu_n14908));
INVX1 exu_U35525(.A(div_z_in[40]), .Y(exu_n14909));
INVX1 exu_U35526(.A(div_z_in[38]), .Y(exu_n14910));
INVX1 exu_U35527(.A(div_z_in[36]), .Y(exu_n14911));
INVX1 exu_U35528(.A(div_z_in[34]), .Y(exu_n14912));
INVX1 exu_U35529(.A(div_z_in[32]), .Y(exu_n14913));
INVX1 exu_U35530(.A(div_z_in[31]), .Y(exu_n14914));
INVX1 exu_U35531(.A(div_z_in[2]), .Y(exu_n14915));
INVX1 exu_U35532(.A(div_z_in[28]), .Y(exu_n14916));
INVX1 exu_U35533(.A(div_z_in[26]), .Y(exu_n14917));
INVX1 exu_U35534(.A(div_z_in[24]), .Y(exu_n14918));
INVX1 exu_U35535(.A(div_z_in[22]), .Y(exu_n14919));
INVX1 exu_U35536(.A(div_z_in[20]), .Y(exu_n14920));
INVX1 exu_U35537(.A(div_z_in[19]), .Y(exu_n14921));
INVX1 exu_U35538(.A(div_z_in[17]), .Y(exu_n14922));
INVX1 exu_U35539(.A(div_z_in[15]), .Y(exu_n14923));
INVX1 exu_U35540(.A(div_z_in[13]), .Y(exu_n14924));
INVX1 exu_U35541(.A(div_z_in[11]), .Y(exu_n14925));
INVX1 exu_U35542(.A(div_z_in[0]), .Y(exu_n14926));
INVX1 exu_U35543(.A(exu_n31621), .Y(exu_n14927));
INVX1 exu_U35544(.A(exu_n31627), .Y(exu_n14928));
INVX1 exu_U35545(.A(exu_n31635), .Y(exu_n14929));
INVX1 exu_U35546(.A(exu_n31641), .Y(exu_n14930));
INVX1 exu_U35547(.A(exu_n31651), .Y(exu_n14931));
INVX1 exu_U35548(.A(exu_n31657), .Y(exu_n14932));
INVX1 exu_U35549(.A(exu_n31665), .Y(exu_n14933));
INVX1 exu_U35550(.A(exu_n31671), .Y(exu_n14934));
INVX1 exu_U35551(.A(exu_n31681), .Y(exu_n14935));
INVX1 exu_U35552(.A(exu_n31687), .Y(exu_n14936));
INVX1 exu_U35553(.A(exu_n31694), .Y(exu_n14937));
INVX1 exu_U35554(.A(exu_n31700), .Y(exu_n14938));
INVX1 exu_U35555(.A(ecl_divcntl_n89), .Y(exu_n14939));
AND2X1 exu_U35556(.A(ecl_divcntl_cntr[1]), .B(ecl_divcntl_cntr[0]), .Y(ecl_divcntl_n89));
AND2X1 exu_U35557(.A(ecl_byplog_rs1_w_comp7_n5), .B(ecl_byplog_rs1_w_comp7_n6), .Y(ecl_byplog_rs1_w_comp7_n4));
INVX1 exu_U35558(.A(ecl_byplog_rs1_w_comp7_n4), .Y(exu_n14940));
AND2X1 exu_U35559(.A(ecl_byplog_rs1_w_comp7_n11), .B(ecl_byplog_rs1_w_comp7_n12), .Y(ecl_byplog_rs1_w_comp7_n10));
INVX1 exu_U35560(.A(ecl_byplog_rs1_w_comp7_n10), .Y(exu_n14941));
AND2X1 exu_U35561(.A(rml_cwp_swap_tid[0]), .B(rml_cwp_swap_tid[1]), .Y(rml_cwp_n48));
INVX1 exu_U35562(.A(rml_cwp_n48), .Y(exu_n14942));
AND2X1 exu_U35563(.A(rml_cwp_swap_tid[1]), .B(exu_n16619), .Y(rml_cwp_n49));
INVX1 exu_U35564(.A(rml_cwp_n49), .Y(exu_n14943));
AND2X1 exu_U35565(.A(rml_cwp_swap_tid[0]), .B(exu_n16620), .Y(rml_cwp_n50));
INVX1 exu_U35566(.A(rml_cwp_n50), .Y(exu_n14944));
AND2X1 exu_U35567(.A(exu_n16619), .B(exu_n16620), .Y(rml_cwp_n51));
INVX1 exu_U35568(.A(rml_cwp_n51), .Y(exu_n14945));
AND2X1 exu_U35569(.A(rml_cwp_n99), .B(rml_cwp_n100), .Y(rml_cwp_n98));
INVX1 exu_U35570(.A(rml_cwp_n98), .Y(exu_n14946));
OR2X1 exu_U35571(.A(rml_ecl_wstate_d[3]), .B(exu_n16572), .Y(rml_wtype_mux_n8));
INVX1 exu_U35572(.A(rml_wtype_mux_n8), .Y(exu_n14947));
OR2X1 exu_U35573(.A(rml_ecl_wstate_d[4]), .B(exu_n16572), .Y(rml_wtype_mux_n10));
INVX1 exu_U35574(.A(rml_wtype_mux_n10), .Y(exu_n14948));
OR2X1 exu_U35575(.A(rml_ecl_wstate_d[5]), .B(exu_n16572), .Y(rml_wtype_mux_n12));
INVX1 exu_U35576(.A(rml_wtype_mux_n12), .Y(exu_n14949));
INVX1 exu_U35577(.A(div_low32or_n6), .Y(exu_n14950));
INVX1 exu_U35578(.A(div_low32or_n12), .Y(exu_n14951));
INVX1 exu_U35579(.A(div_low32or_n20), .Y(exu_n14952));
INVX1 exu_U35580(.A(div_low32or_n26), .Y(exu_n14953));
INVX1 exu_U35581(.A(alu_chk_mem_addr_n2), .Y(exu_n14954));
AND2X1 exu_U35582(.A(alu_chk_mem_addr_n7), .B(alu_chk_mem_addr_n8), .Y(alu_chk_mem_addr_n6));
INVX1 exu_U35583(.A(alu_chk_mem_addr_n6), .Y(exu_n14955));
AND2X1 exu_U35584(.A(alu_chk_mem_addr_n13), .B(alu_chk_mem_addr_n14), .Y(alu_chk_mem_addr_n12));
INVX1 exu_U35585(.A(alu_chk_mem_addr_n12), .Y(exu_n14956));
AND2X1 exu_U35586(.A(alu_chk_mem_addr_n21), .B(alu_chk_mem_addr_n22), .Y(alu_chk_mem_addr_n20));
INVX1 exu_U35587(.A(alu_chk_mem_addr_n20), .Y(exu_n14957));
AND2X1 exu_U35588(.A(alu_chk_mem_addr_n27), .B(alu_chk_mem_addr_n28), .Y(alu_chk_mem_addr_n26));
INVX1 exu_U35589(.A(alu_chk_mem_addr_n26), .Y(exu_n14958));
AND2X1 exu_U35590(.A(mul_exu_ack), .B(ecl_mdqctl_n22), .Y(ecl_mdqctl_n25));
INVX1 exu_U35591(.A(ecl_mdqctl_n25), .Y(exu_n14959));
INVX1 exu_U35592(.A(ecl_divcntl_n54), .Y(exu_n14960));
AND2X1 exu_U35593(.A(exu_n15206), .B(exu_n15204), .Y(ecl_divcntl_n54));
AND2X1 exu_U35594(.A(exu_n15471), .B(ecl_divcntl_div_state_1), .Y(ecl_divcntl_n29));
INVX1 exu_U35595(.A(ecl_divcntl_n29), .Y(exu_n14961));
AND2X1 exu_U35596(.A(ecl_wb_e), .B(ecl_restore_e), .Y(ecl_writeback_n60));
INVX1 exu_U35597(.A(ecl_writeback_n60), .Y(exu_n14962));
AND2X1 exu_U35598(.A(ecl_wb_e), .B(exu_n16598), .Y(ecl_writeback_n64));
INVX1 exu_U35599(.A(ecl_writeback_n64), .Y(exu_n14963));
OR2X1 exu_U35600(.A(exu_n15768), .B(exu_n14965), .Y(ecl_writeback_n94));
INVX1 exu_U35601(.A(ecl_writeback_n94), .Y(exu_n14964));
AND2X1 exu_U35602(.A(exu_n15742), .B(exu_n15739), .Y(ecl_writeback_n96));
INVX1 exu_U35603(.A(ecl_writeback_n96), .Y(exu_n14965));
OR2X1 exu_U35604(.A(exu_n15742), .B(exu_n14967), .Y(ecl_writeback_n105));
INVX1 exu_U35605(.A(ecl_writeback_n105), .Y(exu_n14966));
AND2X1 exu_U35606(.A(ecl_mdqctl_n63), .B(exu_n15739), .Y(ecl_writeback_n106));
INVX1 exu_U35607(.A(ecl_writeback_n106), .Y(exu_n14967));
OR2X1 exu_U35608(.A(exu_n15739), .B(exu_n14969), .Y(ecl_writeback_n113));
INVX1 exu_U35609(.A(ecl_writeback_n113), .Y(exu_n14968));
AND2X1 exu_U35610(.A(ecl_mdqctl_n63), .B(exu_n15742), .Y(ecl_writeback_n114));
INVX1 exu_U35611(.A(ecl_writeback_n114), .Y(exu_n14969));
OR2X1 exu_U35612(.A(exu_n15739), .B(ecl_writeback_n121), .Y(ecl_writeback_n120));
INVX1 exu_U35613(.A(ecl_writeback_n120), .Y(exu_n14970));
AND2X1 exu_U35614(.A(ecl_writeback_sraddr_w[1]), .B(exu_n16553), .Y(ecl_writeback_n132));
INVX1 exu_U35615(.A(ecl_writeback_n132), .Y(exu_n14971));
AND2X1 exu_U35616(.A(exu_n16553), .B(exu_n16554), .Y(ecl_writeback_n140));
INVX1 exu_U35617(.A(ecl_writeback_n140), .Y(exu_n14972));
OR2X1 exu_U35618(.A(ecl_writeback_n157), .B(exu_n14974), .Y(ecl_writeback_n156));
INVX1 exu_U35619(.A(ecl_writeback_n156), .Y(exu_n14973));
AND2X1 exu_U35620(.A(ecl_writeback_n159), .B(ecl_flush_w1), .Y(ecl_writeback_n158));
INVX1 exu_U35621(.A(ecl_writeback_n158), .Y(exu_n14974));
AND2X1 exu_U35622(.A(ifu_exu_inst_vld_w), .B(exu_n15414), .Y(ecl_ccr_n23));
INVX1 exu_U35623(.A(ecl_ccr_n23), .Y(exu_n14975));
OR2X1 exu_U35624(.A(rml_win_trap_w), .B(exu_n16608), .Y(rml_n108));
INVX1 exu_U35625(.A(rml_n108), .Y(exu_n14976));
AND2X1 exu_U35626(.A(rml_save_e), .B(rml_exu_tlu_spill_e), .Y(rml_n118));
INVX1 exu_U35627(.A(rml_n118), .Y(exu_n14977));
INVX1 exu_U35628(.A(div_n42), .Y(exu_n14978));
INVX1 exu_U35629(.A(div_n48), .Y(exu_n14979));
INVX1 exu_U35630(.A(div_n56), .Y(exu_n14980));
INVX1 exu_U35631(.A(div_n62), .Y(exu_n14981));
INVX1 exu_U35632(.A(div_n72), .Y(exu_n14982));
INVX1 exu_U35633(.A(div_n78), .Y(exu_n14983));
INVX1 exu_U35634(.A(div_n86), .Y(exu_n14984));
INVX1 exu_U35635(.A(div_n92), .Y(exu_n14985));
INVX1 exu_U35636(.A(alu_n74), .Y(exu_n14986));
INVX1 exu_U35637(.A(alu_n80), .Y(exu_n14987));
INVX1 exu_U35638(.A(alu_n88), .Y(exu_n14988));
INVX1 exu_U35639(.A(alu_n94), .Y(exu_n14989));
INVX1 exu_U35640(.A(alu_n100), .Y(exu_n14990));
INVX1 exu_U35641(.A(alu_n104), .Y(exu_n14991));
INVX1 exu_U35642(.A(alu_n110), .Y(exu_n14992));
INVX1 exu_U35643(.A(alu_n118), .Y(exu_n14993));
INVX1 exu_U35644(.A(alu_n124), .Y(exu_n14994));
OR2X1 exu_U35645(.A(ecl_n91), .B(exu_n14996), .Y(ecl_n90));
INVX1 exu_U35646(.A(ecl_n90), .Y(exu_n14995));
INVX1 exu_U35647(.A(ecl_n92), .Y(exu_n14996));
OR2X1 exu_U35648(.A(exu_n16512), .B(ecl_n143), .Y(ecl_n142));
INVX1 exu_U35649(.A(ecl_n142), .Y(exu_n14997));
AND2X1 exu_U35650(.A(rml_cwp_next_slot1_state[1]), .B(exu_n15941), .Y(exu_n17460));
AND2X1 exu_U35651(.A(rml_cwp_next_slot1_state[0]), .B(exu_n15941), .Y(exu_n17461));
AND2X1 exu_U35652(.A(rml_cwp_next_slot2_state[1]), .B(exu_n15942), .Y(exu_n17475));
AND2X1 exu_U35653(.A(rml_cwp_next_slot2_state[0]), .B(exu_n15942), .Y(exu_n17477));
AND2X1 exu_U35654(.A(rml_cwp_next_slot3_state[1]), .B(exu_n15943), .Y(exu_n17491));
AND2X1 exu_U35655(.A(rml_cwp_next_slot3_state[0]), .B(exu_n15943), .Y(exu_n17492));
AND2X1 exu_U35656(.A(ecl_divcntl_cnt6_next_cntr[1]), .B(exu_n17619), .Y(exu_n17624));
AND2X1 exu_U35657(.A(ecl_divcntl_cnt6_n30), .B(exu_n17619), .Y(exu_n17625));
AND2X1 exu_U35658(.A(rml_ecl_wstate_d[5]), .B(exu_n15824), .Y(exu_n18013));
AND2X1 exu_U35659(.A(exu_ifu_cc_d[5]), .B(exu_n16373), .Y(exu_n18014));
AND2X1 exu_U35660(.A(rml_ecl_wstate_d[4]), .B(exu_n15824), .Y(exu_n18015));
AND2X1 exu_U35661(.A(exu_ifu_cc_d[4]), .B(exu_n16373), .Y(exu_n18016));
AND2X1 exu_U35662(.A(rml_ecl_wstate_d[3]), .B(exu_n15824), .Y(exu_n18017));
AND2X1 exu_U35663(.A(exu_ifu_cc_d[3]), .B(exu_n16373), .Y(exu_n18018));
AND2X1 exu_U35664(.A(rml_cwp_next_swap_thr[3]), .B(exu_n18407), .Y(exu_n18408));
AND2X1 exu_U35665(.A(rml_cwp_next_swap_thr[2]), .B(exu_n18407), .Y(exu_n18409));
AND2X1 exu_U35666(.A(rml_cwp_next_swap_thr[1]), .B(exu_n18407), .Y(exu_n18410));
AND2X1 exu_U35667(.A(exu_n15234), .B(exu_n18407), .Y(exu_n18411));
AND2X1 exu_U35668(.A(rml_cwp_cwp_cmplt_next), .B(exu_n18417), .Y(exu_n18418));
AND2X1 exu_U35669(.A(rml_cwp_swap_tid[1]), .B(exu_n18417), .Y(exu_n18419));
AND2X1 exu_U35670(.A(rml_cwp_swap_tid[0]), .B(exu_n18417), .Y(exu_n18420));
AND2X1 exu_U35671(.A(rml_cwp_swap_data_12), .B(exu_n18417), .Y(exu_n18421));
AND2X1 exu_U35672(.A(ecl_dff_sel_sum_d2e_din[0]), .B(exu_n19255), .Y(exu_n19256));
AND2X1 exu_U35673(.A(ifu_exu_tv_d), .B(exu_n19257), .Y(exu_n19258));
AND2X1 exu_U35674(.A(ifu_exu_tagop_d), .B(exu_n19259), .Y(exu_n19260));
AND2X1 exu_U35675(.A(ifu_exu_ialign_d), .B(exu_n19261), .Y(exu_n19262));
AND2X1 exu_U35676(.A(ecl_ialign_e), .B(exu_n19263), .Y(exu_n19264));
AND2X1 exu_U35677(.A(lsu_exu_ldxa_m), .B(exu_n19265), .Y(exu_n19266));
AND2X1 exu_U35678(.A(ifu_exu_sethi_inst_d), .B(exu_n19267), .Y(exu_n19268));
AND2X1 exu_U35679(.A(ifu_exu_rs1_vld_d), .B(exu_n19269), .Y(exu_n19270));
AND2X1 exu_U35680(.A(ifu_exu_rs2_vld_d), .B(exu_n19271), .Y(exu_n19272));
AND2X1 exu_U35681(.A(ecl_rs3_vld_d), .B(exu_n19273), .Y(exu_n19274));
AND2X1 exu_U35682(.A(ifu_exu_casa_d), .B(exu_n19275), .Y(exu_n19276));
AND2X1 exu_U35683(.A(ifu_exu_invert_d), .B(exu_n19279), .Y(exu_n19280));
INVX1 exu_U35684(.A(exu_n19280), .Y(exu_n14998));
INVX1 exu_U35685(.A(exu_n14998), .Y(exu_n16320));
AND2X1 exu_U35686(.A(ecl_c_used_dff_din[0]), .B(exu_n19281), .Y(exu_n19282));
AND2X1 exu_U35687(.A(ifu_exu_muls_d), .B(exu_n19283), .Y(exu_n19284));
AND2X1 exu_U35688(.A(ecl_div_muls_rs1_31_e_l), .B(exu_n19287), .Y(exu_n19288));
AND2X1 exu_U35689(.A(div_input_data_e[95]), .B(exu_n19289), .Y(exu_n19290));
AND2X1 exu_U35690(.A(ifu_exu_save_d), .B(exu_n19291), .Y(exu_n19292));
AND2X1 exu_U35691(.A(ifu_exu_restore_d), .B(exu_n19293), .Y(exu_n19294));
AND2X1 exu_U35692(.A(ifu_exu_addr_mask_d), .B(exu_n19295), .Y(exu_n19296));
AND2X1 exu_U35693(.A(ecl_misalign_addr_e), .B(exu_n19299), .Y(exu_n19300));
AND2X1 exu_U35694(.A(ifu_exu_range_check_jlret_d), .B(exu_n19301), .Y(exu_n19302));
AND2X1 exu_U35695(.A(ifu_exu_range_check_other_d), .B(exu_n19305), .Y(exu_n19306));
AND2X1 exu_U35696(.A(ecl_ifu_exu_range_check_other_e), .B(exu_n19307), .Y(exu_n19308));
AND2X1 exu_U35697(.A(ifu_exu_inst_vld_w), .B(exu_n19309), .Y(exu_n19310));
AND2X1 exu_U35698(.A(tlu_exu_priv_trap_m), .B(exu_n19311), .Y(exu_n19312));
AND2X1 exu_U35699(.A(ifu_tlu_flush_m), .B(exu_n19315), .Y(exu_n19316));
AND2X1 exu_U35700(.A(ecl_flush_w), .B(exu_n19317), .Y(exu_n19318));
AND2X1 exu_U35701(.A(ecl_std_d), .B(exu_n19323), .Y(exu_n19324));
AND2X1 exu_U35702(.A(ecl_early_ttype_vld_e), .B(exu_n19325), .Y(exu_n19326));
AND2X1 exu_U35703(.A(exu_n15030), .B(exu_n19327), .Y(exu_n19328));
AND2X1 exu_U35704(.A(ifu_exu_invert_d), .B(exu_n19337), .Y(exu_n19338));
INVX1 exu_U35705(.A(exu_n19338), .Y(exu_n14999));
INVX1 exu_U35706(.A(exu_n14999), .Y(exu_n16321));
AND2X1 exu_U35707(.A(rml_save_e), .B(exu_n19339), .Y(exu_n19340));
AND2X1 exu_U35708(.A(rml_win_trap_e), .B(exu_n19341), .Y(exu_n19342));
AND2X1 exu_U35709(.A(rml_win_trap_m), .B(exu_n19343), .Y(exu_n19344));
AND2X1 exu_U35710(.A(exu_n15940), .B(exu_n19345), .Y(exu_n19346));
AND2X1 exu_U35711(.A(rml_rml_ecl_kill_e), .B(exu_n19347), .Y(exu_n19348));
AND2X1 exu_U35712(.A(rml_rml_ecl_other_d), .B(exu_n19349), .Y(exu_n19350));
AND2X1 exu_U35713(.A(exu_n15346), .B(exu_n19351), .Y(exu_n19352));
AND2X1 exu_U35714(.A(rml_did_restore_m), .B(exu_n19353), .Y(exu_n19354));
AND2X1 exu_U35715(.A(rml_rml_cwp_wen_m), .B(exu_n19359), .Y(exu_n19360));
AND2X1 exu_U35716(.A(rml_cansave_wen_e), .B(exu_n19361), .Y(exu_n19362));
AND2X1 exu_U35717(.A(rml_cansave_wen_m), .B(exu_n19363), .Y(exu_n19364));
AND2X1 exu_U35718(.A(rml_canrestore_wen_e), .B(exu_n19365), .Y(exu_n19366));
AND2X1 exu_U35719(.A(rml_canrestore_wen_m), .B(exu_n19367), .Y(exu_n19368));
AND2X1 exu_U35720(.A(rml_n130), .B(exu_n19369), .Y(exu_n19370));
AND2X1 exu_U35721(.A(rml_otherwin_wen_m), .B(exu_n19371), .Y(exu_n19372));
AND2X1 exu_U35722(.A(rml_n131), .B(exu_n19373), .Y(exu_n19374));
AND2X1 exu_U35723(.A(rml_cleanwin_wen_m), .B(exu_n19375), .Y(exu_n19376));
AND2X1 exu_U35724(.A(exu_n15335), .B(exu_n19377), .Y(exu_n19378));
AND2X1 exu_U35725(.A(exu_n15336), .B(exu_n19379), .Y(exu_n19380));
AND2X1 exu_U35726(.A(bypass_w1_eccgen_p0_g[7]), .B(exu_n19381), .Y(exu_n19382));
AND2X1 exu_U35727(.A(bypass_w1_eccgen_p0_g[6]), .B(exu_n19383), .Y(exu_n19384));
AND2X1 exu_U35728(.A(bypass_w1_eccgen_p0_g[5]), .B(exu_n19385), .Y(exu_n19386));
AND2X1 exu_U35729(.A(bypass_w1_eccgen_p0_g[4]), .B(exu_n19387), .Y(exu_n19388));
AND2X1 exu_U35730(.A(bypass_w1_eccgen_p0_g[3]), .B(exu_n19389), .Y(exu_n19390));
AND2X1 exu_U35731(.A(bypass_w1_eccgen_p0_g[2]), .B(exu_n19391), .Y(exu_n19392));
AND2X1 exu_U35732(.A(bypass_w1_eccgen_p0_g[1]), .B(exu_n19393), .Y(exu_n19394));
AND2X1 exu_U35733(.A(bypass_w1_eccgen_p0_g[0]), .B(exu_n19395), .Y(exu_n19396));
AND2X1 exu_U35734(.A(bypass_w1_eccgen_p1_g[7]), .B(exu_n19397), .Y(exu_n19398));
AND2X1 exu_U35735(.A(bypass_w1_eccgen_p1_g[6]), .B(exu_n19399), .Y(exu_n19400));
AND2X1 exu_U35736(.A(bypass_w1_eccgen_p1_g[5]), .B(exu_n19401), .Y(exu_n19402));
AND2X1 exu_U35737(.A(bypass_w1_eccgen_p1_g[4]), .B(exu_n19403), .Y(exu_n19404));
AND2X1 exu_U35738(.A(bypass_w1_eccgen_p1_g[3]), .B(exu_n19405), .Y(exu_n19406));
AND2X1 exu_U35739(.A(bypass_w1_eccgen_p1_g[2]), .B(exu_n19407), .Y(exu_n19408));
AND2X1 exu_U35740(.A(bypass_w1_eccgen_p1_g[1]), .B(exu_n19409), .Y(exu_n19410));
AND2X1 exu_U35741(.A(bypass_w1_eccgen_p1_g[0]), .B(exu_n19411), .Y(exu_n19412));
AND2X1 exu_U35742(.A(bypass_w1_eccgen_p2_g[7]), .B(exu_n19413), .Y(exu_n19414));
AND2X1 exu_U35743(.A(bypass_w1_eccgen_p2_g[6]), .B(exu_n19415), .Y(exu_n19416));
AND2X1 exu_U35744(.A(bypass_w1_eccgen_p2_g[5]), .B(exu_n19417), .Y(exu_n19418));
AND2X1 exu_U35745(.A(bypass_w1_eccgen_p2_g[4]), .B(exu_n19419), .Y(exu_n19420));
AND2X1 exu_U35746(.A(bypass_w1_eccgen_p2_g[3]), .B(exu_n19421), .Y(exu_n19422));
AND2X1 exu_U35747(.A(bypass_w1_eccgen_p2_g[2]), .B(exu_n19423), .Y(exu_n19424));
AND2X1 exu_U35748(.A(bypass_w1_eccgen_p2_g[1]), .B(exu_n19425), .Y(exu_n19426));
AND2X1 exu_U35749(.A(bypass_w1_eccgen_p2_g[0]), .B(exu_n19427), .Y(exu_n19428));
AND2X1 exu_U35750(.A(bypass_w1_eccgen_p3_g[7]), .B(exu_n19429), .Y(exu_n19430));
AND2X1 exu_U35751(.A(bypass_w1_eccgen_p3_g[6]), .B(exu_n19431), .Y(exu_n19432));
AND2X1 exu_U35752(.A(bypass_w1_eccgen_p3_g[5]), .B(exu_n19433), .Y(exu_n19434));
AND2X1 exu_U35753(.A(bypass_w1_eccgen_p3_g[4]), .B(exu_n19435), .Y(exu_n19436));
AND2X1 exu_U35754(.A(bypass_w1_eccgen_p3_g[3]), .B(exu_n19437), .Y(exu_n19438));
AND2X1 exu_U35755(.A(bypass_w1_eccgen_p3_g[2]), .B(exu_n19439), .Y(exu_n19440));
AND2X1 exu_U35756(.A(bypass_w1_eccgen_p3_g[1]), .B(exu_n19441), .Y(exu_n19442));
AND2X1 exu_U35757(.A(bypass_w1_eccgen_p3_g[0]), .B(exu_n19443), .Y(exu_n19444));
AND2X1 exu_U35758(.A(bypass_w1_eccgen_p4_g[3]), .B(exu_n19445), .Y(exu_n19446));
AND2X1 exu_U35759(.A(bypass_w1_eccgen_p4_g[2]), .B(exu_n19447), .Y(exu_n19448));
AND2X1 exu_U35760(.A(bypass_w1_eccgen_p4_g[1]), .B(exu_n19449), .Y(exu_n19450));
AND2X1 exu_U35761(.A(bypass_w1_eccgen_p4_g[0]), .B(exu_n19451), .Y(exu_n19452));
AND2X1 exu_U35762(.A(bypass_w1_eccgen_p5_g[1]), .B(exu_n19453), .Y(exu_n19454));
AND2X1 exu_U35763(.A(bypass_w1_eccgen_p5_g[0]), .B(exu_n19455), .Y(exu_n19456));
AND2X1 exu_U35764(.A(bypass_w1_eccgen_p6_g[1]), .B(exu_n19457), .Y(exu_n19458));
AND2X1 exu_U35765(.A(bypass_w1_eccgen_p6_g[0]), .B(exu_n19459), .Y(exu_n19460));
AND2X1 exu_U35766(.A(bypass_w1_eccgen_p7_g[7]), .B(exu_n19461), .Y(exu_n19462));
AND2X1 exu_U35767(.A(bypass_w1_eccgen_p7_g[6]), .B(exu_n19463), .Y(exu_n19464));
AND2X1 exu_U35768(.A(bypass_w1_eccgen_p7_g[5]), .B(exu_n19465), .Y(exu_n19466));
AND2X1 exu_U35769(.A(bypass_w1_eccgen_p7_g[4]), .B(exu_n19467), .Y(exu_n19468));
AND2X1 exu_U35770(.A(bypass_w1_eccgen_p7_g[3]), .B(exu_n19469), .Y(exu_n19470));
AND2X1 exu_U35771(.A(bypass_w1_eccgen_p7_g[2]), .B(exu_n19471), .Y(exu_n19472));
AND2X1 exu_U35772(.A(bypass_w1_eccgen_p7_g[1]), .B(exu_n19473), .Y(exu_n19474));
AND2X1 exu_U35773(.A(bypass_w1_eccgen_p7_g[0]), .B(exu_n19475), .Y(exu_n19476));
AND2X1 exu_U35774(.A(bypass_w2_eccgen_p0_g[7]), .B(exu_n19477), .Y(exu_n19478));
AND2X1 exu_U35775(.A(bypass_w2_eccgen_p0_g[6]), .B(exu_n19479), .Y(exu_n19480));
AND2X1 exu_U35776(.A(bypass_w2_eccgen_p0_g[5]), .B(exu_n19481), .Y(exu_n19482));
AND2X1 exu_U35777(.A(bypass_w2_eccgen_p0_g[4]), .B(exu_n19483), .Y(exu_n19484));
AND2X1 exu_U35778(.A(bypass_w2_eccgen_p0_g[3]), .B(exu_n19485), .Y(exu_n19486));
AND2X1 exu_U35779(.A(bypass_w2_eccgen_p0_g[2]), .B(exu_n19487), .Y(exu_n19488));
AND2X1 exu_U35780(.A(bypass_w2_eccgen_p0_g[1]), .B(exu_n19489), .Y(exu_n19490));
AND2X1 exu_U35781(.A(bypass_w2_eccgen_p0_g[0]), .B(exu_n19491), .Y(exu_n19492));
AND2X1 exu_U35782(.A(bypass_w2_eccgen_p1_g[7]), .B(exu_n19493), .Y(exu_n19494));
AND2X1 exu_U35783(.A(bypass_w2_eccgen_p1_g[6]), .B(exu_n19495), .Y(exu_n19496));
AND2X1 exu_U35784(.A(bypass_w2_eccgen_p1_g[5]), .B(exu_n19497), .Y(exu_n19498));
AND2X1 exu_U35785(.A(bypass_w2_eccgen_p1_g[4]), .B(exu_n19499), .Y(exu_n19500));
AND2X1 exu_U35786(.A(bypass_w2_eccgen_p1_g[3]), .B(exu_n19501), .Y(exu_n19502));
AND2X1 exu_U35787(.A(bypass_w2_eccgen_p1_g[2]), .B(exu_n19503), .Y(exu_n19504));
AND2X1 exu_U35788(.A(bypass_w2_eccgen_p1_g[1]), .B(exu_n19505), .Y(exu_n19506));
AND2X1 exu_U35789(.A(bypass_w2_eccgen_p1_g[0]), .B(exu_n19507), .Y(exu_n19508));
AND2X1 exu_U35790(.A(bypass_w2_eccgen_p2_g[7]), .B(exu_n19509), .Y(exu_n19510));
AND2X1 exu_U35791(.A(bypass_w2_eccgen_p2_g[6]), .B(exu_n19511), .Y(exu_n19512));
AND2X1 exu_U35792(.A(bypass_w2_eccgen_p2_g[5]), .B(exu_n19513), .Y(exu_n19514));
AND2X1 exu_U35793(.A(bypass_w2_eccgen_p2_g[4]), .B(exu_n19515), .Y(exu_n19516));
AND2X1 exu_U35794(.A(bypass_w2_eccgen_p2_g[3]), .B(exu_n19517), .Y(exu_n19518));
AND2X1 exu_U35795(.A(bypass_w2_eccgen_p2_g[2]), .B(exu_n19519), .Y(exu_n19520));
AND2X1 exu_U35796(.A(bypass_w2_eccgen_p2_g[1]), .B(exu_n19521), .Y(exu_n19522));
AND2X1 exu_U35797(.A(bypass_w2_eccgen_p2_g[0]), .B(exu_n19523), .Y(exu_n19524));
AND2X1 exu_U35798(.A(bypass_w2_eccgen_p3_g[7]), .B(exu_n19525), .Y(exu_n19526));
AND2X1 exu_U35799(.A(bypass_w2_eccgen_p3_g[6]), .B(exu_n19527), .Y(exu_n19528));
AND2X1 exu_U35800(.A(bypass_w2_eccgen_p3_g[5]), .B(exu_n19529), .Y(exu_n19530));
AND2X1 exu_U35801(.A(bypass_w2_eccgen_p3_g[4]), .B(exu_n19531), .Y(exu_n19532));
AND2X1 exu_U35802(.A(bypass_w2_eccgen_p3_g[3]), .B(exu_n19533), .Y(exu_n19534));
AND2X1 exu_U35803(.A(bypass_w2_eccgen_p3_g[2]), .B(exu_n19535), .Y(exu_n19536));
AND2X1 exu_U35804(.A(bypass_w2_eccgen_p3_g[1]), .B(exu_n19537), .Y(exu_n19538));
AND2X1 exu_U35805(.A(bypass_w2_eccgen_p3_g[0]), .B(exu_n19539), .Y(exu_n19540));
AND2X1 exu_U35806(.A(bypass_w2_eccgen_p4_g[3]), .B(exu_n19541), .Y(exu_n19542));
AND2X1 exu_U35807(.A(bypass_w2_eccgen_p4_g[2]), .B(exu_n19543), .Y(exu_n19544));
AND2X1 exu_U35808(.A(bypass_w2_eccgen_p4_g[1]), .B(exu_n19545), .Y(exu_n19546));
AND2X1 exu_U35809(.A(bypass_w2_eccgen_p4_g[0]), .B(exu_n19547), .Y(exu_n19548));
AND2X1 exu_U35810(.A(bypass_w2_eccgen_p5_g[1]), .B(exu_n19549), .Y(exu_n19550));
AND2X1 exu_U35811(.A(bypass_w2_eccgen_p5_g[0]), .B(exu_n19551), .Y(exu_n19552));
AND2X1 exu_U35812(.A(bypass_w2_eccgen_p6_g[1]), .B(exu_n19553), .Y(exu_n19554));
AND2X1 exu_U35813(.A(bypass_w2_eccgen_p6_g[0]), .B(exu_n19555), .Y(exu_n19556));
AND2X1 exu_U35814(.A(bypass_w2_eccgen_p7_g[7]), .B(exu_n19557), .Y(exu_n19558));
AND2X1 exu_U35815(.A(bypass_w2_eccgen_p7_g[6]), .B(exu_n19559), .Y(exu_n19560));
AND2X1 exu_U35816(.A(bypass_w2_eccgen_p7_g[5]), .B(exu_n19561), .Y(exu_n19562));
AND2X1 exu_U35817(.A(bypass_w2_eccgen_p7_g[4]), .B(exu_n19563), .Y(exu_n19564));
AND2X1 exu_U35818(.A(bypass_w2_eccgen_p7_g[3]), .B(exu_n19565), .Y(exu_n19566));
AND2X1 exu_U35819(.A(bypass_w2_eccgen_p7_g[2]), .B(exu_n19567), .Y(exu_n19568));
AND2X1 exu_U35820(.A(bypass_w2_eccgen_p7_g[1]), .B(exu_n19569), .Y(exu_n19570));
AND2X1 exu_U35821(.A(bypass_w2_eccgen_p7_g[0]), .B(exu_n19571), .Y(exu_n19572));
AND2X1 exu_U35822(.A(ifu_exu_setcc_d), .B(exu_n19573), .Y(exu_n19574));
AND2X1 exu_U35823(.A(exu_n15235), .B(exu_n19575), .Y(exu_n19576));
AND2X1 exu_U35824(.A(ecl_ccr_valid_setcc_m), .B(exu_n19577), .Y(exu_n19578));
AND2X1 exu_U35825(.A(ecl_writeback_ld_g), .B(exu_n19579), .Y(exu_n19580));
AND2X1 exu_U35826(.A(ifu_exu_wen_d), .B(exu_n19587), .Y(exu_n19588));
AND2X1 exu_U35827(.A(ifu_tlu_wsr_inst_d), .B(exu_n19591), .Y(exu_n19592));
AND2X1 exu_U35828(.A(exu_ffu_wsr_inst_e), .B(exu_n19593), .Y(exu_n19594));
AND2X1 exu_U35829(.A(ecl_writeback_wrsr_m), .B(exu_n19595), .Y(exu_n19596));
AND2X1 exu_U35830(.A(ecl_writeback_yreg_wen_w), .B(exu_n19597), .Y(exu_n19598));
AND2X1 exu_U35831(.A(ifu_exu_return_d), .B(exu_n19599), .Y(exu_n19600));
AND2X1 exu_U35832(.A(ecl_byp_restore_m), .B(exu_n19603), .Y(exu_n19604));
AND2X1 exu_U35833(.A(ecl_writeback_short_longop_done_e), .B(exu_n19607), .Y(exu_n19608));
AND2X1 exu_U35834(.A(exu_n16305), .B(exu_n19609), .Y(exu_n19610));
AND2X1 exu_U35835(.A(ecl_byp_rs2_mux2_sel_rf), .B(exu_n19611), .Y(exu_n19612));
AND2X1 exu_U35836(.A(exu_n16004), .B(exu_n19613), .Y(exu_n19614));
AND2X1 exu_U35837(.A(ifu_exu_nceen_e), .B(exu_n19619), .Y(exu_n19620));
AND2X1 exu_U35838(.A(ecc_ecl_rs1_ce), .B(exu_n19621), .Y(exu_n19622));
AND2X1 exu_U35839(.A(ecl_eccctl_sel_rs2_e), .B(exu_n19623), .Y(exu_n19624));
AND2X1 exu_U35840(.A(exu_n15205), .B(exu_n19625), .Y(exu_n19626));
AND2X1 exu_U35841(.A(ecl_eccctl_inj_irferr_m), .B(exu_n19627), .Y(exu_n19628));
AND2X1 exu_U35842(.A(ecc_ecl_rs1_ue), .B(exu_n19629), .Y(exu_n19630));
AND2X1 exu_U35843(.A(ecc_ecl_rs2_ue), .B(exu_n19631), .Y(exu_n19632));
AND2X1 exu_U35844(.A(ecc_ecl_rs2_ce), .B(exu_n19633), .Y(exu_n19634));
AND2X1 exu_U35845(.A(ecl_eccctl_n14), .B(exu_n19635), .Y(exu_n19636));
AND2X1 exu_U35846(.A(ecl_divcntl_n23), .B(exu_n19640), .Y(exu_n19641));
AND2X1 exu_U35847(.A(ecl_mdqctl_new_div_vld), .B(exu_n19650), .Y(exu_n19651));
AND2X1 exu_U35848(.A(ecl_mdqctl_isdiv_e_valid), .B(exu_n19652), .Y(exu_n19653));
AND2X1 exu_U35849(.A(ecl_mdqctl_isdiv_m_valid), .B(exu_n19654), .Y(exu_n19655));
AND2X1 exu_U35850(.A(ifu_exu_muldivop_d[4]), .B(exu_n19656), .Y(exu_n19657));
AND2X1 exu_U35851(.A(ecl_mdqctl_n16), .B(exu_n19281), .Y(exu_n19658));
AND2X1 exu_U35852(.A(ecl_mdqctl_ismul_m_valid), .B(exu_n19279), .Y(exu_n19659));
AND2X1 exu_U35853(.A(ecl_mdqctl_mul_done_valid_c0), .B(exu_n19271), .Y(exu_n19662));
AND2X1 exu_U35854(.A(ecl_mdqctl_mul_done_valid_c1), .B(exu_n19269), .Y(exu_n19663));
AND2X1 exu_U35855(.A(ecl_mdqctl_mul_done_c2), .B(exu_n19267), .Y(exu_n19664));
AND2X1 exu_U35856(.A(ecl_mdqctl_mul_done_c3), .B(exu_n19265), .Y(exu_n19665));
AND2X1 exu_U35857(.A(ecl_mdqctl_next_mul_done), .B(exu_n19263), .Y(exu_n19666));
AND2X1 exu_U35858(.A(exu_n15925), .B(exu_n19261), .Y(exu_n19667));
AND2X1 exu_U35859(.A(rml_cwp_full_swap_m), .B(exu_n19259), .Y(exu_n19668));
AND2X1 exu_U35860(.A(ecl_shiftop_d[2]), .B(exu_n19670), .Y(exu_n19671));
AND2X1 exu_U35861(.A(ecl_shiftop_d[1]), .B(exu_n19670), .Y(exu_n19672));
AND2X1 exu_U35862(.A(ecl_shiftop_d[0]), .B(exu_n19670), .Y(exu_n19673));
AND2X1 exu_U35863(.A(exu_n15851), .B(exu_n19678), .Y(exu_n19679));
AND2X1 exu_U35864(.A(exu_n15852), .B(exu_n19678), .Y(exu_n19680));
AND2X1 exu_U35865(.A(exu_n15853), .B(exu_n19678), .Y(exu_n19681));
AND2X1 exu_U35866(.A(rml_next_cwp_m[2]), .B(exu_n19682), .Y(exu_n19683));
AND2X1 exu_U35867(.A(rml_next_cwp_m[1]), .B(exu_n19682), .Y(exu_n19684));
AND2X1 exu_U35868(.A(rml_next_cwp_m[0]), .B(exu_n19682), .Y(exu_n19685));
AND2X1 exu_U35869(.A(rml_next_cansave_m[2]), .B(exu_n19690), .Y(exu_n19691));
AND2X1 exu_U35870(.A(rml_next_cansave_m[1]), .B(exu_n19690), .Y(exu_n19692));
AND2X1 exu_U35871(.A(rml_next_cansave_m[0]), .B(exu_n19690), .Y(exu_n19693));
AND2X1 exu_U35872(.A(rml_next_canrestore_m[2]), .B(exu_n19698), .Y(exu_n19699));
AND2X1 exu_U35873(.A(rml_next_canrestore_m[1]), .B(exu_n19698), .Y(exu_n19700));
AND2X1 exu_U35874(.A(rml_next_canrestore_m[0]), .B(exu_n19698), .Y(exu_n19701));
AND2X1 exu_U35875(.A(rml_next_otherwin_m[2]), .B(exu_n19706), .Y(exu_n19707));
AND2X1 exu_U35876(.A(rml_next_otherwin_m[1]), .B(exu_n19706), .Y(exu_n19708));
AND2X1 exu_U35877(.A(rml_next_otherwin_m[0]), .B(exu_n19706), .Y(exu_n19709));
AND2X1 exu_U35878(.A(rml_next_cleanwin_m[2]), .B(exu_n19714), .Y(exu_n19715));
AND2X1 exu_U35879(.A(rml_next_cleanwin_m[1]), .B(exu_n19714), .Y(exu_n19716));
AND2X1 exu_U35880(.A(rml_next_cleanwin_m[0]), .B(exu_n19714), .Y(exu_n19717));
AND2X1 exu_U35881(.A(rml_ecl_cansave_d[2]), .B(exu_n19718), .Y(exu_n19719));
AND2X1 exu_U35882(.A(rml_ecl_cansave_d[1]), .B(exu_n19718), .Y(exu_n19720));
AND2X1 exu_U35883(.A(rml_ecl_cansave_d[0]), .B(exu_n19718), .Y(exu_n19721));
AND2X1 exu_U35884(.A(rml_ecl_canrestore_d[2]), .B(exu_n19722), .Y(exu_n19723));
AND2X1 exu_U35885(.A(rml_ecl_canrestore_d[1]), .B(exu_n19722), .Y(exu_n19724));
AND2X1 exu_U35886(.A(rml_ecl_canrestore_d[0]), .B(exu_n19722), .Y(exu_n19725));
AND2X1 exu_U35887(.A(rml_ecl_otherwin_d[2]), .B(exu_n19726), .Y(exu_n19727));
AND2X1 exu_U35888(.A(rml_ecl_otherwin_d[1]), .B(exu_n19726), .Y(exu_n19728));
AND2X1 exu_U35889(.A(rml_ecl_otherwin_d[0]), .B(exu_n19726), .Y(exu_n19729));
AND2X1 exu_U35890(.A(rml_ecl_cleanwin_d[2]), .B(exu_n19730), .Y(exu_n19731));
AND2X1 exu_U35891(.A(rml_ecl_cleanwin_d[1]), .B(exu_n19730), .Y(exu_n19732));
AND2X1 exu_U35892(.A(rml_ecl_cleanwin_d[0]), .B(exu_n19730), .Y(exu_n19733));
AND2X1 exu_U35893(.A(ecl_wb_ccr_setcc_g), .B(exu_n19734), .Y(exu_n19735));
AND2X1 exu_U35894(.A(ecl_irf_tid_g[1]), .B(exu_n19734), .Y(exu_n19736));
AND2X1 exu_U35895(.A(ecl_irf_tid_g[0]), .B(exu_n19734), .Y(exu_n19737));
AND2X1 exu_U35896(.A(rml_ecl_cwp_d[2]), .B(exu_n19738), .Y(exu_n19739));
AND2X1 exu_U35897(.A(rml_ecl_cwp_d[1]), .B(exu_n19738), .Y(exu_n19740));
AND2X1 exu_U35898(.A(rml_ecl_cwp_d[0]), .B(exu_n19738), .Y(exu_n19741));
AND2X1 exu_U35899(.A(ecl_eccctl_cwp_e[2]), .B(exu_n19742), .Y(exu_n19743));
AND2X1 exu_U35900(.A(ecl_eccctl_cwp_e[1]), .B(exu_n19742), .Y(exu_n19744));
AND2X1 exu_U35901(.A(ecl_eccctl_cwp_e[0]), .B(exu_n19742), .Y(exu_n19745));
AND2X1 exu_U35902(.A(exu_n16612), .B(exu_n19746), .Y(exu_n19747));
AND2X1 exu_U35903(.A(ecl_rs2_data_31_m), .B(exu_n19746), .Y(exu_n19748));
AND2X1 exu_U35904(.A(div_ecl_adder_out_31), .B(exu_n19746), .Y(exu_n19749));
AND2X1 exu_U35905(.A(rml_cwp_cwp_thr0_next[2]), .B(exu_n19750), .Y(exu_n19751));
AND2X1 exu_U35906(.A(rml_cwp_cwp_thr0_next[1]), .B(exu_n19750), .Y(exu_n19752));
AND2X1 exu_U35907(.A(rml_oddwin_w[0]), .B(exu_n19750), .Y(exu_n19753));
AND2X1 exu_U35908(.A(rml_cwp_cwp_thr1_next[2]), .B(exu_n19754), .Y(exu_n19755));
AND2X1 exu_U35909(.A(rml_cwp_cwp_thr1_next[1]), .B(exu_n19754), .Y(exu_n19756));
AND2X1 exu_U35910(.A(rml_oddwin_w[1]), .B(exu_n19754), .Y(exu_n19757));
AND2X1 exu_U35911(.A(rml_cwp_cwp_thr2_next[2]), .B(exu_n19758), .Y(exu_n19759));
AND2X1 exu_U35912(.A(rml_cwp_cwp_thr2_next[1]), .B(exu_n19758), .Y(exu_n19760));
AND2X1 exu_U35913(.A(rml_oddwin_w[2]), .B(exu_n19758), .Y(exu_n19761));
AND2X1 exu_U35914(.A(rml_cwp_cwp_thr3_next[2]), .B(exu_n19762), .Y(exu_n19763));
AND2X1 exu_U35915(.A(rml_cwp_cwp_thr3_next[1]), .B(exu_n19762), .Y(exu_n19764));
AND2X1 exu_U35916(.A(rml_oddwin_w[3]), .B(exu_n19762), .Y(exu_n19765));
AND2X1 exu_U35917(.A(ecl_read_ffusr_e), .B(exu_n19782), .Y(exu_n19783));
AND2X1 exu_U35918(.A(ecl_read_tlusr_e), .B(exu_n19782), .Y(exu_n19784));
AND2X1 exu_U35919(.A(exu_ifu_cc_d[3]), .B(exu_n19785), .Y(exu_n19786));
AND2X1 exu_U35920(.A(exu_ifu_cc_d[1]), .B(exu_n19785), .Y(exu_n19787));
AND2X1 exu_U35921(.A(ifu_exu_tid_s2[1]), .B(exu_n19788), .Y(exu_n19789));
AND2X1 exu_U35922(.A(ifu_exu_tid_s2[0]), .B(exu_n19788), .Y(exu_n19790));
AND2X1 exu_U35923(.A(ecl_tid_d[1]), .B(exu_n19791), .Y(exu_n19792));
AND2X1 exu_U35924(.A(ecl_tid_d[0]), .B(exu_n19791), .Y(exu_n19793));
AND2X1 exu_U35925(.A(ecl_tid_e[1]), .B(exu_n19794), .Y(exu_n19795));
AND2X1 exu_U35926(.A(ecl_tid_e[0]), .B(exu_n19794), .Y(exu_n19796));
AND2X1 exu_U35927(.A(ecl_tid_w[1]), .B(exu_n19797), .Y(exu_n19798));
AND2X1 exu_U35928(.A(ecl_tid_w[0]), .B(exu_n19797), .Y(exu_n19799));
AND2X1 exu_U35929(.A(exu_n15034), .B(exu_n19800), .Y(exu_n19801));
AND2X1 exu_U35930(.A(exu_n15035), .B(exu_n19800), .Y(exu_n19802));
AND2X1 exu_U35931(.A(rml_tid_d[1]), .B(exu_n19803), .Y(exu_n19804));
AND2X1 exu_U35932(.A(rml_tid_d[0]), .B(exu_n19803), .Y(exu_n19805));
AND2X1 exu_U35933(.A(ecl_ld_tid_g[1]), .B(exu_n19818), .Y(exu_n19819));
AND2X1 exu_U35934(.A(ecl_ld_tid_g[0]), .B(exu_n19818), .Y(exu_n19820));
AND2X1 exu_U35935(.A(rml_ecl_gl_e[1]), .B(exu_n19821), .Y(exu_n19822));
AND2X1 exu_U35936(.A(rml_ecl_gl_e[0]), .B(exu_n19821), .Y(exu_n19823));
AND2X1 exu_U35937(.A(ifu_exu_rs2_s[4]), .B(exu_n19824), .Y(exu_n19825));
AND2X1 exu_U35938(.A(ifu_exu_rs2_s[3]), .B(exu_n19824), .Y(exu_n19826));
AND2X1 exu_U35939(.A(ifu_exu_rs2_s[2]), .B(exu_n19824), .Y(exu_n19827));
AND2X1 exu_U35940(.A(ifu_exu_rs2_s[1]), .B(exu_n19824), .Y(exu_n19828));
AND2X1 exu_U35941(.A(ifu_exu_rs2_s[0]), .B(exu_n19824), .Y(exu_n19829));
AND2X1 exu_U35942(.A(ifu_exu_rs3_s[4]), .B(exu_n19830), .Y(exu_n19831));
AND2X1 exu_U35943(.A(ifu_exu_rs3_s[3]), .B(exu_n19830), .Y(exu_n19832));
AND2X1 exu_U35944(.A(ifu_exu_rs3_s[2]), .B(exu_n19830), .Y(exu_n19833));
AND2X1 exu_U35945(.A(ifu_exu_rs3_s[1]), .B(exu_n19830), .Y(exu_n19834));
AND2X1 exu_U35946(.A(ifu_exu_rs3_s[0]), .B(exu_n19830), .Y(exu_n19835));
AND2X1 exu_U35947(.A(ecl_ifu_exu_rs1_d[4]), .B(exu_n19836), .Y(exu_n19837));
AND2X1 exu_U35948(.A(ecl_ifu_exu_rs1_d[3]), .B(exu_n19836), .Y(exu_n19838));
AND2X1 exu_U35949(.A(ecl_ifu_exu_rs1_d[2]), .B(exu_n19836), .Y(exu_n19839));
AND2X1 exu_U35950(.A(ecl_ifu_exu_rs1_d[1]), .B(exu_n19836), .Y(exu_n19840));
AND2X1 exu_U35951(.A(ecl_ifu_exu_rs1_d[0]), .B(exu_n19836), .Y(exu_n19841));
AND2X1 exu_U35952(.A(ecl_ifu_exu_rs2_d[4]), .B(exu_n19842), .Y(exu_n19843));
AND2X1 exu_U35953(.A(ecl_ifu_exu_rs2_d[3]), .B(exu_n19842), .Y(exu_n19844));
AND2X1 exu_U35954(.A(ecl_ifu_exu_rs2_d[2]), .B(exu_n19842), .Y(exu_n19845));
AND2X1 exu_U35955(.A(ecl_ifu_exu_rs2_d[1]), .B(exu_n19842), .Y(exu_n19846));
AND2X1 exu_U35956(.A(ecl_ifu_exu_rs2_d[0]), .B(exu_n19842), .Y(exu_n19847));
AND2X1 exu_U35957(.A(ecl_ifu_exu_rs3_d[4]), .B(exu_n19848), .Y(exu_n19849));
AND2X1 exu_U35958(.A(ecl_ifu_exu_rs3_d[3]), .B(exu_n19848), .Y(exu_n19850));
AND2X1 exu_U35959(.A(ecl_ifu_exu_rs3_d[2]), .B(exu_n19848), .Y(exu_n19851));
AND2X1 exu_U35960(.A(ecl_ifu_exu_rs3_d[1]), .B(exu_n19848), .Y(exu_n19852));
AND2X1 exu_U35961(.A(ecl_ifu_exu_rs3_d[0]), .B(exu_n19848), .Y(exu_n19853));
AND2X1 exu_U35962(.A(ecl_ifu_exu_rs1_e[4]), .B(exu_n19854), .Y(exu_n19855));
AND2X1 exu_U35963(.A(ecl_ifu_exu_rs1_e[3]), .B(exu_n19854), .Y(exu_n19856));
AND2X1 exu_U35964(.A(ecl_ifu_exu_rs1_e[2]), .B(exu_n19854), .Y(exu_n19857));
AND2X1 exu_U35965(.A(ecl_ifu_exu_rs1_e[1]), .B(exu_n19854), .Y(exu_n19858));
AND2X1 exu_U35966(.A(ecl_ifu_exu_rs1_e[0]), .B(exu_n19854), .Y(exu_n19859));
AND2X1 exu_U35967(.A(ecl_ifu_exu_rs2_e[4]), .B(exu_n19860), .Y(exu_n19861));
AND2X1 exu_U35968(.A(ecl_ifu_exu_rs2_e[3]), .B(exu_n19860), .Y(exu_n19862));
AND2X1 exu_U35969(.A(ecl_ifu_exu_rs2_e[2]), .B(exu_n19860), .Y(exu_n19863));
AND2X1 exu_U35970(.A(ecl_ifu_exu_rs2_e[1]), .B(exu_n19860), .Y(exu_n19864));
AND2X1 exu_U35971(.A(ecl_ifu_exu_rs2_e[0]), .B(exu_n19860), .Y(exu_n19865));
AND2X1 exu_U35972(.A(ecl_ifu_exu_rs3_e[4]), .B(exu_n19866), .Y(exu_n19867));
AND2X1 exu_U35973(.A(ecl_ifu_exu_rs3_e[3]), .B(exu_n19866), .Y(exu_n19868));
AND2X1 exu_U35974(.A(ecl_ifu_exu_rs3_e[2]), .B(exu_n19866), .Y(exu_n19869));
AND2X1 exu_U35975(.A(ecl_ifu_exu_rs3_e[1]), .B(exu_n19866), .Y(exu_n19870));
AND2X1 exu_U35976(.A(ecl_ifu_exu_rs3_e[0]), .B(exu_n19866), .Y(exu_n19871));
AND2X1 exu_U35977(.A(lsu_exu_rd_m[4]), .B(exu_n19872), .Y(exu_n19873));
AND2X1 exu_U35978(.A(lsu_exu_rd_m[3]), .B(exu_n19872), .Y(exu_n19874));
AND2X1 exu_U35979(.A(lsu_exu_rd_m[2]), .B(exu_n19872), .Y(exu_n19875));
AND2X1 exu_U35980(.A(lsu_exu_rd_m[1]), .B(exu_n19872), .Y(exu_n19876));
AND2X1 exu_U35981(.A(lsu_exu_rd_m[0]), .B(exu_n19872), .Y(exu_n19877));
AND2X1 exu_U35982(.A(ifu_exu_rd_d[4]), .B(exu_n19878), .Y(exu_n19879));
AND2X1 exu_U35983(.A(ifu_exu_rd_d[3]), .B(exu_n19878), .Y(exu_n19880));
AND2X1 exu_U35984(.A(ifu_exu_rd_d[2]), .B(exu_n19878), .Y(exu_n19881));
AND2X1 exu_U35985(.A(ifu_exu_rd_d[1]), .B(exu_n19878), .Y(exu_n19882));
AND2X1 exu_U35986(.A(ifu_exu_rd_d[0]), .B(exu_n19878), .Y(exu_n19883));
AND2X1 exu_U35987(.A(ecl_real_rd_e[4]), .B(exu_n19884), .Y(exu_n19885));
AND2X1 exu_U35988(.A(ecl_rd_e[3]), .B(exu_n19884), .Y(exu_n19886));
AND2X1 exu_U35989(.A(ecl_rd_e[2]), .B(exu_n19884), .Y(exu_n19887));
AND2X1 exu_U35990(.A(ecl_rd_e[1]), .B(exu_n19884), .Y(exu_n19888));
AND2X1 exu_U35991(.A(ecl_rd_e[0]), .B(exu_n19884), .Y(exu_n19889));
AND2X1 exu_U35992(.A(ecl_irf_rd_m[4]), .B(exu_n19890), .Y(exu_n19891));
AND2X1 exu_U35993(.A(ecl_irf_rd_m[3]), .B(exu_n19890), .Y(exu_n19892));
AND2X1 exu_U35994(.A(ecl_irf_rd_m[2]), .B(exu_n19890), .Y(exu_n19893));
AND2X1 exu_U35995(.A(ecl_irf_rd_m[1]), .B(exu_n19890), .Y(exu_n19894));
AND2X1 exu_U35996(.A(ecl_irf_rd_m[0]), .B(exu_n19890), .Y(exu_n19895));
AND2X1 exu_U35997(.A(ecl_ld_rd_g[4]), .B(exu_n19896), .Y(exu_n19897));
AND2X1 exu_U35998(.A(ecl_ld_rd_g[3]), .B(exu_n19896), .Y(exu_n19898));
AND2X1 exu_U35999(.A(ecl_ld_rd_g[2]), .B(exu_n19896), .Y(exu_n19899));
AND2X1 exu_U36000(.A(ecl_ld_rd_g[1]), .B(exu_n19896), .Y(exu_n19900));
AND2X1 exu_U36001(.A(ecl_ld_rd_g[0]), .B(exu_n19896), .Y(exu_n19901));
AND2X1 exu_U36002(.A(ecl_irf_rd_g[4]), .B(exu_n19902), .Y(exu_n19903));
AND2X1 exu_U36003(.A(ecl_irf_rd_g[3]), .B(exu_n19902), .Y(exu_n19904));
AND2X1 exu_U36004(.A(ecl_irf_rd_g[2]), .B(exu_n19902), .Y(exu_n19905));
AND2X1 exu_U36005(.A(ecl_irf_rd_g[1]), .B(exu_n19902), .Y(exu_n19906));
AND2X1 exu_U36006(.A(ecl_irf_rd_g[0]), .B(exu_n19902), .Y(exu_n19907));
AND2X1 exu_U36007(.A(exu_n16436), .B(exu_n19908), .Y(exu_n19909));
AND2X1 exu_U36008(.A(div_gencc_in[63]), .B(exu_n19908), .Y(exu_n19910));
AND2X1 exu_U36009(.A(exu_n15352), .B(exu_n19908), .Y(exu_n19911));
AND2X1 exu_U36010(.A(exu_n16197), .B(exu_n19908), .Y(exu_n19912));
AND2X1 exu_U36011(.A(div_ecl_low32_nonzero), .B(exu_n19908), .Y(exu_n19913));
AND2X1 exu_U36012(.A(tlu_exu_cwpccr_update_m), .B(exu_n19914), .Y(exu_n19915));
AND2X1 exu_U36013(.A(tlu_exu_cwp_m[2]), .B(exu_n19914), .Y(exu_n19916));
AND2X1 exu_U36014(.A(tlu_exu_cwp_m[1]), .B(exu_n19914), .Y(exu_n19917));
AND2X1 exu_U36015(.A(tlu_exu_cwp_m[0]), .B(exu_n19914), .Y(exu_n19918));
AND2X1 exu_U36016(.A(tlu_exu_cwp_retry_m), .B(exu_n19914), .Y(exu_n19919));
AND2X1 exu_U36017(.A(grst_l), .B(exu_n19257), .Y(exu_n19921));
AND2X1 exu_U36018(.A(ecc_rs2_err_e[6]), .B(exu_n19950), .Y(exu_n19951));
AND2X1 exu_U36019(.A(ecc_rs2_err_e[5]), .B(exu_n19950), .Y(exu_n19952));
AND2X1 exu_U36020(.A(ecc_rs2_err_e[4]), .B(exu_n19950), .Y(exu_n19953));
AND2X1 exu_U36021(.A(ecc_rs2_err_e[3]), .B(exu_n19950), .Y(exu_n19954));
AND2X1 exu_U36022(.A(ecc_rs2_err_e[2]), .B(exu_n19950), .Y(exu_n19955));
AND2X1 exu_U36023(.A(ecc_rs2_err_e[1]), .B(exu_n19950), .Y(exu_n19956));
AND2X1 exu_U36024(.A(ecc_rs2_err_e[0]), .B(exu_n19950), .Y(exu_n19957));
AND2X1 exu_U36025(.A(ecc_rs3_err_e[6]), .B(exu_n19958), .Y(exu_n19959));
AND2X1 exu_U36026(.A(ecc_rs3_err_e[5]), .B(exu_n19958), .Y(exu_n19960));
AND2X1 exu_U36027(.A(ecc_rs3_err_e[4]), .B(exu_n19958), .Y(exu_n19961));
AND2X1 exu_U36028(.A(ecc_rs3_err_e[3]), .B(exu_n19958), .Y(exu_n19962));
AND2X1 exu_U36029(.A(ecc_rs3_err_e[2]), .B(exu_n19958), .Y(exu_n19963));
AND2X1 exu_U36030(.A(ecc_rs3_err_e[1]), .B(exu_n19958), .Y(exu_n19964));
AND2X1 exu_U36031(.A(ecc_rs3_err_e[0]), .B(exu_n19958), .Y(exu_n19965));
AND2X1 exu_U36032(.A(ifu_tlu_sraddr_d[6]), .B(exu_n19966), .Y(exu_n19967));
AND2X1 exu_U36033(.A(ifu_tlu_sraddr_d[5]), .B(exu_n19966), .Y(exu_n19968));
AND2X1 exu_U36034(.A(ifu_tlu_sraddr_d[4]), .B(exu_n19966), .Y(exu_n19969));
AND2X1 exu_U36035(.A(ifu_tlu_sraddr_d[3]), .B(exu_n19966), .Y(exu_n19970));
AND2X1 exu_U36036(.A(ifu_tlu_sraddr_d[2]), .B(exu_n19966), .Y(exu_n19971));
AND2X1 exu_U36037(.A(ifu_tlu_sraddr_d[1]), .B(exu_n19966), .Y(exu_n19972));
AND2X1 exu_U36038(.A(ifu_tlu_sraddr_d[0]), .B(exu_n19966), .Y(exu_n19973));
AND2X1 exu_U36039(.A(ecl_writeback_sraddr_e[6]), .B(exu_n19974), .Y(exu_n19975));
AND2X1 exu_U36040(.A(ecl_writeback_sraddr_e[5]), .B(exu_n19974), .Y(exu_n19976));
AND2X1 exu_U36041(.A(ecl_writeback_sraddr_e[4]), .B(exu_n19974), .Y(exu_n19977));
AND2X1 exu_U36042(.A(ecl_writeback_sraddr_e[3]), .B(exu_n19974), .Y(exu_n19978));
AND2X1 exu_U36043(.A(ecl_writeback_sraddr_e[2]), .B(exu_n19974), .Y(exu_n19979));
AND2X1 exu_U36044(.A(ecl_writeback_sraddr_e[1]), .B(exu_n19974), .Y(exu_n19980));
AND2X1 exu_U36045(.A(ecl_writeback_sraddr_e[0]), .B(exu_n19974), .Y(exu_n19981));
AND2X1 exu_U36046(.A(ecl_writeback_sraddr_m[6]), .B(exu_n19982), .Y(exu_n19983));
AND2X1 exu_U36047(.A(ecl_writeback_sraddr_m[5]), .B(exu_n19982), .Y(exu_n19984));
AND2X1 exu_U36048(.A(ecl_writeback_sraddr_m[4]), .B(exu_n19982), .Y(exu_n19985));
AND2X1 exu_U36049(.A(ecl_writeback_sraddr_m[3]), .B(exu_n19982), .Y(exu_n19986));
AND2X1 exu_U36050(.A(ecl_writeback_sraddr_m[2]), .B(exu_n19982), .Y(exu_n19987));
AND2X1 exu_U36051(.A(ecl_writeback_sraddr_m[1]), .B(exu_n19982), .Y(exu_n19988));
AND2X1 exu_U36052(.A(ecl_writeback_sraddr_m[0]), .B(exu_n19982), .Y(exu_n19989));
AND2X1 exu_U36053(.A(rml_cwp_spill_next), .B(exu_n19990), .Y(exu_n19991));
AND2X1 exu_U36054(.A(rml_cwp_swap_data[8]), .B(exu_n19990), .Y(exu_n19992));
AND2X1 exu_U36055(.A(rml_cwp_spill_wtype_next[2]), .B(exu_n19990), .Y(exu_n19993));
AND2X1 exu_U36056(.A(rml_cwp_spill_wtype_next[1]), .B(exu_n19990), .Y(exu_n19994));
AND2X1 exu_U36057(.A(rml_cwp_spill_wtype_next[0]), .B(exu_n19990), .Y(exu_n19995));
AND2X1 exu_U36058(.A(byp_ecc_rs2_synd_d[6]), .B(exu_n20268), .Y(exu_n20269));
AND2X1 exu_U36059(.A(byp_ecc_rs2_synd_d[5]), .B(exu_n20268), .Y(exu_n20270));
AND2X1 exu_U36060(.A(byp_ecc_rs2_synd_d[4]), .B(exu_n20268), .Y(exu_n20271));
AND2X1 exu_U36061(.A(byp_ecc_rs2_synd_d[3]), .B(exu_n20268), .Y(exu_n20272));
AND2X1 exu_U36062(.A(byp_ecc_rs2_synd_d[2]), .B(exu_n20268), .Y(exu_n20273));
AND2X1 exu_U36063(.A(byp_ecc_rs2_synd_d[1]), .B(exu_n20268), .Y(exu_n20274));
AND2X1 exu_U36064(.A(byp_ecc_rs2_synd_d[0]), .B(exu_n20268), .Y(exu_n20275));
AND2X1 exu_U36065(.A(byp_ecc_rs2_synd_d[7]), .B(exu_n20268), .Y(exu_n20276));
AND2X1 exu_U36066(.A(byp_ecc_rs3_synd_d[6]), .B(exu_n20277), .Y(exu_n20278));
AND2X1 exu_U36067(.A(byp_ecc_rs3_synd_d[5]), .B(exu_n20277), .Y(exu_n20279));
AND2X1 exu_U36068(.A(byp_ecc_rs3_synd_d[4]), .B(exu_n20277), .Y(exu_n20280));
AND2X1 exu_U36069(.A(byp_ecc_rs3_synd_d[3]), .B(exu_n20277), .Y(exu_n20281));
AND2X1 exu_U36070(.A(byp_ecc_rs3_synd_d[2]), .B(exu_n20277), .Y(exu_n20282));
AND2X1 exu_U36071(.A(byp_ecc_rs3_synd_d[1]), .B(exu_n20277), .Y(exu_n20283));
AND2X1 exu_U36072(.A(byp_ecc_rs3_synd_d[0]), .B(exu_n20277), .Y(exu_n20284));
AND2X1 exu_U36073(.A(byp_ecc_rs3_synd_d[7]), .B(exu_n20277), .Y(exu_n20285));
AND2X1 exu_U36074(.A(ecl_alu_xcc_e[2]), .B(exu_n20286), .Y(exu_n20287));
AND2X1 exu_U36075(.A(ecl_adder_xcc[1]), .B(exu_n20286), .Y(exu_n20288));
AND2X1 exu_U36076(.A(ecl_adder_xcc[0]), .B(exu_n20286), .Y(exu_n20289));
AND2X1 exu_U36077(.A(exu_n15339), .B(exu_n20286), .Y(exu_n20290));
AND2X1 exu_U36078(.A(exu_n15426), .B(exu_n20286), .Y(exu_n20291));
AND2X1 exu_U36079(.A(ecl_adder_icc[1]), .B(exu_n20286), .Y(exu_n20292));
AND2X1 exu_U36080(.A(ecl_adder_icc[0]), .B(exu_n20286), .Y(exu_n20293));
AND2X1 exu_U36081(.A(exu_n15338), .B(exu_n20286), .Y(exu_n20294));
AND2X1 exu_U36082(.A(exu_n18012), .B(exu_n20340), .Y(exu_n20341));
AND2X1 exu_U36083(.A(ecl_writeback_rdpr_mux2_out[5]), .B(exu_n20340), .Y(exu_n20342));
AND2X1 exu_U36084(.A(ecl_writeback_rdpr_mux2_out[4]), .B(exu_n20340), .Y(exu_n20343));
AND2X1 exu_U36085(.A(ecl_writeback_rdpr_mux2_out[3]), .B(exu_n20340), .Y(exu_n20344));
AND2X1 exu_U36086(.A(ecl_writeback_rdpr_mux2_out[2]), .B(exu_n20340), .Y(exu_n20345));
AND2X1 exu_U36087(.A(ecl_writeback_rdpr_mux2_out[1]), .B(exu_n20340), .Y(exu_n20346));
AND2X1 exu_U36088(.A(ecl_writeback_rdpr_mux2_out[0]), .B(exu_n20340), .Y(exu_n20347));
AND2X1 exu_U36089(.A(exu_n18011), .B(exu_n20340), .Y(exu_n20348));
AND2X1 exu_U36090(.A(byp_irf_rd_data_w[6]), .B(exu_n16008), .Y(exu_n21629));
AND2X1 exu_U36091(.A(byp_irf_rd_data_w[5]), .B(exu_n16008), .Y(exu_n21630));
AND2X1 exu_U36092(.A(byp_irf_rd_data_w[4]), .B(exu_n16008), .Y(exu_n21631));
AND2X1 exu_U36093(.A(byp_irf_rd_data_w[3]), .B(exu_n16008), .Y(exu_n21632));
AND2X1 exu_U36094(.A(byp_irf_rd_data_w[2]), .B(exu_n16008), .Y(exu_n21633));
AND2X1 exu_U36095(.A(byp_irf_rd_data_w[1]), .B(exu_n16008), .Y(exu_n21634));
AND2X1 exu_U36096(.A(byp_irf_rd_data_w[31]), .B(exu_n16007), .Y(exu_n21635));
AND2X1 exu_U36097(.A(byp_irf_rd_data_w[30]), .B(exu_n16007), .Y(exu_n21636));
AND2X1 exu_U36098(.A(byp_irf_rd_data_w[29]), .B(exu_n16007), .Y(exu_n21637));
AND2X1 exu_U36099(.A(byp_irf_rd_data_w[28]), .B(exu_n16007), .Y(exu_n21638));
AND2X1 exu_U36100(.A(byp_irf_rd_data_w[27]), .B(exu_n16007), .Y(exu_n21639));
AND2X1 exu_U36101(.A(byp_irf_rd_data_w[0]), .B(exu_n16007), .Y(exu_n21640));
AND2X1 exu_U36102(.A(byp_irf_rd_data_w[26]), .B(exu_n16007), .Y(exu_n21641));
AND2X1 exu_U36103(.A(byp_irf_rd_data_w[25]), .B(exu_n16007), .Y(exu_n21642));
AND2X1 exu_U36104(.A(byp_irf_rd_data_w[24]), .B(exu_n16007), .Y(exu_n21643));
AND2X1 exu_U36105(.A(byp_irf_rd_data_w[23]), .B(exu_n16007), .Y(exu_n21644));
AND2X1 exu_U36106(.A(byp_irf_rd_data_w[22]), .B(exu_n16007), .Y(exu_n21645));
AND2X1 exu_U36107(.A(byp_irf_rd_data_w[21]), .B(exu_n16007), .Y(exu_n21646));
AND2X1 exu_U36108(.A(byp_irf_rd_data_w[20]), .B(exu_n16007), .Y(exu_n21647));
AND2X1 exu_U36109(.A(byp_irf_rd_data_w[19]), .B(exu_n16006), .Y(exu_n21648));
AND2X1 exu_U36110(.A(byp_irf_rd_data_w[18]), .B(exu_n16006), .Y(exu_n21649));
AND2X1 exu_U36111(.A(byp_irf_rd_data_w[17]), .B(exu_n16006), .Y(exu_n21650));
AND2X1 exu_U36112(.A(byp_irf_rd_data_w[16]), .B(exu_n16006), .Y(exu_n21651));
AND2X1 exu_U36113(.A(byp_irf_rd_data_w[15]), .B(exu_n16006), .Y(exu_n21652));
AND2X1 exu_U36114(.A(byp_irf_rd_data_w[14]), .B(exu_n16006), .Y(exu_n21653));
AND2X1 exu_U36115(.A(byp_irf_rd_data_w[13]), .B(exu_n16006), .Y(exu_n21654));
AND2X1 exu_U36116(.A(byp_irf_rd_data_w[12]), .B(exu_n16006), .Y(exu_n21655));
AND2X1 exu_U36117(.A(byp_irf_rd_data_w[11]), .B(exu_n16006), .Y(exu_n21656));
AND2X1 exu_U36118(.A(byp_irf_rd_data_w[10]), .B(exu_n16006), .Y(exu_n21657));
AND2X1 exu_U36119(.A(byp_irf_rd_data_w[9]), .B(exu_n16006), .Y(exu_n21658));
AND2X1 exu_U36120(.A(byp_irf_rd_data_w[8]), .B(exu_n16006), .Y(exu_n21659));
AND2X1 exu_U36121(.A(byp_irf_rd_data_w[7]), .B(exu_n16006), .Y(exu_n21660));
AND2X1 exu_U36122(.A(div_yreg_next_yreg_thr0[6]), .B(exu_n16012), .Y(exu_n21662));
AND2X1 exu_U36123(.A(div_yreg_next_yreg_thr0[5]), .B(exu_n16012), .Y(exu_n21663));
AND2X1 exu_U36124(.A(div_yreg_next_yreg_thr0[4]), .B(exu_n16012), .Y(exu_n21664));
AND2X1 exu_U36125(.A(div_yreg_next_yreg_thr0[3]), .B(exu_n16012), .Y(exu_n21665));
AND2X1 exu_U36126(.A(div_yreg_next_yreg_thr0[2]), .B(exu_n16012), .Y(exu_n21666));
AND2X1 exu_U36127(.A(div_yreg_next_yreg_thr0[1]), .B(exu_n16012), .Y(exu_n21667));
AND2X1 exu_U36128(.A(div_yreg_next_yreg_thr0[31]), .B(exu_n16011), .Y(exu_n21668));
AND2X1 exu_U36129(.A(div_yreg_next_yreg_thr0[30]), .B(exu_n16011), .Y(exu_n21669));
AND2X1 exu_U36130(.A(div_yreg_next_yreg_thr0[29]), .B(exu_n16011), .Y(exu_n21670));
AND2X1 exu_U36131(.A(div_yreg_next_yreg_thr0[28]), .B(exu_n16011), .Y(exu_n21671));
AND2X1 exu_U36132(.A(div_yreg_next_yreg_thr0[27]), .B(exu_n16011), .Y(exu_n21672));
AND2X1 exu_U36133(.A(div_yreg_next_yreg_thr0[0]), .B(exu_n16011), .Y(exu_n21673));
AND2X1 exu_U36134(.A(div_yreg_next_yreg_thr0[26]), .B(exu_n16011), .Y(exu_n21674));
AND2X1 exu_U36135(.A(div_yreg_next_yreg_thr0[25]), .B(exu_n16011), .Y(exu_n21675));
AND2X1 exu_U36136(.A(div_yreg_next_yreg_thr0[24]), .B(exu_n16011), .Y(exu_n21676));
AND2X1 exu_U36137(.A(div_yreg_next_yreg_thr0[23]), .B(exu_n16011), .Y(exu_n21677));
AND2X1 exu_U36138(.A(div_yreg_next_yreg_thr0[22]), .B(exu_n16011), .Y(exu_n21678));
AND2X1 exu_U36139(.A(div_yreg_next_yreg_thr0[21]), .B(exu_n16011), .Y(exu_n21679));
AND2X1 exu_U36140(.A(div_yreg_next_yreg_thr0[20]), .B(exu_n16011), .Y(exu_n21680));
AND2X1 exu_U36141(.A(div_yreg_next_yreg_thr0[19]), .B(exu_n16010), .Y(exu_n21681));
AND2X1 exu_U36142(.A(div_yreg_next_yreg_thr0[18]), .B(exu_n16010), .Y(exu_n21682));
AND2X1 exu_U36143(.A(div_yreg_next_yreg_thr0[17]), .B(exu_n16010), .Y(exu_n21683));
AND2X1 exu_U36144(.A(div_yreg_next_yreg_thr0[16]), .B(exu_n16010), .Y(exu_n21684));
AND2X1 exu_U36145(.A(div_yreg_next_yreg_thr0[15]), .B(exu_n16010), .Y(exu_n21685));
AND2X1 exu_U36146(.A(div_yreg_next_yreg_thr0[14]), .B(exu_n16010), .Y(exu_n21686));
AND2X1 exu_U36147(.A(div_yreg_next_yreg_thr0[13]), .B(exu_n16010), .Y(exu_n21687));
AND2X1 exu_U36148(.A(div_yreg_next_yreg_thr0[12]), .B(exu_n16010), .Y(exu_n21688));
AND2X1 exu_U36149(.A(div_yreg_next_yreg_thr0[11]), .B(exu_n16010), .Y(exu_n21689));
AND2X1 exu_U36150(.A(div_yreg_next_yreg_thr0[10]), .B(exu_n16010), .Y(exu_n21690));
AND2X1 exu_U36151(.A(div_yreg_next_yreg_thr0[9]), .B(exu_n16010), .Y(exu_n21691));
AND2X1 exu_U36152(.A(div_yreg_next_yreg_thr0[8]), .B(exu_n16010), .Y(exu_n21692));
AND2X1 exu_U36153(.A(div_yreg_next_yreg_thr0[7]), .B(exu_n16010), .Y(exu_n21693));
AND2X1 exu_U36154(.A(div_yreg_next_yreg_thr1[6]), .B(exu_n16016), .Y(exu_n21695));
AND2X1 exu_U36155(.A(div_yreg_next_yreg_thr1[5]), .B(exu_n16016), .Y(exu_n21696));
AND2X1 exu_U36156(.A(div_yreg_next_yreg_thr1[4]), .B(exu_n16016), .Y(exu_n21697));
AND2X1 exu_U36157(.A(div_yreg_next_yreg_thr1[3]), .B(exu_n16016), .Y(exu_n21698));
AND2X1 exu_U36158(.A(div_yreg_next_yreg_thr1[2]), .B(exu_n16016), .Y(exu_n21699));
AND2X1 exu_U36159(.A(div_yreg_next_yreg_thr1[1]), .B(exu_n16016), .Y(exu_n21700));
AND2X1 exu_U36160(.A(div_yreg_next_yreg_thr1[31]), .B(exu_n16015), .Y(exu_n21701));
AND2X1 exu_U36161(.A(div_yreg_next_yreg_thr1[30]), .B(exu_n16015), .Y(exu_n21702));
AND2X1 exu_U36162(.A(div_yreg_next_yreg_thr1[29]), .B(exu_n16015), .Y(exu_n21703));
AND2X1 exu_U36163(.A(div_yreg_next_yreg_thr1[28]), .B(exu_n16015), .Y(exu_n21704));
AND2X1 exu_U36164(.A(div_yreg_next_yreg_thr1[27]), .B(exu_n16015), .Y(exu_n21705));
AND2X1 exu_U36165(.A(div_yreg_next_yreg_thr1[0]), .B(exu_n16015), .Y(exu_n21706));
AND2X1 exu_U36166(.A(div_yreg_next_yreg_thr1[26]), .B(exu_n16015), .Y(exu_n21707));
AND2X1 exu_U36167(.A(div_yreg_next_yreg_thr1[25]), .B(exu_n16015), .Y(exu_n21708));
AND2X1 exu_U36168(.A(div_yreg_next_yreg_thr1[24]), .B(exu_n16015), .Y(exu_n21709));
AND2X1 exu_U36169(.A(div_yreg_next_yreg_thr1[23]), .B(exu_n16015), .Y(exu_n21710));
AND2X1 exu_U36170(.A(div_yreg_next_yreg_thr1[22]), .B(exu_n16015), .Y(exu_n21711));
AND2X1 exu_U36171(.A(div_yreg_next_yreg_thr1[21]), .B(exu_n16015), .Y(exu_n21712));
AND2X1 exu_U36172(.A(div_yreg_next_yreg_thr1[20]), .B(exu_n16015), .Y(exu_n21713));
AND2X1 exu_U36173(.A(div_yreg_next_yreg_thr1[19]), .B(exu_n16014), .Y(exu_n21714));
AND2X1 exu_U36174(.A(div_yreg_next_yreg_thr1[18]), .B(exu_n16014), .Y(exu_n21715));
AND2X1 exu_U36175(.A(div_yreg_next_yreg_thr1[17]), .B(exu_n16014), .Y(exu_n21716));
AND2X1 exu_U36176(.A(div_yreg_next_yreg_thr1[16]), .B(exu_n16014), .Y(exu_n21717));
AND2X1 exu_U36177(.A(div_yreg_next_yreg_thr1[15]), .B(exu_n16014), .Y(exu_n21718));
AND2X1 exu_U36178(.A(div_yreg_next_yreg_thr1[14]), .B(exu_n16014), .Y(exu_n21719));
AND2X1 exu_U36179(.A(div_yreg_next_yreg_thr1[13]), .B(exu_n16014), .Y(exu_n21720));
AND2X1 exu_U36180(.A(div_yreg_next_yreg_thr1[12]), .B(exu_n16014), .Y(exu_n21721));
AND2X1 exu_U36181(.A(div_yreg_next_yreg_thr1[11]), .B(exu_n16014), .Y(exu_n21722));
AND2X1 exu_U36182(.A(div_yreg_next_yreg_thr1[10]), .B(exu_n16014), .Y(exu_n21723));
AND2X1 exu_U36183(.A(div_yreg_next_yreg_thr1[9]), .B(exu_n16014), .Y(exu_n21724));
AND2X1 exu_U36184(.A(div_yreg_next_yreg_thr1[8]), .B(exu_n16014), .Y(exu_n21725));
AND2X1 exu_U36185(.A(div_yreg_next_yreg_thr1[7]), .B(exu_n16014), .Y(exu_n21726));
AND2X1 exu_U36186(.A(div_yreg_next_yreg_thr2[6]), .B(exu_n16020), .Y(exu_n21728));
AND2X1 exu_U36187(.A(div_yreg_next_yreg_thr2[5]), .B(exu_n16020), .Y(exu_n21729));
AND2X1 exu_U36188(.A(div_yreg_next_yreg_thr2[4]), .B(exu_n16020), .Y(exu_n21730));
AND2X1 exu_U36189(.A(div_yreg_next_yreg_thr2[3]), .B(exu_n16020), .Y(exu_n21731));
AND2X1 exu_U36190(.A(div_yreg_next_yreg_thr2[2]), .B(exu_n16020), .Y(exu_n21732));
AND2X1 exu_U36191(.A(div_yreg_next_yreg_thr2[1]), .B(exu_n16020), .Y(exu_n21733));
AND2X1 exu_U36192(.A(div_yreg_next_yreg_thr2[31]), .B(exu_n16019), .Y(exu_n21734));
AND2X1 exu_U36193(.A(div_yreg_next_yreg_thr2[30]), .B(exu_n16019), .Y(exu_n21735));
AND2X1 exu_U36194(.A(div_yreg_next_yreg_thr2[29]), .B(exu_n16019), .Y(exu_n21736));
AND2X1 exu_U36195(.A(div_yreg_next_yreg_thr2[28]), .B(exu_n16019), .Y(exu_n21737));
AND2X1 exu_U36196(.A(div_yreg_next_yreg_thr2[27]), .B(exu_n16019), .Y(exu_n21738));
AND2X1 exu_U36197(.A(div_yreg_next_yreg_thr2[0]), .B(exu_n16019), .Y(exu_n21739));
AND2X1 exu_U36198(.A(div_yreg_next_yreg_thr2[26]), .B(exu_n16019), .Y(exu_n21740));
AND2X1 exu_U36199(.A(div_yreg_next_yreg_thr2[25]), .B(exu_n16019), .Y(exu_n21741));
AND2X1 exu_U36200(.A(div_yreg_next_yreg_thr2[24]), .B(exu_n16019), .Y(exu_n21742));
AND2X1 exu_U36201(.A(div_yreg_next_yreg_thr2[23]), .B(exu_n16019), .Y(exu_n21743));
AND2X1 exu_U36202(.A(div_yreg_next_yreg_thr2[22]), .B(exu_n16019), .Y(exu_n21744));
AND2X1 exu_U36203(.A(div_yreg_next_yreg_thr2[21]), .B(exu_n16019), .Y(exu_n21745));
AND2X1 exu_U36204(.A(div_yreg_next_yreg_thr2[20]), .B(exu_n16019), .Y(exu_n21746));
AND2X1 exu_U36205(.A(div_yreg_next_yreg_thr2[19]), .B(exu_n16018), .Y(exu_n21747));
AND2X1 exu_U36206(.A(div_yreg_next_yreg_thr2[18]), .B(exu_n16018), .Y(exu_n21748));
AND2X1 exu_U36207(.A(div_yreg_next_yreg_thr2[17]), .B(exu_n16018), .Y(exu_n21749));
AND2X1 exu_U36208(.A(div_yreg_next_yreg_thr2[16]), .B(exu_n16018), .Y(exu_n21750));
AND2X1 exu_U36209(.A(div_yreg_next_yreg_thr2[15]), .B(exu_n16018), .Y(exu_n21751));
AND2X1 exu_U36210(.A(div_yreg_next_yreg_thr2[14]), .B(exu_n16018), .Y(exu_n21752));
AND2X1 exu_U36211(.A(div_yreg_next_yreg_thr2[13]), .B(exu_n16018), .Y(exu_n21753));
AND2X1 exu_U36212(.A(div_yreg_next_yreg_thr2[12]), .B(exu_n16018), .Y(exu_n21754));
AND2X1 exu_U36213(.A(div_yreg_next_yreg_thr2[11]), .B(exu_n16018), .Y(exu_n21755));
AND2X1 exu_U36214(.A(div_yreg_next_yreg_thr2[10]), .B(exu_n16018), .Y(exu_n21756));
AND2X1 exu_U36215(.A(div_yreg_next_yreg_thr2[9]), .B(exu_n16018), .Y(exu_n21757));
AND2X1 exu_U36216(.A(div_yreg_next_yreg_thr2[8]), .B(exu_n16018), .Y(exu_n21758));
AND2X1 exu_U36217(.A(div_yreg_next_yreg_thr2[7]), .B(exu_n16018), .Y(exu_n21759));
AND2X1 exu_U36218(.A(div_yreg_next_yreg_thr3[6]), .B(exu_n16024), .Y(exu_n21761));
AND2X1 exu_U36219(.A(div_yreg_next_yreg_thr3[5]), .B(exu_n16024), .Y(exu_n21762));
AND2X1 exu_U36220(.A(div_yreg_next_yreg_thr3[4]), .B(exu_n16024), .Y(exu_n21763));
AND2X1 exu_U36221(.A(div_yreg_next_yreg_thr3[3]), .B(exu_n16024), .Y(exu_n21764));
AND2X1 exu_U36222(.A(div_yreg_next_yreg_thr3[2]), .B(exu_n16024), .Y(exu_n21765));
AND2X1 exu_U36223(.A(div_yreg_next_yreg_thr3[1]), .B(exu_n16024), .Y(exu_n21766));
AND2X1 exu_U36224(.A(div_yreg_next_yreg_thr3[31]), .B(exu_n16023), .Y(exu_n21767));
AND2X1 exu_U36225(.A(div_yreg_next_yreg_thr3[30]), .B(exu_n16023), .Y(exu_n21768));
AND2X1 exu_U36226(.A(div_yreg_next_yreg_thr3[29]), .B(exu_n16023), .Y(exu_n21769));
AND2X1 exu_U36227(.A(div_yreg_next_yreg_thr3[28]), .B(exu_n16023), .Y(exu_n21770));
AND2X1 exu_U36228(.A(div_yreg_next_yreg_thr3[27]), .B(exu_n16023), .Y(exu_n21771));
AND2X1 exu_U36229(.A(div_yreg_next_yreg_thr3[0]), .B(exu_n16023), .Y(exu_n21772));
AND2X1 exu_U36230(.A(div_yreg_next_yreg_thr3[26]), .B(exu_n16023), .Y(exu_n21773));
AND2X1 exu_U36231(.A(div_yreg_next_yreg_thr3[25]), .B(exu_n16023), .Y(exu_n21774));
AND2X1 exu_U36232(.A(div_yreg_next_yreg_thr3[24]), .B(exu_n16023), .Y(exu_n21775));
AND2X1 exu_U36233(.A(div_yreg_next_yreg_thr3[23]), .B(exu_n16023), .Y(exu_n21776));
AND2X1 exu_U36234(.A(div_yreg_next_yreg_thr3[22]), .B(exu_n16023), .Y(exu_n21777));
AND2X1 exu_U36235(.A(div_yreg_next_yreg_thr3[21]), .B(exu_n16023), .Y(exu_n21778));
AND2X1 exu_U36236(.A(div_yreg_next_yreg_thr3[20]), .B(exu_n16023), .Y(exu_n21779));
AND2X1 exu_U36237(.A(div_yreg_next_yreg_thr3[19]), .B(exu_n16022), .Y(exu_n21780));
AND2X1 exu_U36238(.A(div_yreg_next_yreg_thr3[18]), .B(exu_n16022), .Y(exu_n21781));
AND2X1 exu_U36239(.A(div_yreg_next_yreg_thr3[17]), .B(exu_n16022), .Y(exu_n21782));
AND2X1 exu_U36240(.A(div_yreg_next_yreg_thr3[16]), .B(exu_n16022), .Y(exu_n21783));
AND2X1 exu_U36241(.A(div_yreg_next_yreg_thr3[15]), .B(exu_n16022), .Y(exu_n21784));
AND2X1 exu_U36242(.A(div_yreg_next_yreg_thr3[14]), .B(exu_n16022), .Y(exu_n21785));
AND2X1 exu_U36243(.A(div_yreg_next_yreg_thr3[13]), .B(exu_n16022), .Y(exu_n21786));
AND2X1 exu_U36244(.A(div_yreg_next_yreg_thr3[12]), .B(exu_n16022), .Y(exu_n21787));
AND2X1 exu_U36245(.A(div_yreg_next_yreg_thr3[11]), .B(exu_n16022), .Y(exu_n21788));
AND2X1 exu_U36246(.A(div_yreg_next_yreg_thr3[10]), .B(exu_n16022), .Y(exu_n21789));
AND2X1 exu_U36247(.A(div_yreg_next_yreg_thr3[9]), .B(exu_n16022), .Y(exu_n21790));
AND2X1 exu_U36248(.A(div_yreg_next_yreg_thr3[8]), .B(exu_n16022), .Y(exu_n21791));
AND2X1 exu_U36249(.A(div_yreg_next_yreg_thr3[7]), .B(exu_n16022), .Y(exu_n21792));
AND2X1 exu_U36250(.A(exu_n16300), .B(exu_n15211), .Y(exu_n24338));
AND2X1 exu_U36251(.A(exu_n15271), .B(exu_n16300), .Y(exu_n24342));
AND2X1 exu_U36252(.A(exu_n15272), .B(exu_n16300), .Y(exu_n24346));
AND2X1 exu_U36253(.A(exu_n15273), .B(exu_n16300), .Y(exu_n24350));
AND2X1 exu_U36254(.A(exu_n15274), .B(exu_n16300), .Y(exu_n24354));
AND2X1 exu_U36255(.A(exu_n15275), .B(exu_n16300), .Y(exu_n24358));
AND2X1 exu_U36256(.A(exu_n15276), .B(exu_n16300), .Y(exu_n24362));
AND2X1 exu_U36257(.A(exu_n15277), .B(exu_n16300), .Y(exu_n24366));
AND2X1 exu_U36258(.A(exu_n15278), .B(exu_n16300), .Y(exu_n24370));
AND2X1 exu_U36259(.A(exu_n15279), .B(exu_n16300), .Y(exu_n24374));
AND2X1 exu_U36260(.A(exu_n15280), .B(exu_n16300), .Y(exu_n24378));
AND2X1 exu_U36261(.A(exu_n15281), .B(exu_n16300), .Y(exu_n24382));
AND2X1 exu_U36262(.A(exu_n15282), .B(exu_n16300), .Y(exu_n24386));
AND2X1 exu_U36263(.A(exu_n15283), .B(exu_n16300), .Y(exu_n24390));
AND2X1 exu_U36264(.A(exu_n15284), .B(exu_n16300), .Y(exu_n24394));
AND2X1 exu_U36265(.A(exu_n15285), .B(exu_n16300), .Y(exu_n24398));
AND2X1 exu_U36266(.A(exu_n15286), .B(exu_n16300), .Y(exu_n24402));
AND2X1 exu_U36267(.A(exu_n15287), .B(exu_n16300), .Y(exu_n24406));
AND2X1 exu_U36268(.A(exu_n15288), .B(exu_n16300), .Y(exu_n24410));
AND2X1 exu_U36269(.A(exu_n15289), .B(exu_n16300), .Y(exu_n24414));
AND2X1 exu_U36270(.A(exu_n15290), .B(exu_n16300), .Y(exu_n24418));
AND2X1 exu_U36271(.A(exu_n15291), .B(exu_n16300), .Y(exu_n24422));
AND2X1 exu_U36272(.A(exu_n15292), .B(exu_n16300), .Y(exu_n24426));
AND2X1 exu_U36273(.A(exu_n15293), .B(exu_n16300), .Y(exu_n24430));
AND2X1 exu_U36274(.A(exu_n15294), .B(exu_n16300), .Y(exu_n24434));
AND2X1 exu_U36275(.A(exu_n15295), .B(exu_n16300), .Y(exu_n24438));
AND2X1 exu_U36276(.A(exu_n15296), .B(exu_n16300), .Y(exu_n24442));
AND2X1 exu_U36277(.A(exu_n15297), .B(exu_n16300), .Y(exu_n24446));
AND2X1 exu_U36278(.A(exu_n15298), .B(exu_n16300), .Y(exu_n24450));
AND2X1 exu_U36279(.A(exu_n15299), .B(exu_n16300), .Y(exu_n24454));
AND2X1 exu_U36280(.A(exu_n15300), .B(exu_n16300), .Y(exu_n24458));
AND2X1 exu_U36281(.A(exu_n15301), .B(exu_n16300), .Y(exu_n24462));
AND2X1 exu_U36282(.A(exu_n15302), .B(exu_n16300), .Y(exu_n24466));
AND2X1 exu_U36283(.A(exu_n15303), .B(exu_n16300), .Y(exu_n24470));
AND2X1 exu_U36284(.A(exu_n15304), .B(exu_n16300), .Y(exu_n24474));
AND2X1 exu_U36285(.A(exu_n15305), .B(exu_n16300), .Y(exu_n24478));
AND2X1 exu_U36286(.A(exu_n15306), .B(exu_n16300), .Y(exu_n24482));
AND2X1 exu_U36287(.A(exu_n15307), .B(exu_n16300), .Y(exu_n24486));
AND2X1 exu_U36288(.A(exu_n15308), .B(exu_n16300), .Y(exu_n24490));
AND2X1 exu_U36289(.A(exu_n15309), .B(exu_n16300), .Y(exu_n24494));
AND2X1 exu_U36290(.A(exu_n15310), .B(exu_n16300), .Y(exu_n24498));
AND2X1 exu_U36291(.A(exu_n15311), .B(exu_n16300), .Y(exu_n24502));
AND2X1 exu_U36292(.A(exu_n15312), .B(exu_n16300), .Y(exu_n24506));
AND2X1 exu_U36293(.A(exu_n15313), .B(exu_n16300), .Y(exu_n24510));
AND2X1 exu_U36294(.A(exu_n15314), .B(exu_n16300), .Y(exu_n24514));
AND2X1 exu_U36295(.A(exu_n15315), .B(exu_n16300), .Y(exu_n24518));
AND2X1 exu_U36296(.A(exu_n15316), .B(exu_n16300), .Y(exu_n24522));
AND2X1 exu_U36297(.A(exu_n15317), .B(exu_n16300), .Y(exu_n24526));
AND2X1 exu_U36298(.A(exu_n15318), .B(exu_n16300), .Y(exu_n24530));
AND2X1 exu_U36299(.A(exu_n15319), .B(exu_n16300), .Y(exu_n24534));
AND2X1 exu_U36300(.A(exu_n15320), .B(exu_n16300), .Y(exu_n24538));
AND2X1 exu_U36301(.A(exu_n15321), .B(exu_n16300), .Y(exu_n24542));
AND2X1 exu_U36302(.A(exu_n15322), .B(exu_n16300), .Y(exu_n24546));
AND2X1 exu_U36303(.A(exu_n15323), .B(exu_n16300), .Y(exu_n24550));
AND2X1 exu_U36304(.A(exu_n15324), .B(exu_n16300), .Y(exu_n24554));
AND2X1 exu_U36305(.A(exu_n15325), .B(exu_n16300), .Y(exu_n24558));
AND2X1 exu_U36306(.A(exu_n15326), .B(exu_n16300), .Y(exu_n24562));
AND2X1 exu_U36307(.A(exu_n15327), .B(exu_n16300), .Y(exu_n24566));
AND2X1 exu_U36308(.A(exu_n15328), .B(exu_n16300), .Y(exu_n24570));
AND2X1 exu_U36309(.A(exu_n15329), .B(exu_n16300), .Y(exu_n24574));
AND2X1 exu_U36310(.A(exu_n15330), .B(exu_n16300), .Y(exu_n24578));
AND2X1 exu_U36311(.A(exu_n15331), .B(exu_n16300), .Y(exu_n24582));
AND2X1 exu_U36312(.A(exu_n15332), .B(exu_n16300), .Y(exu_n24586));
AND2X1 exu_U36313(.A(exu_n15333), .B(exu_n16300), .Y(exu_n24590));
AND2X1 exu_U36314(.A(shft_shift16_e[0]), .B(shft_rshifterinput_b1[9]), .Y(exu_n27754));
INVX1 exu_U36315(.A(exu_n27754), .Y(exu_n15000));
AND2X1 exu_U36316(.A(shft_rshifterinput_b1[8]), .B(exu_n16148), .Y(exu_n27755));
INVX1 exu_U36317(.A(exu_n27755), .Y(exu_n15001));
AND2X1 exu_U36318(.A(shft_rshifterinput_b1[7]), .B(exu_n16148), .Y(exu_n27756));
INVX1 exu_U36319(.A(exu_n27756), .Y(exu_n15002));
AND2X1 exu_U36320(.A(shft_rshifterinput_b1[6]), .B(shft_shift16_e[0]), .Y(exu_n27757));
INVX1 exu_U36321(.A(exu_n27757), .Y(exu_n15003));
AND2X1 exu_U36322(.A(shft_rshifterinput_b1[5]), .B(exu_n16148), .Y(exu_n27782));
INVX1 exu_U36323(.A(exu_n27782), .Y(exu_n15004));
AND2X1 exu_U36324(.A(shft_rshifterinput_b1[4]), .B(shft_shift16_e[0]), .Y(exu_n27843));
INVX1 exu_U36325(.A(exu_n27843), .Y(exu_n15005));
AND2X1 exu_U36326(.A(shft_rshifterinput_b1[15]), .B(exu_n16145), .Y(exu_n27859));
AND2X1 exu_U36327(.A(shft_rshifterinput_b1[14]), .B(exu_n16145), .Y(exu_n27863));
AND2X1 exu_U36328(.A(shft_rshifterinput_b1[13]), .B(exu_n16145), .Y(exu_n27867));
AND2X1 exu_U36329(.A(shft_rshifterinput_b1[12]), .B(exu_n16145), .Y(exu_n27871));
AND2X1 exu_U36330(.A(shft_rshifterinput_b1[11]), .B(exu_n16145), .Y(exu_n27875));
AND2X1 exu_U36331(.A(shft_rshifterinput_b1[10]), .B(exu_n16145), .Y(exu_n27879));
AND2X1 exu_U36332(.A(shft_rshifterinput_b1[9]), .B(exu_n16145), .Y(exu_n27883));
AND2X1 exu_U36333(.A(shft_rshifterinput_b1[8]), .B(exu_n16145), .Y(exu_n27887));
AND2X1 exu_U36334(.A(shft_rshifterinput_b1[7]), .B(exu_n16145), .Y(exu_n27892));
AND2X1 exu_U36335(.A(shft_rshifterinput_b1[6]), .B(exu_n16145), .Y(exu_n27896));
AND2X1 exu_U36336(.A(shft_rshifterinput_b1[5]), .B(exu_n16145), .Y(exu_n27900));
AND2X1 exu_U36337(.A(shft_rshifterinput_b1[4]), .B(exu_n16145), .Y(exu_n27904));
AND2X1 exu_U36338(.A(shft_rshifterinput_b1[3]), .B(exu_n16145), .Y(exu_n27908));
AND2X1 exu_U36339(.A(shft_rshifterinput_b1[2]), .B(exu_n16145), .Y(exu_n27912));
AND2X1 exu_U36340(.A(shft_rshifterinput_b1[1]), .B(exu_n16145), .Y(exu_n27916));
AND2X1 exu_U36341(.A(shft_rshifterinput_b1[0]), .B(exu_n16145), .Y(exu_n27920));
AND2X1 exu_U36342(.A(shft_rshifterinput_b1[15]), .B(exu_n16148), .Y(exu_n27971));
INVX1 exu_U36343(.A(exu_n27971), .Y(exu_n15006));
AND2X1 exu_U36344(.A(shft_rshifterinput_b1[14]), .B(shft_shift16_e[0]), .Y(exu_n27972));
INVX1 exu_U36345(.A(exu_n27972), .Y(exu_n15007));
AND2X1 exu_U36346(.A(shft_rshifterinput_b1[13]), .B(shft_shift16_e[0]), .Y(exu_n27973));
INVX1 exu_U36347(.A(exu_n27973), .Y(exu_n15008));
AND2X1 exu_U36348(.A(shft_rshifterinput_b1[12]), .B(exu_n16148), .Y(exu_n27974));
INVX1 exu_U36349(.A(exu_n27974), .Y(exu_n15009));
AND2X1 exu_U36350(.A(shft_rshifterinput_b1[11]), .B(exu_n16148), .Y(exu_n27975));
INVX1 exu_U36351(.A(exu_n27975), .Y(exu_n15010));
AND2X1 exu_U36352(.A(shft_rshifterinput_b1[10]), .B(shft_shift16_e[0]), .Y(exu_n27976));
INVX1 exu_U36353(.A(exu_n27976), .Y(exu_n15011));
AND2X1 exu_U36354(.A(exu_n16233), .B(exu_n27958), .Y(exu_n27981));
AND2X1 exu_U36355(.A(exu_n27977), .B(exu_n16232), .Y(exu_n27985));
AND2X1 exu_U36356(.A(exu_n27888), .B(exu_n16230), .Y(exu_n28142));
AND2X1 exu_U36357(.A(exu_n27927), .B(exu_n16230), .Y(exu_n28203));
AND2X1 exu_U36358(.A(exu_n27958), .B(exu_n15401), .Y(exu_n28264));
AND2X1 exu_U36359(.A(exu_n27888), .B(exu_n16233), .Y(exu_n28316));
AND2X1 exu_U36360(.A(exu_n27927), .B(exu_n16233), .Y(exu_n28320));
AND2X1 exu_U36361(.A(exu_n28321), .B(exu_n15402), .Y(exu_n28571));
AND2X1 exu_U36362(.A(exu_n28321), .B(exu_n16223), .Y(exu_n28695));
AND2X1 exu_U36363(.A(div_ecl_d_msb), .B(ecl_div_sel_64b), .Y(exu_n28720));
AND2X1 exu_U36364(.A(div_curr_q[62]), .B(exu_n16252), .Y(exu_n28721));
AND2X1 exu_U36365(.A(div_curr_q[61]), .B(ecl_div_sel_64b), .Y(exu_n28722));
AND2X1 exu_U36366(.A(div_curr_q[60]), .B(ecl_div_sel_64b), .Y(exu_n28723));
AND2X1 exu_U36367(.A(div_curr_q[59]), .B(ecl_div_sel_64b), .Y(exu_n28730));
AND2X1 exu_U36368(.A(div_curr_q[58]), .B(exu_n16252), .Y(exu_n28731));
AND2X1 exu_U36369(.A(div_curr_q[57]), .B(exu_n16252), .Y(exu_n28732));
AND2X1 exu_U36370(.A(div_curr_q[56]), .B(exu_n16252), .Y(exu_n28733));
AND2X1 exu_U36371(.A(div_curr_q[55]), .B(exu_n16252), .Y(exu_n28734));
AND2X1 exu_U36372(.A(div_curr_q[54]), .B(exu_n16252), .Y(exu_n28735));
AND2X1 exu_U36373(.A(div_curr_q[53]), .B(exu_n16252), .Y(exu_n28736));
AND2X1 exu_U36374(.A(div_curr_q[52]), .B(exu_n16252), .Y(exu_n28737));
AND2X1 exu_U36375(.A(div_curr_q[51]), .B(exu_n16252), .Y(exu_n28738));
AND2X1 exu_U36376(.A(div_curr_q[50]), .B(exu_n16252), .Y(exu_n28739));
AND2X1 exu_U36377(.A(div_curr_q[49]), .B(exu_n16252), .Y(exu_n28746));
AND2X1 exu_U36378(.A(div_curr_q[48]), .B(exu_n16252), .Y(exu_n28747));
AND2X1 exu_U36379(.A(div_curr_q[47]), .B(exu_n16252), .Y(exu_n28748));
AND2X1 exu_U36380(.A(div_curr_q[46]), .B(exu_n16252), .Y(exu_n28749));
AND2X1 exu_U36381(.A(div_curr_q[45]), .B(exu_n16252), .Y(exu_n28750));
AND2X1 exu_U36382(.A(div_curr_q[44]), .B(exu_n16252), .Y(exu_n28751));
AND2X1 exu_U36383(.A(div_curr_q[43]), .B(exu_n16252), .Y(exu_n28752));
AND2X1 exu_U36384(.A(div_curr_q[42]), .B(ecl_div_sel_64b), .Y(exu_n28753));
AND2X1 exu_U36385(.A(div_curr_q[41]), .B(exu_n16252), .Y(exu_n28754));
AND2X1 exu_U36386(.A(div_curr_q[40]), .B(exu_n16252), .Y(exu_n28755));
AND2X1 exu_U36387(.A(div_curr_q[39]), .B(ecl_div_sel_64b), .Y(exu_n28762));
AND2X1 exu_U36388(.A(div_curr_q[38]), .B(exu_n16252), .Y(exu_n28763));
AND2X1 exu_U36389(.A(div_curr_q[37]), .B(ecl_div_sel_64b), .Y(exu_n28764));
AND2X1 exu_U36390(.A(div_curr_q[36]), .B(ecl_div_sel_64b), .Y(exu_n28765));
AND2X1 exu_U36391(.A(div_curr_q[35]), .B(exu_n16252), .Y(exu_n28766));
AND2X1 exu_U36392(.A(div_curr_q[34]), .B(exu_n16252), .Y(exu_n28767));
AND2X1 exu_U36393(.A(div_curr_q[33]), .B(ecl_div_sel_64b), .Y(exu_n28768));
AND2X1 exu_U36394(.A(div_curr_q[32]), .B(exu_n16252), .Y(exu_n28769));
AND2X1 exu_U36395(.A(bypass_rd_data_e[6]), .B(exu_n16030), .Y(exu_n29302));
AND2X1 exu_U36396(.A(bypass_rd_data_e[5]), .B(exu_n16030), .Y(exu_n29303));
AND2X1 exu_U36397(.A(bypass_rd_data_e[4]), .B(exu_n16030), .Y(exu_n29304));
AND2X1 exu_U36398(.A(bypass_rd_data_e[3]), .B(exu_n16030), .Y(exu_n29312));
AND2X1 exu_U36399(.A(bypass_rd_data_e[2]), .B(exu_n16029), .Y(exu_n29323));
AND2X1 exu_U36400(.A(bypass_rd_data_e[1]), .B(exu_n16028), .Y(exu_n29334));
AND2X1 exu_U36401(.A(bypass_rd_data_e[31]), .B(exu_n16027), .Y(exu_n29340));
AND2X1 exu_U36402(.A(bypass_rd_data_e[30]), .B(exu_n16027), .Y(exu_n29341));
AND2X1 exu_U36403(.A(bypass_rd_data_e[29]), .B(exu_n16027), .Y(exu_n29342));
AND2X1 exu_U36404(.A(bypass_rd_data_e[28]), .B(exu_n16027), .Y(exu_n29343));
AND2X1 exu_U36405(.A(bypass_rd_data_e[27]), .B(exu_n16027), .Y(exu_n29344));
AND2X1 exu_U36406(.A(bypass_rd_data_e[0]), .B(exu_n16027), .Y(exu_n29345));
AND2X1 exu_U36407(.A(bypass_rd_data_e[26]), .B(exu_n16027), .Y(exu_n29346));
AND2X1 exu_U36408(.A(bypass_rd_data_e[25]), .B(exu_n16027), .Y(exu_n29347));
AND2X1 exu_U36409(.A(bypass_rd_data_e[24]), .B(exu_n16027), .Y(exu_n29348));
AND2X1 exu_U36410(.A(bypass_rd_data_e[23]), .B(exu_n16027), .Y(exu_n29349));
AND2X1 exu_U36411(.A(bypass_rd_data_e[22]), .B(exu_n16027), .Y(exu_n29350));
AND2X1 exu_U36412(.A(bypass_rd_data_e[21]), .B(exu_n16027), .Y(exu_n29351));
AND2X1 exu_U36413(.A(bypass_rd_data_e[20]), .B(exu_n16027), .Y(exu_n29352));
AND2X1 exu_U36414(.A(bypass_rd_data_e[19]), .B(exu_n16026), .Y(exu_n29353));
AND2X1 exu_U36415(.A(bypass_rd_data_e[18]), .B(exu_n16026), .Y(exu_n29354));
AND2X1 exu_U36416(.A(bypass_rd_data_e[17]), .B(exu_n16026), .Y(exu_n29355));
AND2X1 exu_U36417(.A(bypass_rd_data_e[16]), .B(exu_n16026), .Y(exu_n29356));
AND2X1 exu_U36418(.A(bypass_rd_data_e[15]), .B(exu_n16026), .Y(exu_n29357));
AND2X1 exu_U36419(.A(bypass_rd_data_e[14]), .B(exu_n16026), .Y(exu_n29358));
AND2X1 exu_U36420(.A(bypass_rd_data_e[13]), .B(exu_n16026), .Y(exu_n29359));
AND2X1 exu_U36421(.A(bypass_rd_data_e[12]), .B(exu_n16026), .Y(exu_n29360));
AND2X1 exu_U36422(.A(bypass_rd_data_e[11]), .B(exu_n16026), .Y(exu_n29361));
AND2X1 exu_U36423(.A(bypass_rd_data_e[10]), .B(exu_n16026), .Y(exu_n29362));
AND2X1 exu_U36424(.A(bypass_rd_data_e[9]), .B(exu_n16026), .Y(exu_n29363));
AND2X1 exu_U36425(.A(bypass_rd_data_e[8]), .B(exu_n16026), .Y(exu_n29364));
AND2X1 exu_U36426(.A(bypass_rd_data_e[7]), .B(exu_n16026), .Y(exu_n29365));
AND2X1 exu_U36427(.A(bypass_byp_irf_rd_data_m[6]), .B(exu_n16044), .Y(exu_n29432));
AND2X1 exu_U36428(.A(bypass_byp_irf_rd_data_m[5]), .B(exu_n16044), .Y(exu_n29433));
AND2X1 exu_U36429(.A(bypass_byp_irf_rd_data_m[4]), .B(exu_n16044), .Y(exu_n29434));
AND2X1 exu_U36430(.A(bypass_byp_irf_rd_data_m[63]), .B(exu_n16044), .Y(exu_n29435));
AND2X1 exu_U36431(.A(bypass_byp_irf_rd_data_m[62]), .B(exu_n16044), .Y(exu_n29436));
AND2X1 exu_U36432(.A(bypass_byp_irf_rd_data_m[61]), .B(exu_n16044), .Y(exu_n29437));
AND2X1 exu_U36433(.A(bypass_byp_irf_rd_data_m[60]), .B(exu_n16044), .Y(exu_n29438));
AND2X1 exu_U36434(.A(bypass_byp_irf_rd_data_m[59]), .B(exu_n16044), .Y(exu_n29439));
AND2X1 exu_U36435(.A(bypass_byp_irf_rd_data_m[58]), .B(exu_n16044), .Y(exu_n29440));
AND2X1 exu_U36436(.A(bypass_byp_irf_rd_data_m[57]), .B(exu_n16044), .Y(exu_n29441));
AND2X1 exu_U36437(.A(bypass_byp_irf_rd_data_m[3]), .B(exu_n16044), .Y(exu_n29442));
AND2X1 exu_U36438(.A(bypass_byp_irf_rd_data_m[56]), .B(exu_n16044), .Y(exu_n29443));
AND2X1 exu_U36439(.A(bypass_byp_irf_rd_data_m[55]), .B(exu_n16043), .Y(exu_n29444));
AND2X1 exu_U36440(.A(bypass_byp_irf_rd_data_m[54]), .B(exu_n16043), .Y(exu_n29445));
AND2X1 exu_U36441(.A(bypass_byp_irf_rd_data_m[53]), .B(exu_n16043), .Y(exu_n29446));
AND2X1 exu_U36442(.A(bypass_byp_irf_rd_data_m[52]), .B(exu_n16043), .Y(exu_n29447));
AND2X1 exu_U36443(.A(bypass_byp_irf_rd_data_m[51]), .B(exu_n16043), .Y(exu_n29448));
AND2X1 exu_U36444(.A(bypass_byp_irf_rd_data_m[50]), .B(exu_n16043), .Y(exu_n29449));
AND2X1 exu_U36445(.A(bypass_byp_irf_rd_data_m[49]), .B(exu_n16043), .Y(exu_n29450));
AND2X1 exu_U36446(.A(bypass_byp_irf_rd_data_m[48]), .B(exu_n16043), .Y(exu_n29451));
AND2X1 exu_U36447(.A(bypass_byp_irf_rd_data_m[47]), .B(exu_n16043), .Y(exu_n29452));
AND2X1 exu_U36448(.A(bypass_byp_irf_rd_data_m[2]), .B(exu_n16043), .Y(exu_n29453));
AND2X1 exu_U36449(.A(bypass_byp_irf_rd_data_m[46]), .B(exu_n16043), .Y(exu_n29454));
AND2X1 exu_U36450(.A(bypass_byp_irf_rd_data_m[45]), .B(exu_n16043), .Y(exu_n29455));
AND2X1 exu_U36451(.A(bypass_byp_irf_rd_data_m[44]), .B(exu_n16043), .Y(exu_n29456));
AND2X1 exu_U36452(.A(bypass_byp_irf_rd_data_m[43]), .B(exu_n16042), .Y(exu_n29457));
AND2X1 exu_U36453(.A(bypass_byp_irf_rd_data_m[42]), .B(exu_n16042), .Y(exu_n29458));
AND2X1 exu_U36454(.A(bypass_byp_irf_rd_data_m[41]), .B(exu_n16042), .Y(exu_n29459));
AND2X1 exu_U36455(.A(bypass_byp_irf_rd_data_m[40]), .B(exu_n16042), .Y(exu_n29460));
AND2X1 exu_U36456(.A(bypass_byp_irf_rd_data_m[39]), .B(exu_n16042), .Y(exu_n29461));
AND2X1 exu_U36457(.A(bypass_byp_irf_rd_data_m[38]), .B(exu_n16042), .Y(exu_n29462));
AND2X1 exu_U36458(.A(bypass_byp_irf_rd_data_m[37]), .B(exu_n16042), .Y(exu_n29463));
AND2X1 exu_U36459(.A(bypass_byp_irf_rd_data_m[1]), .B(exu_n16042), .Y(exu_n29464));
AND2X1 exu_U36460(.A(bypass_byp_irf_rd_data_m[36]), .B(exu_n16042), .Y(exu_n29465));
AND2X1 exu_U36461(.A(bypass_byp_irf_rd_data_m[35]), .B(exu_n16042), .Y(exu_n29466));
AND2X1 exu_U36462(.A(bypass_byp_irf_rd_data_m[34]), .B(exu_n16042), .Y(exu_n29467));
AND2X1 exu_U36463(.A(bypass_byp_irf_rd_data_m[33]), .B(exu_n16042), .Y(exu_n29468));
AND2X1 exu_U36464(.A(bypass_byp_irf_rd_data_m[32]), .B(exu_n16042), .Y(exu_n29469));
AND2X1 exu_U36465(.A(bypass_byp_irf_rd_data_m[31]), .B(exu_n16041), .Y(exu_n29470));
AND2X1 exu_U36466(.A(bypass_byp_irf_rd_data_m[30]), .B(exu_n16041), .Y(exu_n29471));
AND2X1 exu_U36467(.A(bypass_byp_irf_rd_data_m[29]), .B(exu_n16041), .Y(exu_n29472));
AND2X1 exu_U36468(.A(bypass_byp_irf_rd_data_m[28]), .B(exu_n16041), .Y(exu_n29473));
AND2X1 exu_U36469(.A(bypass_byp_irf_rd_data_m[27]), .B(exu_n16041), .Y(exu_n29474));
AND2X1 exu_U36470(.A(bypass_byp_irf_rd_data_m[0]), .B(exu_n16041), .Y(exu_n29475));
AND2X1 exu_U36471(.A(bypass_byp_irf_rd_data_m[26]), .B(exu_n16041), .Y(exu_n29476));
AND2X1 exu_U36472(.A(bypass_byp_irf_rd_data_m[25]), .B(exu_n16041), .Y(exu_n29477));
AND2X1 exu_U36473(.A(bypass_byp_irf_rd_data_m[24]), .B(exu_n16041), .Y(exu_n29478));
AND2X1 exu_U36474(.A(bypass_byp_irf_rd_data_m[23]), .B(exu_n16041), .Y(exu_n29479));
AND2X1 exu_U36475(.A(bypass_byp_irf_rd_data_m[22]), .B(exu_n16041), .Y(exu_n29480));
AND2X1 exu_U36476(.A(bypass_byp_irf_rd_data_m[21]), .B(exu_n16041), .Y(exu_n29481));
AND2X1 exu_U36477(.A(bypass_byp_irf_rd_data_m[20]), .B(exu_n16041), .Y(exu_n29482));
AND2X1 exu_U36478(.A(bypass_byp_irf_rd_data_m[19]), .B(exu_n16040), .Y(exu_n29483));
AND2X1 exu_U36479(.A(bypass_byp_irf_rd_data_m[18]), .B(exu_n16040), .Y(exu_n29484));
AND2X1 exu_U36480(.A(bypass_byp_irf_rd_data_m[17]), .B(exu_n16040), .Y(exu_n29485));
AND2X1 exu_U36481(.A(bypass_byp_irf_rd_data_m[16]), .B(exu_n16040), .Y(exu_n29486));
AND2X1 exu_U36482(.A(bypass_byp_irf_rd_data_m[15]), .B(exu_n16040), .Y(exu_n29487));
AND2X1 exu_U36483(.A(bypass_byp_irf_rd_data_m[14]), .B(exu_n16040), .Y(exu_n29488));
AND2X1 exu_U36484(.A(bypass_byp_irf_rd_data_m[13]), .B(exu_n16040), .Y(exu_n29489));
AND2X1 exu_U36485(.A(bypass_byp_irf_rd_data_m[12]), .B(exu_n16040), .Y(exu_n29490));
AND2X1 exu_U36486(.A(bypass_byp_irf_rd_data_m[11]), .B(exu_n16040), .Y(exu_n29491));
AND2X1 exu_U36487(.A(bypass_byp_irf_rd_data_m[10]), .B(exu_n16040), .Y(exu_n29492));
AND2X1 exu_U36488(.A(bypass_byp_irf_rd_data_m[9]), .B(exu_n16040), .Y(exu_n29493));
AND2X1 exu_U36489(.A(bypass_byp_irf_rd_data_m[8]), .B(exu_n16040), .Y(exu_n29494));
AND2X1 exu_U36490(.A(bypass_byp_irf_rd_data_m[7]), .B(exu_n16040), .Y(exu_n29495));
AND2X1 exu_U36491(.A(exu_n15854), .B(exu_n16051), .Y(exu_n29497));
AND2X1 exu_U36492(.A(exu_n15833), .B(exu_n16051), .Y(exu_n29498));
AND2X1 exu_U36493(.A(exu_n15801), .B(exu_n16051), .Y(exu_n29499));
AND2X1 exu_U36494(.A(exu_n15826), .B(exu_n16051), .Y(exu_n29500));
AND2X1 exu_U36495(.A(exu_n15796), .B(exu_n16051), .Y(exu_n29501));
AND2X1 exu_U36496(.A(exu_n15779), .B(exu_n16051), .Y(exu_n29502));
AND2X1 exu_U36497(.A(exu_n15780), .B(exu_n16051), .Y(exu_n29503));
AND2X1 exu_U36498(.A(exu_n15797), .B(exu_n16051), .Y(exu_n29504));
AND2X1 exu_U36499(.A(exu_n15811), .B(exu_n16051), .Y(exu_n29505));
AND2X1 exu_U36500(.A(exu_n15798), .B(exu_n16051), .Y(exu_n29506));
AND2X1 exu_U36501(.A(exu_n15843), .B(exu_n16051), .Y(exu_n29507));
AND2X1 exu_U36502(.A(exu_n15834), .B(exu_n16051), .Y(exu_n29508));
AND2X1 exu_U36503(.A(exu_n15799), .B(exu_n16050), .Y(exu_n29509));
AND2X1 exu_U36504(.A(exu_n15781), .B(exu_n16050), .Y(exu_n29510));
AND2X1 exu_U36505(.A(exu_n15827), .B(exu_n16050), .Y(exu_n29511));
AND2X1 exu_U36506(.A(exu_n15812), .B(exu_n16050), .Y(exu_n29512));
AND2X1 exu_U36507(.A(exu_n15835), .B(exu_n16050), .Y(exu_n29513));
AND2X1 exu_U36508(.A(exu_n15800), .B(exu_n16050), .Y(exu_n29514));
AND2X1 exu_U36509(.A(exu_n15782), .B(exu_n16050), .Y(exu_n29515));
AND2X1 exu_U36510(.A(exu_n15783), .B(exu_n16050), .Y(exu_n29516));
AND2X1 exu_U36511(.A(exu_n15802), .B(exu_n16050), .Y(exu_n29517));
AND2X1 exu_U36512(.A(exu_n15831), .B(exu_n16050), .Y(exu_n29518));
AND2X1 exu_U36513(.A(exu_n15855), .B(exu_n16050), .Y(exu_n29519));
AND2X1 exu_U36514(.A(exu_n15784), .B(exu_n16050), .Y(exu_n29520));
AND2X1 exu_U36515(.A(exu_n15841), .B(exu_n16050), .Y(exu_n29521));
AND2X1 exu_U36516(.A(exu_n15785), .B(exu_n16049), .Y(exu_n29522));
AND2X1 exu_U36517(.A(exu_n15803), .B(exu_n16049), .Y(exu_n29523));
AND2X1 exu_U36518(.A(exu_n15828), .B(exu_n16049), .Y(exu_n29524));
AND2X1 exu_U36519(.A(exu_n15842), .B(exu_n16049), .Y(exu_n29525));
AND2X1 exu_U36520(.A(exu_n15844), .B(exu_n16049), .Y(exu_n29526));
AND2X1 exu_U36521(.A(exu_n15829), .B(exu_n16049), .Y(exu_n29527));
AND2X1 exu_U36522(.A(exu_n15786), .B(exu_n16049), .Y(exu_n29528));
AND2X1 exu_U36523(.A(exu_n15813), .B(exu_n16049), .Y(exu_n29529));
AND2X1 exu_U36524(.A(exu_n15927), .B(exu_n16049), .Y(exu_n29530));
AND2X1 exu_U36525(.A(exu_n15787), .B(exu_n16049), .Y(exu_n29531));
AND2X1 exu_U36526(.A(exu_n15804), .B(exu_n16049), .Y(exu_n29532));
AND2X1 exu_U36527(.A(exu_n15788), .B(exu_n16049), .Y(exu_n29533));
AND2X1 exu_U36528(.A(exu_n15928), .B(exu_n16049), .Y(exu_n29534));
AND2X1 exu_U36529(.A(exu_n15830), .B(exu_n16048), .Y(exu_n29535));
AND2X1 exu_U36530(.A(exu_n15845), .B(exu_n16048), .Y(exu_n29536));
AND2X1 exu_U36531(.A(exu_n15789), .B(exu_n16048), .Y(exu_n29537));
AND2X1 exu_U36532(.A(exu_n15846), .B(exu_n16048), .Y(exu_n29538));
AND2X1 exu_U36533(.A(exu_n15805), .B(exu_n16048), .Y(exu_n29539));
AND2X1 exu_U36534(.A(exu_n15810), .B(exu_n16048), .Y(exu_n29540));
AND2X1 exu_U36535(.A(exu_n15806), .B(exu_n16048), .Y(exu_n29541));
AND2X1 exu_U36536(.A(exu_n15836), .B(exu_n16048), .Y(exu_n29542));
AND2X1 exu_U36537(.A(exu_n15837), .B(exu_n16048), .Y(exu_n29543));
AND2X1 exu_U36538(.A(exu_n15807), .B(exu_n16048), .Y(exu_n29544));
AND2X1 exu_U36539(.A(exu_n15790), .B(exu_n16048), .Y(exu_n29545));
AND2X1 exu_U36540(.A(exu_n15847), .B(exu_n16048), .Y(exu_n29546));
AND2X1 exu_U36541(.A(exu_n15791), .B(exu_n16048), .Y(exu_n29547));
AND2X1 exu_U36542(.A(exu_n15808), .B(exu_n16047), .Y(exu_n29548));
AND2X1 exu_U36543(.A(exu_n15792), .B(exu_n16047), .Y(exu_n29549));
AND2X1 exu_U36544(.A(exu_n15929), .B(exu_n16047), .Y(exu_n29550));
AND2X1 exu_U36545(.A(exu_n15832), .B(exu_n16047), .Y(exu_n29551));
AND2X1 exu_U36546(.A(exu_n15848), .B(exu_n16047), .Y(exu_n29552));
AND2X1 exu_U36547(.A(exu_n15793), .B(exu_n16047), .Y(exu_n29553));
AND2X1 exu_U36548(.A(exu_n15849), .B(exu_n16047), .Y(exu_n29554));
AND2X1 exu_U36549(.A(exu_n15809), .B(exu_n16047), .Y(exu_n29555));
AND2X1 exu_U36550(.A(exu_n15838), .B(exu_n16047), .Y(exu_n29556));
AND2X1 exu_U36551(.A(exu_n15850), .B(exu_n16047), .Y(exu_n29557));
AND2X1 exu_U36552(.A(exu_n15418), .B(exu_n16047), .Y(exu_n29558));
AND2X1 exu_U36553(.A(exu_n15840), .B(exu_n16047), .Y(exu_n29559));
AND2X1 exu_U36554(.A(exu_n15825), .B(exu_n16047), .Y(exu_n29560));
AND2X1 exu_U36555(.A(bypass_byp_alu_rs1_data_d[6]), .B(exu_n16058), .Y(exu_n29562));
AND2X1 exu_U36556(.A(bypass_byp_alu_rs1_data_d[5]), .B(exu_n16058), .Y(exu_n29563));
AND2X1 exu_U36557(.A(bypass_byp_alu_rs1_data_d[4]), .B(exu_n16058), .Y(exu_n29564));
AND2X1 exu_U36558(.A(bypass_byp_alu_rs1_data_d[63]), .B(exu_n16058), .Y(exu_n29565));
AND2X1 exu_U36559(.A(bypass_byp_alu_rs1_data_d[62]), .B(exu_n16058), .Y(exu_n29566));
AND2X1 exu_U36560(.A(bypass_byp_alu_rs1_data_d[61]), .B(exu_n16058), .Y(exu_n29567));
AND2X1 exu_U36561(.A(bypass_byp_alu_rs1_data_d[60]), .B(exu_n16058), .Y(exu_n29568));
AND2X1 exu_U36562(.A(bypass_byp_alu_rs1_data_d[59]), .B(exu_n16058), .Y(exu_n29569));
AND2X1 exu_U36563(.A(bypass_byp_alu_rs1_data_d[58]), .B(exu_n16058), .Y(exu_n29570));
AND2X1 exu_U36564(.A(bypass_byp_alu_rs1_data_d[57]), .B(exu_n16058), .Y(exu_n29571));
AND2X1 exu_U36565(.A(bypass_byp_alu_rs1_data_d[3]), .B(exu_n16058), .Y(exu_n29572));
AND2X1 exu_U36566(.A(bypass_byp_alu_rs1_data_d[56]), .B(exu_n16058), .Y(exu_n29573));
AND2X1 exu_U36567(.A(bypass_byp_alu_rs1_data_d[55]), .B(exu_n16057), .Y(exu_n29574));
AND2X1 exu_U36568(.A(bypass_byp_alu_rs1_data_d[54]), .B(exu_n16057), .Y(exu_n29575));
AND2X1 exu_U36569(.A(bypass_byp_alu_rs1_data_d[53]), .B(exu_n16057), .Y(exu_n29576));
AND2X1 exu_U36570(.A(bypass_byp_alu_rs1_data_d[52]), .B(exu_n16057), .Y(exu_n29577));
AND2X1 exu_U36571(.A(bypass_byp_alu_rs1_data_d[51]), .B(exu_n16057), .Y(exu_n29578));
AND2X1 exu_U36572(.A(bypass_byp_alu_rs1_data_d[50]), .B(exu_n16057), .Y(exu_n29579));
AND2X1 exu_U36573(.A(bypass_byp_alu_rs1_data_d[49]), .B(exu_n16057), .Y(exu_n29580));
AND2X1 exu_U36574(.A(bypass_byp_alu_rs1_data_d[48]), .B(exu_n16057), .Y(exu_n29581));
AND2X1 exu_U36575(.A(bypass_byp_alu_rs1_data_d[47]), .B(exu_n16057), .Y(exu_n29582));
AND2X1 exu_U36576(.A(bypass_byp_alu_rs1_data_d[2]), .B(exu_n16057), .Y(exu_n29583));
AND2X1 exu_U36577(.A(bypass_byp_alu_rs1_data_d[46]), .B(exu_n16057), .Y(exu_n29584));
AND2X1 exu_U36578(.A(bypass_byp_alu_rs1_data_d[45]), .B(exu_n16057), .Y(exu_n29585));
AND2X1 exu_U36579(.A(bypass_byp_alu_rs1_data_d[44]), .B(exu_n16057), .Y(exu_n29586));
AND2X1 exu_U36580(.A(bypass_byp_alu_rs1_data_d[43]), .B(exu_n16056), .Y(exu_n29587));
AND2X1 exu_U36581(.A(bypass_byp_alu_rs1_data_d[42]), .B(exu_n16056), .Y(exu_n29588));
AND2X1 exu_U36582(.A(bypass_byp_alu_rs1_data_d[41]), .B(exu_n16056), .Y(exu_n29589));
AND2X1 exu_U36583(.A(bypass_byp_alu_rs1_data_d[40]), .B(exu_n16056), .Y(exu_n29590));
AND2X1 exu_U36584(.A(bypass_byp_alu_rs1_data_d[39]), .B(exu_n16056), .Y(exu_n29591));
AND2X1 exu_U36585(.A(bypass_byp_alu_rs1_data_d[38]), .B(exu_n16056), .Y(exu_n29592));
AND2X1 exu_U36586(.A(bypass_byp_alu_rs1_data_d[37]), .B(exu_n16056), .Y(exu_n29593));
AND2X1 exu_U36587(.A(bypass_byp_alu_rs1_data_d[1]), .B(exu_n16056), .Y(exu_n29594));
AND2X1 exu_U36588(.A(bypass_byp_alu_rs1_data_d[36]), .B(exu_n16056), .Y(exu_n29595));
AND2X1 exu_U36589(.A(bypass_byp_alu_rs1_data_d[35]), .B(exu_n16056), .Y(exu_n29596));
AND2X1 exu_U36590(.A(bypass_byp_alu_rs1_data_d[34]), .B(exu_n16056), .Y(exu_n29597));
AND2X1 exu_U36591(.A(bypass_byp_alu_rs1_data_d[33]), .B(exu_n16056), .Y(exu_n29598));
AND2X1 exu_U36592(.A(bypass_byp_alu_rs1_data_d[32]), .B(exu_n16056), .Y(exu_n29599));
AND2X1 exu_U36593(.A(bypass_byp_alu_rs1_data_d[31]), .B(exu_n16055), .Y(exu_n29600));
AND2X1 exu_U36594(.A(bypass_byp_alu_rs1_data_d[30]), .B(exu_n16055), .Y(exu_n29601));
AND2X1 exu_U36595(.A(bypass_byp_alu_rs1_data_d[29]), .B(exu_n16055), .Y(exu_n29602));
AND2X1 exu_U36596(.A(bypass_byp_alu_rs1_data_d[28]), .B(exu_n16055), .Y(exu_n29603));
AND2X1 exu_U36597(.A(bypass_byp_alu_rs1_data_d[27]), .B(exu_n16055), .Y(exu_n29604));
AND2X1 exu_U36598(.A(bypass_byp_alu_rs1_data_d[0]), .B(exu_n16055), .Y(exu_n29605));
AND2X1 exu_U36599(.A(bypass_byp_alu_rs1_data_d[26]), .B(exu_n16055), .Y(exu_n29606));
AND2X1 exu_U36600(.A(bypass_byp_alu_rs1_data_d[25]), .B(exu_n16055), .Y(exu_n29607));
AND2X1 exu_U36601(.A(bypass_byp_alu_rs1_data_d[24]), .B(exu_n16055), .Y(exu_n29608));
AND2X1 exu_U36602(.A(bypass_byp_alu_rs1_data_d[23]), .B(exu_n16055), .Y(exu_n29609));
AND2X1 exu_U36603(.A(bypass_byp_alu_rs1_data_d[22]), .B(exu_n16055), .Y(exu_n29610));
AND2X1 exu_U36604(.A(bypass_byp_alu_rs1_data_d[21]), .B(exu_n16055), .Y(exu_n29611));
AND2X1 exu_U36605(.A(bypass_byp_alu_rs1_data_d[20]), .B(exu_n16055), .Y(exu_n29612));
AND2X1 exu_U36606(.A(bypass_byp_alu_rs1_data_d[19]), .B(exu_n16054), .Y(exu_n29613));
AND2X1 exu_U36607(.A(bypass_byp_alu_rs1_data_d[18]), .B(exu_n16054), .Y(exu_n29614));
AND2X1 exu_U36608(.A(bypass_byp_alu_rs1_data_d[17]), .B(exu_n16054), .Y(exu_n29615));
AND2X1 exu_U36609(.A(bypass_byp_alu_rs1_data_d[16]), .B(exu_n16054), .Y(exu_n29616));
AND2X1 exu_U36610(.A(bypass_byp_alu_rs1_data_d[15]), .B(exu_n16054), .Y(exu_n29617));
AND2X1 exu_U36611(.A(bypass_byp_alu_rs1_data_d[14]), .B(exu_n16054), .Y(exu_n29618));
AND2X1 exu_U36612(.A(bypass_byp_alu_rs1_data_d[13]), .B(exu_n16054), .Y(exu_n29619));
AND2X1 exu_U36613(.A(bypass_byp_alu_rs1_data_d[12]), .B(exu_n16054), .Y(exu_n29620));
AND2X1 exu_U36614(.A(bypass_byp_alu_rs1_data_d[11]), .B(exu_n16054), .Y(exu_n29621));
AND2X1 exu_U36615(.A(bypass_byp_alu_rs1_data_d[10]), .B(exu_n16054), .Y(exu_n29622));
AND2X1 exu_U36616(.A(bypass_byp_alu_rs1_data_d[9]), .B(exu_n16054), .Y(exu_n29623));
AND2X1 exu_U36617(.A(bypass_byp_alu_rs1_data_d[8]), .B(exu_n16054), .Y(exu_n29624));
AND2X1 exu_U36618(.A(bypass_byp_alu_rs1_data_d[7]), .B(exu_n16054), .Y(exu_n29625));
AND2X1 exu_U36619(.A(bypass_byp_alu_rs2_data_d[6]), .B(exu_n16065), .Y(exu_n29627));
AND2X1 exu_U36620(.A(bypass_byp_alu_rs2_data_d[5]), .B(exu_n16065), .Y(exu_n29628));
AND2X1 exu_U36621(.A(bypass_byp_alu_rs2_data_d[4]), .B(exu_n16065), .Y(exu_n29629));
AND2X1 exu_U36622(.A(bypass_byp_alu_rs2_data_d[63]), .B(exu_n16065), .Y(exu_n29630));
AND2X1 exu_U36623(.A(bypass_byp_alu_rs2_data_d[62]), .B(exu_n16065), .Y(exu_n29631));
AND2X1 exu_U36624(.A(bypass_byp_alu_rs2_data_d[61]), .B(exu_n16065), .Y(exu_n29632));
AND2X1 exu_U36625(.A(bypass_byp_alu_rs2_data_d[60]), .B(exu_n16065), .Y(exu_n29633));
AND2X1 exu_U36626(.A(bypass_byp_alu_rs2_data_d[59]), .B(exu_n16065), .Y(exu_n29634));
AND2X1 exu_U36627(.A(bypass_byp_alu_rs2_data_d[58]), .B(exu_n16065), .Y(exu_n29635));
AND2X1 exu_U36628(.A(bypass_byp_alu_rs2_data_d[57]), .B(exu_n16065), .Y(exu_n29636));
AND2X1 exu_U36629(.A(bypass_byp_alu_rs2_data_d[3]), .B(exu_n16065), .Y(exu_n29637));
AND2X1 exu_U36630(.A(bypass_byp_alu_rs2_data_d[56]), .B(exu_n16065), .Y(exu_n29638));
AND2X1 exu_U36631(.A(bypass_byp_alu_rs2_data_d[55]), .B(exu_n16064), .Y(exu_n29639));
AND2X1 exu_U36632(.A(bypass_byp_alu_rs2_data_d[54]), .B(exu_n16064), .Y(exu_n29640));
AND2X1 exu_U36633(.A(bypass_byp_alu_rs2_data_d[53]), .B(exu_n16064), .Y(exu_n29641));
AND2X1 exu_U36634(.A(bypass_byp_alu_rs2_data_d[52]), .B(exu_n16064), .Y(exu_n29642));
AND2X1 exu_U36635(.A(bypass_byp_alu_rs2_data_d[51]), .B(exu_n16064), .Y(exu_n29643));
AND2X1 exu_U36636(.A(bypass_byp_alu_rs2_data_d[50]), .B(exu_n16064), .Y(exu_n29644));
AND2X1 exu_U36637(.A(bypass_byp_alu_rs2_data_d[49]), .B(exu_n16064), .Y(exu_n29645));
AND2X1 exu_U36638(.A(bypass_byp_alu_rs2_data_d[48]), .B(exu_n16064), .Y(exu_n29646));
AND2X1 exu_U36639(.A(bypass_byp_alu_rs2_data_d[47]), .B(exu_n16064), .Y(exu_n29647));
AND2X1 exu_U36640(.A(bypass_byp_alu_rs2_data_d[2]), .B(exu_n16064), .Y(exu_n29648));
AND2X1 exu_U36641(.A(bypass_byp_alu_rs2_data_d[46]), .B(exu_n16064), .Y(exu_n29649));
AND2X1 exu_U36642(.A(bypass_byp_alu_rs2_data_d[45]), .B(exu_n16064), .Y(exu_n29650));
AND2X1 exu_U36643(.A(bypass_byp_alu_rs2_data_d[44]), .B(exu_n16064), .Y(exu_n29651));
AND2X1 exu_U36644(.A(bypass_byp_alu_rs2_data_d[43]), .B(exu_n16063), .Y(exu_n29652));
AND2X1 exu_U36645(.A(bypass_byp_alu_rs2_data_d[42]), .B(exu_n16063), .Y(exu_n29653));
AND2X1 exu_U36646(.A(bypass_byp_alu_rs2_data_d[41]), .B(exu_n16063), .Y(exu_n29654));
AND2X1 exu_U36647(.A(bypass_byp_alu_rs2_data_d[40]), .B(exu_n16063), .Y(exu_n29655));
AND2X1 exu_U36648(.A(bypass_byp_alu_rs2_data_d[39]), .B(exu_n16063), .Y(exu_n29656));
AND2X1 exu_U36649(.A(bypass_byp_alu_rs2_data_d[38]), .B(exu_n16063), .Y(exu_n29657));
AND2X1 exu_U36650(.A(bypass_byp_alu_rs2_data_d[37]), .B(exu_n16063), .Y(exu_n29658));
AND2X1 exu_U36651(.A(bypass_byp_alu_rs2_data_d[1]), .B(exu_n16063), .Y(exu_n29659));
AND2X1 exu_U36652(.A(bypass_byp_alu_rs2_data_d[36]), .B(exu_n16063), .Y(exu_n29660));
AND2X1 exu_U36653(.A(bypass_byp_alu_rs2_data_d[35]), .B(exu_n16063), .Y(exu_n29661));
AND2X1 exu_U36654(.A(bypass_byp_alu_rs2_data_d[34]), .B(exu_n16063), .Y(exu_n29662));
AND2X1 exu_U36655(.A(bypass_byp_alu_rs2_data_d[33]), .B(exu_n16063), .Y(exu_n29663));
AND2X1 exu_U36656(.A(bypass_byp_alu_rs2_data_d[32]), .B(exu_n16063), .Y(exu_n29664));
AND2X1 exu_U36657(.A(bypass_byp_alu_rs2_data_d[31]), .B(exu_n16062), .Y(exu_n29665));
AND2X1 exu_U36658(.A(bypass_byp_alu_rs2_data_d[30]), .B(exu_n16062), .Y(exu_n29666));
AND2X1 exu_U36659(.A(bypass_byp_alu_rs2_data_d[29]), .B(exu_n16062), .Y(exu_n29667));
AND2X1 exu_U36660(.A(bypass_byp_alu_rs2_data_d[28]), .B(exu_n16062), .Y(exu_n29668));
AND2X1 exu_U36661(.A(bypass_byp_alu_rs2_data_d[27]), .B(exu_n16062), .Y(exu_n29669));
AND2X1 exu_U36662(.A(bypass_byp_alu_rs2_data_d[0]), .B(exu_n16062), .Y(exu_n29670));
AND2X1 exu_U36663(.A(bypass_byp_alu_rs2_data_d[26]), .B(exu_n16062), .Y(exu_n29671));
AND2X1 exu_U36664(.A(bypass_byp_alu_rs2_data_d[25]), .B(exu_n16062), .Y(exu_n29672));
AND2X1 exu_U36665(.A(bypass_byp_alu_rs2_data_d[24]), .B(exu_n16062), .Y(exu_n29673));
AND2X1 exu_U36666(.A(bypass_byp_alu_rs2_data_d[23]), .B(exu_n16062), .Y(exu_n29674));
AND2X1 exu_U36667(.A(bypass_byp_alu_rs2_data_d[22]), .B(exu_n16062), .Y(exu_n29675));
AND2X1 exu_U36668(.A(bypass_byp_alu_rs2_data_d[21]), .B(exu_n16062), .Y(exu_n29676));
AND2X1 exu_U36669(.A(bypass_byp_alu_rs2_data_d[20]), .B(exu_n16062), .Y(exu_n29677));
AND2X1 exu_U36670(.A(bypass_byp_alu_rs2_data_d[19]), .B(exu_n16061), .Y(exu_n29678));
AND2X1 exu_U36671(.A(bypass_byp_alu_rs2_data_d[18]), .B(exu_n16061), .Y(exu_n29679));
AND2X1 exu_U36672(.A(bypass_byp_alu_rs2_data_d[17]), .B(exu_n16061), .Y(exu_n29680));
AND2X1 exu_U36673(.A(bypass_byp_alu_rs2_data_d[16]), .B(exu_n16061), .Y(exu_n29681));
AND2X1 exu_U36674(.A(bypass_byp_alu_rs2_data_d[15]), .B(exu_n16061), .Y(exu_n29682));
AND2X1 exu_U36675(.A(bypass_byp_alu_rs2_data_d[14]), .B(exu_n16061), .Y(exu_n29683));
AND2X1 exu_U36676(.A(bypass_byp_alu_rs2_data_d[13]), .B(exu_n16061), .Y(exu_n29684));
AND2X1 exu_U36677(.A(bypass_byp_alu_rs2_data_d[12]), .B(exu_n16061), .Y(exu_n29685));
AND2X1 exu_U36678(.A(bypass_byp_alu_rs2_data_d[11]), .B(exu_n16061), .Y(exu_n29686));
AND2X1 exu_U36679(.A(bypass_byp_alu_rs2_data_d[10]), .B(exu_n16061), .Y(exu_n29687));
AND2X1 exu_U36680(.A(bypass_byp_alu_rs2_data_d[9]), .B(exu_n16061), .Y(exu_n29688));
AND2X1 exu_U36681(.A(bypass_byp_alu_rs2_data_d[8]), .B(exu_n16061), .Y(exu_n29689));
AND2X1 exu_U36682(.A(bypass_byp_alu_rs2_data_d[7]), .B(exu_n16061), .Y(exu_n29690));
AND2X1 exu_U36683(.A(bypass_rs3_data_d[6]), .B(exu_n16072), .Y(exu_n29692));
AND2X1 exu_U36684(.A(bypass_rs3_data_d[5]), .B(exu_n16072), .Y(exu_n29693));
AND2X1 exu_U36685(.A(bypass_rs3_data_d[4]), .B(exu_n16072), .Y(exu_n29694));
AND2X1 exu_U36686(.A(bypass_rs3_data_d[63]), .B(exu_n16072), .Y(exu_n29695));
AND2X1 exu_U36687(.A(bypass_rs3_data_d[62]), .B(exu_n16072), .Y(exu_n29696));
AND2X1 exu_U36688(.A(bypass_rs3_data_d[61]), .B(exu_n16072), .Y(exu_n29697));
AND2X1 exu_U36689(.A(bypass_rs3_data_d[60]), .B(exu_n16072), .Y(exu_n29698));
AND2X1 exu_U36690(.A(bypass_rs3_data_d[59]), .B(exu_n16072), .Y(exu_n29699));
AND2X1 exu_U36691(.A(bypass_rs3_data_d[58]), .B(exu_n16072), .Y(exu_n29700));
AND2X1 exu_U36692(.A(bypass_rs3_data_d[57]), .B(exu_n16072), .Y(exu_n29701));
AND2X1 exu_U36693(.A(bypass_rs3_data_d[3]), .B(exu_n16072), .Y(exu_n29702));
AND2X1 exu_U36694(.A(bypass_rs3_data_d[56]), .B(exu_n16072), .Y(exu_n29703));
AND2X1 exu_U36695(.A(bypass_rs3_data_d[55]), .B(exu_n16071), .Y(exu_n29704));
AND2X1 exu_U36696(.A(bypass_rs3_data_d[54]), .B(exu_n16071), .Y(exu_n29705));
AND2X1 exu_U36697(.A(bypass_rs3_data_d[53]), .B(exu_n16071), .Y(exu_n29706));
AND2X1 exu_U36698(.A(bypass_rs3_data_d[52]), .B(exu_n16071), .Y(exu_n29707));
AND2X1 exu_U36699(.A(bypass_rs3_data_d[51]), .B(exu_n16071), .Y(exu_n29708));
AND2X1 exu_U36700(.A(bypass_rs3_data_d[50]), .B(exu_n16071), .Y(exu_n29709));
AND2X1 exu_U36701(.A(bypass_rs3_data_d[49]), .B(exu_n16071), .Y(exu_n29710));
AND2X1 exu_U36702(.A(bypass_rs3_data_d[48]), .B(exu_n16071), .Y(exu_n29711));
AND2X1 exu_U36703(.A(bypass_rs3_data_d[47]), .B(exu_n16071), .Y(exu_n29712));
AND2X1 exu_U36704(.A(bypass_rs3_data_d[2]), .B(exu_n16071), .Y(exu_n29713));
AND2X1 exu_U36705(.A(bypass_rs3_data_d[46]), .B(exu_n16071), .Y(exu_n29714));
AND2X1 exu_U36706(.A(bypass_rs3_data_d[45]), .B(exu_n16071), .Y(exu_n29715));
AND2X1 exu_U36707(.A(bypass_rs3_data_d[44]), .B(exu_n16071), .Y(exu_n29716));
AND2X1 exu_U36708(.A(bypass_rs3_data_d[43]), .B(exu_n16070), .Y(exu_n29717));
AND2X1 exu_U36709(.A(bypass_rs3_data_d[42]), .B(exu_n16070), .Y(exu_n29718));
AND2X1 exu_U36710(.A(bypass_rs3_data_d[41]), .B(exu_n16070), .Y(exu_n29719));
AND2X1 exu_U36711(.A(bypass_rs3_data_d[40]), .B(exu_n16070), .Y(exu_n29720));
AND2X1 exu_U36712(.A(bypass_rs3_data_d[39]), .B(exu_n16070), .Y(exu_n29721));
AND2X1 exu_U36713(.A(bypass_rs3_data_d[38]), .B(exu_n16070), .Y(exu_n29722));
AND2X1 exu_U36714(.A(bypass_rs3_data_d[37]), .B(exu_n16070), .Y(exu_n29723));
AND2X1 exu_U36715(.A(bypass_rs3_data_d[1]), .B(exu_n16070), .Y(exu_n29724));
AND2X1 exu_U36716(.A(bypass_rs3_data_d[36]), .B(exu_n16070), .Y(exu_n29725));
AND2X1 exu_U36717(.A(bypass_rs3_data_d[35]), .B(exu_n16070), .Y(exu_n29726));
AND2X1 exu_U36718(.A(bypass_rs3_data_d[34]), .B(exu_n16070), .Y(exu_n29727));
AND2X1 exu_U36719(.A(bypass_rs3_data_d[33]), .B(exu_n16070), .Y(exu_n29728));
AND2X1 exu_U36720(.A(bypass_rs3_data_d[32]), .B(exu_n16070), .Y(exu_n29729));
AND2X1 exu_U36721(.A(bypass_rs3_data_d[31]), .B(exu_n16069), .Y(exu_n29730));
AND2X1 exu_U36722(.A(bypass_rs3_data_d[30]), .B(exu_n16069), .Y(exu_n29731));
AND2X1 exu_U36723(.A(bypass_rs3_data_d[29]), .B(exu_n16069), .Y(exu_n29732));
AND2X1 exu_U36724(.A(bypass_rs3_data_d[28]), .B(exu_n16069), .Y(exu_n29733));
AND2X1 exu_U36725(.A(bypass_rs3_data_d[27]), .B(exu_n16069), .Y(exu_n29734));
AND2X1 exu_U36726(.A(bypass_rs3_data_d[0]), .B(exu_n16069), .Y(exu_n29735));
AND2X1 exu_U36727(.A(bypass_rs3_data_d[26]), .B(exu_n16069), .Y(exu_n29736));
AND2X1 exu_U36728(.A(bypass_rs3_data_d[25]), .B(exu_n16069), .Y(exu_n29737));
AND2X1 exu_U36729(.A(bypass_rs3_data_d[24]), .B(exu_n16069), .Y(exu_n29738));
AND2X1 exu_U36730(.A(bypass_rs3_data_d[23]), .B(exu_n16069), .Y(exu_n29739));
AND2X1 exu_U36731(.A(bypass_rs3_data_d[22]), .B(exu_n16069), .Y(exu_n29740));
AND2X1 exu_U36732(.A(bypass_rs3_data_d[21]), .B(exu_n16069), .Y(exu_n29741));
AND2X1 exu_U36733(.A(bypass_rs3_data_d[20]), .B(exu_n16069), .Y(exu_n29742));
AND2X1 exu_U36734(.A(bypass_rs3_data_d[19]), .B(exu_n16068), .Y(exu_n29743));
AND2X1 exu_U36735(.A(bypass_rs3_data_d[18]), .B(exu_n16068), .Y(exu_n29744));
AND2X1 exu_U36736(.A(bypass_rs3_data_d[17]), .B(exu_n16068), .Y(exu_n29745));
AND2X1 exu_U36737(.A(bypass_rs3_data_d[16]), .B(exu_n16068), .Y(exu_n29746));
AND2X1 exu_U36738(.A(bypass_rs3_data_d[15]), .B(exu_n16068), .Y(exu_n29747));
AND2X1 exu_U36739(.A(bypass_rs3_data_d[14]), .B(exu_n16068), .Y(exu_n29748));
AND2X1 exu_U36740(.A(bypass_rs3_data_d[13]), .B(exu_n16068), .Y(exu_n29749));
AND2X1 exu_U36741(.A(bypass_rs3_data_d[12]), .B(exu_n16068), .Y(exu_n29750));
AND2X1 exu_U36742(.A(bypass_rs3_data_d[11]), .B(exu_n16068), .Y(exu_n29751));
AND2X1 exu_U36743(.A(bypass_rs3_data_d[10]), .B(exu_n16068), .Y(exu_n29752));
AND2X1 exu_U36744(.A(bypass_rs3_data_d[9]), .B(exu_n16068), .Y(exu_n29753));
AND2X1 exu_U36745(.A(bypass_rs3_data_d[8]), .B(exu_n16068), .Y(exu_n29754));
AND2X1 exu_U36746(.A(bypass_rs3_data_d[7]), .B(exu_n16068), .Y(exu_n29755));
AND2X1 exu_U36747(.A(bypass_byp_alu_rcc_data_d[6]), .B(exu_n16079), .Y(exu_n29757));
AND2X1 exu_U36748(.A(bypass_byp_alu_rcc_data_d[5]), .B(exu_n16079), .Y(exu_n29758));
AND2X1 exu_U36749(.A(bypass_byp_alu_rcc_data_d[4]), .B(exu_n16079), .Y(exu_n29759));
AND2X1 exu_U36750(.A(bypass_byp_alu_rcc_data_d[63]), .B(exu_n16079), .Y(exu_n29760));
AND2X1 exu_U36751(.A(bypass_byp_alu_rcc_data_d[62]), .B(exu_n16079), .Y(exu_n29761));
AND2X1 exu_U36752(.A(bypass_byp_alu_rcc_data_d[61]), .B(exu_n16079), .Y(exu_n29762));
AND2X1 exu_U36753(.A(bypass_byp_alu_rcc_data_d[60]), .B(exu_n16079), .Y(exu_n29763));
AND2X1 exu_U36754(.A(bypass_byp_alu_rcc_data_d[59]), .B(exu_n16079), .Y(exu_n29764));
AND2X1 exu_U36755(.A(bypass_byp_alu_rcc_data_d[58]), .B(exu_n16079), .Y(exu_n29765));
AND2X1 exu_U36756(.A(bypass_byp_alu_rcc_data_d[57]), .B(exu_n16079), .Y(exu_n29766));
AND2X1 exu_U36757(.A(bypass_byp_alu_rcc_data_d[3]), .B(exu_n16079), .Y(exu_n29767));
AND2X1 exu_U36758(.A(bypass_byp_alu_rcc_data_d[56]), .B(exu_n16079), .Y(exu_n29768));
AND2X1 exu_U36759(.A(bypass_byp_alu_rcc_data_d[55]), .B(exu_n16078), .Y(exu_n29769));
AND2X1 exu_U36760(.A(bypass_byp_alu_rcc_data_d[54]), .B(exu_n16078), .Y(exu_n29770));
AND2X1 exu_U36761(.A(bypass_byp_alu_rcc_data_d[53]), .B(exu_n16078), .Y(exu_n29771));
AND2X1 exu_U36762(.A(bypass_byp_alu_rcc_data_d[52]), .B(exu_n16078), .Y(exu_n29772));
AND2X1 exu_U36763(.A(bypass_byp_alu_rcc_data_d[51]), .B(exu_n16078), .Y(exu_n29773));
AND2X1 exu_U36764(.A(bypass_byp_alu_rcc_data_d[50]), .B(exu_n16078), .Y(exu_n29774));
AND2X1 exu_U36765(.A(bypass_byp_alu_rcc_data_d[49]), .B(exu_n16078), .Y(exu_n29775));
AND2X1 exu_U36766(.A(bypass_byp_alu_rcc_data_d[48]), .B(exu_n16078), .Y(exu_n29776));
AND2X1 exu_U36767(.A(bypass_byp_alu_rcc_data_d[47]), .B(exu_n16078), .Y(exu_n29777));
AND2X1 exu_U36768(.A(bypass_byp_alu_rcc_data_d[2]), .B(exu_n16078), .Y(exu_n29778));
AND2X1 exu_U36769(.A(bypass_byp_alu_rcc_data_d[46]), .B(exu_n16078), .Y(exu_n29779));
AND2X1 exu_U36770(.A(bypass_byp_alu_rcc_data_d[45]), .B(exu_n16078), .Y(exu_n29780));
AND2X1 exu_U36771(.A(bypass_byp_alu_rcc_data_d[44]), .B(exu_n16078), .Y(exu_n29781));
AND2X1 exu_U36772(.A(bypass_byp_alu_rcc_data_d[43]), .B(exu_n16077), .Y(exu_n29782));
AND2X1 exu_U36773(.A(bypass_byp_alu_rcc_data_d[42]), .B(exu_n16077), .Y(exu_n29783));
AND2X1 exu_U36774(.A(bypass_byp_alu_rcc_data_d[41]), .B(exu_n16077), .Y(exu_n29784));
AND2X1 exu_U36775(.A(bypass_byp_alu_rcc_data_d[40]), .B(exu_n16077), .Y(exu_n29785));
AND2X1 exu_U36776(.A(bypass_byp_alu_rcc_data_d[39]), .B(exu_n16077), .Y(exu_n29786));
AND2X1 exu_U36777(.A(bypass_byp_alu_rcc_data_d[38]), .B(exu_n16077), .Y(exu_n29787));
AND2X1 exu_U36778(.A(bypass_byp_alu_rcc_data_d[37]), .B(exu_n16077), .Y(exu_n29788));
AND2X1 exu_U36779(.A(bypass_byp_alu_rcc_data_d[1]), .B(exu_n16077), .Y(exu_n29789));
AND2X1 exu_U36780(.A(bypass_byp_alu_rcc_data_d[36]), .B(exu_n16077), .Y(exu_n29790));
AND2X1 exu_U36781(.A(bypass_byp_alu_rcc_data_d[35]), .B(exu_n16077), .Y(exu_n29791));
AND2X1 exu_U36782(.A(bypass_byp_alu_rcc_data_d[34]), .B(exu_n16077), .Y(exu_n29792));
AND2X1 exu_U36783(.A(bypass_byp_alu_rcc_data_d[33]), .B(exu_n16077), .Y(exu_n29793));
AND2X1 exu_U36784(.A(bypass_byp_alu_rcc_data_d[32]), .B(exu_n16077), .Y(exu_n29794));
AND2X1 exu_U36785(.A(bypass_byp_alu_rcc_data_d[31]), .B(exu_n16076), .Y(exu_n29795));
AND2X1 exu_U36786(.A(bypass_byp_alu_rcc_data_d[30]), .B(exu_n16076), .Y(exu_n29796));
AND2X1 exu_U36787(.A(bypass_byp_alu_rcc_data_d[29]), .B(exu_n16076), .Y(exu_n29797));
AND2X1 exu_U36788(.A(bypass_byp_alu_rcc_data_d[28]), .B(exu_n16076), .Y(exu_n29798));
AND2X1 exu_U36789(.A(bypass_byp_alu_rcc_data_d[27]), .B(exu_n16076), .Y(exu_n29799));
AND2X1 exu_U36790(.A(bypass_byp_alu_rcc_data_d[0]), .B(exu_n16076), .Y(exu_n29800));
AND2X1 exu_U36791(.A(bypass_byp_alu_rcc_data_d[26]), .B(exu_n16076), .Y(exu_n29801));
AND2X1 exu_U36792(.A(bypass_byp_alu_rcc_data_d[25]), .B(exu_n16076), .Y(exu_n29802));
AND2X1 exu_U36793(.A(bypass_byp_alu_rcc_data_d[24]), .B(exu_n16076), .Y(exu_n29803));
AND2X1 exu_U36794(.A(bypass_byp_alu_rcc_data_d[23]), .B(exu_n16076), .Y(exu_n29804));
AND2X1 exu_U36795(.A(bypass_byp_alu_rcc_data_d[22]), .B(exu_n16076), .Y(exu_n29805));
AND2X1 exu_U36796(.A(bypass_byp_alu_rcc_data_d[21]), .B(exu_n16076), .Y(exu_n29806));
AND2X1 exu_U36797(.A(bypass_byp_alu_rcc_data_d[20]), .B(exu_n16076), .Y(exu_n29807));
AND2X1 exu_U36798(.A(bypass_byp_alu_rcc_data_d[19]), .B(exu_n16075), .Y(exu_n29808));
AND2X1 exu_U36799(.A(bypass_byp_alu_rcc_data_d[18]), .B(exu_n16075), .Y(exu_n29809));
AND2X1 exu_U36800(.A(bypass_byp_alu_rcc_data_d[17]), .B(exu_n16075), .Y(exu_n29810));
AND2X1 exu_U36801(.A(bypass_byp_alu_rcc_data_d[16]), .B(exu_n16075), .Y(exu_n29811));
AND2X1 exu_U36802(.A(bypass_byp_alu_rcc_data_d[15]), .B(exu_n16075), .Y(exu_n29812));
AND2X1 exu_U36803(.A(bypass_byp_alu_rcc_data_d[14]), .B(exu_n16075), .Y(exu_n29813));
AND2X1 exu_U36804(.A(bypass_byp_alu_rcc_data_d[13]), .B(exu_n16075), .Y(exu_n29814));
AND2X1 exu_U36805(.A(bypass_byp_alu_rcc_data_d[12]), .B(exu_n16075), .Y(exu_n29815));
AND2X1 exu_U36806(.A(bypass_byp_alu_rcc_data_d[11]), .B(exu_n16075), .Y(exu_n29816));
AND2X1 exu_U36807(.A(bypass_byp_alu_rcc_data_d[10]), .B(exu_n16075), .Y(exu_n29817));
AND2X1 exu_U36808(.A(bypass_byp_alu_rcc_data_d[9]), .B(exu_n16075), .Y(exu_n29818));
AND2X1 exu_U36809(.A(bypass_byp_alu_rcc_data_d[8]), .B(exu_n16075), .Y(exu_n29819));
AND2X1 exu_U36810(.A(bypass_byp_alu_rcc_data_d[7]), .B(exu_n16075), .Y(exu_n29820));
AND2X1 exu_U36811(.A(byp_alu_rcc_data_e[6]), .B(exu_n16086), .Y(exu_n29822));
AND2X1 exu_U36812(.A(byp_alu_rcc_data_e[5]), .B(exu_n16086), .Y(exu_n29823));
AND2X1 exu_U36813(.A(byp_alu_rcc_data_e[4]), .B(exu_n16086), .Y(exu_n29824));
AND2X1 exu_U36814(.A(exu_ifu_regn_e), .B(exu_n16086), .Y(exu_n29825));
AND2X1 exu_U36815(.A(byp_alu_rcc_data_e[62]), .B(exu_n16086), .Y(exu_n29826));
AND2X1 exu_U36816(.A(byp_alu_rcc_data_e[61]), .B(exu_n16086), .Y(exu_n29827));
AND2X1 exu_U36817(.A(byp_alu_rcc_data_e[60]), .B(exu_n16086), .Y(exu_n29828));
AND2X1 exu_U36818(.A(byp_alu_rcc_data_e[59]), .B(exu_n16086), .Y(exu_n29829));
AND2X1 exu_U36819(.A(byp_alu_rcc_data_e[58]), .B(exu_n16086), .Y(exu_n29830));
AND2X1 exu_U36820(.A(byp_alu_rcc_data_e[57]), .B(exu_n16086), .Y(exu_n29831));
AND2X1 exu_U36821(.A(byp_alu_rcc_data_e[3]), .B(exu_n16086), .Y(exu_n29832));
AND2X1 exu_U36822(.A(byp_alu_rcc_data_e[56]), .B(exu_n16086), .Y(exu_n29833));
AND2X1 exu_U36823(.A(byp_alu_rcc_data_e[55]), .B(exu_n16085), .Y(exu_n29834));
AND2X1 exu_U36824(.A(byp_alu_rcc_data_e[54]), .B(exu_n16085), .Y(exu_n29835));
AND2X1 exu_U36825(.A(byp_alu_rcc_data_e[53]), .B(exu_n16085), .Y(exu_n29836));
AND2X1 exu_U36826(.A(byp_alu_rcc_data_e[52]), .B(exu_n16085), .Y(exu_n29837));
AND2X1 exu_U36827(.A(byp_alu_rcc_data_e[51]), .B(exu_n16085), .Y(exu_n29838));
AND2X1 exu_U36828(.A(byp_alu_rcc_data_e[50]), .B(exu_n16085), .Y(exu_n29839));
AND2X1 exu_U36829(.A(byp_alu_rcc_data_e[49]), .B(exu_n16085), .Y(exu_n29840));
AND2X1 exu_U36830(.A(byp_alu_rcc_data_e[48]), .B(exu_n16085), .Y(exu_n29841));
AND2X1 exu_U36831(.A(byp_alu_rcc_data_e[47]), .B(exu_n16085), .Y(exu_n29842));
AND2X1 exu_U36832(.A(byp_alu_rcc_data_e[2]), .B(exu_n16085), .Y(exu_n29843));
AND2X1 exu_U36833(.A(byp_alu_rcc_data_e[46]), .B(exu_n16085), .Y(exu_n29844));
AND2X1 exu_U36834(.A(byp_alu_rcc_data_e[45]), .B(exu_n16085), .Y(exu_n29845));
AND2X1 exu_U36835(.A(byp_alu_rcc_data_e[44]), .B(exu_n16085), .Y(exu_n29846));
AND2X1 exu_U36836(.A(byp_alu_rcc_data_e[43]), .B(exu_n16084), .Y(exu_n29847));
AND2X1 exu_U36837(.A(byp_alu_rcc_data_e[42]), .B(exu_n16084), .Y(exu_n29848));
AND2X1 exu_U36838(.A(byp_alu_rcc_data_e[41]), .B(exu_n16084), .Y(exu_n29849));
AND2X1 exu_U36839(.A(byp_alu_rcc_data_e[40]), .B(exu_n16084), .Y(exu_n29850));
AND2X1 exu_U36840(.A(byp_alu_rcc_data_e[39]), .B(exu_n16084), .Y(exu_n29851));
AND2X1 exu_U36841(.A(byp_alu_rcc_data_e[38]), .B(exu_n16084), .Y(exu_n29852));
AND2X1 exu_U36842(.A(byp_alu_rcc_data_e[37]), .B(exu_n16084), .Y(exu_n29853));
AND2X1 exu_U36843(.A(byp_alu_rcc_data_e[1]), .B(exu_n16084), .Y(exu_n29854));
AND2X1 exu_U36844(.A(byp_alu_rcc_data_e[36]), .B(exu_n16084), .Y(exu_n29855));
AND2X1 exu_U36845(.A(byp_alu_rcc_data_e[35]), .B(exu_n16084), .Y(exu_n29856));
AND2X1 exu_U36846(.A(byp_alu_rcc_data_e[34]), .B(exu_n16084), .Y(exu_n29857));
AND2X1 exu_U36847(.A(byp_alu_rcc_data_e[33]), .B(exu_n16084), .Y(exu_n29858));
AND2X1 exu_U36848(.A(byp_alu_rcc_data_e[32]), .B(exu_n16084), .Y(exu_n29859));
AND2X1 exu_U36849(.A(byp_alu_rcc_data_e[31]), .B(exu_n16083), .Y(exu_n29860));
AND2X1 exu_U36850(.A(byp_alu_rcc_data_e[30]), .B(exu_n16083), .Y(exu_n29861));
AND2X1 exu_U36851(.A(byp_alu_rcc_data_e[29]), .B(exu_n16083), .Y(exu_n29862));
AND2X1 exu_U36852(.A(byp_alu_rcc_data_e[28]), .B(exu_n16083), .Y(exu_n29863));
AND2X1 exu_U36853(.A(byp_alu_rcc_data_e[27]), .B(exu_n16083), .Y(exu_n29864));
AND2X1 exu_U36854(.A(byp_alu_rcc_data_e[0]), .B(exu_n16083), .Y(exu_n29865));
AND2X1 exu_U36855(.A(byp_alu_rcc_data_e[26]), .B(exu_n16083), .Y(exu_n29866));
AND2X1 exu_U36856(.A(byp_alu_rcc_data_e[25]), .B(exu_n16083), .Y(exu_n29867));
AND2X1 exu_U36857(.A(byp_alu_rcc_data_e[24]), .B(exu_n16083), .Y(exu_n29868));
AND2X1 exu_U36858(.A(byp_alu_rcc_data_e[23]), .B(exu_n16083), .Y(exu_n29869));
AND2X1 exu_U36859(.A(byp_alu_rcc_data_e[22]), .B(exu_n16083), .Y(exu_n29870));
AND2X1 exu_U36860(.A(byp_alu_rcc_data_e[21]), .B(exu_n16083), .Y(exu_n29871));
AND2X1 exu_U36861(.A(byp_alu_rcc_data_e[20]), .B(exu_n16083), .Y(exu_n29872));
AND2X1 exu_U36862(.A(byp_alu_rcc_data_e[19]), .B(exu_n16082), .Y(exu_n29873));
AND2X1 exu_U36863(.A(byp_alu_rcc_data_e[18]), .B(exu_n16082), .Y(exu_n29874));
AND2X1 exu_U36864(.A(byp_alu_rcc_data_e[17]), .B(exu_n16082), .Y(exu_n29875));
AND2X1 exu_U36865(.A(byp_alu_rcc_data_e[16]), .B(exu_n16082), .Y(exu_n29876));
AND2X1 exu_U36866(.A(byp_alu_rcc_data_e[15]), .B(exu_n16082), .Y(exu_n29877));
AND2X1 exu_U36867(.A(byp_alu_rcc_data_e[14]), .B(exu_n16082), .Y(exu_n29878));
AND2X1 exu_U36868(.A(byp_alu_rcc_data_e[13]), .B(exu_n16082), .Y(exu_n29879));
AND2X1 exu_U36869(.A(byp_alu_rcc_data_e[12]), .B(exu_n16082), .Y(exu_n29880));
AND2X1 exu_U36870(.A(byp_alu_rcc_data_e[11]), .B(exu_n16082), .Y(exu_n29881));
AND2X1 exu_U36871(.A(byp_alu_rcc_data_e[10]), .B(exu_n16082), .Y(exu_n29882));
AND2X1 exu_U36872(.A(byp_alu_rcc_data_e[9]), .B(exu_n16082), .Y(exu_n29883));
AND2X1 exu_U36873(.A(byp_alu_rcc_data_e[8]), .B(exu_n16082), .Y(exu_n29884));
AND2X1 exu_U36874(.A(byp_alu_rcc_data_e[7]), .B(exu_n16082), .Y(exu_n29885));
AND2X1 exu_U36875(.A(div_input_data_e[70]), .B(exu_n16093), .Y(exu_n29887));
AND2X1 exu_U36876(.A(div_input_data_e[69]), .B(exu_n16093), .Y(exu_n29888));
AND2X1 exu_U36877(.A(div_input_data_e[68]), .B(exu_n16093), .Y(exu_n29889));
AND2X1 exu_U36878(.A(div_input_data_e[127]), .B(exu_n16093), .Y(exu_n29890));
AND2X1 exu_U36879(.A(div_input_data_e[126]), .B(exu_n16093), .Y(exu_n29891));
AND2X1 exu_U36880(.A(div_input_data_e[125]), .B(exu_n16093), .Y(exu_n29892));
AND2X1 exu_U36881(.A(div_input_data_e[124]), .B(exu_n16093), .Y(exu_n29893));
AND2X1 exu_U36882(.A(div_input_data_e[123]), .B(exu_n16093), .Y(exu_n29894));
AND2X1 exu_U36883(.A(div_input_data_e[122]), .B(exu_n16093), .Y(exu_n29895));
AND2X1 exu_U36884(.A(div_input_data_e[121]), .B(exu_n16093), .Y(exu_n29896));
AND2X1 exu_U36885(.A(div_input_data_e[67]), .B(exu_n16093), .Y(exu_n29897));
AND2X1 exu_U36886(.A(div_input_data_e[120]), .B(exu_n16093), .Y(exu_n29898));
AND2X1 exu_U36887(.A(div_input_data_e[119]), .B(exu_n16092), .Y(exu_n29899));
AND2X1 exu_U36888(.A(div_input_data_e[118]), .B(exu_n16092), .Y(exu_n29900));
AND2X1 exu_U36889(.A(div_input_data_e[117]), .B(exu_n16092), .Y(exu_n29901));
AND2X1 exu_U36890(.A(div_input_data_e[116]), .B(exu_n16092), .Y(exu_n29902));
AND2X1 exu_U36891(.A(div_input_data_e[115]), .B(exu_n16092), .Y(exu_n29903));
AND2X1 exu_U36892(.A(div_input_data_e[114]), .B(exu_n16092), .Y(exu_n29904));
AND2X1 exu_U36893(.A(div_input_data_e[113]), .B(exu_n16092), .Y(exu_n29905));
AND2X1 exu_U36894(.A(div_input_data_e[112]), .B(exu_n16092), .Y(exu_n29906));
AND2X1 exu_U36895(.A(div_input_data_e[111]), .B(exu_n16092), .Y(exu_n29907));
AND2X1 exu_U36896(.A(div_input_data_e[66]), .B(exu_n16092), .Y(exu_n29908));
AND2X1 exu_U36897(.A(div_input_data_e[110]), .B(exu_n16092), .Y(exu_n29909));
AND2X1 exu_U36898(.A(div_input_data_e[109]), .B(exu_n16092), .Y(exu_n29910));
AND2X1 exu_U36899(.A(div_input_data_e[108]), .B(exu_n16092), .Y(exu_n29911));
AND2X1 exu_U36900(.A(div_input_data_e[107]), .B(exu_n16091), .Y(exu_n29912));
AND2X1 exu_U36901(.A(div_input_data_e[106]), .B(exu_n16091), .Y(exu_n29913));
AND2X1 exu_U36902(.A(div_input_data_e[105]), .B(exu_n16091), .Y(exu_n29914));
AND2X1 exu_U36903(.A(div_input_data_e[104]), .B(exu_n16091), .Y(exu_n29915));
AND2X1 exu_U36904(.A(div_input_data_e[103]), .B(exu_n16091), .Y(exu_n29916));
AND2X1 exu_U36905(.A(div_input_data_e[102]), .B(exu_n16091), .Y(exu_n29917));
AND2X1 exu_U36906(.A(div_input_data_e[101]), .B(exu_n16091), .Y(exu_n29918));
AND2X1 exu_U36907(.A(div_input_data_e[65]), .B(exu_n16091), .Y(exu_n29919));
AND2X1 exu_U36908(.A(div_input_data_e[100]), .B(exu_n16091), .Y(exu_n29920));
AND2X1 exu_U36909(.A(div_input_data_e[99]), .B(exu_n16091), .Y(exu_n29921));
AND2X1 exu_U36910(.A(div_input_data_e[98]), .B(exu_n16091), .Y(exu_n29922));
AND2X1 exu_U36911(.A(div_input_data_e[97]), .B(exu_n16091), .Y(exu_n29923));
AND2X1 exu_U36912(.A(div_input_data_e[96]), .B(exu_n16091), .Y(exu_n29924));
AND2X1 exu_U36913(.A(div_input_data_e[94]), .B(exu_n16090), .Y(exu_n29925));
AND2X1 exu_U36914(.A(div_input_data_e[93]), .B(exu_n16090), .Y(exu_n29926));
AND2X1 exu_U36915(.A(div_input_data_e[92]), .B(exu_n16090), .Y(exu_n29927));
AND2X1 exu_U36916(.A(div_input_data_e[91]), .B(exu_n16090), .Y(exu_n29928));
AND2X1 exu_U36917(.A(div_input_data_e[64]), .B(exu_n16090), .Y(exu_n29929));
AND2X1 exu_U36918(.A(div_input_data_e[90]), .B(exu_n16090), .Y(exu_n29930));
AND2X1 exu_U36919(.A(div_input_data_e[89]), .B(exu_n16090), .Y(exu_n29931));
AND2X1 exu_U36920(.A(div_input_data_e[88]), .B(exu_n16090), .Y(exu_n29932));
AND2X1 exu_U36921(.A(div_input_data_e[87]), .B(exu_n16090), .Y(exu_n29933));
AND2X1 exu_U36922(.A(div_input_data_e[86]), .B(exu_n16090), .Y(exu_n29934));
AND2X1 exu_U36923(.A(div_input_data_e[85]), .B(exu_n16090), .Y(exu_n29935));
AND2X1 exu_U36924(.A(div_input_data_e[84]), .B(exu_n16090), .Y(exu_n29936));
AND2X1 exu_U36925(.A(div_input_data_e[83]), .B(exu_n16089), .Y(exu_n29937));
AND2X1 exu_U36926(.A(div_input_data_e[82]), .B(exu_n16089), .Y(exu_n29938));
AND2X1 exu_U36927(.A(div_input_data_e[81]), .B(exu_n16089), .Y(exu_n29939));
AND2X1 exu_U36928(.A(div_input_data_e[80]), .B(exu_n16089), .Y(exu_n29940));
AND2X1 exu_U36929(.A(div_input_data_e[79]), .B(exu_n16089), .Y(exu_n29941));
AND2X1 exu_U36930(.A(div_input_data_e[78]), .B(exu_n16089), .Y(exu_n29942));
AND2X1 exu_U36931(.A(div_input_data_e[77]), .B(exu_n16089), .Y(exu_n29943));
AND2X1 exu_U36932(.A(div_input_data_e[76]), .B(exu_n16089), .Y(exu_n29944));
AND2X1 exu_U36933(.A(div_input_data_e[75]), .B(exu_n16089), .Y(exu_n29945));
AND2X1 exu_U36934(.A(div_input_data_e[74]), .B(exu_n16089), .Y(exu_n29946));
AND2X1 exu_U36935(.A(div_input_data_e[73]), .B(exu_n16089), .Y(exu_n29947));
AND2X1 exu_U36936(.A(div_input_data_e[72]), .B(exu_n16089), .Y(exu_n29948));
AND2X1 exu_U36937(.A(div_input_data_e[71]), .B(exu_n16089), .Y(exu_n29949));
AND2X1 exu_U36938(.A(exu_spu_rs3_data_e[6]), .B(exu_n16100), .Y(exu_n29951));
AND2X1 exu_U36939(.A(exu_spu_rs3_data_e[5]), .B(exu_n16100), .Y(exu_n29952));
AND2X1 exu_U36940(.A(exu_spu_rs3_data_e[4]), .B(exu_n16100), .Y(exu_n29953));
AND2X1 exu_U36941(.A(exu_spu_rs3_data_e[63]), .B(exu_n16100), .Y(exu_n29954));
AND2X1 exu_U36942(.A(exu_spu_rs3_data_e[62]), .B(exu_n16100), .Y(exu_n29955));
AND2X1 exu_U36943(.A(exu_spu_rs3_data_e[61]), .B(exu_n16100), .Y(exu_n29956));
AND2X1 exu_U36944(.A(exu_spu_rs3_data_e[60]), .B(exu_n16100), .Y(exu_n29957));
AND2X1 exu_U36945(.A(exu_spu_rs3_data_e[59]), .B(exu_n16100), .Y(exu_n29958));
AND2X1 exu_U36946(.A(exu_spu_rs3_data_e[58]), .B(exu_n16100), .Y(exu_n29959));
AND2X1 exu_U36947(.A(exu_spu_rs3_data_e[57]), .B(exu_n16100), .Y(exu_n29960));
AND2X1 exu_U36948(.A(exu_spu_rs3_data_e[3]), .B(exu_n16100), .Y(exu_n29961));
AND2X1 exu_U36949(.A(exu_spu_rs3_data_e[56]), .B(exu_n16100), .Y(exu_n29962));
AND2X1 exu_U36950(.A(exu_spu_rs3_data_e[55]), .B(exu_n16099), .Y(exu_n29963));
AND2X1 exu_U36951(.A(exu_spu_rs3_data_e[54]), .B(exu_n16099), .Y(exu_n29964));
AND2X1 exu_U36952(.A(exu_spu_rs3_data_e[53]), .B(exu_n16099), .Y(exu_n29965));
AND2X1 exu_U36953(.A(exu_spu_rs3_data_e[52]), .B(exu_n16099), .Y(exu_n29966));
AND2X1 exu_U36954(.A(exu_spu_rs3_data_e[51]), .B(exu_n16099), .Y(exu_n29967));
AND2X1 exu_U36955(.A(exu_spu_rs3_data_e[50]), .B(exu_n16099), .Y(exu_n29968));
AND2X1 exu_U36956(.A(exu_spu_rs3_data_e[49]), .B(exu_n16099), .Y(exu_n29969));
AND2X1 exu_U36957(.A(exu_spu_rs3_data_e[48]), .B(exu_n16099), .Y(exu_n29970));
AND2X1 exu_U36958(.A(exu_spu_rs3_data_e[47]), .B(exu_n16099), .Y(exu_n29971));
AND2X1 exu_U36959(.A(exu_spu_rs3_data_e[2]), .B(exu_n16099), .Y(exu_n29972));
AND2X1 exu_U36960(.A(exu_spu_rs3_data_e[46]), .B(exu_n16099), .Y(exu_n29973));
AND2X1 exu_U36961(.A(exu_spu_rs3_data_e[45]), .B(exu_n16099), .Y(exu_n29974));
AND2X1 exu_U36962(.A(exu_spu_rs3_data_e[44]), .B(exu_n16099), .Y(exu_n29975));
AND2X1 exu_U36963(.A(exu_spu_rs3_data_e[43]), .B(exu_n16098), .Y(exu_n29976));
AND2X1 exu_U36964(.A(exu_spu_rs3_data_e[42]), .B(exu_n16098), .Y(exu_n29977));
AND2X1 exu_U36965(.A(exu_spu_rs3_data_e[41]), .B(exu_n16098), .Y(exu_n29978));
AND2X1 exu_U36966(.A(exu_spu_rs3_data_e[40]), .B(exu_n16098), .Y(exu_n29979));
AND2X1 exu_U36967(.A(exu_spu_rs3_data_e[39]), .B(exu_n16098), .Y(exu_n29980));
AND2X1 exu_U36968(.A(exu_spu_rs3_data_e[38]), .B(exu_n16098), .Y(exu_n29981));
AND2X1 exu_U36969(.A(exu_spu_rs3_data_e[37]), .B(exu_n16098), .Y(exu_n29982));
AND2X1 exu_U36970(.A(exu_spu_rs3_data_e[1]), .B(exu_n16098), .Y(exu_n29983));
AND2X1 exu_U36971(.A(exu_spu_rs3_data_e[36]), .B(exu_n16098), .Y(exu_n29984));
AND2X1 exu_U36972(.A(exu_spu_rs3_data_e[35]), .B(exu_n16098), .Y(exu_n29985));
AND2X1 exu_U36973(.A(exu_spu_rs3_data_e[34]), .B(exu_n16098), .Y(exu_n29986));
AND2X1 exu_U36974(.A(exu_spu_rs3_data_e[33]), .B(exu_n16098), .Y(exu_n29987));
AND2X1 exu_U36975(.A(exu_spu_rs3_data_e[32]), .B(exu_n16098), .Y(exu_n29988));
AND2X1 exu_U36976(.A(exu_spu_rs3_data_e[31]), .B(exu_n16097), .Y(exu_n29989));
AND2X1 exu_U36977(.A(exu_spu_rs3_data_e[30]), .B(exu_n16097), .Y(exu_n29990));
AND2X1 exu_U36978(.A(exu_spu_rs3_data_e[29]), .B(exu_n16097), .Y(exu_n29991));
AND2X1 exu_U36979(.A(exu_spu_rs3_data_e[28]), .B(exu_n16097), .Y(exu_n29992));
AND2X1 exu_U36980(.A(exu_spu_rs3_data_e[27]), .B(exu_n16097), .Y(exu_n29993));
AND2X1 exu_U36981(.A(exu_spu_rs3_data_e[0]), .B(exu_n16097), .Y(exu_n29994));
AND2X1 exu_U36982(.A(exu_spu_rs3_data_e[26]), .B(exu_n16097), .Y(exu_n29995));
AND2X1 exu_U36983(.A(exu_spu_rs3_data_e[25]), .B(exu_n16097), .Y(exu_n29996));
AND2X1 exu_U36984(.A(exu_spu_rs3_data_e[24]), .B(exu_n16097), .Y(exu_n29997));
AND2X1 exu_U36985(.A(exu_spu_rs3_data_e[23]), .B(exu_n16097), .Y(exu_n29998));
AND2X1 exu_U36986(.A(exu_spu_rs3_data_e[22]), .B(exu_n16097), .Y(exu_n29999));
AND2X1 exu_U36987(.A(exu_spu_rs3_data_e[21]), .B(exu_n16097), .Y(exu_n30000));
AND2X1 exu_U36988(.A(exu_spu_rs3_data_e[20]), .B(exu_n16097), .Y(exu_n30001));
AND2X1 exu_U36989(.A(exu_spu_rs3_data_e[19]), .B(exu_n16096), .Y(exu_n30002));
AND2X1 exu_U36990(.A(exu_spu_rs3_data_e[18]), .B(exu_n16096), .Y(exu_n30003));
AND2X1 exu_U36991(.A(exu_spu_rs3_data_e[17]), .B(exu_n16096), .Y(exu_n30004));
AND2X1 exu_U36992(.A(exu_spu_rs3_data_e[16]), .B(exu_n16096), .Y(exu_n30005));
AND2X1 exu_U36993(.A(exu_spu_rs3_data_e[15]), .B(exu_n16096), .Y(exu_n30006));
AND2X1 exu_U36994(.A(exu_spu_rs3_data_e[14]), .B(exu_n16096), .Y(exu_n30007));
AND2X1 exu_U36995(.A(exu_spu_rs3_data_e[13]), .B(exu_n16096), .Y(exu_n30008));
AND2X1 exu_U36996(.A(exu_spu_rs3_data_e[12]), .B(exu_n16096), .Y(exu_n30009));
AND2X1 exu_U36997(.A(exu_spu_rs3_data_e[11]), .B(exu_n16096), .Y(exu_n30010));
AND2X1 exu_U36998(.A(exu_spu_rs3_data_e[10]), .B(exu_n16096), .Y(exu_n30011));
AND2X1 exu_U36999(.A(exu_spu_rs3_data_e[9]), .B(exu_n16096), .Y(exu_n30012));
AND2X1 exu_U37000(.A(exu_spu_rs3_data_e[8]), .B(exu_n16096), .Y(exu_n30013));
AND2X1 exu_U37001(.A(exu_spu_rs3_data_e[7]), .B(exu_n16096), .Y(exu_n30014));
AND2X1 exu_U37002(.A(exu_n16442), .B(exu_n16107), .Y(exu_n30016));
AND2X1 exu_U37003(.A(exu_n16447), .B(exu_n16107), .Y(exu_n30017));
AND2X1 exu_U37004(.A(exu_n16458), .B(exu_n16107), .Y(exu_n30018));
AND2X1 exu_U37005(.A(exu_n16443), .B(exu_n16107), .Y(exu_n30019));
AND2X1 exu_U37006(.A(exu_n16444), .B(exu_n16107), .Y(exu_n30020));
AND2X1 exu_U37007(.A(exu_n16445), .B(exu_n16107), .Y(exu_n30021));
AND2X1 exu_U37008(.A(exu_n16446), .B(exu_n16107), .Y(exu_n30022));
AND2X1 exu_U37009(.A(exu_n16448), .B(exu_n16107), .Y(exu_n30023));
AND2X1 exu_U37010(.A(exu_n16449), .B(exu_n16107), .Y(exu_n30024));
AND2X1 exu_U37011(.A(exu_n16450), .B(exu_n16107), .Y(exu_n30025));
AND2X1 exu_U37012(.A(exu_n16469), .B(exu_n16107), .Y(exu_n30026));
AND2X1 exu_U37013(.A(exu_n16451), .B(exu_n16107), .Y(exu_n30027));
AND2X1 exu_U37014(.A(exu_n16452), .B(exu_n16106), .Y(exu_n30028));
AND2X1 exu_U37015(.A(exu_n16453), .B(exu_n16106), .Y(exu_n30029));
AND2X1 exu_U37016(.A(exu_n16454), .B(exu_n16106), .Y(exu_n30030));
AND2X1 exu_U37017(.A(exu_n16455), .B(exu_n16106), .Y(exu_n30031));
AND2X1 exu_U37018(.A(exu_n16456), .B(exu_n16106), .Y(exu_n30032));
AND2X1 exu_U37019(.A(exu_n16457), .B(exu_n16106), .Y(exu_n30033));
AND2X1 exu_U37020(.A(exu_n16459), .B(exu_n16106), .Y(exu_n30034));
AND2X1 exu_U37021(.A(exu_n16460), .B(exu_n16106), .Y(exu_n30035));
AND2X1 exu_U37022(.A(exu_n16461), .B(exu_n16106), .Y(exu_n30036));
AND2X1 exu_U37023(.A(exu_n16480), .B(exu_n16106), .Y(exu_n30037));
AND2X1 exu_U37024(.A(exu_n16462), .B(exu_n16106), .Y(exu_n30038));
AND2X1 exu_U37025(.A(exu_n16463), .B(exu_n16106), .Y(exu_n30039));
AND2X1 exu_U37026(.A(exu_n16464), .B(exu_n16106), .Y(exu_n30040));
AND2X1 exu_U37027(.A(exu_n16465), .B(exu_n16105), .Y(exu_n30041));
AND2X1 exu_U37028(.A(exu_n16466), .B(exu_n16105), .Y(exu_n30042));
AND2X1 exu_U37029(.A(exu_n16467), .B(exu_n16105), .Y(exu_n30043));
AND2X1 exu_U37030(.A(exu_n16468), .B(exu_n16105), .Y(exu_n30044));
AND2X1 exu_U37031(.A(exu_n16470), .B(exu_n16105), .Y(exu_n30045));
AND2X1 exu_U37032(.A(exu_n16471), .B(exu_n16105), .Y(exu_n30046));
AND2X1 exu_U37033(.A(exu_n16472), .B(exu_n16105), .Y(exu_n30047));
AND2X1 exu_U37034(.A(exu_n16491), .B(exu_n16105), .Y(exu_n30048));
AND2X1 exu_U37035(.A(exu_n16473), .B(exu_n16105), .Y(exu_n30049));
AND2X1 exu_U37036(.A(exu_n16474), .B(exu_n16105), .Y(exu_n30050));
AND2X1 exu_U37037(.A(exu_n16475), .B(exu_n16105), .Y(exu_n30051));
AND2X1 exu_U37038(.A(exu_n16476), .B(exu_n16105), .Y(exu_n30052));
AND2X1 exu_U37039(.A(exu_n16477), .B(exu_n16105), .Y(exu_n30053));
AND2X1 exu_U37040(.A(exu_n16478), .B(exu_n16104), .Y(exu_n30054));
AND2X1 exu_U37041(.A(exu_n16479), .B(exu_n16104), .Y(exu_n30055));
AND2X1 exu_U37042(.A(exu_n16481), .B(exu_n16104), .Y(exu_n30056));
AND2X1 exu_U37043(.A(exu_n16482), .B(exu_n16104), .Y(exu_n30057));
AND2X1 exu_U37044(.A(exu_n16483), .B(exu_n16104), .Y(exu_n30058));
AND2X1 exu_U37045(.A(exu_n16502), .B(exu_n16104), .Y(exu_n30059));
AND2X1 exu_U37046(.A(exu_n16484), .B(exu_n16104), .Y(exu_n30060));
AND2X1 exu_U37047(.A(exu_n16485), .B(exu_n16104), .Y(exu_n30061));
AND2X1 exu_U37048(.A(exu_n16486), .B(exu_n16104), .Y(exu_n30062));
AND2X1 exu_U37049(.A(exu_n16487), .B(exu_n16104), .Y(exu_n30063));
AND2X1 exu_U37050(.A(exu_n16488), .B(exu_n16104), .Y(exu_n30064));
AND2X1 exu_U37051(.A(exu_n16489), .B(exu_n16104), .Y(exu_n30065));
AND2X1 exu_U37052(.A(exu_n16490), .B(exu_n16104), .Y(exu_n30066));
AND2X1 exu_U37053(.A(exu_n16492), .B(exu_n16103), .Y(exu_n30067));
AND2X1 exu_U37054(.A(exu_n16493), .B(exu_n16103), .Y(exu_n30068));
AND2X1 exu_U37055(.A(exu_n16494), .B(exu_n16103), .Y(exu_n30069));
AND2X1 exu_U37056(.A(exu_n16495), .B(exu_n16103), .Y(exu_n30070));
AND2X1 exu_U37057(.A(exu_n16496), .B(exu_n16103), .Y(exu_n30071));
AND2X1 exu_U37058(.A(exu_n16497), .B(exu_n16103), .Y(exu_n30072));
AND2X1 exu_U37059(.A(exu_n16498), .B(exu_n16103), .Y(exu_n30073));
AND2X1 exu_U37060(.A(exu_n16499), .B(exu_n16103), .Y(exu_n30074));
AND2X1 exu_U37061(.A(exu_n16500), .B(exu_n16103), .Y(exu_n30075));
AND2X1 exu_U37062(.A(exu_n16501), .B(exu_n16103), .Y(exu_n30076));
AND2X1 exu_U37063(.A(exu_n16439), .B(exu_n16103), .Y(exu_n30077));
AND2X1 exu_U37064(.A(exu_n16440), .B(exu_n16103), .Y(exu_n30078));
AND2X1 exu_U37065(.A(exu_n16441), .B(exu_n16103), .Y(exu_n30079));
INVX1 exu_U37066(.A(exu_n15012), .Y(exu_n16322));
INVX1 exu_U37067(.A(exu_n15013), .Y(exu_n16325));
INVX1 exu_U37068(.A(exu_n15012), .Y(exu_n16326));
INVX1 exu_U37069(.A(exu_n15013), .Y(exu_n16327));
INVX1 exu_U37070(.A(exu_n15012), .Y(exu_n16328));
INVX1 exu_U37071(.A(exu_n15013), .Y(exu_n16329));
INVX1 exu_U37072(.A(exu_n15012), .Y(exu_n16330));
INVX1 exu_U37073(.A(exu_n15013), .Y(exu_n16331));
INVX1 exu_U37074(.A(exu_n16324), .Y(exu_n15012));
INVX1 exu_U37075(.A(exu_n15012), .Y(exu_n16332));
INVX1 exu_U37076(.A(exu_n15013), .Y(exu_n16324));
INVX1 exu_U37077(.A(exu_n16323), .Y(exu_n15013));
INVX1 exu_U37078(.A(exu_n14998), .Y(exu_n16323));
INVX1 exu_U37079(.A(exu_n15015), .Y(exu_n16333));
INVX1 exu_U37080(.A(exu_n15014), .Y(exu_n16334));
INVX1 exu_U37081(.A(exu_n15015), .Y(exu_n16335));
INVX1 exu_U37082(.A(exu_n15014), .Y(exu_n16336));
INVX1 exu_U37083(.A(exu_n15015), .Y(exu_n16337));
INVX1 exu_U37084(.A(exu_n15014), .Y(exu_n16338));
INVX1 exu_U37085(.A(exu_n15015), .Y(exu_n16339));
INVX1 exu_U37086(.A(exu_n15015), .Y(exu_n16340));
INVX1 exu_U37087(.A(exu_n16341), .Y(exu_n15014));
INVX1 exu_U37088(.A(exu_n14999), .Y(exu_n16341));
INVX1 exu_U37089(.A(exu_n16342), .Y(exu_n15015));
INVX1 exu_U37090(.A(exu_n15014), .Y(exu_n16342));
INVX1 exu_U37091(.A(exu_n15017), .Y(exu_n16343));
INVX1 exu_U37092(.A(exu_n15016), .Y(exu_n16344));
INVX1 exu_U37093(.A(exu_n15017), .Y(exu_n16345));
INVX1 exu_U37094(.A(exu_n15016), .Y(exu_n16346));
INVX1 exu_U37095(.A(exu_n15017), .Y(exu_n16347));
INVX1 exu_U37096(.A(exu_n15016), .Y(exu_n16348));
INVX1 exu_U37097(.A(exu_n15017), .Y(exu_n16349));
INVX1 exu_U37098(.A(exu_n16350), .Y(exu_n15016));
INVX1 exu_U37099(.A(exu_n14998), .Y(exu_n16350));
INVX1 exu_U37100(.A(exu_n16351), .Y(exu_n15017));
INVX1 exu_U37101(.A(exu_n15016), .Y(exu_n16351));
INVX1 exu_U37102(.A(exu_n15019), .Y(exu_n16352));
INVX1 exu_U37103(.A(exu_n15018), .Y(exu_n16353));
INVX1 exu_U37104(.A(exu_n15019), .Y(exu_n16354));
INVX1 exu_U37105(.A(exu_n15018), .Y(exu_n16355));
INVX1 exu_U37106(.A(exu_n15019), .Y(exu_n16356));
INVX1 exu_U37107(.A(exu_n15018), .Y(exu_n16358));
INVX1 exu_U37108(.A(exu_n15019), .Y(exu_n16359));
INVX1 exu_U37109(.A(exu_n16357), .Y(exu_n15018));
INVX1 exu_U37110(.A(exu_n14999), .Y(exu_n16357));
INVX1 exu_U37111(.A(exu_n16360), .Y(exu_n15019));
INVX1 exu_U37112(.A(exu_n15018), .Y(exu_n16360));
INVX1 exu_U37113(.A(exu_n15021), .Y(exu_n16361));
INVX1 exu_U37114(.A(exu_n15020), .Y(exu_n16362));
INVX1 exu_U37115(.A(exu_n15021), .Y(exu_n16363));
INVX1 exu_U37116(.A(exu_n15020), .Y(exu_n16364));
INVX1 exu_U37117(.A(exu_n15021), .Y(exu_n16365));
INVX1 exu_U37118(.A(exu_n15020), .Y(exu_n16366));
INVX1 exu_U37119(.A(exu_n15020), .Y(exu_n16367));
INVX1 exu_U37120(.A(exu_n16369), .Y(exu_n15020));
INVX1 exu_U37121(.A(exu_n15021), .Y(exu_n16369));
INVX1 exu_U37122(.A(exu_n16368), .Y(exu_n15021));
INVX1 exu_U37123(.A(exu_n14998), .Y(exu_n16368));
AND2X1 exu_U37124(.A(exu_spu_rs3_data_e[63]), .B(exu_n16167), .Y(exu_lsu_rs3_data_e[63]));
AND2X1 exu_U37125(.A(exu_spu_rs3_data_e[62]), .B(exu_n16167), .Y(exu_lsu_rs3_data_e[62]));
AND2X1 exu_U37126(.A(exu_spu_rs3_data_e[61]), .B(exu_n16169), .Y(exu_lsu_rs3_data_e[61]));
AND2X1 exu_U37127(.A(exu_spu_rs3_data_e[60]), .B(exu_n16167), .Y(exu_lsu_rs3_data_e[60]));
AND2X1 exu_U37128(.A(exu_spu_rs3_data_e[59]), .B(exu_n16168), .Y(exu_lsu_rs3_data_e[59]));
AND2X1 exu_U37129(.A(exu_spu_rs3_data_e[58]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[58]));
AND2X1 exu_U37130(.A(exu_spu_rs3_data_e[57]), .B(exu_n16168), .Y(exu_lsu_rs3_data_e[57]));
AND2X1 exu_U37131(.A(exu_spu_rs3_data_e[56]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[56]));
AND2X1 exu_U37132(.A(exu_spu_rs3_data_e[55]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[55]));
AND2X1 exu_U37133(.A(exu_spu_rs3_data_e[54]), .B(exu_n16169), .Y(exu_lsu_rs3_data_e[54]));
AND2X1 exu_U37134(.A(exu_spu_rs3_data_e[53]), .B(exu_n16167), .Y(exu_lsu_rs3_data_e[53]));
AND2X1 exu_U37135(.A(exu_spu_rs3_data_e[52]), .B(exu_n16168), .Y(exu_lsu_rs3_data_e[52]));
AND2X1 exu_U37136(.A(exu_spu_rs3_data_e[51]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[51]));
AND2X1 exu_U37137(.A(exu_spu_rs3_data_e[50]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[50]));
AND2X1 exu_U37138(.A(exu_spu_rs3_data_e[49]), .B(exu_n16169), .Y(exu_lsu_rs3_data_e[49]));
AND2X1 exu_U37139(.A(exu_spu_rs3_data_e[48]), .B(exu_n16167), .Y(exu_lsu_rs3_data_e[48]));
AND2X1 exu_U37140(.A(exu_spu_rs3_data_e[47]), .B(exu_n16168), .Y(exu_lsu_rs3_data_e[47]));
AND2X1 exu_U37141(.A(exu_spu_rs3_data_e[46]), .B(exu_n16169), .Y(exu_lsu_rs3_data_e[46]));
AND2X1 exu_U37142(.A(exu_spu_rs3_data_e[45]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[45]));
AND2X1 exu_U37143(.A(exu_spu_rs3_data_e[44]), .B(exu_n16169), .Y(exu_lsu_rs3_data_e[44]));
AND2X1 exu_U37144(.A(exu_spu_rs3_data_e[43]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[43]));
AND2X1 exu_U37145(.A(exu_spu_rs3_data_e[42]), .B(exu_n16169), .Y(exu_lsu_rs3_data_e[42]));
AND2X1 exu_U37146(.A(exu_spu_rs3_data_e[41]), .B(exu_n16167), .Y(exu_lsu_rs3_data_e[41]));
AND2X1 exu_U37147(.A(exu_spu_rs3_data_e[40]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[40]));
AND2X1 exu_U37148(.A(exu_spu_rs3_data_e[39]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[39]));
AND2X1 exu_U37149(.A(exu_spu_rs3_data_e[38]), .B(exu_n16169), .Y(exu_lsu_rs3_data_e[38]));
AND2X1 exu_U37150(.A(exu_spu_rs3_data_e[37]), .B(exu_n16167), .Y(exu_lsu_rs3_data_e[37]));
AND2X1 exu_U37151(.A(exu_spu_rs3_data_e[36]), .B(exu_n16167), .Y(exu_lsu_rs3_data_e[36]));
AND2X1 exu_U37152(.A(exu_spu_rs3_data_e[35]), .B(exu_n16170), .Y(exu_lsu_rs3_data_e[35]));
AND2X1 exu_U37153(.A(exu_spu_rs3_data_e[34]), .B(exu_n16169), .Y(exu_lsu_rs3_data_e[34]));
AND2X1 exu_U37154(.A(exu_spu_rs3_data_e[33]), .B(exu_n16167), .Y(exu_lsu_rs3_data_e[33]));
AND2X1 exu_U37155(.A(exu_spu_rs3_data_e[32]), .B(exu_n16168), .Y(exu_lsu_rs3_data_e[32]));
AND2X1 exu_U37156(.A(rml_cwp_swap_slot0_state_valid[0]), .B(rml_cwp_swap_keep_state[0]), .Y(exu_n31472));
AND2X1 exu_U37157(.A(rml_cwp_valid_tlu_swap_w), .B(rml_cwp_swap_sel_tlu[0]), .Y(exu_n31473));
AND2X1 exu_U37158(.A(rml_cwp_swap_slot1_state_valid[0]), .B(rml_cwp_swap_keep_state[1]), .Y(exu_n31477));
AND2X1 exu_U37159(.A(rml_cwp_valid_tlu_swap_w), .B(rml_cwp_n34), .Y(exu_n31478));
AND2X1 exu_U37160(.A(rml_cwp_swap_slot2_state_valid[0]), .B(rml_cwp_swap_keep_state[2]), .Y(exu_n31482));
AND2X1 exu_U37161(.A(rml_cwp_valid_tlu_swap_w), .B(rml_cwp_n33), .Y(exu_n31483));
AND2X1 exu_U37162(.A(rml_cwp_swap_slot3_state_valid[0]), .B(rml_cwp_swap_keep_state[3]), .Y(exu_n31487));
AND2X1 exu_U37163(.A(rml_cwp_valid_tlu_swap_w), .B(rml_cwp_n32), .Y(exu_n31488));
AND2X1 exu_U37164(.A(rml_cwp_next_slot0_state[1]), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n2));
AND2X1 exu_U37165(.A(rml_cwp_next_slot0_state[0]), .B(exu_n15946), .Y(rml_cwp_slot0_data_dff_n5));
AND2X1 exu_U37166(.A(ecl_divcntl_inputs_neg_d), .B(exu_n19255), .Y(ecl_divcntl_inputs_neg_dff_n8));
AND2X1 exu_U37167(.A(ecl_divcntl_next_state[5]), .B(ecl_divcntl_divstate_dff_n1), .Y(ecl_divcntl_divstate_dff_n3));
AND2X1 exu_U37168(.A(ecl_divcntl_next_state[4]), .B(ecl_divcntl_divstate_dff_n1), .Y(ecl_divcntl_divstate_dff_n5));
AND2X1 exu_U37169(.A(ecl_divcntl_next_state[1]), .B(ecl_divcntl_divstate_dff_n1), .Y(ecl_divcntl_divstate_dff_n11));
AND2X1 exu_U37170(.A(ecl_tid_m[0]), .B(ecl_writeback_restore_tid_dff_n2), .Y(ecl_writeback_restore_tid_dff_n8));
AND2X1 exu_U37171(.A(ecl_tid_m[1]), .B(ecl_writeback_restore_tid_dff_n2), .Y(ecl_writeback_restore_tid_dff_n13));
OR2X1 exu_U37172(.A(mux_drive_disable), .B(ecl_eccctl_sel_rs1_m), .Y(ecl_ecc_sel_rs1_m_l));
AND2X1 exu_U37173(.A(ecl_eccctl_sel_rs2_m), .B(exu_n16396), .Y(ecl_ecc_sel_rs2_m_l));
INVX1 exu_U37174(.A(ecl_ecc_sel_rs2_m_l), .Y(exu_n15022));
AND2X1 exu_U37175(.A(ecl_eccctl_sel_rs3_m), .B(exu_n16396), .Y(ecl_ecc_sel_rs3_m_l));
INVX1 exu_U37176(.A(ecl_ecc_sel_rs3_m_l), .Y(exu_n15023));
AND2X1 exu_U37177(.A(exu_n16379), .B(ecl_ttype_e2m_n1), .Y(ecl_ttype_e2m_n3));
AND2X1 exu_U37178(.A(exu_n16378), .B(ecl_ttype_e2m_n1), .Y(ecl_ttype_e2m_n9));
AND2X1 exu_U37179(.A(exu_n16377), .B(ecl_ttype_e2m_n1), .Y(ecl_ttype_e2m_n13));
AND2X1 exu_U37180(.A(exu_n16376), .B(ecl_ttype_e2m_n1), .Y(ecl_ttype_e2m_n15));
AND2X1 exu_U37181(.A(ifu_exu_tcc_e), .B(ecl_ttype_e2m_n1), .Y(ecl_ttype_e2m_n17));
AND2X1 exu_U37182(.A(exu_n16380), .B(ecl_ttype_e2m_n1), .Y(ecl_ttype_e2m_n19));
AND2X1 exu_U37183(.A(ifu_exu_enshift_d), .B(bypass_irf_write_clkbuf_tmb_l), .Y(ecl_dff_enshift_d2e_n3));
AND2X1 exu_U37184(.A(ifu_exu_aluop_d[2]), .B(ecl_dff_aluop_d2e_n1), .Y(ecl_dff_aluop_d2e_n3));
AND2X1 exu_U37185(.A(ifu_exu_aluop_d[1]), .B(ecl_dff_aluop_d2e_n1), .Y(ecl_dff_aluop_d2e_n5));
AND2X1 exu_U37186(.A(ifu_exu_aluop_d[0]), .B(ecl_dff_aluop_d2e_n1), .Y(ecl_dff_aluop_d2e_n7));
AND2X1 exu_U37187(.A(lsu_exu_thr_m[1]), .B(ecl_dff_ld_tid_m2g_n1), .Y(ecl_dff_ld_tid_m2g_n3));
AND2X1 exu_U37188(.A(lsu_exu_thr_m[0]), .B(ecl_dff_ld_tid_m2g_n1), .Y(ecl_dff_ld_tid_m2g_n5));
AND2X1 exu_U37189(.A(ifu_exu_rs1_s[4]), .B(ecl_dff_rs1_s2d_n1), .Y(ecl_dff_rs1_s2d_n3));
AND2X1 exu_U37190(.A(ifu_exu_rs1_s[3]), .B(ecl_dff_rs1_s2d_n1), .Y(ecl_dff_rs1_s2d_n5));
AND2X1 exu_U37191(.A(ifu_exu_rs1_s[2]), .B(ecl_dff_rs1_s2d_n1), .Y(ecl_dff_rs1_s2d_n7));
AND2X1 exu_U37192(.A(ifu_exu_rs1_s[1]), .B(ecl_dff_rs1_s2d_n1), .Y(ecl_dff_rs1_s2d_n9));
AND2X1 exu_U37193(.A(ifu_exu_rs1_s[0]), .B(ecl_dff_rs1_s2d_n1), .Y(ecl_dff_rs1_s2d_n11));
AND2X1 exu_U37194(.A(ecc_rs1_err_e[6]), .B(ecc_rs1_err_e2m_n1), .Y(ecc_rs1_err_e2m_n3));
AND2X1 exu_U37195(.A(ecc_rs1_err_e[5]), .B(ecc_rs1_err_e2m_n1), .Y(ecc_rs1_err_e2m_n5));
AND2X1 exu_U37196(.A(ecc_rs1_err_e[4]), .B(ecc_rs1_err_e2m_n1), .Y(ecc_rs1_err_e2m_n7));
AND2X1 exu_U37197(.A(ecc_rs1_err_e[3]), .B(ecc_rs1_err_e2m_n1), .Y(ecc_rs1_err_e2m_n9));
AND2X1 exu_U37198(.A(ecc_rs1_err_e[2]), .B(ecc_rs1_err_e2m_n1), .Y(ecc_rs1_err_e2m_n11));
AND2X1 exu_U37199(.A(ecc_rs1_err_e[1]), .B(ecc_rs1_err_e2m_n1), .Y(ecc_rs1_err_e2m_n13));
AND2X1 exu_U37200(.A(ecc_rs1_err_e[0]), .B(ecc_rs1_err_e2m_n1), .Y(ecc_rs1_err_e2m_n15));
AND2X1 exu_U37201(.A(byp_ecc_rs1_synd_d[6]), .B(ecc_rs1_ecc_d2e_n1), .Y(ecc_rs1_ecc_d2e_n3));
AND2X1 exu_U37202(.A(byp_ecc_rs1_synd_d[5]), .B(ecc_rs1_ecc_d2e_n1), .Y(ecc_rs1_ecc_d2e_n5));
AND2X1 exu_U37203(.A(byp_ecc_rs1_synd_d[4]), .B(ecc_rs1_ecc_d2e_n1), .Y(ecc_rs1_ecc_d2e_n7));
AND2X1 exu_U37204(.A(byp_ecc_rs1_synd_d[3]), .B(ecc_rs1_ecc_d2e_n1), .Y(ecc_rs1_ecc_d2e_n9));
AND2X1 exu_U37205(.A(byp_ecc_rs1_synd_d[2]), .B(ecc_rs1_ecc_d2e_n1), .Y(ecc_rs1_ecc_d2e_n11));
AND2X1 exu_U37206(.A(byp_ecc_rs1_synd_d[1]), .B(ecc_rs1_ecc_d2e_n1), .Y(ecc_rs1_ecc_d2e_n13));
AND2X1 exu_U37207(.A(byp_ecc_rs1_synd_d[0]), .B(ecc_rs1_ecc_d2e_n1), .Y(ecc_rs1_ecc_d2e_n15));
AND2X1 exu_U37208(.A(byp_ecc_rs1_synd_d[7]), .B(ecc_rs1_ecc_d2e_n1), .Y(ecc_rs1_ecc_d2e_n17));
AND2X1 exu_U37209(.A(bypass_rs3h_data_d[6]), .B(exu_n16133), .Y(bypass_rs3h_data_dff_n3));
AND2X1 exu_U37210(.A(bypass_rs3h_data_d[5]), .B(exu_n16133), .Y(bypass_rs3h_data_dff_n5));
AND2X1 exu_U37211(.A(bypass_rs3h_data_d[4]), .B(exu_n16133), .Y(bypass_rs3h_data_dff_n7));
AND2X1 exu_U37212(.A(bypass_rs3h_data_d[3]), .B(exu_n16133), .Y(bypass_rs3h_data_dff_n9));
AND2X1 exu_U37213(.A(bypass_rs3h_data_d[2]), .B(exu_n16133), .Y(bypass_rs3h_data_dff_n11));
AND2X1 exu_U37214(.A(bypass_rs3h_data_d[1]), .B(exu_n16133), .Y(bypass_rs3h_data_dff_n13));
AND2X1 exu_U37215(.A(bypass_rs3h_data_d[31]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n15));
AND2X1 exu_U37216(.A(bypass_rs3h_data_d[30]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n17));
AND2X1 exu_U37217(.A(bypass_rs3h_data_d[29]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n19));
AND2X1 exu_U37218(.A(bypass_rs3h_data_d[28]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n21));
AND2X1 exu_U37219(.A(bypass_rs3h_data_d[27]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n23));
AND2X1 exu_U37220(.A(bypass_rs3h_data_d[0]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n25));
AND2X1 exu_U37221(.A(bypass_rs3h_data_d[26]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n27));
AND2X1 exu_U37222(.A(bypass_rs3h_data_d[25]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n29));
AND2X1 exu_U37223(.A(bypass_rs3h_data_d[24]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n31));
AND2X1 exu_U37224(.A(bypass_rs3h_data_d[23]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n33));
AND2X1 exu_U37225(.A(bypass_rs3h_data_d[22]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n35));
AND2X1 exu_U37226(.A(bypass_rs3h_data_d[21]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n37));
AND2X1 exu_U37227(.A(bypass_rs3h_data_d[20]), .B(exu_n16132), .Y(bypass_rs3h_data_dff_n39));
AND2X1 exu_U37228(.A(bypass_rs3h_data_d[19]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n41));
AND2X1 exu_U37229(.A(bypass_rs3h_data_d[18]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n43));
AND2X1 exu_U37230(.A(bypass_rs3h_data_d[17]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n45));
AND2X1 exu_U37231(.A(bypass_rs3h_data_d[16]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n47));
AND2X1 exu_U37232(.A(bypass_rs3h_data_d[15]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n49));
AND2X1 exu_U37233(.A(bypass_rs3h_data_d[14]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n51));
AND2X1 exu_U37234(.A(bypass_rs3h_data_d[13]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n53));
AND2X1 exu_U37235(.A(bypass_rs3h_data_d[12]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n55));
AND2X1 exu_U37236(.A(bypass_rs3h_data_d[11]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n57));
AND2X1 exu_U37237(.A(bypass_rs3h_data_d[10]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n59));
AND2X1 exu_U37238(.A(bypass_rs3h_data_d[9]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n61));
AND2X1 exu_U37239(.A(bypass_rs3h_data_d[8]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n63));
AND2X1 exu_U37240(.A(bypass_rs3h_data_d[7]), .B(exu_n16131), .Y(bypass_rs3h_data_dff_n65));
AND2X1 exu_U37241(.A(ecl_byp_sel_yreg_e), .B(div_byp_yreg_e[9]), .Y(bypass_ifu_exu_sr_mux_n6));
AND2X1 exu_U37242(.A(div_byp_yreg_e[8]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n12));
AND2X1 exu_U37243(.A(div_byp_yreg_e[31]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n240));
AND2X1 exu_U37244(.A(div_byp_yreg_e[30]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n246));
AND2X1 exu_U37245(.A(div_byp_yreg_e[29]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n258));
AND2X1 exu_U37246(.A(div_byp_yreg_e[28]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n264));
AND2X1 exu_U37247(.A(div_byp_yreg_e[27]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n270));
AND2X1 exu_U37248(.A(div_byp_yreg_e[26]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n276));
AND2X1 exu_U37249(.A(div_byp_yreg_e[25]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n282));
AND2X1 exu_U37250(.A(div_byp_yreg_e[24]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n288));
AND2X1 exu_U37251(.A(div_byp_yreg_e[23]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n294));
AND2X1 exu_U37252(.A(div_byp_yreg_e[22]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n300));
AND2X1 exu_U37253(.A(div_byp_yreg_e[21]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n306));
AND2X1 exu_U37254(.A(div_byp_yreg_e[20]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n312));
AND2X1 exu_U37255(.A(div_byp_yreg_e[19]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n324));
AND2X1 exu_U37256(.A(div_byp_yreg_e[18]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n330));
AND2X1 exu_U37257(.A(div_byp_yreg_e[17]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n336));
AND2X1 exu_U37258(.A(div_byp_yreg_e[16]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n342));
AND2X1 exu_U37259(.A(div_byp_yreg_e[15]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n348));
AND2X1 exu_U37260(.A(div_byp_yreg_e[14]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n354));
AND2X1 exu_U37261(.A(div_byp_yreg_e[13]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n360));
AND2X1 exu_U37262(.A(div_byp_yreg_e[12]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n366));
AND2X1 exu_U37263(.A(div_byp_yreg_e[11]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n372));
AND2X1 exu_U37264(.A(div_byp_yreg_e[10]), .B(ecl_byp_sel_yreg_e), .Y(bypass_ifu_exu_sr_mux_n378));
AND2X1 exu_U37265(.A(ecl_cancel_rs3_ecc_e), .B(exu_n16159), .Y(ecl_alu_out_sel_logic_e_l));
BUFX2 exu_U37266(.A(exu_n15024), .Y(exu_n15941));
OR2X1 exu_U37267(.A(se), .B(exu_n16556), .Y(exu_n17476));
INVX1 exu_U37268(.A(exu_n17476), .Y(exu_n15024));
BUFX2 exu_U37269(.A(exu_n15024), .Y(exu_n15942));
BUFX2 exu_U37270(.A(exu_n15024), .Y(exu_n15943));
BUFX2 exu_U37271(.A(exu_n15024), .Y(exu_n15946));
BUFX2 exu_U37272(.A(exu_n15688), .Y(exu_n15947));
AND2X1 exu_U37273(.A(exu_n16396), .B(rml_cwp_n38), .Y(rml_cwp_swap_sel[0]));
INVX1 exu_U37274(.A(rml_cwp_swap_sel[0]), .Y(exu_n15025));
OR2X1 exu_U37275(.A(rml_cwp_n74), .B(rml_cwp_swap_sel_tlu[0]), .Y(rml_cwp_slot0_data_mux_sel2));
INVX1 exu_U37276(.A(rml_cwp_slot0_data_mux_sel2), .Y(exu_n15026));
INVX1 exu_U37277(.A(rml_cwp_N99), .Y(exu_n15027));
INVX1 exu_U37278(.A(ecl_ecc_log_rs1_m), .Y(exu_n15028));
AND2X1 exu_U37279(.A(ecl_thr_match_de), .B(exu_n15235), .Y(ecl_ccr_n40));
INVX1 exu_U37280(.A(ecl_ccr_n40), .Y(exu_n15029));
OR2X1 exu_U37281(.A(exu_n16604), .B(exu_n15344), .Y(rml_ecl_fill_e));
INVX1 exu_U37282(.A(rml_ecl_fill_e), .Y(exu_n15030));
BUFX2 exu_U37283(.A(ecl_irf_wen_w), .Y(exu_n15031));
INVX1 exu_U37284(.A(exu_n31727), .Y(exu_lsu_rs3_data_e[9]));
INVX1 exu_U37285(.A(exu_n31741), .Y(exu_ifu_cc_d[7]));
BUFX2 exu_U37286(.A(ecl_irf_tid_m[1]), .Y(exu_n15034));
BUFX2 exu_U37287(.A(ecl_irf_tid_m[0]), .Y(exu_n15035));
INVX1 exu_U37288(.A(exu_n31728), .Y(exu_lsu_rs3_data_e[8]));
INVX1 exu_U37289(.A(exu_n31729), .Y(exu_lsu_rs3_data_e[7]));
INVX1 exu_U37290(.A(exu_n31730), .Y(exu_lsu_rs3_data_e[6]));
INVX1 exu_U37291(.A(exu_n31731), .Y(exu_lsu_rs3_data_e[5]));
INVX1 exu_U37292(.A(exu_n31732), .Y(exu_lsu_rs3_data_e[4]));
INVX1 exu_U37293(.A(exu_n31733), .Y(exu_lsu_rs3_data_e[3]));
INVX1 exu_U37294(.A(exu_n31705), .Y(exu_lsu_rs3_data_e[31]));
INVX1 exu_U37295(.A(exu_n31706), .Y(exu_lsu_rs3_data_e[30]));
INVX1 exu_U37296(.A(exu_n31734), .Y(exu_lsu_rs3_data_e[2]));
INVX1 exu_U37297(.A(exu_n31707), .Y(exu_lsu_rs3_data_e[29]));
INVX1 exu_U37298(.A(exu_n31708), .Y(exu_lsu_rs3_data_e[28]));
INVX1 exu_U37299(.A(exu_n31709), .Y(exu_lsu_rs3_data_e[27]));
INVX1 exu_U37300(.A(exu_n31710), .Y(exu_lsu_rs3_data_e[26]));
INVX1 exu_U37301(.A(exu_n31711), .Y(exu_lsu_rs3_data_e[25]));
INVX1 exu_U37302(.A(exu_n31712), .Y(exu_lsu_rs3_data_e[24]));
INVX1 exu_U37303(.A(exu_n31713), .Y(exu_lsu_rs3_data_e[23]));
INVX1 exu_U37304(.A(exu_n31714), .Y(exu_lsu_rs3_data_e[22]));
INVX1 exu_U37305(.A(exu_n31715), .Y(exu_lsu_rs3_data_e[21]));
INVX1 exu_U37306(.A(exu_n31716), .Y(exu_lsu_rs3_data_e[20]));
INVX1 exu_U37307(.A(exu_n31735), .Y(exu_lsu_rs3_data_e[1]));
INVX1 exu_U37308(.A(exu_n31717), .Y(exu_lsu_rs3_data_e[19]));
INVX1 exu_U37309(.A(exu_n31718), .Y(exu_lsu_rs3_data_e[18]));
INVX1 exu_U37310(.A(exu_n31719), .Y(exu_lsu_rs3_data_e[17]));
INVX1 exu_U37311(.A(exu_n31720), .Y(exu_lsu_rs3_data_e[16]));
INVX1 exu_U37312(.A(exu_n31721), .Y(exu_lsu_rs3_data_e[15]));
INVX1 exu_U37313(.A(exu_n31722), .Y(exu_lsu_rs3_data_e[14]));
INVX1 exu_U37314(.A(exu_n31723), .Y(exu_lsu_rs3_data_e[13]));
INVX1 exu_U37315(.A(exu_n31724), .Y(exu_lsu_rs3_data_e[12]));
INVX1 exu_U37316(.A(exu_n31725), .Y(exu_lsu_rs3_data_e[11]));
INVX1 exu_U37317(.A(exu_n31726), .Y(exu_lsu_rs3_data_e[10]));
INVX1 exu_U37318(.A(exu_n31736), .Y(exu_lsu_rs3_data_e[0]));
INVX1 exu_U37319(.A(exu_n31742), .Y(exu_ifu_cc_d[6]));
INVX1 exu_U37320(.A(exu_n31743), .Y(exu_ifu_cc_d[5]));
INVX1 exu_U37321(.A(exu_n31744), .Y(exu_ifu_cc_d[4]));
INVX1 exu_U37322(.A(exu_n31746), .Y(exu_ifu_cc_d[2]));
INVX1 exu_U37323(.A(exu_n31739), .Y(exu_ifu_err_reg_m[4]));
INVX1 exu_U37324(.A(exu_n31740), .Y(exu_ifu_err_reg_m[3]));
INVX1 exu_U37325(.A(exu_n18423), .Y(exu_n15073));
INVX1 exu_U37326(.A(exu_n18428), .Y(exu_n15074));
INVX1 exu_U37327(.A(ecl_divcntl_cnt6_n10), .Y(exu_n15075));
INVX1 exu_U37328(.A(rml_cwp_inc_n3), .Y(exu_n15076));
AND2X1 exu_U37329(.A(div_ecl_d_62), .B(exu_n15372), .Y(ecl_divcntl_n51));
INVX1 exu_U37330(.A(ecl_divcntl_n51), .Y(exu_n15077));
OR2X1 exu_U37331(.A(exu_n15510), .B(exu_n15774), .Y(ecc_error_data_m[63]));
INVX1 exu_U37332(.A(ecc_error_data_m[63]), .Y(exu_n15078));
OR2X1 exu_U37333(.A(exu_n15510), .B(exu_n15506), .Y(ecc_error_data_m[62]));
INVX1 exu_U37334(.A(ecc_error_data_m[62]), .Y(exu_n15079));
OR2X1 exu_U37335(.A(exu_n15509), .B(exu_n15774), .Y(ecc_error_data_m[61]));
INVX1 exu_U37336(.A(ecc_error_data_m[61]), .Y(exu_n15080));
OR2X1 exu_U37337(.A(exu_n15509), .B(exu_n15506), .Y(ecc_error_data_m[60]));
INVX1 exu_U37338(.A(ecc_error_data_m[60]), .Y(exu_n15081));
OR2X1 exu_U37339(.A(exu_n15511), .B(exu_n15774), .Y(ecc_error_data_m[59]));
INVX1 exu_U37340(.A(ecc_error_data_m[59]), .Y(exu_n15082));
OR2X1 exu_U37341(.A(exu_n15511), .B(exu_n15506), .Y(ecc_error_data_m[58]));
INVX1 exu_U37342(.A(ecc_error_data_m[58]), .Y(exu_n15083));
OR2X1 exu_U37343(.A(exu_n15774), .B(exu_n15516), .Y(ecc_error_data_m[57]));
INVX1 exu_U37344(.A(ecc_error_data_m[57]), .Y(exu_n15084));
OR2X1 exu_U37345(.A(exu_n15937), .B(exu_n15770), .Y(ecc_error_data_m[56]));
INVX1 exu_U37346(.A(ecc_error_data_m[56]), .Y(exu_n15085));
OR2X1 exu_U37347(.A(exu_n15936), .B(exu_n15770), .Y(ecc_error_data_m[55]));
INVX1 exu_U37348(.A(ecc_error_data_m[55]), .Y(exu_n15086));
OR2X1 exu_U37349(.A(exu_n15937), .B(exu_n15771), .Y(ecc_error_data_m[54]));
INVX1 exu_U37350(.A(ecc_error_data_m[54]), .Y(exu_n15087));
OR2X1 exu_U37351(.A(exu_n15936), .B(exu_n15771), .Y(ecc_error_data_m[53]));
INVX1 exu_U37352(.A(ecc_error_data_m[53]), .Y(exu_n15088));
OR2X1 exu_U37353(.A(exu_n15937), .B(exu_n15772), .Y(ecc_error_data_m[52]));
INVX1 exu_U37354(.A(ecc_error_data_m[52]), .Y(exu_n15089));
OR2X1 exu_U37355(.A(exu_n15936), .B(exu_n15772), .Y(ecc_error_data_m[51]));
INVX1 exu_U37356(.A(ecc_error_data_m[51]), .Y(exu_n15090));
OR2X1 exu_U37357(.A(exu_n15937), .B(exu_n15773), .Y(ecc_error_data_m[50]));
INVX1 exu_U37358(.A(ecc_error_data_m[50]), .Y(exu_n15091));
INVX1 exu_U37359(.A(ecc_error_data_m[4]), .Y(exu_n15092));
OR2X1 exu_U37360(.A(exu_n15936), .B(exu_n15773), .Y(ecc_error_data_m[49]));
INVX1 exu_U37361(.A(ecc_error_data_m[49]), .Y(exu_n15093));
OR2X1 exu_U37362(.A(exu_n15770), .B(exu_n15938), .Y(ecc_error_data_m[48]));
INVX1 exu_U37363(.A(ecc_error_data_m[48]), .Y(exu_n15094));
OR2X1 exu_U37364(.A(exu_n15770), .B(exu_n15932), .Y(ecc_error_data_m[47]));
INVX1 exu_U37365(.A(ecc_error_data_m[47]), .Y(exu_n15095));
OR2X1 exu_U37366(.A(exu_n15771), .B(exu_n15938), .Y(ecc_error_data_m[46]));
INVX1 exu_U37367(.A(ecc_error_data_m[46]), .Y(exu_n15096));
OR2X1 exu_U37368(.A(exu_n15771), .B(exu_n15932), .Y(ecc_error_data_m[45]));
INVX1 exu_U37369(.A(ecc_error_data_m[45]), .Y(exu_n15097));
OR2X1 exu_U37370(.A(exu_n15772), .B(exu_n15938), .Y(ecc_error_data_m[44]));
INVX1 exu_U37371(.A(ecc_error_data_m[44]), .Y(exu_n15098));
OR2X1 exu_U37372(.A(exu_n15772), .B(exu_n15932), .Y(ecc_error_data_m[43]));
INVX1 exu_U37373(.A(ecc_error_data_m[43]), .Y(exu_n15099));
OR2X1 exu_U37374(.A(exu_n15773), .B(exu_n15938), .Y(ecc_error_data_m[42]));
INVX1 exu_U37375(.A(ecc_error_data_m[42]), .Y(exu_n15100));
OR2X1 exu_U37376(.A(exu_n15773), .B(exu_n15932), .Y(ecc_error_data_m[41]));
INVX1 exu_U37377(.A(ecc_error_data_m[41]), .Y(exu_n15101));
OR2X1 exu_U37378(.A(exu_n15937), .B(exu_n15776), .Y(ecc_error_data_m[40]));
INVX1 exu_U37379(.A(ecc_error_data_m[40]), .Y(exu_n15102));
OR2X1 exu_U37380(.A(exu_n15936), .B(exu_n15776), .Y(ecc_error_data_m[39]));
INVX1 exu_U37381(.A(ecc_error_data_m[39]), .Y(exu_n15103));
OR2X1 exu_U37382(.A(exu_n15937), .B(exu_n15777), .Y(ecc_error_data_m[38]));
INVX1 exu_U37383(.A(ecc_error_data_m[38]), .Y(exu_n15104));
OR2X1 exu_U37384(.A(exu_n15936), .B(exu_n15777), .Y(ecc_error_data_m[37]));
INVX1 exu_U37385(.A(ecc_error_data_m[37]), .Y(exu_n15105));
OR2X1 exu_U37386(.A(exu_n15937), .B(exu_n15778), .Y(ecc_error_data_m[36]));
INVX1 exu_U37387(.A(ecc_error_data_m[36]), .Y(exu_n15106));
OR2X1 exu_U37388(.A(exu_n15936), .B(exu_n15778), .Y(ecc_error_data_m[35]));
INVX1 exu_U37389(.A(ecc_error_data_m[35]), .Y(exu_n15107));
OR2X1 exu_U37390(.A(exu_n15937), .B(exu_n15507), .Y(ecc_error_data_m[34]));
INVX1 exu_U37391(.A(ecc_error_data_m[34]), .Y(exu_n15108));
OR2X1 exu_U37392(.A(exu_n15936), .B(exu_n15507), .Y(ecc_error_data_m[33]));
INVX1 exu_U37393(.A(ecc_error_data_m[33]), .Y(exu_n15109));
OR2X1 exu_U37394(.A(exu_n15938), .B(exu_n15776), .Y(ecc_error_data_m[32]));
INVX1 exu_U37395(.A(ecc_error_data_m[32]), .Y(exu_n15110));
OR2X1 exu_U37396(.A(exu_n15932), .B(exu_n15776), .Y(ecc_error_data_m[31]));
INVX1 exu_U37397(.A(ecc_error_data_m[31]), .Y(exu_n15111));
OR2X1 exu_U37398(.A(exu_n15938), .B(exu_n15777), .Y(ecc_error_data_m[30]));
INVX1 exu_U37399(.A(ecc_error_data_m[30]), .Y(exu_n15112));
OR2X1 exu_U37400(.A(exu_n15932), .B(exu_n15777), .Y(ecc_error_data_m[29]));
INVX1 exu_U37401(.A(ecc_error_data_m[29]), .Y(exu_n15113));
OR2X1 exu_U37402(.A(exu_n15938), .B(exu_n15778), .Y(ecc_error_data_m[28]));
INVX1 exu_U37403(.A(ecc_error_data_m[28]), .Y(exu_n15114));
OR2X1 exu_U37404(.A(exu_n15932), .B(exu_n15778), .Y(ecc_error_data_m[27]));
INVX1 exu_U37405(.A(ecc_error_data_m[27]), .Y(exu_n15115));
OR2X1 exu_U37406(.A(exu_n15938), .B(exu_n15507), .Y(ecc_error_data_m[26]));
INVX1 exu_U37407(.A(ecc_error_data_m[26]), .Y(exu_n15116));
INVX1 exu_U37408(.A(rml_n36), .Y(exu_n15117));
INVX1 exu_U37409(.A(alu_va_e[63]), .Y(exu_n15118));
AND2X1 exu_U37410(.A(exu_n15547), .B(exu_n15857), .Y(rml_n57));
INVX1 exu_U37411(.A(rml_n57), .Y(exu_n15119));
AND2X1 exu_U37412(.A(exu_n15548), .B(exu_n15553), .Y(rml_n58));
INVX1 exu_U37413(.A(rml_n58), .Y(exu_n15120));
AND2X1 exu_U37414(.A(ecl_rd_e[3]), .B(ecl_n44), .Y(ecl_n43));
INVX1 exu_U37415(.A(ecl_n43), .Y(exu_n15121));
AND2X1 exu_U37416(.A(ifu_exu_usecin_d), .B(exu_ifu_cc_d[0]), .Y(ecl_n76));
INVX1 exu_U37417(.A(ecl_n76), .Y(exu_n15122));
INVX1 exu_U37418(.A(ecc_ecc_datain_m[9]), .Y(exu_n15123));
INVX1 exu_U37419(.A(ecc_ecc_datain_m[8]), .Y(exu_n15124));
INVX1 exu_U37420(.A(ecc_ecc_datain_m[7]), .Y(exu_n15125));
INVX1 exu_U37421(.A(ecc_ecc_datain_m[6]), .Y(exu_n15126));
INVX1 exu_U37422(.A(ecc_ecc_datain_m[63]), .Y(exu_n15127));
INVX1 exu_U37423(.A(ecc_ecc_datain_m[62]), .Y(exu_n15128));
INVX1 exu_U37424(.A(ecc_ecc_datain_m[61]), .Y(exu_n15129));
INVX1 exu_U37425(.A(ecc_ecc_datain_m[60]), .Y(exu_n15130));
INVX1 exu_U37426(.A(ecc_ecc_datain_m[5]), .Y(exu_n15131));
INVX1 exu_U37427(.A(ecc_ecc_datain_m[59]), .Y(exu_n15132));
INVX1 exu_U37428(.A(ecc_ecc_datain_m[58]), .Y(exu_n15133));
INVX1 exu_U37429(.A(ecc_ecc_datain_m[57]), .Y(exu_n15134));
INVX1 exu_U37430(.A(ecc_ecc_datain_m[56]), .Y(exu_n15135));
INVX1 exu_U37431(.A(ecc_ecc_datain_m[55]), .Y(exu_n15136));
INVX1 exu_U37432(.A(ecc_ecc_datain_m[54]), .Y(exu_n15137));
INVX1 exu_U37433(.A(ecc_ecc_datain_m[53]), .Y(exu_n15138));
INVX1 exu_U37434(.A(ecc_ecc_datain_m[52]), .Y(exu_n15139));
INVX1 exu_U37435(.A(ecc_ecc_datain_m[51]), .Y(exu_n15140));
INVX1 exu_U37436(.A(ecc_ecc_datain_m[50]), .Y(exu_n15141));
INVX1 exu_U37437(.A(ecc_ecc_datain_m[4]), .Y(exu_n15142));
INVX1 exu_U37438(.A(ecc_ecc_datain_m[49]), .Y(exu_n15143));
INVX1 exu_U37439(.A(ecc_ecc_datain_m[48]), .Y(exu_n15144));
INVX1 exu_U37440(.A(ecc_ecc_datain_m[47]), .Y(exu_n15145));
INVX1 exu_U37441(.A(ecc_ecc_datain_m[46]), .Y(exu_n15146));
INVX1 exu_U37442(.A(ecc_ecc_datain_m[45]), .Y(exu_n15147));
INVX1 exu_U37443(.A(ecc_ecc_datain_m[44]), .Y(exu_n15148));
INVX1 exu_U37444(.A(ecc_ecc_datain_m[43]), .Y(exu_n15149));
INVX1 exu_U37445(.A(ecc_ecc_datain_m[42]), .Y(exu_n15150));
INVX1 exu_U37446(.A(ecc_ecc_datain_m[41]), .Y(exu_n15151));
INVX1 exu_U37447(.A(ecc_ecc_datain_m[40]), .Y(exu_n15152));
INVX1 exu_U37448(.A(ecc_ecc_datain_m[3]), .Y(exu_n15153));
INVX1 exu_U37449(.A(ecc_ecc_datain_m[39]), .Y(exu_n15154));
INVX1 exu_U37450(.A(ecc_ecc_datain_m[38]), .Y(exu_n15155));
INVX1 exu_U37451(.A(ecc_ecc_datain_m[37]), .Y(exu_n15156));
INVX1 exu_U37452(.A(ecc_ecc_datain_m[36]), .Y(exu_n15157));
INVX1 exu_U37453(.A(ecc_ecc_datain_m[35]), .Y(exu_n15158));
INVX1 exu_U37454(.A(ecc_ecc_datain_m[34]), .Y(exu_n15159));
INVX1 exu_U37455(.A(ecc_ecc_datain_m[33]), .Y(exu_n15160));
INVX1 exu_U37456(.A(ecc_ecc_datain_m[32]), .Y(exu_n15161));
INVX1 exu_U37457(.A(ecc_ecc_datain_m[31]), .Y(exu_n15162));
INVX1 exu_U37458(.A(ecc_ecc_datain_m[30]), .Y(exu_n15163));
INVX1 exu_U37459(.A(ecc_ecc_datain_m[2]), .Y(exu_n15164));
INVX1 exu_U37460(.A(ecc_ecc_datain_m[29]), .Y(exu_n15165));
INVX1 exu_U37461(.A(ecc_ecc_datain_m[28]), .Y(exu_n15166));
INVX1 exu_U37462(.A(ecc_ecc_datain_m[27]), .Y(exu_n15167));
INVX1 exu_U37463(.A(ecc_ecc_datain_m[26]), .Y(exu_n15168));
INVX1 exu_U37464(.A(ecc_ecc_datain_m[25]), .Y(exu_n15169));
INVX1 exu_U37465(.A(ecc_ecc_datain_m[24]), .Y(exu_n15170));
INVX1 exu_U37466(.A(ecc_ecc_datain_m[23]), .Y(exu_n15171));
INVX1 exu_U37467(.A(ecc_ecc_datain_m[22]), .Y(exu_n15172));
INVX1 exu_U37468(.A(ecc_ecc_datain_m[21]), .Y(exu_n15173));
INVX1 exu_U37469(.A(ecc_ecc_datain_m[20]), .Y(exu_n15174));
INVX1 exu_U37470(.A(ecc_ecc_datain_m[1]), .Y(exu_n15175));
INVX1 exu_U37471(.A(ecc_ecc_datain_m[19]), .Y(exu_n15176));
INVX1 exu_U37472(.A(ecc_ecc_datain_m[18]), .Y(exu_n15177));
INVX1 exu_U37473(.A(ecc_ecc_datain_m[17]), .Y(exu_n15178));
INVX1 exu_U37474(.A(ecc_ecc_datain_m[16]), .Y(exu_n15179));
INVX1 exu_U37475(.A(ecc_ecc_datain_m[15]), .Y(exu_n15180));
INVX1 exu_U37476(.A(ecc_ecc_datain_m[14]), .Y(exu_n15181));
INVX1 exu_U37477(.A(ecc_ecc_datain_m[13]), .Y(exu_n15182));
INVX1 exu_U37478(.A(ecc_ecc_datain_m[12]), .Y(exu_n15183));
INVX1 exu_U37479(.A(ecc_ecc_datain_m[11]), .Y(exu_n15184));
INVX1 exu_U37480(.A(ecc_ecc_datain_m[10]), .Y(exu_n15185));
INVX1 exu_U37481(.A(ecc_ecc_datain_m[0]), .Y(exu_n15186));
INVX1 exu_U37482(.A(div_gencc_in[32]), .Y(exu_n15187));
INVX1 exu_U37483(.A(exu_n15189), .Y(exu_n15188));
INVX1 exu_U37484(.A(exu_n15191), .Y(exu_n15190));
INVX1 exu_U37485(.A(exu_n15193), .Y(exu_n15192));
AND2X1 exu_U37486(.A(rml_wstate_wen_w), .B(ecl_rml_thr_w[3]), .Y(exu_n18323));
INVX1 exu_U37487(.A(exu_n18323), .Y(exu_n15194));
AND2X1 exu_U37488(.A(ecl_rml_thr_w[2]), .B(rml_wstate_wen_w), .Y(exu_n18324));
INVX1 exu_U37489(.A(exu_n18324), .Y(exu_n15195));
AND2X1 exu_U37490(.A(exu_n15957), .B(rml_wstate_wen_w), .Y(exu_n18325));
INVX1 exu_U37491(.A(exu_n18325), .Y(exu_n15196));
AND2X1 exu_U37492(.A(exu_n15959), .B(rml_wstate_wen_w), .Y(exu_n18326));
INVX1 exu_U37493(.A(exu_n18326), .Y(exu_n15197));
AND2X1 exu_U37494(.A(ecl_divcntl_n80), .B(exu_n16247), .Y(ecl_divcntl_n67));
INVX1 exu_U37495(.A(ecl_divcntl_n67), .Y(exu_n15198));
INVX1 exu_U37496(.A(ecc_decode_n23), .Y(exu_n15199));
OR2X1 exu_U37497(.A(exu_n15480), .B(exu_n15396), .Y(ecc_decode_n49));
INVX1 exu_U37498(.A(ecc_decode_n49), .Y(exu_n15200));
AND2X1 exu_U37499(.A(ifu_exu_useimm_d), .B(ecl_writeback_n19), .Y(ecl_byplog_rs2_n12));
INVX1 exu_U37500(.A(ecl_byplog_rs2_n12), .Y(exu_n15201));
OR2X1 exu_U37501(.A(ecc_err_m[5]), .B(exu_n15480), .Y(ecc_decode_n38));
INVX1 exu_U37502(.A(ecc_decode_n38), .Y(exu_n15202));
INVX1 exu_U37503(.A(ecl_byplog_rs1_n38), .Y(exu_n15203));
INVX1 exu_U37504(.A(div_ecl_detect_zero_high), .Y(exu_n15204));
OR2X1 exu_U37505(.A(ecc_ecl_rs1_ce), .B(ecc_ecl_rs2_ce), .Y(ecl_eccctl_ecc_sel_rs3_dff_din[0]));
INVX1 exu_U37506(.A(ecl_eccctl_ecc_sel_rs3_dff_din[0]), .Y(exu_n15205));
INVX1 exu_U37507(.A(div_ecl_detect_zero_low), .Y(exu_n15206));
INVX1 exu_U37508(.A(ecl_byplog_rs1_N2), .Y(exu_n15207));
INVX1 exu_U37509(.A(ecl_byplog_rs2_N2), .Y(exu_n15208));
INVX1 exu_U37510(.A(ecl_byplog_rs3h_N2), .Y(exu_n15209));
INVX1 exu_U37511(.A(ecl_byplog_rs3_N2), .Y(exu_n15210));
INVX1 exu_U37512(.A(bypass_rs1_data_w2[9]), .Y(exu_n15211));
INVX1 exu_U37513(.A(ecl_n62), .Y(exu_n15212));
AND2X1 exu_U37514(.A(rml_cwp_valid_tlu_swap_w), .B(ecl_rml_thr_w[3]), .Y(rml_cwp_n71));
INVX1 exu_U37515(.A(rml_cwp_n71), .Y(exu_n15213));
AND2X1 exu_U37516(.A(rml_cwp_valid_tlu_swap_w), .B(ecl_rml_thr_w[2]), .Y(rml_cwp_n69));
INVX1 exu_U37517(.A(rml_cwp_n69), .Y(exu_n15214));
AND2X1 exu_U37518(.A(rml_cwp_valid_tlu_swap_w), .B(exu_n15958), .Y(rml_cwp_n67));
INVX1 exu_U37519(.A(rml_cwp_n67), .Y(exu_n15215));
AND2X1 exu_U37520(.A(rml_cwp_valid_tlu_swap_w), .B(exu_n15960), .Y(rml_cwp_n65));
INVX1 exu_U37521(.A(rml_cwp_n65), .Y(exu_n15216));
INVX1 exu_U37522(.A(ecl_writeback_n74), .Y(exu_n15217));
INVX1 exu_U37523(.A(ecl_writeback_n78), .Y(exu_n15218));
OR2X1 exu_U37524(.A(exu_n15775), .B(ecl_writeback_n181), .Y(ecl_writeback_n82));
INVX1 exu_U37525(.A(ecl_writeback_n82), .Y(exu_n15219));
INVX1 exu_U37526(.A(ecl_writeback_n86), .Y(exu_n15220));
OR2X1 exu_U37527(.A(ecl_divcntl_gencc_in_msb_l_d1), .B(ecl_divcntl_inputs_neg_q), .Y(ecl_divcntl_n78));
INVX1 exu_U37528(.A(ecl_divcntl_n78), .Y(exu_n15221));
AND2X1 exu_U37529(.A(ecl_ifu_exu_rs1_d[0]), .B(exu_n16559), .Y(exu_n16630));
INVX1 exu_U37530(.A(exu_n16630), .Y(exu_n15222));
AND2X1 exu_U37531(.A(ecl_ifu_exu_rs1_d[0]), .B(exu_n16565), .Y(exu_n16644));
INVX1 exu_U37532(.A(exu_n16644), .Y(exu_n15223));
AND2X1 exu_U37533(.A(ecl_ifu_exu_rs1_d[0]), .B(exu_n16561), .Y(exu_n16658));
INVX1 exu_U37534(.A(exu_n16658), .Y(exu_n15224));
AND2X1 exu_U37535(.A(ecl_ifu_exu_rs1_d[0]), .B(exu_n16563), .Y(exu_n16672));
INVX1 exu_U37536(.A(exu_n16672), .Y(exu_n15225));
AND2X1 exu_U37537(.A(ecl_ifu_exu_rs2_d[0]), .B(exu_n16559), .Y(exu_n16686));
INVX1 exu_U37538(.A(exu_n16686), .Y(exu_n15226));
AND2X1 exu_U37539(.A(ecl_ifu_exu_rs2_d[0]), .B(exu_n16565), .Y(exu_n16700));
INVX1 exu_U37540(.A(exu_n16700), .Y(exu_n15227));
AND2X1 exu_U37541(.A(ecl_ifu_exu_rs2_d[0]), .B(exu_n16561), .Y(exu_n16714));
INVX1 exu_U37542(.A(exu_n16714), .Y(exu_n15228));
AND2X1 exu_U37543(.A(ecl_ifu_exu_rs2_d[0]), .B(exu_n16563), .Y(exu_n16728));
INVX1 exu_U37544(.A(exu_n16728), .Y(exu_n15229));
AND2X1 exu_U37545(.A(ecl_ifu_exu_rs3_d[0]), .B(exu_n16559), .Y(exu_n17406));
INVX1 exu_U37546(.A(exu_n17406), .Y(exu_n15230));
AND2X1 exu_U37547(.A(ecl_ifu_exu_rs3_d[0]), .B(exu_n16565), .Y(exu_n17420));
INVX1 exu_U37548(.A(exu_n17420), .Y(exu_n15231));
AND2X1 exu_U37549(.A(ecl_ifu_exu_rs3_d[0]), .B(exu_n16561), .Y(exu_n17434));
INVX1 exu_U37550(.A(exu_n17434), .Y(exu_n15232));
AND2X1 exu_U37551(.A(ecl_ifu_exu_rs3_d[0]), .B(exu_n16563), .Y(exu_n17448));
INVX1 exu_U37552(.A(exu_n17448), .Y(exu_n15233));
INVX1 exu_U37553(.A(rml_cwp_next_swap_thr[0]), .Y(exu_n15234));
OR2X1 exu_U37554(.A(exu_n16602), .B(ecl_rml_kill_e), .Y(ecl_ccr_valid_setcc_e));
INVX1 exu_U37555(.A(ecl_ccr_valid_setcc_e), .Y(exu_n15235));
INVX1 exu_U37556(.A(ecl_divcntl_wb_req_g), .Y(exu_n15236));
OR2X1 exu_U37557(.A(ecl_bypass_m), .B(ecl_writeback_wrsr_m), .Y(ecl_writeback_n199));
INVX1 exu_U37558(.A(ecl_writeback_n199), .Y(exu_n15237));
AND2X1 exu_U37559(.A(exu_n15382), .B(exu_n15761), .Y(ecl_writeback_n73));
INVX1 exu_U37560(.A(ecl_writeback_n73), .Y(exu_n15238));
AND2X1 exu_U37561(.A(ecl_ifu_exu_tv_e), .B(ecl_adder_icc[1]), .Y(ecl_n120));
INVX1 exu_U37562(.A(ecl_n120), .Y(exu_n15239));
INVX1 exu_U37563(.A(div_xin[41]), .Y(exu_n15240));
INVX1 exu_U37564(.A(div_xin[40]), .Y(exu_n15241));
INVX1 exu_U37565(.A(div_xin[39]), .Y(exu_n15242));
INVX1 exu_U37566(.A(div_xin[38]), .Y(exu_n15243));
INVX1 exu_U37567(.A(div_xin[37]), .Y(exu_n15244));
INVX1 exu_U37568(.A(div_xin[36]), .Y(exu_n15245));
INVX1 exu_U37569(.A(div_xin[35]), .Y(exu_n15246));
INVX1 exu_U37570(.A(div_xin[62]), .Y(exu_n15247));
INVX1 exu_U37571(.A(div_xin[34]), .Y(exu_n15248));
INVX1 exu_U37572(.A(div_xin[61]), .Y(exu_n15249));
INVX1 exu_U37573(.A(div_xin[60]), .Y(exu_n15250));
INVX1 exu_U37574(.A(div_xin[59]), .Y(exu_n15251));
INVX1 exu_U37575(.A(div_xin[58]), .Y(exu_n15252));
INVX1 exu_U37576(.A(div_xin[57]), .Y(exu_n15253));
INVX1 exu_U37577(.A(div_xin[56]), .Y(exu_n15254));
INVX1 exu_U37578(.A(div_xin[55]), .Y(exu_n15255));
INVX1 exu_U37579(.A(div_xin[54]), .Y(exu_n15256));
INVX1 exu_U37580(.A(div_xin[53]), .Y(exu_n15257));
INVX1 exu_U37581(.A(div_xin[52]), .Y(exu_n15258));
INVX1 exu_U37582(.A(div_xin[33]), .Y(exu_n15259));
INVX1 exu_U37583(.A(div_xin[51]), .Y(exu_n15260));
INVX1 exu_U37584(.A(div_xin[50]), .Y(exu_n15261));
INVX1 exu_U37585(.A(div_xin[49]), .Y(exu_n15262));
INVX1 exu_U37586(.A(div_xin[48]), .Y(exu_n15263));
INVX1 exu_U37587(.A(div_xin[47]), .Y(exu_n15264));
INVX1 exu_U37588(.A(div_xin[46]), .Y(exu_n15265));
INVX1 exu_U37589(.A(div_xin[45]), .Y(exu_n15266));
INVX1 exu_U37590(.A(div_xin[44]), .Y(exu_n15267));
INVX1 exu_U37591(.A(div_xin[43]), .Y(exu_n15268));
INVX1 exu_U37592(.A(div_xin[42]), .Y(exu_n15269));
INVX1 exu_U37593(.A(div_xin[32]), .Y(exu_n15270));
INVX1 exu_U37594(.A(bypass_rs1_data_w2[8]), .Y(exu_n15271));
INVX1 exu_U37595(.A(bypass_rs1_data_w2[7]), .Y(exu_n15272));
INVX1 exu_U37596(.A(bypass_rs1_data_w2[6]), .Y(exu_n15273));
INVX1 exu_U37597(.A(bypass_rs1_data_w2[63]), .Y(exu_n15274));
INVX1 exu_U37598(.A(bypass_rs1_data_w2[62]), .Y(exu_n15275));
INVX1 exu_U37599(.A(bypass_rs1_data_w2[61]), .Y(exu_n15276));
INVX1 exu_U37600(.A(bypass_rs1_data_w2[60]), .Y(exu_n15277));
INVX1 exu_U37601(.A(bypass_rs1_data_w2[5]), .Y(exu_n15278));
INVX1 exu_U37602(.A(bypass_rs1_data_w2[59]), .Y(exu_n15279));
INVX1 exu_U37603(.A(bypass_rs1_data_w2[58]), .Y(exu_n15280));
INVX1 exu_U37604(.A(bypass_rs1_data_w2[57]), .Y(exu_n15281));
INVX1 exu_U37605(.A(bypass_rs1_data_w2[56]), .Y(exu_n15282));
INVX1 exu_U37606(.A(bypass_rs1_data_w2[55]), .Y(exu_n15283));
INVX1 exu_U37607(.A(bypass_rs1_data_w2[54]), .Y(exu_n15284));
INVX1 exu_U37608(.A(bypass_rs1_data_w2[53]), .Y(exu_n15285));
INVX1 exu_U37609(.A(bypass_rs1_data_w2[52]), .Y(exu_n15286));
INVX1 exu_U37610(.A(bypass_rs1_data_w2[51]), .Y(exu_n15287));
INVX1 exu_U37611(.A(bypass_rs1_data_w2[50]), .Y(exu_n15288));
INVX1 exu_U37612(.A(bypass_rs1_data_w2[4]), .Y(exu_n15289));
INVX1 exu_U37613(.A(bypass_rs1_data_w2[49]), .Y(exu_n15290));
INVX1 exu_U37614(.A(bypass_rs1_data_w2[48]), .Y(exu_n15291));
INVX1 exu_U37615(.A(bypass_rs1_data_w2[47]), .Y(exu_n15292));
INVX1 exu_U37616(.A(bypass_rs1_data_w2[46]), .Y(exu_n15293));
INVX1 exu_U37617(.A(bypass_rs1_data_w2[45]), .Y(exu_n15294));
INVX1 exu_U37618(.A(bypass_rs1_data_w2[44]), .Y(exu_n15295));
INVX1 exu_U37619(.A(bypass_rs1_data_w2[43]), .Y(exu_n15296));
INVX1 exu_U37620(.A(bypass_rs1_data_w2[42]), .Y(exu_n15297));
INVX1 exu_U37621(.A(bypass_rs1_data_w2[41]), .Y(exu_n15298));
INVX1 exu_U37622(.A(bypass_rs1_data_w2[40]), .Y(exu_n15299));
INVX1 exu_U37623(.A(bypass_rs1_data_w2[3]), .Y(exu_n15300));
INVX1 exu_U37624(.A(bypass_rs1_data_w2[39]), .Y(exu_n15301));
INVX1 exu_U37625(.A(bypass_rs1_data_w2[38]), .Y(exu_n15302));
INVX1 exu_U37626(.A(bypass_rs1_data_w2[37]), .Y(exu_n15303));
INVX1 exu_U37627(.A(bypass_rs1_data_w2[36]), .Y(exu_n15304));
INVX1 exu_U37628(.A(bypass_rs1_data_w2[35]), .Y(exu_n15305));
INVX1 exu_U37629(.A(bypass_rs1_data_w2[34]), .Y(exu_n15306));
INVX1 exu_U37630(.A(bypass_rs1_data_w2[33]), .Y(exu_n15307));
INVX1 exu_U37631(.A(bypass_rs1_data_w2[32]), .Y(exu_n15308));
INVX1 exu_U37632(.A(bypass_rs1_data_w2[31]), .Y(exu_n15309));
INVX1 exu_U37633(.A(bypass_rs1_data_w2[30]), .Y(exu_n15310));
INVX1 exu_U37634(.A(bypass_rs1_data_w2[2]), .Y(exu_n15311));
INVX1 exu_U37635(.A(bypass_rs1_data_w2[29]), .Y(exu_n15312));
INVX1 exu_U37636(.A(bypass_rs1_data_w2[28]), .Y(exu_n15313));
INVX1 exu_U37637(.A(bypass_rs1_data_w2[27]), .Y(exu_n15314));
INVX1 exu_U37638(.A(bypass_rs1_data_w2[26]), .Y(exu_n15315));
INVX1 exu_U37639(.A(bypass_rs1_data_w2[25]), .Y(exu_n15316));
INVX1 exu_U37640(.A(bypass_rs1_data_w2[24]), .Y(exu_n15317));
INVX1 exu_U37641(.A(bypass_rs1_data_w2[23]), .Y(exu_n15318));
INVX1 exu_U37642(.A(bypass_rs1_data_w2[22]), .Y(exu_n15319));
INVX1 exu_U37643(.A(bypass_rs1_data_w2[21]), .Y(exu_n15320));
INVX1 exu_U37644(.A(bypass_rs1_data_w2[20]), .Y(exu_n15321));
INVX1 exu_U37645(.A(bypass_rs1_data_w2[1]), .Y(exu_n15322));
INVX1 exu_U37646(.A(bypass_rs1_data_w2[19]), .Y(exu_n15323));
INVX1 exu_U37647(.A(bypass_rs1_data_w2[18]), .Y(exu_n15324));
INVX1 exu_U37648(.A(bypass_rs1_data_w2[17]), .Y(exu_n15325));
INVX1 exu_U37649(.A(bypass_rs1_data_w2[16]), .Y(exu_n15326));
INVX1 exu_U37650(.A(bypass_rs1_data_w2[15]), .Y(exu_n15327));
INVX1 exu_U37651(.A(bypass_rs1_data_w2[14]), .Y(exu_n15328));
INVX1 exu_U37652(.A(bypass_rs1_data_w2[13]), .Y(exu_n15329));
INVX1 exu_U37653(.A(bypass_rs1_data_w2[12]), .Y(exu_n15330));
INVX1 exu_U37654(.A(bypass_rs1_data_w2[11]), .Y(exu_n15331));
INVX1 exu_U37655(.A(bypass_rs1_data_w2[10]), .Y(exu_n15332));
INVX1 exu_U37656(.A(bypass_rs1_data_w2[0]), .Y(exu_n15333));
INVX1 exu_U37657(.A(ecl_divcntl_firstlast_sub), .Y(exu_n15334));
AND2X1 exu_U37658(.A(ifu_exu_ecc_mask[5]), .B(ecl_eccctl_inj_irferr_m), .Y(ecl_byp_ecc_mask_m_l[5]));
INVX1 exu_U37659(.A(ecl_byp_ecc_mask_m_l[5]), .Y(exu_n15335));
AND2X1 exu_U37660(.A(ifu_exu_ecc_mask[4]), .B(ecl_eccctl_inj_irferr_m), .Y(ecl_byp_ecc_mask_m_l[4]));
INVX1 exu_U37661(.A(ecl_byp_ecc_mask_m_l[4]), .Y(exu_n15336));
INVX1 exu_U37662(.A(ecl_early1_ttype_e[1]), .Y(exu_n15337));
INVX1 exu_U37663(.A(ecl_alu_xcc_e[3]), .Y(exu_n15338));
INVX1 exu_U37664(.A(ecl_alu_icc_e[3]), .Y(exu_n15339));
AND2X1 exu_U37665(.A(rml_cwp_swap_thr[3]), .B(rml_cwp_N99), .Y(rml_cwp_n40));
INVX1 exu_U37666(.A(rml_cwp_n40), .Y(exu_n15340));
AND2X1 exu_U37667(.A(rml_cwp_swap_thr[2]), .B(rml_cwp_N99), .Y(rml_cwp_n42));
INVX1 exu_U37668(.A(rml_cwp_n42), .Y(exu_n15341));
AND2X1 exu_U37669(.A(rml_cwp_swap_thr[1]), .B(rml_cwp_N99), .Y(rml_cwp_n44));
INVX1 exu_U37670(.A(rml_cwp_n44), .Y(exu_n15342));
OR2X1 exu_U37671(.A(rml_n121), .B(rml_rml_ecl_cansave_e[0]), .Y(rml_n114));
INVX1 exu_U37672(.A(rml_n114), .Y(exu_n15343));
INVX1 exu_U37673(.A(rml_n79), .Y(exu_n15344));
INVX1 exu_U37674(.A(ecl_byplog_rs1_n29), .Y(exu_n15345));
AND2X1 exu_U37675(.A(rml_n50), .B(rml_n51), .Y(rml_swap_e));
INVX1 exu_U37676(.A(rml_swap_e), .Y(exu_n15346));
AND2X1 exu_U37677(.A(ecl_divcntl_n79), .B(ecl_divcntl_gencc_in_31_d1), .Y(ecl_divcntl_n60));
INVX1 exu_U37678(.A(ecl_divcntl_n60), .Y(exu_n15347));
OR2X1 exu_U37679(.A(ecl_writeback_sraddr_e[3]), .B(ecl_writeback_sraddr_e[1]), .Y(ecl_read_yreg_e));
INVX1 exu_U37680(.A(ecl_read_yreg_e), .Y(exu_n15348));
INVX1 exu_U37681(.A(exu_ifu_spill_e), .Y(exu_n15349));
INVX1 exu_U37682(.A(exu_n15351), .Y(exu_n15350));
AND2X1 exu_U37683(.A(ecl_n105), .B(ecl_shiftop_e_0), .Y(ecl_shft_extend32bit_e_l));
INVX1 exu_U37684(.A(ecl_shft_extend32bit_e_l), .Y(exu_n15351));
INVX1 exu_U37685(.A(div_ecl_gencc_in_31), .Y(exu_n15352));
AND2X1 exu_U37686(.A(ecc_ecl_rs3_ue), .B(exu_n16394), .Y(ecl_eccctl_n14));
INVX1 exu_U37687(.A(ecl_eccctl_n14), .Y(exu_n15353));
AND2X1 exu_U37688(.A(ifu_tlu_sraddr_d[0]), .B(ifu_tlu_sraddr_d[1]), .Y(ecl_writeback_n72));
INVX1 exu_U37689(.A(ecl_writeback_n72), .Y(exu_n15354));
AND2X1 exu_U37690(.A(exu_n16571), .B(exu_n16570), .Y(rml_n77));
INVX1 exu_U37691(.A(rml_n77), .Y(exu_n15355));
INVX1 exu_U37692(.A(ecl_writeback_n44), .Y(exu_n15356));
AND2X1 exu_U37693(.A(exu_n19203), .B(exu_n19199), .Y(exu_n19201));
INVX1 exu_U37694(.A(exu_n19201), .Y(exu_n15357));
AND2X1 exu_U37695(.A(exu_n19239), .B(exu_n19235), .Y(exu_n19237));
INVX1 exu_U37696(.A(exu_n19237), .Y(exu_n15358));
AND2X1 exu_U37697(.A(ecl_byplog_rs2_n33), .B(ecl_byplog_rs2_n29), .Y(ecl_byplog_rs2_n31));
INVX1 exu_U37698(.A(ecl_byplog_rs2_n31), .Y(exu_n15359));
INVX1 exu_U37699(.A(rml_n103), .Y(exu_n15360));
AND2X1 exu_U37700(.A(ecl_writeback_n144), .B(ecl_writeback_sraddr_w[5]), .Y(ecl_writeback_n141));
INVX1 exu_U37701(.A(ecl_writeback_n141), .Y(exu_n15361));
AND2X1 exu_U37702(.A(exu_n16392), .B(rml_ecl_fill_e), .Y(ecl_n47));
INVX1 exu_U37703(.A(ecl_n47), .Y(exu_n15362));
AND2X1 exu_U37704(.A(ecl_mdqctl_div_data[11]), .B(ecl_mdqctl_n51), .Y(ecl_mdqctl_divcntl_reset_div));
INVX1 exu_U37705(.A(ecl_mdqctl_divcntl_reset_div), .Y(exu_n15363));
AND2X1 exu_U37706(.A(exu_n15457), .B(ecl_mdqctl_wb_multhr_g[1]), .Y(ecl_writeback_n185));
INVX1 exu_U37707(.A(ecl_writeback_n185), .Y(exu_n15364));
INVX1 exu_U37708(.A(rml_cwp_cwp_output_queue_n22), .Y(exu_n15365));
INVX1 exu_U37709(.A(ecl_divcntl_cnt6_n20), .Y(exu_n15366));
AND2X1 exu_U37710(.A(exu_n15378), .B(ecl_divcntl_cnt6_n31), .Y(ecl_divcntl_cnt6_n26));
INVX1 exu_U37711(.A(ecl_divcntl_cnt6_n26), .Y(exu_n15367));
AND2X1 exu_U37712(.A(rml_cwp_n91), .B(rml_cwp_wen_w), .Y(rml_cwp_n80));
INVX1 exu_U37713(.A(rml_cwp_n80), .Y(exu_n15368));
AND2X1 exu_U37714(.A(rml_cwp_n92), .B(rml_cwp_wen_w), .Y(rml_cwp_n83));
INVX1 exu_U37715(.A(rml_cwp_n83), .Y(exu_n15369));
AND2X1 exu_U37716(.A(rml_cwp_n93), .B(rml_cwp_wen_w), .Y(rml_cwp_n86));
INVX1 exu_U37717(.A(rml_cwp_n86), .Y(exu_n15370));
AND2X1 exu_U37718(.A(rml_cwp_n94), .B(rml_cwp_wen_w), .Y(rml_cwp_n89));
INVX1 exu_U37719(.A(rml_cwp_n89), .Y(exu_n15371));
AND2X1 exu_U37720(.A(ecl_divcntl_n52), .B(ecl_divcntl_n53), .Y(ecl_divcntl_n23));
INVX1 exu_U37721(.A(ecl_divcntl_n23), .Y(exu_n15372));
INVX1 exu_U37722(.A(ecl_eccctl_n21), .Y(exu_n15373));
INVX1 exu_U37723(.A(ecl_writeback_n191), .Y(exu_n15374));
INVX1 exu_U37724(.A(exu_n15376), .Y(exu_n15375));
INVX1 exu_U37725(.A(exu_n19200), .Y(exu_n15376));
INVX1 exu_U37726(.A(exu_n19236), .Y(exu_n15377));
INVX1 exu_U37727(.A(ecl_divcntl_cnt6_n30), .Y(exu_n15378));
AND2X1 exu_U37728(.A(exu_n16621), .B(ecl_divcntl_div_state_1), .Y(ecl_divcntl_cnt6_n30));
AND2X1 exu_U37729(.A(ecl_mdqctl_n20), .B(ecl_mdqctl_ismul_e), .Y(ecl_mdqctl_n16));
INVX1 exu_U37730(.A(ecl_mdqctl_n16), .Y(exu_n15379));
INVX1 exu_U37731(.A(ecl_byplog_rs2_n14), .Y(exu_n15380));
INVX1 exu_U37732(.A(ecl_byplog_rs2_n30), .Y(exu_n15381));
INVX1 exu_U37733(.A(ecl_writeback_n129), .Y(exu_n15382));
AND2X1 exu_U37734(.A(exu_n16606), .B(exu_n16604), .Y(rml_n51));
INVX1 exu_U37735(.A(rml_n51), .Y(exu_n15383));
AND2X1 exu_U37736(.A(rml_cwp_swap_state[1]), .B(rml_cwp_N99), .Y(rml_cwp_n96));
INVX1 exu_U37737(.A(rml_cwp_n96), .Y(exu_n15384));
INVX1 exu_U37738(.A(exu_n19199), .Y(exu_n15385));
INVX1 exu_U37739(.A(exu_n19235), .Y(exu_n15386));
INVX1 exu_U37740(.A(ecl_divcntl_cnt6_n23), .Y(exu_n15387));
INVX1 exu_U37741(.A(ecl_divcntl_n72), .Y(exu_n15388));
INVX1 exu_U37742(.A(ecl_byplog_rs2_n29), .Y(exu_n15389));
AND2X1 exu_U37743(.A(ifu_tlu_sraddr_d[0]), .B(exu_n16375), .Y(ecl_writeback_n70));
INVX1 exu_U37744(.A(ecl_writeback_n70), .Y(exu_n15390));
BUFX2 exu_U37745(.A(rml_irf_old_lo_cwp_e[2]), .Y(exu_n15391));
BUFX2 exu_U37746(.A(rml_irf_new_lo_cwp_e[2]), .Y(exu_n15392));
INVX1 exu_U37747(.A(ecl_pick_not_aligned), .Y(exu_n15393));
INVX1 exu_U37748(.A(ecl_divcntl_n61), .Y(exu_n15394));
INVX1 exu_U37749(.A(ecl_writeback_n149), .Y(exu_n15395));
INVX1 exu_U37750(.A(ecc_err_m[5]), .Y(exu_n15396));
OR2X1 exu_U37751(.A(exu_n15965), .B(exu_n15462), .Y(ecl_byp_rs3_longmux_sel_g2));
OR2X1 exu_U37752(.A(exu_n19227), .B(exu_n15463), .Y(ecl_byp_rs3h_longmux_sel_g2));
OR2X1 exu_U37753(.A(ecl_mdqctl_mul_data[9]), .B(exu_n15986), .Y(ecl_div_mul_get_32bit_data));
OR2X1 exu_U37754(.A(ecl_div_sel_64b), .B(ecl_ecl_div_signed_div), .Y(ecl_div_sel_u32));
OR2X1 exu_U37755(.A(exu_n15487), .B(ecl_divcntl_gencc_in_31_d1), .Y(ecl_div_upper33_zero));
OR2X1 exu_U37756(.A(exu_n15966), .B(exu_n15464), .Y(ecl_byp_rs2_longmux_sel_g2));
OR2X1 exu_U37757(.A(exu_n15508), .B(ecl_byplog_rs1_n21), .Y(ecl_byp_rs1_mux2_sel_ld));
OR2X1 exu_U37758(.A(exu_n15508), .B(ecl_byp_rcc_mux1_sel_w2), .Y(ecl_byp_rs1_mux1_sel_w2));
OR2X1 exu_U37759(.A(exu_n15967), .B(exu_n15465), .Y(ecl_byp_rs1_longmux_sel_g2));
AND2X1 exu_U37760(.A(ecl_byplog_rs1_n20), .B(exu_n15767), .Y(ecl_byp_rs1_mux1_sel_other));
INVX1 exu_U37761(.A(ecl_byp_rs1_mux1_sel_other), .Y(exu_n15397));
AND2X1 exu_U37762(.A(exu_n15476), .B(ecl_byplog_rs1_n19), .Y(ecl_byp_rcc_mux2_sel_rf));
OR2X1 exu_U37763(.A(ecl_byplog_rs1_n26), .B(ecl_byplog_rs1_n21), .Y(ecl_byp_rcc_mux2_sel_ld));
OR2X1 exu_U37764(.A(ecl_byplog_rs1_n17), .B(ecl_byplog_rs1_n26), .Y(ecl_byp_rcc_mux2_sel_e));
OR2X1 exu_U37765(.A(exu_n15437), .B(exu_n16300), .Y(ecl_byp_rcc_mux1_sel_w));
OR2X1 exu_U37766(.A(ecl_byplog_rs1_n32), .B(exu_n16300), .Y(ecl_byp_rcc_mux1_sel_m));
OR2X1 exu_U37767(.A(ecl_writeback_n129), .B(exu_n16271), .Y(ecl_byp_sel_muldiv_g));
INVX1 exu_U37768(.A(ecl_byp_sel_muldiv_g), .Y(exu_n15398));
OR2X1 exu_U37769(.A(exu_n15690), .B(exu_n16519), .Y(shft_shift16_e[3]));
INVX1 exu_U37770(.A(shft_shift16_e[3]), .Y(exu_n15399));
OR2X1 exu_U37771(.A(div_input_data_e[68]), .B(exu_n15690), .Y(shft_shift16_e[2]));
OR2X1 exu_U37772(.A(div_input_data_e[66]), .B(exu_n16518), .Y(ecl_shft_shift4_e[2]));
OR2X1 exu_U37773(.A(div_input_data_e[67]), .B(exu_n16517), .Y(ecl_shft_shift4_e[1]));
INVX1 exu_U37774(.A(ecl_shft_shift4_e[1]), .Y(exu_n15400));
OR2X1 exu_U37775(.A(div_input_data_e[67]), .B(div_input_data_e[66]), .Y(ecl_shft_shift4_e[0]));
INVX1 exu_U37776(.A(ecl_shft_shift4_e[0]), .Y(exu_n15401));
OR2X1 exu_U37777(.A(div_input_data_e[64]), .B(exu_n16516), .Y(ecl_shft_shift1_e[2]));
INVX1 exu_U37778(.A(ecl_shft_shift1_e[2]), .Y(exu_n15402));
OR2X1 exu_U37779(.A(div_input_data_e[65]), .B(exu_n16514), .Y(ecl_shft_shift1_e[1]));
INVX1 exu_U37780(.A(ecl_shft_extendbit_e), .Y(exu_n15403));
OR2X1 exu_U37781(.A(ecl_tid_e[0]), .B(exu_n16580), .Y(ecl_div_thr_e[2]));
OR2X1 exu_U37782(.A(ecl_tid_e[1]), .B(exu_n16579), .Y(ecl_div_thr_e[1]));
OR2X1 exu_U37783(.A(ecl_tid_e[1]), .B(ecl_tid_e[0]), .Y(ecl_div_thr_e[0]));
OR2X1 exu_U37784(.A(ecl_byp_sel_ffusr_m), .B(exu_n16582), .Y(ecl_byp_sel_tlusr_m));
OR2X1 exu_U37785(.A(ecl_read_tlusr_m), .B(ecl_byp_sel_ffusr_m), .Y(ecl_byp_sel_ifex_m));
OR2X1 exu_U37786(.A(div_input_data_e[64]), .B(div_input_data_e[65]), .Y(ecl_shft_shift1_e[0]));
OR2X1 exu_U37787(.A(exu_n16576), .B(ecl_tid_w[1]), .Y(ecl_rml_thr_w[1]));
INVX1 exu_U37788(.A(ecl_rml_thr_w[1]), .Y(exu_n15404));
OR2X1 exu_U37789(.A(ecl_tid_w[0]), .B(ecl_tid_w[1]), .Y(ecl_rml_thr_w[0]));
INVX1 exu_U37790(.A(ecl_rml_thr_w[0]), .Y(exu_n15405));
INVX1 exu_U37791(.A(exu_n31737), .Y(exu_lsu_ldst_va_e[47]));
INVX1 exu_U37792(.A(exu_n31748), .Y(exu_ifu_cc_d[0]));
INVX1 exu_U37793(.A(exu_n31745), .Y(exu_ifu_cc_d[3]));
INVX1 exu_U37794(.A(exu_n31747), .Y(exu_ifu_cc_d[1]));
AND2X1 exu_U37795(.A(exu_n15691), .B(exu_n15925), .Y(rml_cwp_n74));
INVX1 exu_U37796(.A(rml_cwp_n74), .Y(exu_n15410));
OR2X1 exu_U37797(.A(alu_regzcmp_low_nonzero), .B(alu_regzcmp_high_nonzero), .Y(exu_n31738));
INVX1 exu_U37798(.A(exu_n31738), .Y(exu_ifu_regz_e));
AND2X1 exu_U37799(.A(exu_n16604), .B(exu_n16383), .Y(rml_cansave_inc_e));
INVX1 exu_U37800(.A(rml_cansave_inc_e), .Y(exu_n15412));
AND2X1 exu_U37801(.A(exu_n16606), .B(exu_n16385), .Y(rml_canrestore_inc_e));
INVX1 exu_U37802(.A(rml_canrestore_inc_e), .Y(exu_n15413));
AND2X1 exu_U37803(.A(ecl_thr_match_dm), .B(ecl_ccr_setcc_m), .Y(ecl_ccr_n24));
INVX1 exu_U37804(.A(ecl_ccr_n24), .Y(exu_n15414));
AND2X1 exu_U37805(.A(exu_n15554), .B(exu_n15488), .Y(rml_cwp_n43));
INVX1 exu_U37806(.A(rml_cwp_n43), .Y(exu_n15415));
AND2X1 exu_U37807(.A(exu_n15555), .B(exu_n15489), .Y(rml_cwp_n41));
INVX1 exu_U37808(.A(rml_cwp_n41), .Y(exu_n15416));
AND2X1 exu_U37809(.A(exu_n15556), .B(exu_n15490), .Y(rml_cwp_n39));
INVX1 exu_U37810(.A(rml_cwp_n39), .Y(exu_n15417));
INVX1 exu_U37811(.A(bypass_rd_data_g[9]), .Y(exu_n15418));
INVX1 exu_U37812(.A(div_gencc_in[63]), .Y(exu_n15419));
OR2X1 exu_U37813(.A(ecl_byp_sel_alu_e), .B(ifu_exu_rd_ifusr_e), .Y(ecl_n46));
INVX1 exu_U37814(.A(ecl_n46), .Y(exu_n15420));
INVX1 exu_U37815(.A(exu_n19197), .Y(exu_n15421));
INVX1 exu_U37816(.A(exu_n19233), .Y(exu_n15422));
INVX1 exu_U37817(.A(ecl_byplog_rs2_n26), .Y(exu_n15423));
AND2X1 exu_U37818(.A(ecl_divcntl_n85), .B(exu_n15471), .Y(ecl_divcntl_n56));
INVX1 exu_U37819(.A(ecl_divcntl_n56), .Y(exu_n15424));
AND2X1 exu_U37820(.A(ecl_mdqctl_ismul_w), .B(exu_n16390), .Y(ecl_mdqctl_n21));
INVX1 exu_U37821(.A(ecl_mdqctl_n21), .Y(exu_n15425));
INVX1 exu_U37822(.A(alu_ecl_zlow_e), .Y(exu_n15426));
INVX1 exu_U37823(.A(ecl_writeback_sel_cwp_d), .Y(exu_n15427));
INVX1 exu_U37824(.A(rml_cwp_cwp_wen_tlu_w[3]), .Y(exu_n15428));
INVX1 exu_U37825(.A(rml_cwp_cwp_wen_tlu_w[2]), .Y(exu_n15429));
INVX1 exu_U37826(.A(rml_cwp_cwp_wen_tlu_w[1]), .Y(exu_n15430));
INVX1 exu_U37827(.A(rml_cwp_cwp_wen_tlu_w[0]), .Y(exu_n15431));
OR2X1 exu_U37828(.A(ifu_tlu_sraddr_d[1]), .B(ifu_tlu_sraddr_d[0]), .Y(ecl_writeback_sel_cleanwin_d));
INVX1 exu_U37829(.A(ecl_writeback_sel_cleanwin_d), .Y(exu_n15432));
AND2X1 exu_U37830(.A(exu_n19207), .B(ecl_byplog_rs3_match_w), .Y(exu_n19196));
INVX1 exu_U37831(.A(exu_n19196), .Y(exu_n15433));
AND2X1 exu_U37832(.A(exu_n19243), .B(ecl_byplog_rs3h_match_w), .Y(exu_n19232));
INVX1 exu_U37833(.A(exu_n19232), .Y(exu_n15434));
AND2X1 exu_U37834(.A(ecl_byplog_rs2_n37), .B(ecl_byplog_rs2_match_w), .Y(ecl_byplog_rs2_n25));
INVX1 exu_U37835(.A(ecl_byplog_rs2_n25), .Y(exu_n15435));
INVX1 exu_U37836(.A(ecl_n68), .Y(exu_n15436));
AND2X1 exu_U37837(.A(ecl_byplog_rs1_n42), .B(ecl_byplog_rs1_match_w), .Y(ecl_byplog_rs1_n31));
INVX1 exu_U37838(.A(ecl_byplog_rs1_n31), .Y(exu_n15437));
INVX1 exu_U37839(.A(shft_rshifterinput_b1[41]), .Y(exu_n15438));
OR2X1 exu_U37840(.A(rml_n35), .B(tlu_exu_agp_tid[1]), .Y(rml_agp_thr[1]));
INVX1 exu_U37841(.A(rml_agp_thr[1]), .Y(exu_n15439));
OR2X1 exu_U37842(.A(tlu_exu_agp_tid[0]), .B(tlu_exu_agp_tid[1]), .Y(rml_agp_thr[0]));
INVX1 exu_U37843(.A(rml_agp_thr[0]), .Y(exu_n15440));
INVX1 exu_U37844(.A(ecc_err_m[2]), .Y(exu_n15441));
INVX1 exu_U37845(.A(shft_rshifterinput_b1[40]), .Y(exu_n15442));
INVX1 exu_U37846(.A(shft_rshifterinput_b1[39]), .Y(exu_n15443));
INVX1 exu_U37847(.A(shft_rshifterinput_b1[38]), .Y(exu_n15444));
INVX1 exu_U37848(.A(shft_rshifterinput_b1[37]), .Y(exu_n15445));
INVX1 exu_U37849(.A(shft_rshifterinput_b1[36]), .Y(exu_n15446));
INVX1 exu_U37850(.A(shft_rshifterinput_b1[35]), .Y(exu_n15447));
INVX1 exu_U37851(.A(shft_rshifterinput_b1[34]), .Y(exu_n15448));
INVX1 exu_U37852(.A(shft_rshifterinput_b1[33]), .Y(exu_n15449));
INVX1 exu_U37853(.A(shft_rshifterinput_b1[47]), .Y(exu_n15450));
INVX1 exu_U37854(.A(shft_rshifterinput_b1[46]), .Y(exu_n15451));
INVX1 exu_U37855(.A(shft_rshifterinput_b1[45]), .Y(exu_n15452));
INVX1 exu_U37856(.A(shft_rshifterinput_b1[44]), .Y(exu_n15453));
INVX1 exu_U37857(.A(shft_rshifterinput_b1[43]), .Y(exu_n15454));
INVX1 exu_U37858(.A(shft_rshifterinput_b1[42]), .Y(exu_n15455));
INVX1 exu_U37859(.A(shft_rshifterinput_b1[32]), .Y(exu_n15456));
OR2X1 exu_U37860(.A(ecl_mdqctl_mul_data[9]), .B(exu_n16186), .Y(ecl_mdqctl_wb_yreg_wen_g));
INVX1 exu_U37861(.A(ecl_mdqctl_wb_yreg_wen_g), .Y(exu_n15457));
BUFX2 exu_U37862(.A(ecl_ecl_reset_l), .Y(exu_n15458));
INVX1 exu_U37863(.A(ecc_err_m[4]), .Y(exu_n15459));
INVX1 exu_U37864(.A(ecc_err_m[3]), .Y(exu_n15460));
INVX1 exu_U37865(.A(ecc_err_m[1]), .Y(exu_n15461));
AND2X1 exu_U37866(.A(exu_n19211), .B(ecl_wb_byplog_wen_g2), .Y(exu_n19204));
INVX1 exu_U37867(.A(exu_n19204), .Y(exu_n15462));
AND2X1 exu_U37868(.A(exu_n19247), .B(ecl_wb_byplog_wen_g2), .Y(exu_n19240));
INVX1 exu_U37869(.A(exu_n19240), .Y(exu_n15463));
AND2X1 exu_U37870(.A(ecl_byplog_rs2_n41), .B(ecl_wb_byplog_wen_g2), .Y(ecl_byplog_rs2_n34));
INVX1 exu_U37871(.A(ecl_byplog_rs2_n34), .Y(exu_n15464));
AND2X1 exu_U37872(.A(ecl_byplog_rs1_n45), .B(ecl_wb_byplog_wen_g2), .Y(ecl_byplog_rs1_n23));
INVX1 exu_U37873(.A(ecl_byplog_rs1_n23), .Y(exu_n15465));
AND2X1 exu_U37874(.A(ecl_ccr_n28), .B(ecl_ccr_thr_w2[1]), .Y(ecl_ccr_n12));
INVX1 exu_U37875(.A(ecl_ccr_n12), .Y(exu_n15466));
INVX1 exu_U37876(.A(ecl_ccr_n15), .Y(exu_n15467));
INVX1 exu_U37877(.A(ecl_ccr_n17), .Y(exu_n15468));
INVX1 exu_U37878(.A(ecl_ccr_n19), .Y(exu_n15469));
OR2X1 exu_U37879(.A(exu_n16571), .B(rml_tid_e[0]), .Y(rml_n66));
INVX1 exu_U37880(.A(rml_n66), .Y(exu_n15470));
INVX1 exu_U37881(.A(ecl_divcntl_n30), .Y(exu_n15471));
AND2X1 exu_U37882(.A(rml_cwp_spill_next), .B(rml_cwp_swap_thr[3]), .Y(rml_cwp_n79));
INVX1 exu_U37883(.A(rml_cwp_n79), .Y(exu_n15472));
AND2X1 exu_U37884(.A(rml_cwp_spill_next), .B(rml_cwp_swap_thr[2]), .Y(rml_cwp_n82));
INVX1 exu_U37885(.A(rml_cwp_n82), .Y(exu_n15473));
AND2X1 exu_U37886(.A(rml_cwp_spill_next), .B(rml_cwp_swap_thr[1]), .Y(rml_cwp_n85));
INVX1 exu_U37887(.A(rml_cwp_n85), .Y(exu_n15474));
AND2X1 exu_U37888(.A(rml_cwp_spill_next), .B(rml_cwp_swap_thr[0]), .Y(rml_cwp_n88));
INVX1 exu_U37889(.A(rml_cwp_n88), .Y(exu_n15475));
AND2X1 exu_U37890(.A(ecl_byplog_rs1_n46), .B(ecl_ld_thr_match_dg), .Y(ecl_byplog_rs1_n22));
INVX1 exu_U37891(.A(ecl_byplog_rs1_n26), .Y(exu_n15476));
INVX1 exu_U37892(.A(ecl_writeback_n198), .Y(exu_n15477));
INVX1 exu_U37893(.A(alu_va_e[57]), .Y(exu_n15478));
INVX1 exu_U37894(.A(alu_va_e[48]), .Y(exu_n15479));
INVX1 exu_U37895(.A(ecc_err_m[6]), .Y(exu_n15480));
INVX1 exu_U37896(.A(ecl_eccctl_n25), .Y(exu_n15481));
INVX1 exu_U37897(.A(ecl_writeback_n50), .Y(exu_n15482));
INVX1 exu_U37898(.A(rml_agp_wen_thr3_w), .Y(exu_n15483));
INVX1 exu_U37899(.A(rml_agp_wen_thr2_w), .Y(exu_n15484));
INVX1 exu_U37900(.A(rml_agp_wen_thr1_w), .Y(exu_n15485));
INVX1 exu_U37901(.A(rml_agp_wen_thr0_w), .Y(exu_n15486));
AND2X1 exu_U37902(.A(ecl_divcntl_upper32_equal_d1), .B(ecl_divcntl_gencc_in_msb_l_d1), .Y(ecl_divcntl_n70));
INVX1 exu_U37903(.A(ecl_divcntl_n70), .Y(exu_n15487));
AND2X1 exu_U37904(.A(rml_cwp_n75), .B(exu_n15958), .Y(rml_cwp_n34));
INVX1 exu_U37905(.A(rml_cwp_n34), .Y(exu_n15488));
AND2X1 exu_U37906(.A(rml_cwp_n76), .B(ecl_rml_thr_w[2]), .Y(rml_cwp_n33));
INVX1 exu_U37907(.A(rml_cwp_n33), .Y(exu_n15489));
AND2X1 exu_U37908(.A(rml_cwp_n77), .B(ecl_rml_thr_w[3]), .Y(rml_cwp_n32));
INVX1 exu_U37909(.A(rml_cwp_n32), .Y(exu_n15490));
INVX1 exu_U37910(.A(div_ecl_cout64), .Y(exu_n15491));
INVX1 exu_U37911(.A(div_xin[63]), .Y(exu_n15492));
INVX1 exu_U37912(.A(ecl_n112), .Y(exu_n15493));
INVX1 exu_U37913(.A(alu_va_e[62]), .Y(exu_n15494));
INVX1 exu_U37914(.A(alu_va_e[61]), .Y(exu_n15495));
INVX1 exu_U37915(.A(alu_va_e[60]), .Y(exu_n15496));
INVX1 exu_U37916(.A(alu_va_e[59]), .Y(exu_n15497));
INVX1 exu_U37917(.A(alu_va_e[58]), .Y(exu_n15498));
INVX1 exu_U37918(.A(alu_va_e[55]), .Y(exu_n15499));
INVX1 exu_U37919(.A(alu_va_e[54]), .Y(exu_n15500));
INVX1 exu_U37920(.A(alu_va_e[53]), .Y(exu_n15501));
INVX1 exu_U37921(.A(alu_va_e[52]), .Y(exu_n15502));
INVX1 exu_U37922(.A(alu_va_e[51]), .Y(exu_n15503));
INVX1 exu_U37923(.A(alu_va_e[50]), .Y(exu_n15504));
INVX1 exu_U37924(.A(alu_va_e[49]), .Y(exu_n15505));
INVX1 exu_U37925(.A(ecc_decode_n20), .Y(exu_n15506));
AND2X1 exu_U37926(.A(ecc_decode_n43), .B(ecc_decode_n24), .Y(ecc_decode_n42));
INVX1 exu_U37927(.A(ecc_decode_n42), .Y(exu_n15507));
INVX1 exu_U37928(.A(ecl_byplog_rs1_n20), .Y(exu_n15508));
INVX1 exu_U37929(.A(ecc_decode_n21), .Y(exu_n15509));
INVX1 exu_U37930(.A(ecc_decode_n18), .Y(exu_n15510));
INVX1 exu_U37931(.A(ecc_decode_n22), .Y(exu_n15511));
INVX1 exu_U37932(.A(div_gencc_in[41]), .Y(exu_n15512));
AND2X1 exu_U37933(.A(ifu_exu_ecc_mask[7]), .B(ecl_eccctl_inj_irferr_m), .Y(ecl_byp_ecc_mask_m_l[7]));
INVX1 exu_U37934(.A(ecl_byp_ecc_mask_m_l[7]), .Y(exu_n15513));
AND2X1 exu_U37935(.A(ifu_exu_ecc_mask[6]), .B(ecl_eccctl_inj_irferr_m), .Y(ecl_byp_ecc_mask_m_l[6]));
INVX1 exu_U37936(.A(ecl_byp_ecc_mask_m_l[6]), .Y(exu_n15514));
AND2X1 exu_U37937(.A(ifu_exu_ecc_mask[3]), .B(ecl_eccctl_inj_irferr_m), .Y(ecl_byp_ecc_mask_m_l[3]));
INVX1 exu_U37938(.A(ecl_byp_ecc_mask_m_l[3]), .Y(exu_n15515));
INVX1 exu_U37939(.A(ecc_decode_n24), .Y(exu_n15516));
AND2X1 exu_U37940(.A(ecc_err_m[1]), .B(ecc_err_m[2]), .Y(ecc_decode_n24));
INVX1 exu_U37941(.A(div_gencc_in[62]), .Y(exu_n15517));
INVX1 exu_U37942(.A(div_gencc_in[61]), .Y(exu_n15518));
INVX1 exu_U37943(.A(div_gencc_in[60]), .Y(exu_n15519));
INVX1 exu_U37944(.A(div_gencc_in[59]), .Y(exu_n15520));
INVX1 exu_U37945(.A(div_gencc_in[58]), .Y(exu_n15521));
INVX1 exu_U37946(.A(div_gencc_in[57]), .Y(exu_n15522));
INVX1 exu_U37947(.A(div_gencc_in[56]), .Y(exu_n15523));
INVX1 exu_U37948(.A(div_gencc_in[55]), .Y(exu_n15524));
INVX1 exu_U37949(.A(div_gencc_in[54]), .Y(exu_n15525));
INVX1 exu_U37950(.A(div_gencc_in[53]), .Y(exu_n15526));
INVX1 exu_U37951(.A(div_gencc_in[52]), .Y(exu_n15527));
INVX1 exu_U37952(.A(div_gencc_in[51]), .Y(exu_n15528));
INVX1 exu_U37953(.A(div_gencc_in[50]), .Y(exu_n15529));
INVX1 exu_U37954(.A(div_gencc_in[49]), .Y(exu_n15530));
INVX1 exu_U37955(.A(div_gencc_in[48]), .Y(exu_n15531));
INVX1 exu_U37956(.A(div_gencc_in[47]), .Y(exu_n15532));
INVX1 exu_U37957(.A(div_gencc_in[46]), .Y(exu_n15533));
INVX1 exu_U37958(.A(div_gencc_in[45]), .Y(exu_n15534));
INVX1 exu_U37959(.A(div_gencc_in[44]), .Y(exu_n15535));
INVX1 exu_U37960(.A(div_gencc_in[43]), .Y(exu_n15536));
INVX1 exu_U37961(.A(div_gencc_in[40]), .Y(exu_n15537));
INVX1 exu_U37962(.A(div_gencc_in[39]), .Y(exu_n15538));
INVX1 exu_U37963(.A(div_gencc_in[38]), .Y(exu_n15539));
INVX1 exu_U37964(.A(div_gencc_in[37]), .Y(exu_n15540));
INVX1 exu_U37965(.A(div_gencc_in[36]), .Y(exu_n15541));
INVX1 exu_U37966(.A(div_gencc_in[35]), .Y(exu_n15542));
INVX1 exu_U37967(.A(div_gencc_in[34]), .Y(exu_n15543));
INVX1 exu_U37968(.A(div_gencc_in[33]), .Y(exu_n15544));
INVX1 exu_U37969(.A(ecl_writeback_n110), .Y(exu_n15545));
INVX1 exu_U37970(.A(alu_va_e[56]), .Y(exu_n15546));
BUFX2 exu_U37971(.A(rml_irf_old_lo_cwp_e[1]), .Y(exu_n15547));
BUFX2 exu_U37972(.A(rml_irf_new_lo_cwp_e[1]), .Y(exu_n15548));
INVX1 exu_U37973(.A(div_gencc_in[42]), .Y(exu_n15549));
AND2X1 exu_U37974(.A(ifu_exu_ecc_mask[2]), .B(ecl_eccctl_inj_irferr_m), .Y(ecl_byp_ecc_mask_m_l[2]));
INVX1 exu_U37975(.A(ecl_byp_ecc_mask_m_l[2]), .Y(exu_n15550));
AND2X1 exu_U37976(.A(ifu_exu_ecc_mask[1]), .B(ecl_eccctl_inj_irferr_m), .Y(ecl_byp_ecc_mask_m_l[1]));
INVX1 exu_U37977(.A(ecl_byp_ecc_mask_m_l[1]), .Y(exu_n15551));
AND2X1 exu_U37978(.A(ifu_exu_ecc_mask[0]), .B(ecl_eccctl_inj_irferr_m), .Y(ecl_byp_ecc_mask_m_l[0]));
INVX1 exu_U37979(.A(ecl_byp_ecc_mask_m_l[0]), .Y(exu_n15552));
BUFX2 exu_U37980(.A(rml_irf_new_lo_cwp_e[0]), .Y(exu_n15553));
AND2X1 exu_U37981(.A(exu_n9), .B(exu_n15925), .Y(rml_cwp_n37));
INVX1 exu_U37982(.A(rml_cwp_n37), .Y(exu_n15554));
AND2X1 exu_U37983(.A(rml_cwp_thr_e[2]), .B(exu_n15925), .Y(rml_cwp_n36));
INVX1 exu_U37984(.A(rml_cwp_n36), .Y(exu_n15555));
AND2X1 exu_U37985(.A(exu_n15925), .B(rml_cwp_thr_e[3]), .Y(rml_cwp_n35));
INVX1 exu_U37986(.A(rml_cwp_n35), .Y(exu_n15556));
INVX1 exu_U37987(.A(ecl_bypass_w), .Y(exu_n15557));
INVX1 exu_U37988(.A(div_ecl_cout32), .Y(exu_n15558));
INVX1 exu_U37989(.A(exu_n16817), .Y(exu_n15559));
INVX1 exu_U37990(.A(exu_n16869), .Y(exu_n15560));
INVX1 exu_U37991(.A(exu_n16885), .Y(exu_n15561));
INVX1 exu_U37992(.A(exu_n16887), .Y(exu_n15562));
INVX1 exu_U37993(.A(exu_n16889), .Y(exu_n15563));
INVX1 exu_U37994(.A(exu_n16891), .Y(exu_n15564));
INVX1 exu_U37995(.A(exu_n16893), .Y(exu_n15565));
INVX1 exu_U37996(.A(exu_n16895), .Y(exu_n15566));
INVX1 exu_U37997(.A(exu_n16897), .Y(exu_n15567));
INVX1 exu_U37998(.A(exu_n16976), .Y(exu_n15568));
INVX1 exu_U37999(.A(exu_n17028), .Y(exu_n15569));
INVX1 exu_U38000(.A(exu_n17044), .Y(exu_n15570));
INVX1 exu_U38001(.A(exu_n17046), .Y(exu_n15571));
INVX1 exu_U38002(.A(exu_n17048), .Y(exu_n15572));
INVX1 exu_U38003(.A(exu_n17050), .Y(exu_n15573));
INVX1 exu_U38004(.A(exu_n17052), .Y(exu_n15574));
INVX1 exu_U38005(.A(exu_n17054), .Y(exu_n15575));
INVX1 exu_U38006(.A(exu_n17056), .Y(exu_n15576));
INVX1 exu_U38007(.A(exu_n17135), .Y(exu_n15577));
INVX1 exu_U38008(.A(exu_n17187), .Y(exu_n15578));
INVX1 exu_U38009(.A(exu_n17203), .Y(exu_n15579));
INVX1 exu_U38010(.A(exu_n17205), .Y(exu_n15580));
INVX1 exu_U38011(.A(exu_n17207), .Y(exu_n15581));
INVX1 exu_U38012(.A(exu_n17209), .Y(exu_n15582));
INVX1 exu_U38013(.A(exu_n17211), .Y(exu_n15583));
INVX1 exu_U38014(.A(exu_n17213), .Y(exu_n15584));
INVX1 exu_U38015(.A(exu_n17215), .Y(exu_n15585));
INVX1 exu_U38016(.A(exu_n17294), .Y(exu_n15586));
INVX1 exu_U38017(.A(exu_n17346), .Y(exu_n15587));
INVX1 exu_U38018(.A(exu_n17362), .Y(exu_n15588));
INVX1 exu_U38019(.A(exu_n17364), .Y(exu_n15589));
INVX1 exu_U38020(.A(exu_n17366), .Y(exu_n15590));
INVX1 exu_U38021(.A(exu_n17368), .Y(exu_n15591));
INVX1 exu_U38022(.A(exu_n17370), .Y(exu_n15592));
INVX1 exu_U38023(.A(exu_n17372), .Y(exu_n15593));
INVX1 exu_U38024(.A(exu_n17374), .Y(exu_n15594));
INVX1 exu_U38025(.A(exu_n16771), .Y(exu_n15595));
INVX1 exu_U38026(.A(exu_n16776), .Y(exu_n15596));
INVX1 exu_U38027(.A(exu_n16781), .Y(exu_n15597));
INVX1 exu_U38028(.A(exu_n16786), .Y(exu_n15598));
INVX1 exu_U38029(.A(exu_n16791), .Y(exu_n15599));
INVX1 exu_U38030(.A(exu_n16796), .Y(exu_n15600));
INVX1 exu_U38031(.A(exu_n16801), .Y(exu_n15601));
INVX1 exu_U38032(.A(exu_n16806), .Y(exu_n15602));
INVX1 exu_U38033(.A(exu_n16811), .Y(exu_n15603));
INVX1 exu_U38034(.A(exu_n16818), .Y(exu_n15604));
INVX1 exu_U38035(.A(exu_n16823), .Y(exu_n15605));
INVX1 exu_U38036(.A(exu_n16828), .Y(exu_n15606));
INVX1 exu_U38037(.A(exu_n16833), .Y(exu_n15607));
INVX1 exu_U38038(.A(exu_n16838), .Y(exu_n15608));
INVX1 exu_U38039(.A(exu_n16843), .Y(exu_n15609));
INVX1 exu_U38040(.A(exu_n16848), .Y(exu_n15610));
INVX1 exu_U38041(.A(exu_n16853), .Y(exu_n15611));
INVX1 exu_U38042(.A(exu_n16858), .Y(exu_n15612));
INVX1 exu_U38043(.A(exu_n16863), .Y(exu_n15613));
INVX1 exu_U38044(.A(exu_n16870), .Y(exu_n15614));
INVX1 exu_U38045(.A(exu_n16875), .Y(exu_n15615));
INVX1 exu_U38046(.A(exu_n16880), .Y(exu_n15616));
INVX1 exu_U38047(.A(exu_n16930), .Y(exu_n15617));
INVX1 exu_U38048(.A(exu_n16935), .Y(exu_n15618));
INVX1 exu_U38049(.A(exu_n16940), .Y(exu_n15619));
INVX1 exu_U38050(.A(exu_n16945), .Y(exu_n15620));
INVX1 exu_U38051(.A(exu_n16950), .Y(exu_n15621));
INVX1 exu_U38052(.A(exu_n16955), .Y(exu_n15622));
INVX1 exu_U38053(.A(exu_n16960), .Y(exu_n15623));
INVX1 exu_U38054(.A(exu_n16965), .Y(exu_n15624));
INVX1 exu_U38055(.A(exu_n16970), .Y(exu_n15625));
INVX1 exu_U38056(.A(exu_n16977), .Y(exu_n15626));
INVX1 exu_U38057(.A(exu_n16982), .Y(exu_n15627));
INVX1 exu_U38058(.A(exu_n16987), .Y(exu_n15628));
INVX1 exu_U38059(.A(exu_n16992), .Y(exu_n15629));
INVX1 exu_U38060(.A(exu_n16997), .Y(exu_n15630));
INVX1 exu_U38061(.A(exu_n17002), .Y(exu_n15631));
INVX1 exu_U38062(.A(exu_n17007), .Y(exu_n15632));
INVX1 exu_U38063(.A(exu_n17012), .Y(exu_n15633));
INVX1 exu_U38064(.A(exu_n17017), .Y(exu_n15634));
INVX1 exu_U38065(.A(exu_n17022), .Y(exu_n15635));
INVX1 exu_U38066(.A(exu_n17029), .Y(exu_n15636));
INVX1 exu_U38067(.A(exu_n17034), .Y(exu_n15637));
INVX1 exu_U38068(.A(exu_n17039), .Y(exu_n15638));
INVX1 exu_U38069(.A(exu_n17089), .Y(exu_n15639));
INVX1 exu_U38070(.A(exu_n17094), .Y(exu_n15640));
INVX1 exu_U38071(.A(exu_n17099), .Y(exu_n15641));
INVX1 exu_U38072(.A(exu_n17104), .Y(exu_n15642));
INVX1 exu_U38073(.A(exu_n17109), .Y(exu_n15643));
INVX1 exu_U38074(.A(exu_n17114), .Y(exu_n15644));
INVX1 exu_U38075(.A(exu_n17119), .Y(exu_n15645));
INVX1 exu_U38076(.A(exu_n17124), .Y(exu_n15646));
INVX1 exu_U38077(.A(exu_n17129), .Y(exu_n15647));
INVX1 exu_U38078(.A(exu_n17136), .Y(exu_n15648));
INVX1 exu_U38079(.A(exu_n17141), .Y(exu_n15649));
INVX1 exu_U38080(.A(exu_n17146), .Y(exu_n15650));
INVX1 exu_U38081(.A(exu_n17151), .Y(exu_n15651));
INVX1 exu_U38082(.A(exu_n17156), .Y(exu_n15652));
INVX1 exu_U38083(.A(exu_n17161), .Y(exu_n15653));
INVX1 exu_U38084(.A(exu_n17166), .Y(exu_n15654));
INVX1 exu_U38085(.A(exu_n17171), .Y(exu_n15655));
INVX1 exu_U38086(.A(exu_n17176), .Y(exu_n15656));
INVX1 exu_U38087(.A(exu_n17181), .Y(exu_n15657));
INVX1 exu_U38088(.A(exu_n17188), .Y(exu_n15658));
INVX1 exu_U38089(.A(exu_n17193), .Y(exu_n15659));
INVX1 exu_U38090(.A(exu_n17198), .Y(exu_n15660));
INVX1 exu_U38091(.A(exu_n17248), .Y(exu_n15661));
INVX1 exu_U38092(.A(exu_n17253), .Y(exu_n15662));
INVX1 exu_U38093(.A(exu_n17258), .Y(exu_n15663));
INVX1 exu_U38094(.A(exu_n17263), .Y(exu_n15664));
INVX1 exu_U38095(.A(exu_n17268), .Y(exu_n15665));
INVX1 exu_U38096(.A(exu_n17273), .Y(exu_n15666));
INVX1 exu_U38097(.A(exu_n17278), .Y(exu_n15667));
INVX1 exu_U38098(.A(exu_n17283), .Y(exu_n15668));
INVX1 exu_U38099(.A(exu_n17288), .Y(exu_n15669));
INVX1 exu_U38100(.A(exu_n17295), .Y(exu_n15670));
INVX1 exu_U38101(.A(exu_n17300), .Y(exu_n15671));
INVX1 exu_U38102(.A(exu_n17305), .Y(exu_n15672));
INVX1 exu_U38103(.A(exu_n17310), .Y(exu_n15673));
INVX1 exu_U38104(.A(exu_n17315), .Y(exu_n15674));
INVX1 exu_U38105(.A(exu_n17320), .Y(exu_n15675));
INVX1 exu_U38106(.A(exu_n17325), .Y(exu_n15676));
INVX1 exu_U38107(.A(exu_n17330), .Y(exu_n15677));
INVX1 exu_U38108(.A(exu_n17335), .Y(exu_n15678));
INVX1 exu_U38109(.A(exu_n17340), .Y(exu_n15679));
INVX1 exu_U38110(.A(exu_n17347), .Y(exu_n15680));
INVX1 exu_U38111(.A(exu_n17352), .Y(exu_n15681));
INVX1 exu_U38112(.A(exu_n17357), .Y(exu_n15682));
AND2X1 exu_U38113(.A(rml_rml_ecl_cwp_e[0]), .B(rml_rml_ecl_cansave_e[0]), .Y(rml_n41));
INVX1 exu_U38114(.A(rml_n41), .Y(exu_n15683));
INVX1 exu_U38115(.A(ecl_divcntl_n69), .Y(exu_n15684));
INVX1 exu_U38116(.A(rml_n52), .Y(exu_n15685));
INVX1 exu_U38117(.A(ecl_ccr_exu_ifu_cc_w[7]), .Y(exu_n15686));
OR2X1 exu_U38118(.A(exu_n16596), .B(ecl_ecl_exu_kill_m), .Y(ecl_writeback_n102));
INVX1 exu_U38119(.A(ecl_writeback_n102), .Y(exu_n15687));
OR2X1 exu_U38120(.A(se), .B(exu_n16398), .Y(ecl_perr_dff_n3));
INVX1 exu_U38121(.A(ecl_perr_dff_n3), .Y(exu_n15688));
INVX1 exu_U38122(.A(ecc_err_m[0]), .Y(exu_n15689));
AND2X1 exu_U38123(.A(div_input_data_e[69]), .B(ecl_shiftop_e[2]), .Y(shft_n5));
INVX1 exu_U38124(.A(shft_n5), .Y(exu_n15690));
OR2X1 exu_U38125(.A(rml_tid_e[0]), .B(rml_tid_e[1]), .Y(rml_cwp_thr_e[0]));
INVX1 exu_U38126(.A(rml_cwp_thr_e[0]), .Y(exu_n15691));
INVX1 exu_U38127(.A(rml_tid_e[0]), .Y(exu_n16570));
OR2X1 exu_U38128(.A(exu_n16375), .B(ifu_tlu_sraddr_d[0]), .Y(ecl_writeback_sel_cansave_d));
INVX1 exu_U38129(.A(ecl_writeback_sel_cansave_d), .Y(exu_n15692));
INVX1 exu_U38130(.A(exu_n27986), .Y(exu_n15693));
INVX1 exu_U38131(.A(shft_rshifterinput_b1[57]), .Y(exu_n15694));
INVX1 exu_U38132(.A(exu_n27989), .Y(exu_n15695));
INVX1 exu_U38133(.A(ecl_ccr_exu_ifu_cc_w[0]), .Y(exu_n15696));
INVX1 exu_U38134(.A(ecl_ccr_exu_ifu_cc_w[1]), .Y(exu_n15697));
INVX1 exu_U38135(.A(ecl_ccr_exu_ifu_cc_w[2]), .Y(exu_n15698));
INVX1 exu_U38136(.A(ecl_ccr_exu_ifu_cc_w[3]), .Y(exu_n15699));
INVX1 exu_U38137(.A(ecl_ccr_exu_ifu_cc_w[4]), .Y(exu_n15700));
INVX1 exu_U38138(.A(ecl_ccr_exu_ifu_cc_w[5]), .Y(exu_n15701));
INVX1 exu_U38139(.A(ecl_ccr_exu_ifu_cc_w[6]), .Y(exu_n15702));
INVX1 exu_U38140(.A(exu_n27921), .Y(exu_n15703));
INVX1 exu_U38141(.A(exu_n27924), .Y(exu_n15704));
INVX1 exu_U38142(.A(exu_n27928), .Y(exu_n15705));
INVX1 exu_U38143(.A(exu_n27931), .Y(exu_n15706));
INVX1 exu_U38144(.A(exu_n27934), .Y(exu_n15707));
INVX1 exu_U38145(.A(exu_n27937), .Y(exu_n15708));
INVX1 exu_U38146(.A(exu_n27940), .Y(exu_n15709));
INVX1 exu_U38147(.A(exu_n27943), .Y(exu_n15710));
INVX1 exu_U38148(.A(exu_n27946), .Y(exu_n15711));
INVX1 exu_U38149(.A(exu_n27949), .Y(exu_n15712));
INVX1 exu_U38150(.A(exu_n27952), .Y(exu_n15713));
INVX1 exu_U38151(.A(exu_n27955), .Y(exu_n15714));
INVX1 exu_U38152(.A(exu_n27959), .Y(exu_n15715));
INVX1 exu_U38153(.A(exu_n27962), .Y(exu_n15716));
INVX1 exu_U38154(.A(exu_n27965), .Y(exu_n15717));
INVX1 exu_U38155(.A(exu_n27968), .Y(exu_n15718));
INVX1 exu_U38156(.A(exu_n28016), .Y(exu_n15719));
INVX1 exu_U38157(.A(exu_n28079), .Y(exu_n15720));
INVX1 exu_U38158(.A(shft_rshifterinput_b1[63]), .Y(exu_n15721));
INVX1 exu_U38159(.A(shft_rshifterinput_b1[62]), .Y(exu_n15722));
INVX1 exu_U38160(.A(shft_rshifterinput_b1[61]), .Y(exu_n15723));
INVX1 exu_U38161(.A(shft_rshifterinput_b1[60]), .Y(exu_n15724));
INVX1 exu_U38162(.A(shft_rshifterinput_b1[59]), .Y(exu_n15725));
INVX1 exu_U38163(.A(shft_rshifterinput_b1[58]), .Y(exu_n15726));
INVX1 exu_U38164(.A(shft_rshifterinput_b1[56]), .Y(exu_n15727));
INVX1 exu_U38165(.A(shft_rshifterinput_b1[55]), .Y(exu_n15728));
INVX1 exu_U38166(.A(shft_rshifterinput_b1[54]), .Y(exu_n15729));
INVX1 exu_U38167(.A(shft_rshifterinput_b1[53]), .Y(exu_n15730));
INVX1 exu_U38168(.A(shft_rshifterinput_b1[52]), .Y(exu_n15731));
INVX1 exu_U38169(.A(shft_rshifterinput_b1[51]), .Y(exu_n15732));
INVX1 exu_U38170(.A(shft_rshifterinput_b1[50]), .Y(exu_n15733));
INVX1 exu_U38171(.A(shft_rshifterinput_b1[49]), .Y(exu_n15734));
INVX1 exu_U38172(.A(shft_rshifterinput_b1[48]), .Y(exu_n15735));
INVX1 exu_U38173(.A(ecl_divcntl_ccr_cc_w2[3]), .Y(exu_n15736));
INVX1 exu_U38174(.A(ecl_divcntl_ccr_cc_w2[2]), .Y(exu_n15737));
AND2X1 exu_U38175(.A(ecl_divcntl_n74), .B(ecl_divcntl_n72), .Y(ecl_divcntl_ccr_cc_w2[1]));
INVX1 exu_U38176(.A(ecl_divcntl_ccr_cc_w2[1]), .Y(exu_n15738));
INVX1 exu_U38177(.A(ecl_writeback_n98), .Y(exu_n15739));
INVX1 exu_U38178(.A(rml_rml_kill_w), .Y(exu_n15740));
AND2X1 exu_U38179(.A(ecl_writeback_n192), .B(ecl_mdqctl_wb_yreg_shift_g), .Y(ecl_writeback_n76));
INVX1 exu_U38180(.A(ecl_writeback_n76), .Y(exu_n15741));
INVX1 exu_U38181(.A(ecl_writeback_n97), .Y(exu_n15742));
INVX1 exu_U38182(.A(ecl_writeback_n80), .Y(exu_n15743));
INVX1 exu_U38183(.A(ecl_writeback_n84), .Y(exu_n15744));
INVX1 exu_U38184(.A(exu_n18191), .Y(exu_n15745));
AND2X1 exu_U38185(.A(rml_canrestore_wen_w), .B(ecl_rml_thr_w[3]), .Y(exu_n18191));
INVX1 exu_U38186(.A(exu_n18192), .Y(exu_n15746));
AND2X1 exu_U38187(.A(ecl_rml_thr_w[2]), .B(rml_canrestore_wen_w), .Y(exu_n18192));
INVX1 exu_U38188(.A(exu_n18193), .Y(exu_n15747));
AND2X1 exu_U38189(.A(exu_n15957), .B(rml_canrestore_wen_w), .Y(exu_n18193));
INVX1 exu_U38190(.A(exu_n18194), .Y(exu_n15748));
AND2X1 exu_U38191(.A(exu_n15959), .B(rml_canrestore_wen_w), .Y(exu_n18194));
INVX1 exu_U38192(.A(exu_n18235), .Y(exu_n15749));
AND2X1 exu_U38193(.A(rml_otherwin_wen_w), .B(ecl_rml_thr_w[3]), .Y(exu_n18235));
INVX1 exu_U38194(.A(exu_n18236), .Y(exu_n15750));
AND2X1 exu_U38195(.A(ecl_rml_thr_w[2]), .B(rml_otherwin_wen_w), .Y(exu_n18236));
INVX1 exu_U38196(.A(exu_n18237), .Y(exu_n15751));
AND2X1 exu_U38197(.A(exu_n15957), .B(rml_otherwin_wen_w), .Y(exu_n18237));
INVX1 exu_U38198(.A(exu_n18238), .Y(exu_n15752));
AND2X1 exu_U38199(.A(exu_n15959), .B(rml_otherwin_wen_w), .Y(exu_n18238));
INVX1 exu_U38200(.A(exu_n18279), .Y(exu_n15753));
AND2X1 exu_U38201(.A(rml_cleanwin_wen_w), .B(ecl_rml_thr_w[3]), .Y(exu_n18279));
INVX1 exu_U38202(.A(exu_n18280), .Y(exu_n15754));
AND2X1 exu_U38203(.A(ecl_rml_thr_w[2]), .B(rml_cleanwin_wen_w), .Y(exu_n18280));
INVX1 exu_U38204(.A(exu_n18281), .Y(exu_n15755));
AND2X1 exu_U38205(.A(exu_n15957), .B(rml_cleanwin_wen_w), .Y(exu_n18281));
INVX1 exu_U38206(.A(exu_n18282), .Y(exu_n15756));
AND2X1 exu_U38207(.A(exu_n15959), .B(rml_cleanwin_wen_w), .Y(exu_n18282));
AND2X1 exu_U38208(.A(ecl_tid_w[1]), .B(exu_n16576), .Y(ecl_rml_thr_w[2]));
BUFX2 exu_U38209(.A(exu_n15404), .Y(exu_n15957));
BUFX2 exu_U38210(.A(exu_n15405), .Y(exu_n15959));
INVX1 exu_U38211(.A(rml_cansave_reg_n5), .Y(exu_n15757));
AND2X1 exu_U38212(.A(rml_cansave_wen_w), .B(ecl_rml_thr_w[3]), .Y(rml_cansave_reg_n5));
INVX1 exu_U38213(.A(rml_cansave_reg_n6), .Y(exu_n15758));
AND2X1 exu_U38214(.A(ecl_rml_thr_w[2]), .B(rml_cansave_wen_w), .Y(rml_cansave_reg_n6));
INVX1 exu_U38215(.A(rml_cansave_reg_n7), .Y(exu_n15759));
AND2X1 exu_U38216(.A(exu_n15957), .B(rml_cansave_wen_w), .Y(rml_cansave_reg_n7));
INVX1 exu_U38217(.A(rml_cansave_reg_n8), .Y(exu_n15760));
AND2X1 exu_U38218(.A(exu_n15959), .B(rml_cansave_wen_w), .Y(rml_cansave_reg_n8));
AND2X1 exu_U38219(.A(ecl_writeback_n198), .B(exu_n16600), .Y(ecl_writeback_n130));
INVX1 exu_U38220(.A(ecl_writeback_n130), .Y(exu_n15761));
INVX1 exu_U38221(.A(rml_n130), .Y(exu_n15762));
INVX1 exu_U38222(.A(rml_n131), .Y(exu_n15763));
INVX1 exu_U38223(.A(exu_n15765), .Y(exu_n15764));
AND2X1 exu_U38224(.A(ecl_wb_byplog_wen_g2), .B(ecl_writeback_n198), .Y(ecl_writeback_n167));
INVX1 exu_U38225(.A(ecl_writeback_n167), .Y(exu_n15765));
INVX1 exu_U38226(.A(rml_cwp_n47), .Y(exu_n15766));
INVX1 exu_U38227(.A(ecl_byplog_rs1_n24), .Y(exu_n15767));
INVX1 exu_U38228(.A(ecl_mdqctl_n63), .Y(exu_n15768));
INVX1 exu_U38229(.A(ecl_byplog_rs1_n17), .Y(exu_n15769));
AND2X1 exu_U38230(.A(ecc_decode_n37), .B(ecc_decode_n18), .Y(ecc_decode_n28));
INVX1 exu_U38231(.A(ecc_decode_n28), .Y(exu_n15770));
AND2X1 exu_U38232(.A(ecc_decode_n37), .B(ecc_decode_n21), .Y(ecc_decode_n30));
INVX1 exu_U38233(.A(ecc_decode_n30), .Y(exu_n15771));
AND2X1 exu_U38234(.A(ecc_decode_n37), .B(ecc_decode_n22), .Y(ecc_decode_n31));
INVX1 exu_U38235(.A(ecc_decode_n31), .Y(exu_n15772));
AND2X1 exu_U38236(.A(ecc_decode_n37), .B(ecc_decode_n24), .Y(ecc_decode_n32));
INVX1 exu_U38237(.A(ecc_decode_n32), .Y(exu_n15773));
INVX1 exu_U38238(.A(ecc_decode_n19), .Y(exu_n15774));
INVX1 exu_U38239(.A(ecl_writeback_n176), .Y(exu_n15775));
AND2X1 exu_U38240(.A(ecl_writeback_yreg_wen_w1), .B(exu_n16607), .Y(ecl_writeback_n176));
AND2X1 exu_U38241(.A(ecc_decode_n43), .B(ecc_decode_n18), .Y(ecc_decode_n39));
INVX1 exu_U38242(.A(ecc_decode_n39), .Y(exu_n15776));
AND2X1 exu_U38243(.A(ecc_decode_n43), .B(ecc_decode_n21), .Y(ecc_decode_n40));
INVX1 exu_U38244(.A(ecc_decode_n40), .Y(exu_n15777));
AND2X1 exu_U38245(.A(ecc_decode_n43), .B(ecc_decode_n22), .Y(ecc_decode_n41));
INVX1 exu_U38246(.A(ecc_decode_n41), .Y(exu_n15778));
INVX1 exu_U38247(.A(bypass_rd_data_g[61]), .Y(exu_n15779));
INVX1 exu_U38248(.A(bypass_rd_data_g[60]), .Y(exu_n15780));
INVX1 exu_U38249(.A(bypass_rd_data_g[54]), .Y(exu_n15781));
INVX1 exu_U38250(.A(bypass_rd_data_g[49]), .Y(exu_n15782));
INVX1 exu_U38251(.A(bypass_rd_data_g[48]), .Y(exu_n15783));
INVX1 exu_U38252(.A(bypass_rd_data_g[45]), .Y(exu_n15784));
INVX1 exu_U38253(.A(bypass_rd_data_g[43]), .Y(exu_n15785));
INVX1 exu_U38254(.A(bypass_rd_data_g[37]), .Y(exu_n15786));
INVX1 exu_U38255(.A(bypass_rd_data_g[35]), .Y(exu_n15787));
INVX1 exu_U38256(.A(bypass_rd_data_g[33]), .Y(exu_n15788));
INVX1 exu_U38257(.A(bypass_rd_data_g[29]), .Y(exu_n15789));
INVX1 exu_U38258(.A(bypass_rd_data_g[22]), .Y(exu_n15790));
INVX1 exu_U38259(.A(bypass_rd_data_g[20]), .Y(exu_n15791));
INVX1 exu_U38260(.A(bypass_rd_data_g[18]), .Y(exu_n15792));
INVX1 exu_U38261(.A(bypass_rd_data_g[14]), .Y(exu_n15793));
INVX1 exu_U38262(.A(ecl_div_cin), .Y(exu_n15794));
INVX1 exu_U38263(.A(alu_ecl_cout32_e), .Y(exu_n15795));
INVX1 exu_U38264(.A(bypass_rd_data_g[62]), .Y(exu_n15796));
INVX1 exu_U38265(.A(bypass_rd_data_g[59]), .Y(exu_n15797));
INVX1 exu_U38266(.A(bypass_rd_data_g[57]), .Y(exu_n15798));
INVX1 exu_U38267(.A(bypass_rd_data_g[55]), .Y(exu_n15799));
INVX1 exu_U38268(.A(bypass_rd_data_g[50]), .Y(exu_n15800));
INVX1 exu_U38269(.A(bypass_rd_data_g[4]), .Y(exu_n15801));
INVX1 exu_U38270(.A(bypass_rd_data_g[47]), .Y(exu_n15802));
INVX1 exu_U38271(.A(bypass_rd_data_g[42]), .Y(exu_n15803));
INVX1 exu_U38272(.A(bypass_rd_data_g[34]), .Y(exu_n15804));
INVX1 exu_U38273(.A(bypass_rd_data_g[27]), .Y(exu_n15805));
INVX1 exu_U38274(.A(bypass_rd_data_g[26]), .Y(exu_n15806));
INVX1 exu_U38275(.A(bypass_rd_data_g[23]), .Y(exu_n15807));
INVX1 exu_U38276(.A(bypass_rd_data_g[19]), .Y(exu_n15808));
INVX1 exu_U38277(.A(bypass_rd_data_g[12]), .Y(exu_n15809));
INVX1 exu_U38278(.A(bypass_rd_data_g[0]), .Y(exu_n15810));
INVX1 exu_U38279(.A(bypass_rd_data_g[58]), .Y(exu_n15811));
INVX1 exu_U38280(.A(bypass_rd_data_g[52]), .Y(exu_n15812));
INVX1 exu_U38281(.A(bypass_rd_data_g[1]), .Y(exu_n15813));
INVX1 exu_U38282(.A(div_ecl_dividend_msb), .Y(exu_n15814));
INVX1 exu_U38283(.A(ecl_divcntl_n24), .Y(exu_n15815));
OR2X1 exu_U38284(.A(exu_n15839), .B(se), .Y(ecl_writeback_restore_rd_dff_n6));
INVX1 exu_U38285(.A(ecl_writeback_restore_rd_dff_n6), .Y(exu_n15816));
OR2X1 exu_U38286(.A(exu_n16390), .B(ecl_ifu_tlu_flush_w), .Y(ecl_rml_inst_vld_w));
INVX1 exu_U38287(.A(ecl_rml_inst_vld_w), .Y(exu_n15817));
AND2X1 exu_U38288(.A(exu_n19214), .B(ecl_ld_thr_match_dg), .Y(exu_n19191));
INVX1 exu_U38289(.A(exu_n19191), .Y(exu_n15818));
AND2X1 exu_U38290(.A(exu_n19250), .B(ecl_ld_thr_match_dg), .Y(exu_n19227));
INVX1 exu_U38291(.A(exu_n19227), .Y(exu_n15819));
AND2X1 exu_U38292(.A(ecl_byplog_rs2_n46), .B(ecl_ld_thr_match_dg), .Y(ecl_byplog_rs2_n20));
INVX1 exu_U38293(.A(ecl_byplog_rs2_n20), .Y(exu_n15820));
BUFX2 exu_U38294(.A(rml_rml_reset_l), .Y(exu_n15821));
INVX1 exu_U38295(.A(ecl_rml_cwp_wen_e), .Y(exu_n15822));
INVX1 exu_U38296(.A(div_adderin1[63]), .Y(exu_n15823));
INVX1 exu_U38297(.A(ecl_writeback_sel_wstate_d), .Y(exu_n15824));
INVX1 exu_U38298(.A(bypass_rd_data_g[7]), .Y(exu_n15825));
INVX1 exu_U38299(.A(bypass_rd_data_g[63]), .Y(exu_n15826));
INVX1 exu_U38300(.A(bypass_rd_data_g[53]), .Y(exu_n15827));
INVX1 exu_U38301(.A(bypass_rd_data_g[41]), .Y(exu_n15828));
INVX1 exu_U38302(.A(bypass_rd_data_g[38]), .Y(exu_n15829));
INVX1 exu_U38303(.A(bypass_rd_data_g[31]), .Y(exu_n15830));
INVX1 exu_U38304(.A(bypass_rd_data_g[2]), .Y(exu_n15831));
INVX1 exu_U38305(.A(bypass_rd_data_g[16]), .Y(exu_n15832));
INVX1 exu_U38306(.A(bypass_rd_data_g[5]), .Y(exu_n15833));
INVX1 exu_U38307(.A(bypass_rd_data_g[56]), .Y(exu_n15834));
INVX1 exu_U38308(.A(bypass_rd_data_g[51]), .Y(exu_n15835));
INVX1 exu_U38309(.A(bypass_rd_data_g[25]), .Y(exu_n15836));
INVX1 exu_U38310(.A(bypass_rd_data_g[24]), .Y(exu_n15837));
INVX1 exu_U38311(.A(bypass_rd_data_g[11]), .Y(exu_n15838));
OR2X1 exu_U38312(.A(ecl_byp_restore_m), .B(se), .Y(ecl_writeback_restore_rd_dff_n3));
INVX1 exu_U38313(.A(ecl_writeback_restore_rd_dff_n3), .Y(exu_n15839));
INVX1 exu_U38314(.A(bypass_rd_data_g[8]), .Y(exu_n15840));
INVX1 exu_U38315(.A(bypass_rd_data_g[44]), .Y(exu_n15841));
INVX1 exu_U38316(.A(bypass_rd_data_g[40]), .Y(exu_n15842));
INVX1 exu_U38317(.A(bypass_rd_data_g[3]), .Y(exu_n15843));
INVX1 exu_U38318(.A(bypass_rd_data_g[39]), .Y(exu_n15844));
INVX1 exu_U38319(.A(bypass_rd_data_g[30]), .Y(exu_n15845));
INVX1 exu_U38320(.A(bypass_rd_data_g[28]), .Y(exu_n15846));
INVX1 exu_U38321(.A(bypass_rd_data_g[21]), .Y(exu_n15847));
INVX1 exu_U38322(.A(bypass_rd_data_g[15]), .Y(exu_n15848));
INVX1 exu_U38323(.A(bypass_rd_data_g[13]), .Y(exu_n15849));
INVX1 exu_U38324(.A(bypass_rd_data_g[10]), .Y(exu_n15850));
INVX1 exu_U38325(.A(rml_next_cwp_e[2]), .Y(exu_n15851));
INVX1 exu_U38326(.A(rml_next_cwp_e[1]), .Y(exu_n15852));
INVX1 exu_U38327(.A(rml_next_cwp_e[0]), .Y(exu_n15853));
INVX1 exu_U38328(.A(bypass_rd_data_g[6]), .Y(exu_n15854));
INVX1 exu_U38329(.A(bypass_rd_data_g[46]), .Y(exu_n15855));
INVX1 exu_U38330(.A(exu_n15857), .Y(exu_n15856));
BUFX2 exu_U38331(.A(rml_irf_old_lo_cwp_e[0]), .Y(exu_n15857));
INVX1 exu_U38332(.A(div_adderin1[32]), .Y(exu_n15858));
INVX1 exu_U38333(.A(div_adderin1[0]), .Y(exu_n15859));
INVX1 exu_U38334(.A(div_adderin1[9]), .Y(exu_n15860));
INVX1 exu_U38335(.A(div_adderin1[8]), .Y(exu_n15861));
INVX1 exu_U38336(.A(div_adderin1[7]), .Y(exu_n15862));
INVX1 exu_U38337(.A(div_adderin1[6]), .Y(exu_n15863));
INVX1 exu_U38338(.A(div_adderin1[62]), .Y(exu_n15864));
INVX1 exu_U38339(.A(div_adderin1[61]), .Y(exu_n15865));
INVX1 exu_U38340(.A(div_adderin1[60]), .Y(exu_n15866));
INVX1 exu_U38341(.A(div_adderin1[5]), .Y(exu_n15867));
INVX1 exu_U38342(.A(div_adderin1[59]), .Y(exu_n15868));
INVX1 exu_U38343(.A(div_adderin1[58]), .Y(exu_n15869));
INVX1 exu_U38344(.A(div_adderin1[57]), .Y(exu_n15870));
INVX1 exu_U38345(.A(div_adderin1[56]), .Y(exu_n15871));
INVX1 exu_U38346(.A(div_adderin1[55]), .Y(exu_n15872));
INVX1 exu_U38347(.A(div_adderin1[54]), .Y(exu_n15873));
INVX1 exu_U38348(.A(div_adderin1[53]), .Y(exu_n15874));
INVX1 exu_U38349(.A(div_adderin1[52]), .Y(exu_n15875));
INVX1 exu_U38350(.A(div_adderin1[51]), .Y(exu_n15876));
INVX1 exu_U38351(.A(div_adderin1[50]), .Y(exu_n15877));
INVX1 exu_U38352(.A(div_adderin1[4]), .Y(exu_n15878));
INVX1 exu_U38353(.A(div_adderin1[49]), .Y(exu_n15879));
INVX1 exu_U38354(.A(div_adderin1[48]), .Y(exu_n15880));
INVX1 exu_U38355(.A(div_adderin1[47]), .Y(exu_n15881));
INVX1 exu_U38356(.A(div_adderin1[46]), .Y(exu_n15882));
INVX1 exu_U38357(.A(div_adderin1[45]), .Y(exu_n15883));
INVX1 exu_U38358(.A(div_adderin1[44]), .Y(exu_n15884));
INVX1 exu_U38359(.A(div_adderin1[43]), .Y(exu_n15885));
INVX1 exu_U38360(.A(div_adderin1[42]), .Y(exu_n15886));
INVX1 exu_U38361(.A(div_adderin1[41]), .Y(exu_n15887));
INVX1 exu_U38362(.A(div_adderin1[40]), .Y(exu_n15888));
INVX1 exu_U38363(.A(div_adderin1[3]), .Y(exu_n15889));
INVX1 exu_U38364(.A(div_adderin1[39]), .Y(exu_n15890));
INVX1 exu_U38365(.A(div_adderin1[38]), .Y(exu_n15891));
INVX1 exu_U38366(.A(div_adderin1[37]), .Y(exu_n15892));
INVX1 exu_U38367(.A(div_adderin1[36]), .Y(exu_n15893));
INVX1 exu_U38368(.A(div_adderin1[35]), .Y(exu_n15894));
INVX1 exu_U38369(.A(div_adderin1[34]), .Y(exu_n15895));
INVX1 exu_U38370(.A(div_adderin1[33]), .Y(exu_n15896));
INVX1 exu_U38371(.A(div_adderin1[31]), .Y(exu_n15897));
INVX1 exu_U38372(.A(div_adderin1[30]), .Y(exu_n15898));
INVX1 exu_U38373(.A(div_adderin1[2]), .Y(exu_n15899));
INVX1 exu_U38374(.A(div_adderin1[29]), .Y(exu_n15900));
INVX1 exu_U38375(.A(div_adderin1[28]), .Y(exu_n15901));
INVX1 exu_U38376(.A(div_adderin1[27]), .Y(exu_n15902));
INVX1 exu_U38377(.A(div_adderin1[26]), .Y(exu_n15903));
INVX1 exu_U38378(.A(div_adderin1[25]), .Y(exu_n15904));
INVX1 exu_U38379(.A(div_adderin1[24]), .Y(exu_n15905));
INVX1 exu_U38380(.A(div_adderin1[23]), .Y(exu_n15906));
INVX1 exu_U38381(.A(div_adderin1[22]), .Y(exu_n15907));
INVX1 exu_U38382(.A(div_adderin1[21]), .Y(exu_n15908));
INVX1 exu_U38383(.A(div_adderin1[20]), .Y(exu_n15909));
INVX1 exu_U38384(.A(div_adderin1[1]), .Y(exu_n15910));
INVX1 exu_U38385(.A(div_adderin1[19]), .Y(exu_n15911));
INVX1 exu_U38386(.A(div_adderin1[18]), .Y(exu_n15912));
INVX1 exu_U38387(.A(div_adderin1[17]), .Y(exu_n15913));
INVX1 exu_U38388(.A(div_adderin1[16]), .Y(exu_n15914));
INVX1 exu_U38389(.A(div_adderin1[15]), .Y(exu_n15915));
INVX1 exu_U38390(.A(div_adderin1[14]), .Y(exu_n15916));
INVX1 exu_U38391(.A(div_adderin1[13]), .Y(exu_n15917));
INVX1 exu_U38392(.A(div_adderin1[12]), .Y(exu_n15918));
INVX1 exu_U38393(.A(div_adderin1[11]), .Y(exu_n15919));
INVX1 exu_U38394(.A(div_adderin1[10]), .Y(exu_n15920));
OR2X1 exu_U38395(.A(exu_n16578), .B(exu_n16577), .Y(ecl_rml_thr_m[3]));
INVX1 exu_U38396(.A(ecl_rml_thr_m[3]), .Y(exu_n15921));
OR2X1 exu_U38397(.A(exu_n16578), .B(ecl_tid_m[0]), .Y(ecl_rml_thr_m[2]));
INVX1 exu_U38398(.A(ecl_rml_thr_m[2]), .Y(exu_n15922));
OR2X1 exu_U38399(.A(exu_n16577), .B(ecl_tid_m[1]), .Y(ecl_rml_thr_m[1]));
INVX1 exu_U38400(.A(ecl_rml_thr_m[1]), .Y(exu_n15923));
OR2X1 exu_U38401(.A(ecl_tid_m[0]), .B(ecl_tid_m[1]), .Y(ecl_rml_thr_m[0]));
INVX1 exu_U38402(.A(ecl_rml_thr_m[0]), .Y(exu_n15924));
INVX1 exu_U38403(.A(rml_full_swap_e), .Y(exu_n15925));
AND2X1 exu_U38404(.A(rml_exu_tlu_spill_e), .B(ecl_rml_cwp_wen_e), .Y(rml_full_swap_e));
INVX1 exu_U38405(.A(ecl_ccr_n14), .Y(exu_n15926));
INVX1 exu_U38406(.A(bypass_rd_data_g[36]), .Y(exu_n15927));
INVX1 exu_U38407(.A(bypass_rd_data_g[32]), .Y(exu_n15928));
INVX1 exu_U38408(.A(bypass_rd_data_g[17]), .Y(exu_n15929));
INVX1 exu_U38409(.A(ecl_pick_normal_ttype), .Y(exu_n15930));
OR2X1 exu_U38410(.A(ecl_ccr_n24), .B(ecl_ccr_use_cc_w), .Y(ecl_ccr_mux_ccr_bypass1_sel0));
INVX1 exu_U38411(.A(ecl_ccr_mux_ccr_bypass1_sel0), .Y(exu_n15931));
INVX1 exu_U38412(.A(ecc_decode_n36), .Y(exu_n15932));
AND2X1 exu_U38413(.A(ecc_err_m[0]), .B(ecc_err_m[3]), .Y(ecc_decode_n36));
OR2X1 exu_U38414(.A(ecl_tid_d[0]), .B(exu_n15944), .Y(ecl_thr_d[2]));
INVX1 exu_U38415(.A(ecl_thr_d[2]), .Y(exu_n15933));
OR2X1 exu_U38416(.A(ecl_tid_d[1]), .B(exu_n15945), .Y(ecl_thr_d[1]));
INVX1 exu_U38417(.A(ecl_thr_d[1]), .Y(exu_n15934));
OR2X1 exu_U38418(.A(ecl_tid_d[1]), .B(ecl_tid_d[0]), .Y(ecl_thr_d[0]));
INVX1 exu_U38419(.A(ecl_thr_d[0]), .Y(exu_n15935));
INVX1 exu_U38420(.A(ecc_decode_n29), .Y(exu_n15936));
INVX1 exu_U38421(.A(ecc_decode_n27), .Y(exu_n15937));
INVX1 exu_U38422(.A(ecc_decode_n35), .Y(exu_n15938));
INVX1 exu_U38423(.A(ecl_wb_ccr_wrccr_w), .Y(exu_n15939));
INVX1 exu_U38424(.A(rml_exu_tlu_spill_e), .Y(exu_n15940));
INVX1 exu_U38425(.A(exu_n15189), .Y(exu_n15950));
INVX1 exu_U38426(.A(exu_n15189), .Y(exu_n15951));
INVX1 exu_U38427(.A(exu_n15191), .Y(exu_n15952));
INVX1 exu_U38428(.A(exu_n15191), .Y(exu_n15953));
INVX1 exu_U38429(.A(exu_n15191), .Y(exu_n15954));
INVX1 exu_U38430(.A(exu_n15193), .Y(exu_n15955));
INVX1 exu_U38431(.A(exu_n15193), .Y(exu_n15956));
XNOR2X1 exu_U38432(.A(ecl_wb_byplog_rd_g2[2]), .B(ecl_ifu_exu_rs1_d[2]), .Y(exu_n16635));
XNOR2X1 exu_U38433(.A(ecl_wb_byplog_rd_g2[4]), .B(ecl_ifu_exu_rs1_d[4]), .Y(exu_n16638));
XNOR2X1 exu_U38434(.A(ecl_wb_byplog_rd_g2[3]), .B(ecl_ifu_exu_rs1_d[3]), .Y(exu_n16637));
XNOR2X1 exu_U38435(.A(ecl_ld_rd_g[2]), .B(ecl_ifu_exu_rs1_d[2]), .Y(exu_n16649));
XNOR2X1 exu_U38436(.A(ecl_ld_rd_g[4]), .B(ecl_ifu_exu_rs1_d[4]), .Y(exu_n16652));
XNOR2X1 exu_U38437(.A(ecl_ld_rd_g[3]), .B(ecl_ifu_exu_rs1_d[3]), .Y(exu_n16651));
XNOR2X1 exu_U38438(.A(ecl_rd_m[2]), .B(ecl_ifu_exu_rs1_d[2]), .Y(exu_n16663));
XNOR2X1 exu_U38439(.A(ecl_rd_m[4]), .B(ecl_ifu_exu_rs1_d[4]), .Y(exu_n16666));
XNOR2X1 exu_U38440(.A(ecl_rd_m[3]), .B(ecl_ifu_exu_rs1_d[3]), .Y(exu_n16665));
XNOR2X1 exu_U38441(.A(ecl_rd_e[2]), .B(ecl_ifu_exu_rs1_d[2]), .Y(exu_n16677));
XNOR2X1 exu_U38442(.A(ecl_rd_e[4]), .B(ecl_ifu_exu_rs1_d[4]), .Y(exu_n16680));
XNOR2X1 exu_U38443(.A(ecl_rd_e[3]), .B(ecl_ifu_exu_rs1_d[3]), .Y(exu_n16679));
XNOR2X1 exu_U38444(.A(ecl_wb_byplog_rd_g2[2]), .B(ecl_ifu_exu_rs2_d[2]), .Y(exu_n16691));
XNOR2X1 exu_U38445(.A(ecl_wb_byplog_rd_g2[4]), .B(ecl_ifu_exu_rs2_d[4]), .Y(exu_n16694));
XNOR2X1 exu_U38446(.A(ecl_wb_byplog_rd_g2[3]), .B(ecl_ifu_exu_rs2_d[3]), .Y(exu_n16693));
XNOR2X1 exu_U38447(.A(ecl_ld_rd_g[2]), .B(ecl_ifu_exu_rs2_d[2]), .Y(exu_n16705));
XNOR2X1 exu_U38448(.A(ecl_ld_rd_g[4]), .B(ecl_ifu_exu_rs2_d[4]), .Y(exu_n16708));
XNOR2X1 exu_U38449(.A(ecl_ld_rd_g[3]), .B(ecl_ifu_exu_rs2_d[3]), .Y(exu_n16707));
XNOR2X1 exu_U38450(.A(ecl_rd_m[2]), .B(ecl_ifu_exu_rs2_d[2]), .Y(exu_n16719));
XNOR2X1 exu_U38451(.A(ecl_rd_m[4]), .B(ecl_ifu_exu_rs2_d[4]), .Y(exu_n16722));
XNOR2X1 exu_U38452(.A(ecl_rd_m[3]), .B(ecl_ifu_exu_rs2_d[3]), .Y(exu_n16721));
XNOR2X1 exu_U38453(.A(ecl_rd_e[2]), .B(ecl_ifu_exu_rs2_d[2]), .Y(exu_n16733));
XNOR2X1 exu_U38454(.A(ecl_rd_e[4]), .B(ecl_ifu_exu_rs2_d[4]), .Y(exu_n16736));
XNOR2X1 exu_U38455(.A(ecl_rd_e[3]), .B(ecl_ifu_exu_rs2_d[3]), .Y(exu_n16735));
XOR2X1 exu_U38456(.A(exu_n15794), .B(div_adderin2[0]), .Y(exu_n16739));
XOR2X1 exu_U38457(.A(exu_n15859), .B(exu_n16739), .Y(div_adder_out_0));
XOR2X1 exu_U38458(.A(div_adderin2[10]), .B(exu_n15920), .Y(exu_n16770));
XOR2X1 exu_U38459(.A(exu_n15595), .B(exu_n16770), .Y(div_adder_out_10));
XOR2X1 exu_U38460(.A(div_adderin2[11]), .B(exu_n15919), .Y(exu_n16775));
XOR2X1 exu_U38461(.A(exu_n15596), .B(exu_n16775), .Y(div_adder_out_11));
XOR2X1 exu_U38462(.A(div_adderin2[12]), .B(exu_n15918), .Y(exu_n16780));
XOR2X1 exu_U38463(.A(exu_n15597), .B(exu_n16780), .Y(div_adder_out_12));
XOR2X1 exu_U38464(.A(div_adderin2[13]), .B(exu_n15917), .Y(exu_n16785));
XOR2X1 exu_U38465(.A(exu_n15598), .B(exu_n16785), .Y(div_adder_out_13));
XOR2X1 exu_U38466(.A(div_adderin2[14]), .B(exu_n15916), .Y(exu_n16790));
XOR2X1 exu_U38467(.A(exu_n15599), .B(exu_n16790), .Y(div_adder_out_14));
XOR2X1 exu_U38468(.A(div_adderin2[15]), .B(exu_n15915), .Y(exu_n16795));
XOR2X1 exu_U38469(.A(exu_n15600), .B(exu_n16795), .Y(div_adder_out_15));
XOR2X1 exu_U38470(.A(div_adderin2[16]), .B(exu_n15914), .Y(exu_n16800));
XOR2X1 exu_U38471(.A(exu_n15601), .B(exu_n16800), .Y(div_adder_out_16));
XOR2X1 exu_U38472(.A(div_adderin2[17]), .B(exu_n15913), .Y(exu_n16805));
XOR2X1 exu_U38473(.A(exu_n15602), .B(exu_n16805), .Y(div_adder_out_17));
XOR2X1 exu_U38474(.A(div_adderin2[18]), .B(exu_n15912), .Y(exu_n16810));
XOR2X1 exu_U38475(.A(exu_n15603), .B(exu_n16810), .Y(div_adder_out_18));
XOR2X1 exu_U38476(.A(div_adderin2[19]), .B(exu_n15911), .Y(exu_n16815));
XOR2X1 exu_U38477(.A(exu_n15604), .B(exu_n16815), .Y(div_adder_out_19));
XOR2X1 exu_U38478(.A(div_adderin2[1]), .B(exu_n15910), .Y(exu_n16816));
XOR2X1 exu_U38479(.A(exu_n15559), .B(exu_n16816), .Y(div_adder_out_1));
XOR2X1 exu_U38480(.A(div_adderin2[20]), .B(exu_n15909), .Y(exu_n16822));
XOR2X1 exu_U38481(.A(exu_n15605), .B(exu_n16822), .Y(div_adder_out_20));
XOR2X1 exu_U38482(.A(div_adderin2[21]), .B(exu_n15908), .Y(exu_n16827));
XOR2X1 exu_U38483(.A(exu_n15606), .B(exu_n16827), .Y(div_adder_out_21));
XOR2X1 exu_U38484(.A(div_adderin2[22]), .B(exu_n15907), .Y(exu_n16832));
XOR2X1 exu_U38485(.A(exu_n15607), .B(exu_n16832), .Y(div_adder_out_22));
XOR2X1 exu_U38486(.A(div_adderin2[23]), .B(exu_n15906), .Y(exu_n16837));
XOR2X1 exu_U38487(.A(exu_n15608), .B(exu_n16837), .Y(div_adder_out_23));
XOR2X1 exu_U38488(.A(div_adderin2[24]), .B(exu_n15905), .Y(exu_n16842));
XOR2X1 exu_U38489(.A(exu_n15609), .B(exu_n16842), .Y(div_adder_out_24));
XOR2X1 exu_U38490(.A(div_adderin2[25]), .B(exu_n15904), .Y(exu_n16847));
XOR2X1 exu_U38491(.A(exu_n15610), .B(exu_n16847), .Y(div_adder_out_25));
XOR2X1 exu_U38492(.A(div_adderin2[26]), .B(exu_n15903), .Y(exu_n16852));
XOR2X1 exu_U38493(.A(exu_n15611), .B(exu_n16852), .Y(div_adder_out_26));
XOR2X1 exu_U38494(.A(div_adderin2[27]), .B(exu_n15902), .Y(exu_n16857));
XOR2X1 exu_U38495(.A(exu_n15612), .B(exu_n16857), .Y(div_adder_out_27));
XOR2X1 exu_U38496(.A(div_adderin2[28]), .B(exu_n15901), .Y(exu_n16862));
XOR2X1 exu_U38497(.A(exu_n15613), .B(exu_n16862), .Y(div_adder_out_28));
XOR2X1 exu_U38498(.A(div_adderin2[29]), .B(exu_n15900), .Y(exu_n16867));
XOR2X1 exu_U38499(.A(exu_n15614), .B(exu_n16867), .Y(div_adder_out_29));
XOR2X1 exu_U38500(.A(div_adderin2[2]), .B(exu_n15899), .Y(exu_n16868));
XOR2X1 exu_U38501(.A(exu_n15560), .B(exu_n16868), .Y(div_adder_out_2));
XOR2X1 exu_U38502(.A(div_adderin2[30]), .B(exu_n15898), .Y(exu_n16874));
XOR2X1 exu_U38503(.A(exu_n15615), .B(exu_n16874), .Y(div_adder_out_30));
XOR2X1 exu_U38504(.A(div_adderin2[31]), .B(exu_n15897), .Y(exu_n16879));
XOR2X1 exu_U38505(.A(exu_n15616), .B(exu_n16879), .Y(div_ecl_adder_out_31));
XOR2X1 exu_U38506(.A(div_adderin2[3]), .B(exu_n15889), .Y(exu_n16884));
XOR2X1 exu_U38507(.A(exu_n15561), .B(exu_n16884), .Y(div_adder_out_3));
XOR2X1 exu_U38508(.A(div_adderin2[4]), .B(exu_n15878), .Y(exu_n16886));
XOR2X1 exu_U38509(.A(exu_n15562), .B(exu_n16886), .Y(div_adder_out_4));
XOR2X1 exu_U38510(.A(div_adderin2[5]), .B(exu_n15867), .Y(exu_n16888));
XOR2X1 exu_U38511(.A(exu_n15563), .B(exu_n16888), .Y(div_adder_out_5));
XOR2X1 exu_U38512(.A(div_adderin2[6]), .B(exu_n15863), .Y(exu_n16890));
XOR2X1 exu_U38513(.A(exu_n15564), .B(exu_n16890), .Y(div_adder_out_6));
XOR2X1 exu_U38514(.A(div_adderin2[7]), .B(exu_n15862), .Y(exu_n16892));
XOR2X1 exu_U38515(.A(exu_n15565), .B(exu_n16892), .Y(div_adder_out_7));
XOR2X1 exu_U38516(.A(div_adderin2[8]), .B(exu_n15861), .Y(exu_n16894));
XOR2X1 exu_U38517(.A(exu_n15566), .B(exu_n16894), .Y(div_adder_out_8));
XOR2X1 exu_U38518(.A(div_adderin2[9]), .B(exu_n15860), .Y(exu_n16896));
XOR2X1 exu_U38519(.A(exu_n15567), .B(exu_n16896), .Y(div_adder_out_9));
XOR2X1 exu_U38520(.A(exu_n15558), .B(div_adderin2[32]), .Y(exu_n16898));
XOR2X1 exu_U38521(.A(exu_n15858), .B(exu_n16898), .Y(div_adder_out[32]));
XOR2X1 exu_U38522(.A(div_adderin2[42]), .B(exu_n15886), .Y(exu_n16929));
XOR2X1 exu_U38523(.A(exu_n15617), .B(exu_n16929), .Y(div_adder_out[42]));
XOR2X1 exu_U38524(.A(div_adderin2[43]), .B(exu_n15885), .Y(exu_n16934));
XOR2X1 exu_U38525(.A(exu_n15618), .B(exu_n16934), .Y(div_adder_out[43]));
XOR2X1 exu_U38526(.A(div_adderin2[44]), .B(exu_n15884), .Y(exu_n16939));
XOR2X1 exu_U38527(.A(exu_n15619), .B(exu_n16939), .Y(div_adder_out[44]));
XOR2X1 exu_U38528(.A(div_adderin2[45]), .B(exu_n15883), .Y(exu_n16944));
XOR2X1 exu_U38529(.A(exu_n15620), .B(exu_n16944), .Y(div_adder_out[45]));
XOR2X1 exu_U38530(.A(div_adderin2[46]), .B(exu_n15882), .Y(exu_n16949));
XOR2X1 exu_U38531(.A(exu_n15621), .B(exu_n16949), .Y(div_adder_out[46]));
XOR2X1 exu_U38532(.A(div_adderin2[47]), .B(exu_n15881), .Y(exu_n16954));
XOR2X1 exu_U38533(.A(exu_n15622), .B(exu_n16954), .Y(div_adder_out[47]));
XOR2X1 exu_U38534(.A(div_adderin2[48]), .B(exu_n15880), .Y(exu_n16959));
XOR2X1 exu_U38535(.A(exu_n15623), .B(exu_n16959), .Y(div_adder_out[48]));
XOR2X1 exu_U38536(.A(div_adderin2[49]), .B(exu_n15879), .Y(exu_n16964));
XOR2X1 exu_U38537(.A(exu_n15624), .B(exu_n16964), .Y(div_adder_out[49]));
XOR2X1 exu_U38538(.A(div_adderin2[50]), .B(exu_n15877), .Y(exu_n16969));
XOR2X1 exu_U38539(.A(exu_n15625), .B(exu_n16969), .Y(div_adder_out[50]));
XOR2X1 exu_U38540(.A(div_adderin2[51]), .B(exu_n15876), .Y(exu_n16974));
XOR2X1 exu_U38541(.A(exu_n15626), .B(exu_n16974), .Y(div_adder_out[51]));
XOR2X1 exu_U38542(.A(div_adderin2[33]), .B(exu_n15896), .Y(exu_n16975));
XOR2X1 exu_U38543(.A(exu_n15568), .B(exu_n16975), .Y(div_adder_out[33]));
XOR2X1 exu_U38544(.A(div_adderin2[52]), .B(exu_n15875), .Y(exu_n16981));
XOR2X1 exu_U38545(.A(exu_n15627), .B(exu_n16981), .Y(div_adder_out[52]));
XOR2X1 exu_U38546(.A(div_adderin2[53]), .B(exu_n15874), .Y(exu_n16986));
XOR2X1 exu_U38547(.A(exu_n15628), .B(exu_n16986), .Y(div_adder_out[53]));
XOR2X1 exu_U38548(.A(div_adderin2[54]), .B(exu_n15873), .Y(exu_n16991));
XOR2X1 exu_U38549(.A(exu_n15629), .B(exu_n16991), .Y(div_adder_out[54]));
XOR2X1 exu_U38550(.A(div_adderin2[55]), .B(exu_n15872), .Y(exu_n16996));
XOR2X1 exu_U38551(.A(exu_n15630), .B(exu_n16996), .Y(div_adder_out[55]));
XOR2X1 exu_U38552(.A(div_adderin2[56]), .B(exu_n15871), .Y(exu_n17001));
XOR2X1 exu_U38553(.A(exu_n15631), .B(exu_n17001), .Y(div_adder_out[56]));
XOR2X1 exu_U38554(.A(div_adderin2[57]), .B(exu_n15870), .Y(exu_n17006));
XOR2X1 exu_U38555(.A(exu_n15632), .B(exu_n17006), .Y(div_adder_out[57]));
XOR2X1 exu_U38556(.A(div_adderin2[58]), .B(exu_n15869), .Y(exu_n17011));
XOR2X1 exu_U38557(.A(exu_n15633), .B(exu_n17011), .Y(div_adder_out[58]));
XOR2X1 exu_U38558(.A(div_adderin2[59]), .B(exu_n15868), .Y(exu_n17016));
XOR2X1 exu_U38559(.A(exu_n15634), .B(exu_n17016), .Y(div_adder_out[59]));
XOR2X1 exu_U38560(.A(div_adderin2[60]), .B(exu_n15866), .Y(exu_n17021));
XOR2X1 exu_U38561(.A(exu_n15635), .B(exu_n17021), .Y(div_adder_out[60]));
XOR2X1 exu_U38562(.A(div_adderin2[61]), .B(exu_n15865), .Y(exu_n17026));
XOR2X1 exu_U38563(.A(exu_n15636), .B(exu_n17026), .Y(div_adder_out[61]));
XOR2X1 exu_U38564(.A(div_adderin2[34]), .B(exu_n15895), .Y(exu_n17027));
XOR2X1 exu_U38565(.A(exu_n15569), .B(exu_n17027), .Y(div_adder_out[34]));
XOR2X1 exu_U38566(.A(div_adderin2[62]), .B(exu_n15864), .Y(exu_n17033));
XOR2X1 exu_U38567(.A(exu_n15637), .B(exu_n17033), .Y(div_adder_out[62]));
XOR2X1 exu_U38568(.A(div_adderin2[63]), .B(exu_n15823), .Y(exu_n17038));
XOR2X1 exu_U38569(.A(exu_n15638), .B(exu_n17038), .Y(div_adder_out[63]));
XOR2X1 exu_U38570(.A(div_adderin2[35]), .B(exu_n15894), .Y(exu_n17043));
XOR2X1 exu_U38571(.A(exu_n15570), .B(exu_n17043), .Y(div_adder_out[35]));
XOR2X1 exu_U38572(.A(div_adderin2[36]), .B(exu_n15893), .Y(exu_n17045));
XOR2X1 exu_U38573(.A(exu_n15571), .B(exu_n17045), .Y(div_adder_out[36]));
XOR2X1 exu_U38574(.A(div_adderin2[37]), .B(exu_n15892), .Y(exu_n17047));
XOR2X1 exu_U38575(.A(exu_n15572), .B(exu_n17047), .Y(div_adder_out[37]));
XOR2X1 exu_U38576(.A(div_adderin2[38]), .B(exu_n15891), .Y(exu_n17049));
XOR2X1 exu_U38577(.A(exu_n15573), .B(exu_n17049), .Y(div_adder_out[38]));
XOR2X1 exu_U38578(.A(div_adderin2[39]), .B(exu_n15890), .Y(exu_n17051));
XOR2X1 exu_U38579(.A(exu_n15574), .B(exu_n17051), .Y(div_adder_out[39]));
XOR2X1 exu_U38580(.A(div_adderin2[40]), .B(exu_n15888), .Y(exu_n17053));
XOR2X1 exu_U38581(.A(exu_n15575), .B(exu_n17053), .Y(div_adder_out[40]));
XOR2X1 exu_U38582(.A(div_adderin2[41]), .B(exu_n15887), .Y(exu_n17055));
XOR2X1 exu_U38583(.A(exu_n15576), .B(exu_n17055), .Y(div_adder_out[41]));
XOR2X1 exu_U38584(.A(ecl_alu_cin_e), .B(alu_addsub_rs2_data_0), .Y(exu_n17057));
XOR2X1 exu_U38585(.A(alu_logic_rs1_data_bf1[0]), .B(exu_n17057), .Y(exu_ifu_brpc_e[0]));
XOR2X1 exu_U38586(.A(alu_addsub_rs2_data_10), .B(alu_logic_rs1_data_bf1[10]), .Y(exu_n17088));
XOR2X1 exu_U38587(.A(exu_n15639), .B(exu_n17088), .Y(exu_ifu_brpc_e[10]));
XOR2X1 exu_U38588(.A(alu_addsub_rs2_data_11), .B(alu_logic_rs1_data_bf1[11]), .Y(exu_n17093));
XOR2X1 exu_U38589(.A(exu_n15640), .B(exu_n17093), .Y(exu_ifu_brpc_e[11]));
XOR2X1 exu_U38590(.A(alu_addsub_rs2_data_12), .B(alu_logic_rs1_data_bf1[12]), .Y(exu_n17098));
XOR2X1 exu_U38591(.A(exu_n15641), .B(exu_n17098), .Y(exu_ifu_brpc_e[12]));
XOR2X1 exu_U38592(.A(alu_addsub_rs2_data_13), .B(alu_logic_rs1_data_bf1[13]), .Y(exu_n17103));
XOR2X1 exu_U38593(.A(exu_n15642), .B(exu_n17103), .Y(exu_ifu_brpc_e[13]));
XOR2X1 exu_U38594(.A(alu_addsub_rs2_data_14), .B(alu_logic_rs1_data_bf1[14]), .Y(exu_n17108));
XOR2X1 exu_U38595(.A(exu_n15643), .B(exu_n17108), .Y(exu_ifu_brpc_e[14]));
XOR2X1 exu_U38596(.A(alu_addsub_rs2_data_15), .B(alu_logic_rs1_data_bf1[15]), .Y(exu_n17113));
XOR2X1 exu_U38597(.A(exu_n15644), .B(exu_n17113), .Y(exu_ifu_brpc_e[15]));
XOR2X1 exu_U38598(.A(alu_addsub_rs2_data_16), .B(alu_logic_rs1_data_bf1[16]), .Y(exu_n17118));
XOR2X1 exu_U38599(.A(exu_n15645), .B(exu_n17118), .Y(exu_ifu_brpc_e[16]));
XOR2X1 exu_U38600(.A(alu_addsub_rs2_data_17), .B(alu_logic_rs1_data_bf1[17]), .Y(exu_n17123));
XOR2X1 exu_U38601(.A(exu_n15646), .B(exu_n17123), .Y(exu_ifu_brpc_e[17]));
XOR2X1 exu_U38602(.A(alu_addsub_rs2_data_18), .B(alu_logic_rs1_data_bf1[18]), .Y(exu_n17128));
XOR2X1 exu_U38603(.A(exu_n15647), .B(exu_n17128), .Y(exu_ifu_brpc_e[18]));
XOR2X1 exu_U38604(.A(alu_addsub_rs2_data_19), .B(alu_logic_rs1_data_bf1[19]), .Y(exu_n17133));
XOR2X1 exu_U38605(.A(exu_n15648), .B(exu_n17133), .Y(exu_ifu_brpc_e[19]));
XOR2X1 exu_U38606(.A(alu_addsub_rs2_data_1), .B(alu_logic_rs1_data_bf1[1]), .Y(exu_n17134));
XOR2X1 exu_U38607(.A(exu_n15577), .B(exu_n17134), .Y(exu_ifu_brpc_e[1]));
XOR2X1 exu_U38608(.A(alu_addsub_rs2_data_20), .B(alu_logic_rs1_data_bf1[20]), .Y(exu_n17140));
XOR2X1 exu_U38609(.A(exu_n15649), .B(exu_n17140), .Y(exu_ifu_brpc_e[20]));
XOR2X1 exu_U38610(.A(alu_addsub_rs2_data_21), .B(alu_logic_rs1_data_bf1[21]), .Y(exu_n17145));
XOR2X1 exu_U38611(.A(exu_n15650), .B(exu_n17145), .Y(exu_ifu_brpc_e[21]));
XOR2X1 exu_U38612(.A(alu_addsub_rs2_data_22), .B(alu_logic_rs1_data_bf1[22]), .Y(exu_n17150));
XOR2X1 exu_U38613(.A(exu_n15651), .B(exu_n17150), .Y(exu_ifu_brpc_e[22]));
XOR2X1 exu_U38614(.A(alu_addsub_rs2_data_23), .B(alu_logic_rs1_data_bf1[23]), .Y(exu_n17155));
XOR2X1 exu_U38615(.A(exu_n15652), .B(exu_n17155), .Y(exu_ifu_brpc_e[23]));
XOR2X1 exu_U38616(.A(alu_addsub_rs2_data_24), .B(alu_logic_rs1_data_bf1[24]), .Y(exu_n17160));
XOR2X1 exu_U38617(.A(exu_n15653), .B(exu_n17160), .Y(exu_ifu_brpc_e[24]));
XOR2X1 exu_U38618(.A(alu_addsub_rs2_data_25), .B(alu_logic_rs1_data_bf1[25]), .Y(exu_n17165));
XOR2X1 exu_U38619(.A(exu_n15654), .B(exu_n17165), .Y(exu_ifu_brpc_e[25]));
XOR2X1 exu_U38620(.A(alu_addsub_rs2_data_26), .B(alu_logic_rs1_data_bf1[26]), .Y(exu_n17170));
XOR2X1 exu_U38621(.A(exu_n15655), .B(exu_n17170), .Y(exu_ifu_brpc_e[26]));
XOR2X1 exu_U38622(.A(alu_addsub_rs2_data_27), .B(alu_logic_rs1_data_bf1[27]), .Y(exu_n17175));
XOR2X1 exu_U38623(.A(exu_n15656), .B(exu_n17175), .Y(exu_ifu_brpc_e[27]));
XOR2X1 exu_U38624(.A(alu_addsub_rs2_data_28), .B(alu_logic_rs1_data_bf1[28]), .Y(exu_n17180));
XOR2X1 exu_U38625(.A(exu_n15657), .B(exu_n17180), .Y(exu_ifu_brpc_e[28]));
XOR2X1 exu_U38626(.A(alu_addsub_rs2_data_29), .B(alu_logic_rs1_data_bf1[29]), .Y(exu_n17185));
XOR2X1 exu_U38627(.A(exu_n15658), .B(exu_n17185), .Y(exu_ifu_brpc_e[29]));
XOR2X1 exu_U38628(.A(alu_addsub_rs2_data_2), .B(alu_logic_rs1_data_bf1[2]), .Y(exu_n17186));
XOR2X1 exu_U38629(.A(exu_n15578), .B(exu_n17186), .Y(exu_ifu_brpc_e[2]));
XOR2X1 exu_U38630(.A(alu_addsub_rs2_data_30), .B(alu_logic_rs1_data_bf1[30]), .Y(exu_n17192));
XOR2X1 exu_U38631(.A(exu_n15659), .B(exu_n17192), .Y(exu_ifu_brpc_e[30]));
XOR2X1 exu_U38632(.A(alu_ecl_adderin2_31_e), .B(alu_logic_rs1_data_bf1[31]), .Y(exu_n17197));
XOR2X1 exu_U38633(.A(exu_n15660), .B(exu_n17197), .Y(exu_ifu_brpc_e[31]));
XOR2X1 exu_U38634(.A(alu_addsub_rs2_data_3), .B(alu_logic_rs1_data_bf1[3]), .Y(exu_n17202));
XOR2X1 exu_U38635(.A(exu_n15579), .B(exu_n17202), .Y(exu_ifu_brpc_e[3]));
XOR2X1 exu_U38636(.A(alu_addsub_rs2_data_4), .B(alu_logic_rs1_data_bf1[4]), .Y(exu_n17204));
XOR2X1 exu_U38637(.A(exu_n15580), .B(exu_n17204), .Y(exu_ifu_brpc_e[4]));
XOR2X1 exu_U38638(.A(alu_addsub_rs2_data_5), .B(alu_logic_rs1_data_bf1[5]), .Y(exu_n17206));
XOR2X1 exu_U38639(.A(exu_n15581), .B(exu_n17206), .Y(exu_ifu_brpc_e[5]));
XOR2X1 exu_U38640(.A(alu_addsub_rs2_data_6), .B(alu_logic_rs1_data_bf1[6]), .Y(exu_n17208));
XOR2X1 exu_U38641(.A(exu_n15582), .B(exu_n17208), .Y(exu_ifu_brpc_e[6]));
XOR2X1 exu_U38642(.A(alu_addsub_rs2_data_7), .B(alu_logic_rs1_data_bf1[7]), .Y(exu_n17210));
XOR2X1 exu_U38643(.A(exu_n15583), .B(exu_n17210), .Y(exu_ifu_brpc_e[7]));
XOR2X1 exu_U38644(.A(alu_addsub_rs2_data_8), .B(alu_logic_rs1_data_bf1[8]), .Y(exu_n17212));
XOR2X1 exu_U38645(.A(exu_n15584), .B(exu_n17212), .Y(exu_ifu_brpc_e[8]));
XOR2X1 exu_U38646(.A(alu_addsub_rs2_data_9), .B(alu_logic_rs1_data_bf1[9]), .Y(exu_n17214));
XOR2X1 exu_U38647(.A(exu_n15585), .B(exu_n17214), .Y(exu_ifu_brpc_e[9]));
XOR2X1 exu_U38648(.A(exu_n15795), .B(alu_addsub_rs2_data[32]), .Y(exu_n17216));
XOR2X1 exu_U38649(.A(alu_logic_rs1_data_bf1[32]), .B(exu_n17216), .Y(exu_ifu_brpc_e[32]));
XOR2X1 exu_U38650(.A(alu_addsub_rs2_data[42]), .B(alu_logic_rs1_data_bf1[42]), .Y(exu_n17247));
XOR2X1 exu_U38651(.A(exu_n15661), .B(exu_n17247), .Y(exu_ifu_brpc_e[42]));
XOR2X1 exu_U38652(.A(alu_addsub_rs2_data[43]), .B(alu_logic_rs1_data_bf1[43]), .Y(exu_n17252));
XOR2X1 exu_U38653(.A(exu_n15662), .B(exu_n17252), .Y(exu_ifu_brpc_e[43]));
XOR2X1 exu_U38654(.A(alu_addsub_rs2_data[44]), .B(alu_logic_rs1_data_bf1[44]), .Y(exu_n17257));
XOR2X1 exu_U38655(.A(exu_n15663), .B(exu_n17257), .Y(exu_ifu_brpc_e[44]));
XOR2X1 exu_U38656(.A(alu_addsub_rs2_data[45]), .B(alu_logic_rs1_data_bf1[45]), .Y(exu_n17262));
XOR2X1 exu_U38657(.A(exu_n15664), .B(exu_n17262), .Y(exu_ifu_brpc_e[45]));
XOR2X1 exu_U38658(.A(alu_addsub_rs2_data[46]), .B(alu_logic_rs1_data_bf1[46]), .Y(exu_n17267));
XOR2X1 exu_U38659(.A(exu_n15665), .B(exu_n17267), .Y(exu_ifu_brpc_e[46]));
XOR2X1 exu_U38660(.A(alu_addsub_rs2_data[47]), .B(alu_logic_rs1_data_bf1[47]), .Y(exu_n17272));
XOR2X1 exu_U38661(.A(exu_n15666), .B(exu_n17272), .Y(exu_ifu_brpc_e[47]));
XOR2X1 exu_U38662(.A(alu_addsub_rs2_data[48]), .B(alu_logic_rs1_data_bf1[48]), .Y(exu_n17277));
XOR2X1 exu_U38663(.A(exu_n15667), .B(exu_n17277), .Y(alu_adder_out[48]));
XOR2X1 exu_U38664(.A(alu_addsub_rs2_data[49]), .B(alu_logic_rs1_data_bf1[49]), .Y(exu_n17282));
XOR2X1 exu_U38665(.A(exu_n15668), .B(exu_n17282), .Y(alu_adder_out[49]));
XOR2X1 exu_U38666(.A(alu_addsub_rs2_data[50]), .B(alu_logic_rs1_data_bf1[50]), .Y(exu_n17287));
XOR2X1 exu_U38667(.A(exu_n15669), .B(exu_n17287), .Y(alu_adder_out[50]));
XOR2X1 exu_U38668(.A(alu_addsub_rs2_data[51]), .B(alu_logic_rs1_data_bf1[51]), .Y(exu_n17292));
XOR2X1 exu_U38669(.A(exu_n15670), .B(exu_n17292), .Y(alu_adder_out[51]));
XOR2X1 exu_U38670(.A(alu_addsub_rs2_data[33]), .B(alu_logic_rs1_data_bf1[33]), .Y(exu_n17293));
XOR2X1 exu_U38671(.A(exu_n15586), .B(exu_n17293), .Y(exu_ifu_brpc_e[33]));
XOR2X1 exu_U38672(.A(alu_addsub_rs2_data[52]), .B(alu_logic_rs1_data_bf1[52]), .Y(exu_n17299));
XOR2X1 exu_U38673(.A(exu_n15671), .B(exu_n17299), .Y(alu_adder_out[52]));
XOR2X1 exu_U38674(.A(alu_addsub_rs2_data[53]), .B(alu_logic_rs1_data_bf1[53]), .Y(exu_n17304));
XOR2X1 exu_U38675(.A(exu_n15672), .B(exu_n17304), .Y(alu_adder_out[53]));
XOR2X1 exu_U38676(.A(alu_addsub_rs2_data[54]), .B(alu_logic_rs1_data_bf1[54]), .Y(exu_n17309));
XOR2X1 exu_U38677(.A(exu_n15673), .B(exu_n17309), .Y(alu_adder_out[54]));
XOR2X1 exu_U38678(.A(alu_addsub_rs2_data[55]), .B(alu_logic_rs1_data_bf1[55]), .Y(exu_n17314));
XOR2X1 exu_U38679(.A(exu_n15674), .B(exu_n17314), .Y(alu_adder_out[55]));
XOR2X1 exu_U38680(.A(alu_addsub_rs2_data[56]), .B(alu_logic_rs1_data_bf1[56]), .Y(exu_n17319));
XOR2X1 exu_U38681(.A(exu_n15675), .B(exu_n17319), .Y(alu_adder_out[56]));
XOR2X1 exu_U38682(.A(alu_addsub_rs2_data[57]), .B(alu_logic_rs1_data_bf1[57]), .Y(exu_n17324));
XOR2X1 exu_U38683(.A(exu_n15676), .B(exu_n17324), .Y(alu_adder_out[57]));
XOR2X1 exu_U38684(.A(alu_addsub_rs2_data[58]), .B(alu_logic_rs1_data_bf1[58]), .Y(exu_n17329));
XOR2X1 exu_U38685(.A(exu_n15677), .B(exu_n17329), .Y(alu_adder_out[58]));
XOR2X1 exu_U38686(.A(alu_addsub_rs2_data[59]), .B(alu_logic_rs1_data_bf1[59]), .Y(exu_n17334));
XOR2X1 exu_U38687(.A(exu_n15678), .B(exu_n17334), .Y(alu_adder_out[59]));
XOR2X1 exu_U38688(.A(alu_addsub_rs2_data[60]), .B(alu_logic_rs1_data_bf1[60]), .Y(exu_n17339));
XOR2X1 exu_U38689(.A(exu_n15679), .B(exu_n17339), .Y(alu_adder_out[60]));
XOR2X1 exu_U38690(.A(alu_addsub_rs2_data[61]), .B(alu_logic_rs1_data_bf1[61]), .Y(exu_n17344));
XOR2X1 exu_U38691(.A(exu_n15680), .B(exu_n17344), .Y(alu_adder_out[61]));
XOR2X1 exu_U38692(.A(alu_addsub_rs2_data[34]), .B(alu_logic_rs1_data_bf1[34]), .Y(exu_n17345));
XOR2X1 exu_U38693(.A(exu_n15587), .B(exu_n17345), .Y(exu_ifu_brpc_e[34]));
XOR2X1 exu_U38694(.A(alu_addsub_rs2_data[62]), .B(alu_logic_rs1_data_bf1[62]), .Y(exu_n17351));
XOR2X1 exu_U38695(.A(exu_n15681), .B(exu_n17351), .Y(alu_adder_out[62]));
XOR2X1 exu_U38696(.A(alu_ecl_adderin2_63_e), .B(alu_logic_rs1_data_bf1[63]), .Y(exu_n17356));
XOR2X1 exu_U38697(.A(exu_n15682), .B(exu_n17356), .Y(alu_ecl_add_n64_e));
XOR2X1 exu_U38698(.A(alu_addsub_rs2_data[35]), .B(alu_logic_rs1_data_bf1[35]), .Y(exu_n17361));
XOR2X1 exu_U38699(.A(exu_n15588), .B(exu_n17361), .Y(exu_ifu_brpc_e[35]));
XOR2X1 exu_U38700(.A(alu_addsub_rs2_data[36]), .B(alu_logic_rs1_data_bf1[36]), .Y(exu_n17363));
XOR2X1 exu_U38701(.A(exu_n15589), .B(exu_n17363), .Y(exu_ifu_brpc_e[36]));
XOR2X1 exu_U38702(.A(alu_addsub_rs2_data[37]), .B(alu_logic_rs1_data_bf1[37]), .Y(exu_n17365));
XOR2X1 exu_U38703(.A(exu_n15590), .B(exu_n17365), .Y(exu_ifu_brpc_e[37]));
XOR2X1 exu_U38704(.A(alu_addsub_rs2_data[38]), .B(alu_logic_rs1_data_bf1[38]), .Y(exu_n17367));
XOR2X1 exu_U38705(.A(exu_n15591), .B(exu_n17367), .Y(exu_ifu_brpc_e[38]));
XOR2X1 exu_U38706(.A(alu_addsub_rs2_data[39]), .B(alu_logic_rs1_data_bf1[39]), .Y(exu_n17369));
XOR2X1 exu_U38707(.A(exu_n15592), .B(exu_n17369), .Y(exu_ifu_brpc_e[39]));
XOR2X1 exu_U38708(.A(alu_addsub_rs2_data[40]), .B(alu_logic_rs1_data_bf1[40]), .Y(exu_n17371));
XOR2X1 exu_U38709(.A(exu_n15593), .B(exu_n17371), .Y(exu_ifu_brpc_e[40]));
XOR2X1 exu_U38710(.A(alu_addsub_rs2_data[41]), .B(alu_logic_rs1_data_bf1[41]), .Y(exu_n17373));
XOR2X1 exu_U38711(.A(exu_n15594), .B(exu_n17373), .Y(exu_ifu_brpc_e[41]));
XNOR2X1 exu_U38712(.A(ecl_wb_byplog_rd_g2[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17375));
XNOR2X1 exu_U38713(.A(ecl_wb_byplog_rd_g2[1]), .B(ecl_ifu_exu_rs3_d[1]), .Y(exu_n17376));
XNOR2X1 exu_U38714(.A(ecl_wb_byplog_rd_g2[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17379));
XNOR2X1 exu_U38715(.A(ecl_wb_byplog_rd_g2[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17378));
XNOR2X1 exu_U38716(.A(ecl_ld_rd_g[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17382));
XNOR2X1 exu_U38717(.A(ecl_ld_rd_g[1]), .B(ecl_ifu_exu_rs3_d[1]), .Y(exu_n17383));
XNOR2X1 exu_U38718(.A(ecl_ld_rd_g[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17386));
XNOR2X1 exu_U38719(.A(ecl_ld_rd_g[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17385));
XNOR2X1 exu_U38720(.A(ecl_rd_m[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17389));
XNOR2X1 exu_U38721(.A(ecl_rd_m[1]), .B(ecl_ifu_exu_rs3_d[1]), .Y(exu_n17390));
XNOR2X1 exu_U38722(.A(ecl_rd_m[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17393));
XNOR2X1 exu_U38723(.A(ecl_rd_m[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17392));
XNOR2X1 exu_U38724(.A(ecl_rd_e[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17396));
XNOR2X1 exu_U38725(.A(ecl_rd_e[1]), .B(ecl_ifu_exu_rs3_d[1]), .Y(exu_n17397));
XNOR2X1 exu_U38726(.A(ecl_rd_e[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17400));
XNOR2X1 exu_U38727(.A(ecl_rd_e[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17399));
XNOR2X1 exu_U38728(.A(ecl_wb_byplog_rd_g2[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17411));
XNOR2X1 exu_U38729(.A(ecl_wb_byplog_rd_g2[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17414));
XNOR2X1 exu_U38730(.A(ecl_wb_byplog_rd_g2[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17413));
XNOR2X1 exu_U38731(.A(ecl_ld_rd_g[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17425));
XNOR2X1 exu_U38732(.A(ecl_ld_rd_g[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17428));
XNOR2X1 exu_U38733(.A(ecl_ld_rd_g[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17427));
XNOR2X1 exu_U38734(.A(ecl_rd_m[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17439));
XNOR2X1 exu_U38735(.A(ecl_rd_m[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17442));
XNOR2X1 exu_U38736(.A(ecl_rd_m[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17441));
XNOR2X1 exu_U38737(.A(ecl_rd_e[2]), .B(ecl_ifu_exu_rs3_d[2]), .Y(exu_n17453));
XNOR2X1 exu_U38738(.A(ecl_rd_e[4]), .B(ecl_ifu_exu_rs3_d[4]), .Y(exu_n17456));
XNOR2X1 exu_U38739(.A(ecl_rd_e[3]), .B(ecl_ifu_exu_rs3_d[3]), .Y(exu_n17455));


DFFNEGX1 irf_rst_tri_en_neg_reg(.D(mem_write_disable), .CLK(rclk), .Q(irf_rst_tri_en_neg));

  bw_r_irf irf ( .so(short_scan0_1), .si(short_si0), .reset_l(arst_l), 
        .rst_tri_en(mem_write_disable), .rml_irf_old_e_cwp_e(
        rml_irf_old_e_cwp_e), .rml_irf_new_e_cwp_e(rml_irf_new_e_cwp_e), 
        .irf_byp_rs1_data_d_l(irf_byp_rs1_data_d_l), .irf_byp_rs2_data_d_l(
        irf_byp_rs2_data_d_l), .irf_byp_rs3_data_d_l(irf_byp_rs3_data_d_l), 
        .irf_byp_rs3h_data_d_l(irf_byp_rs3h_data_d_l), .rclk(rclk), .se(se), 
        .sehold(sehold), .ifu_exu_tid_s2(ifu_exu_tid_s2), .ifu_exu_rs1_s(
        ifu_exu_rs1_s), .ifu_exu_rs2_s(ifu_exu_rs2_s), .ifu_exu_rs3_s(
        ifu_exu_rs3_s), .ifu_exu_ren1_s(ifu_exu_ren1_s), .ifu_exu_ren2_s(
        ifu_exu_ren2_s), .ifu_exu_ren3_s(ifu_exu_ren3_s), .ecl_irf_wen_w(
        ecl_irf_wen_w), .ecl_irf_wen_w2(ecl_wb_byplog_wen_w2 ), 
        .ecl_irf_rd_m(ecl_irf_rd_m), .ecl_irf_rd_g(ecl_irf_rd_g), 
        .byp_irf_rd_data_w(byp_irf_rd_data_w), .byp_irf_rd_data_w2(
        byp_irf_rd_data_w2), .ecl_irf_tid_m(ecl_irf_tid_m), .ecl_irf_tid_g(
        ecl_irf_tid_g), .rml_irf_old_lo_cwp_e(rml_irf_old_lo_cwp_e), 
        .rml_irf_new_lo_cwp_e(rml_irf_new_lo_cwp_e), .rml_irf_swap_even_e(
        rml_irf_swap_even_e), .rml_irf_swap_odd_e(rml_irf_swap_odd_e), 
        .rml_irf_swap_local_e(rml_irf_swap_local_e), .rml_irf_kill_restore_w(
        rml_irf_kill_restore_w), .rml_irf_cwpswap_tid_e(rml_irf_cwpswap_tid_e), 
        .rml_irf_old_agp(rml_irf_old_agp), .rml_irf_new_agp(tlu_exu_agp), 
        .rml_irf_swap_global(tlu_exu_agp_swap), .rml_irf_global_tid(
        tlu_exu_agp_tid) );
endmodule
